module top (decrypt_pad, \key1[0]_pad , \key1[10]_pad , \key1[11]_pad , \key1[12]_pad , \key1[13]_pad , \key1[14]_pad , \key1[15]_pad , \key1[16]_pad , \key1[17]_pad , \key1[18]_pad , \key1[19]_pad , \key1[1]_pad , \key1[20]_pad , \key1[21]_pad , \key1[22]_pad , \key1[23]_pad , \key1[24]_pad , \key1[25]_pad , \key1[26]_pad , \key1[27]_pad , \key1[28]_pad , \key1[29]_pad , \key1[2]_pad , \key1[30]_pad , \key1[31]_pad , \key1[32]_pad , \key1[33]_pad , \key1[34]_pad , \key1[35]_pad , \key1[36]_pad , \key1[37]_pad , \key1[38]_pad , \key1[39]_pad , \key1[3]_pad , \key1[40]_pad , \key1[41]_pad , \key1[42]_pad , \key1[43]_pad , \key1[44]_pad , \key1[45]_pad , \key1[46]_pad , \key1[47]_pad , \key1[48]_pad , \key1[49]_pad , \key1[4]_pad , \key1[50]_pad , \key1[51]_pad , \key1[52]_pad , \key1[53]_pad , \key1[54]_pad , \key1[55]_pad , \key1[5]_pad , \key1[6]_pad , \key1[7]_pad , \key1[8]_pad , \key1[9]_pad , \key3[0]_pad , \key3[10]_pad , \key3[11]_pad , \key3[12]_pad , \key3[13]_pad , \key3[14]_pad , \key3[15]_pad , \key3[16]_pad , \key3[17]_pad , \key3[18]_pad , \key3[19]_pad , \key3[1]_pad , \key3[20]_pad , \key3[21]_pad , \key3[22]_pad , \key3[23]_pad , \key3[24]_pad , \key3[25]_pad , \key3[26]_pad , \key3[27]_pad , \key3[28]_pad , \key3[29]_pad , \key3[2]_pad , \key3[30]_pad , \key3[31]_pad , \key3[32]_pad , \key3[33]_pad , \key3[34]_pad , \key3[35]_pad , \key3[36]_pad , \key3[37]_pad , \key3[38]_pad , \key3[39]_pad , \key3[3]_pad , \key3[40]_pad , \key3[41]_pad , \key3[42]_pad , \key3[43]_pad , \key3[44]_pad , \key3[45]_pad , \key3[46]_pad , \key3[47]_pad , \key3[48]_pad , \key3[49]_pad , \key3[4]_pad , \key3[50]_pad , \key3[51]_pad , \key3[52]_pad , \key3[53]_pad , \key3[54]_pad , \key3[55]_pad , \key3[5]_pad , \key3[6]_pad , \key3[7]_pad , \key3[8]_pad , \key3[9]_pad , \u0_L0_reg[10]/NET0131 , \u0_L0_reg[11]/NET0131 , \u0_L0_reg[12]/NET0131 , \u0_L0_reg[13]/NET0131 , \u0_L0_reg[14]/NET0131 , \u0_L0_reg[15]/P0001 , \u0_L0_reg[16]/NET0131 , \u0_L0_reg[17]/NET0131 , \u0_L0_reg[18]/NET0131 , \u0_L0_reg[19]/P0001 , \u0_L0_reg[1]/NET0131 , \u0_L0_reg[20]/NET0131 , \u0_L0_reg[21]/NET0131 , \u0_L0_reg[22]/NET0131 , \u0_L0_reg[23]/NET0131 , \u0_L0_reg[24]/NET0131 , \u0_L0_reg[25]/NET0131 , \u0_L0_reg[26]/NET0131 , \u0_L0_reg[27]/NET0131 , \u0_L0_reg[28]/NET0131 , \u0_L0_reg[29]/NET0131 , \u0_L0_reg[2]/NET0131 , \u0_L0_reg[30]/P0001 , \u0_L0_reg[31]/NET0131 , \u0_L0_reg[32]/NET0131 , \u0_L0_reg[3]/NET0131 , \u0_L0_reg[4]/NET0131 , \u0_L0_reg[5]/NET0131 , \u0_L0_reg[6]/NET0131 , \u0_L0_reg[7]/NET0131 , \u0_L0_reg[8]/NET0131 , \u0_L0_reg[9]/NET0131 , \u0_L10_reg[10]/NET0131 , \u0_L10_reg[11]/NET0131 , \u0_L10_reg[12]/NET0131 , \u0_L10_reg[13]/NET0131 , \u0_L10_reg[14]/NET0131 , \u0_L10_reg[15]/P0001 , \u0_L10_reg[16]/NET0131 , \u0_L10_reg[17]/NET0131 , \u0_L10_reg[18]/NET0131 , \u0_L10_reg[19]/NET0131 , \u0_L10_reg[1]/NET0131 , \u0_L10_reg[20]/NET0131 , \u0_L10_reg[21]/NET0131 , \u0_L10_reg[22]/NET0131 , \u0_L10_reg[23]/NET0131 , \u0_L10_reg[24]/NET0131 , \u0_L10_reg[25]/NET0131 , \u0_L10_reg[26]/NET0131 , \u0_L10_reg[27]/NET0131 , \u0_L10_reg[28]/NET0131 , \u0_L10_reg[29]/NET0131 , \u0_L10_reg[2]/NET0131 , \u0_L10_reg[30]/NET0131 , \u0_L10_reg[31]/NET0131 , \u0_L10_reg[32]/NET0131 , \u0_L10_reg[3]/NET0131 , \u0_L10_reg[4]/NET0131 , \u0_L10_reg[5]/NET0131 , \u0_L10_reg[6]/NET0131 , \u0_L10_reg[7]/NET0131 , \u0_L10_reg[8]/NET0131 , \u0_L10_reg[9]/NET0131 , \u0_L11_reg[10]/NET0131 , \u0_L11_reg[11]/P0001 , \u0_L11_reg[12]/NET0131 , \u0_L11_reg[13]/NET0131 , \u0_L11_reg[14]/NET0131 , \u0_L11_reg[15]/P0001 , \u0_L11_reg[16]/NET0131 , \u0_L11_reg[17]/NET0131 , \u0_L11_reg[18]/NET0131 , \u0_L11_reg[19]/NET0131 , \u0_L11_reg[1]/NET0131 , \u0_L11_reg[20]/NET0131 , \u0_L11_reg[21]/NET0131 , \u0_L11_reg[22]/NET0131 , \u0_L11_reg[23]/NET0131 , \u0_L11_reg[24]/NET0131 , \u0_L11_reg[25]/NET0131 , \u0_L11_reg[26]/NET0131 , \u0_L11_reg[27]/NET0131 , \u0_L11_reg[28]/NET0131 , \u0_L11_reg[29]/NET0131 , \u0_L11_reg[2]/NET0131 , \u0_L11_reg[30]/NET0131 , \u0_L11_reg[31]/NET0131 , \u0_L11_reg[32]/NET0131 , \u0_L11_reg[3]/NET0131 , \u0_L11_reg[4]/NET0131 , \u0_L11_reg[5]/NET0131 , \u0_L11_reg[6]/NET0131 , \u0_L11_reg[7]/NET0131 , \u0_L11_reg[8]/NET0131 , \u0_L11_reg[9]/NET0131 , \u0_L12_reg[10]/NET0131 , \u0_L12_reg[11]/NET0131 , \u0_L12_reg[12]/NET0131 , \u0_L12_reg[13]/NET0131 , \u0_L12_reg[14]/NET0131 , \u0_L12_reg[15]/P0001 , \u0_L12_reg[16]/NET0131 , \u0_L12_reg[17]/NET0131 , \u0_L12_reg[18]/NET0131 , \u0_L12_reg[19]/P0001 , \u0_L12_reg[1]/NET0131 , \u0_L12_reg[20]/NET0131 , \u0_L12_reg[21]/NET0131 , \u0_L12_reg[22]/NET0131 , \u0_L12_reg[23]/NET0131 , \u0_L12_reg[24]/NET0131 , \u0_L12_reg[25]/NET0131 , \u0_L12_reg[26]/NET0131 , \u0_L12_reg[27]/NET0131 , \u0_L12_reg[28]/NET0131 , \u0_L12_reg[29]/NET0131 , \u0_L12_reg[2]/NET0131 , \u0_L12_reg[30]/NET0131 , \u0_L12_reg[31]/NET0131 , \u0_L12_reg[32]/NET0131 , \u0_L12_reg[3]/NET0131 , \u0_L12_reg[4]/NET0131 , \u0_L12_reg[5]/NET0131 , \u0_L12_reg[6]/NET0131 , \u0_L12_reg[7]/NET0131 , \u0_L12_reg[8]/NET0131 , \u0_L12_reg[9]/NET0131 , \u0_L13_reg[10]/NET0131 , \u0_L13_reg[11]/NET0131 , \u0_L13_reg[12]/NET0131 , \u0_L13_reg[13]/NET0131 , \u0_L13_reg[14]/NET0131 , \u0_L13_reg[15]/P0001 , \u0_L13_reg[16]/NET0131 , \u0_L13_reg[17]/NET0131 , \u0_L13_reg[18]/NET0131 , \u0_L13_reg[19]/NET0131 , \u0_L13_reg[1]/NET0131 , \u0_L13_reg[20]/NET0131 , \u0_L13_reg[21]/NET0131 , \u0_L13_reg[22]/NET0131 , \u0_L13_reg[23]/NET0131 , \u0_L13_reg[24]/NET0131 , \u0_L13_reg[25]/NET0131 , \u0_L13_reg[26]/NET0131 , \u0_L13_reg[27]/NET0131 , \u0_L13_reg[28]/NET0131 , \u0_L13_reg[29]/NET0131 , \u0_L13_reg[2]/NET0131 , \u0_L13_reg[30]/NET0131 , \u0_L13_reg[31]/NET0131 , \u0_L13_reg[32]/NET0131 , \u0_L13_reg[3]/NET0131 , \u0_L13_reg[4]/NET0131 , \u0_L13_reg[5]/NET0131 , \u0_L13_reg[6]/NET0131 , \u0_L13_reg[7]/NET0131 , \u0_L13_reg[8]/NET0131 , \u0_L13_reg[9]/NET0131 , \u0_L14_reg[10]/P0001 , \u0_L14_reg[11]/P0001 , \u0_L14_reg[12]/P0001 , \u0_L14_reg[13]/P0001 , \u0_L14_reg[14]/P0001 , \u0_L14_reg[15]/P0001 , \u0_L14_reg[16]/P0001 , \u0_L14_reg[17]/P0001 , \u0_L14_reg[18]/P0001 , \u0_L14_reg[19]/P0001 , \u0_L14_reg[1]/P0001 , \u0_L14_reg[20]/P0001 , \u0_L14_reg[21]/P0001 , \u0_L14_reg[22]/P0001 , \u0_L14_reg[23]/P0001 , \u0_L14_reg[24]/P0001 , \u0_L14_reg[25]/P0001 , \u0_L14_reg[26]/P0001 , \u0_L14_reg[27]/P0001 , \u0_L14_reg[28]/P0001 , \u0_L14_reg[29]/P0001 , \u0_L14_reg[2]/P0001 , \u0_L14_reg[30]/P0001 , \u0_L14_reg[31]/P0001 , \u0_L14_reg[32]/P0001 , \u0_L14_reg[3]/P0001 , \u0_L14_reg[4]/P0001 , \u0_L14_reg[5]/P0001 , \u0_L14_reg[6]/P0001 , \u0_L14_reg[7]/P0001 , \u0_L14_reg[8]/P0001 , \u0_L14_reg[9]/P0001 , \u0_L1_reg[10]/NET0131 , \u0_L1_reg[11]/NET0131 , \u0_L1_reg[12]/NET0131 , \u0_L1_reg[13]/NET0131 , \u0_L1_reg[14]/NET0131 , \u0_L1_reg[15]/P0001 , \u0_L1_reg[16]/NET0131 , \u0_L1_reg[17]/NET0131 , \u0_L1_reg[18]/NET0131 , \u0_L1_reg[19]/NET0131 , \u0_L1_reg[1]/NET0131 , \u0_L1_reg[20]/NET0131 , \u0_L1_reg[21]/NET0131 , \u0_L1_reg[22]/NET0131 , \u0_L1_reg[23]/NET0131 , \u0_L1_reg[24]/NET0131 , \u0_L1_reg[25]/NET0131 , \u0_L1_reg[26]/NET0131 , \u0_L1_reg[27]/NET0131 , \u0_L1_reg[28]/NET0131 , \u0_L1_reg[29]/NET0131 , \u0_L1_reg[2]/NET0131 , \u0_L1_reg[30]/NET0131 , \u0_L1_reg[31]/NET0131 , \u0_L1_reg[32]/NET0131 , \u0_L1_reg[3]/NET0131 , \u0_L1_reg[4]/NET0131 , \u0_L1_reg[5]/NET0131 , \u0_L1_reg[6]/NET0131 , \u0_L1_reg[7]/NET0131 , \u0_L1_reg[8]/NET0131 , \u0_L1_reg[9]/NET0131 , \u0_L2_reg[10]/NET0131 , \u0_L2_reg[11]/NET0131 , \u0_L2_reg[12]/NET0131 , \u0_L2_reg[13]/NET0131 , \u0_L2_reg[14]/NET0131 , \u0_L2_reg[15]/P0001 , \u0_L2_reg[16]/NET0131 , \u0_L2_reg[17]/NET0131 , \u0_L2_reg[18]/NET0131 , \u0_L2_reg[19]/P0001 , \u0_L2_reg[1]/NET0131 , \u0_L2_reg[20]/NET0131 , \u0_L2_reg[21]/NET0131 , \u0_L2_reg[22]/NET0131 , \u0_L2_reg[23]/NET0131 , \u0_L2_reg[24]/NET0131 , \u0_L2_reg[25]/NET0131 , \u0_L2_reg[26]/NET0131 , \u0_L2_reg[27]/NET0131 , \u0_L2_reg[28]/NET0131 , \u0_L2_reg[29]/NET0131 , \u0_L2_reg[2]/NET0131 , \u0_L2_reg[30]/NET0131 , \u0_L2_reg[31]/NET0131 , \u0_L2_reg[32]/NET0131 , \u0_L2_reg[3]/NET0131 , \u0_L2_reg[4]/NET0131 , \u0_L2_reg[5]/NET0131 , \u0_L2_reg[6]/NET0131 , \u0_L2_reg[7]/NET0131 , \u0_L2_reg[8]/NET0131 , \u0_L2_reg[9]/NET0131 , \u0_L3_reg[10]/NET0131 , \u0_L3_reg[11]/NET0131 , \u0_L3_reg[12]/NET0131 , \u0_L3_reg[13]/NET0131 , \u0_L3_reg[14]/NET0131 , \u0_L3_reg[15]/P0001 , \u0_L3_reg[16]/NET0131 , \u0_L3_reg[17]/NET0131 , \u0_L3_reg[18]/NET0131 , \u0_L3_reg[19]/P0001 , \u0_L3_reg[1]/NET0131 , \u0_L3_reg[20]/NET0131 , \u0_L3_reg[21]/NET0131 , \u0_L3_reg[22]/NET0131 , \u0_L3_reg[23]/NET0131 , \u0_L3_reg[24]/NET0131 , \u0_L3_reg[25]/NET0131 , \u0_L3_reg[26]/NET0131 , \u0_L3_reg[27]/NET0131 , \u0_L3_reg[28]/NET0131 , \u0_L3_reg[29]/NET0131 , \u0_L3_reg[2]/NET0131 , \u0_L3_reg[30]/NET0131 , \u0_L3_reg[31]/NET0131 , \u0_L3_reg[32]/NET0131 , \u0_L3_reg[3]/NET0131 , \u0_L3_reg[4]/NET0131 , \u0_L3_reg[5]/NET0131 , \u0_L3_reg[6]/NET0131 , \u0_L3_reg[7]/NET0131 , \u0_L3_reg[8]/NET0131 , \u0_L3_reg[9]/NET0131 , \u0_L4_reg[10]/NET0131 , \u0_L4_reg[11]/NET0131 , \u0_L4_reg[12]/NET0131 , \u0_L4_reg[13]/NET0131 , \u0_L4_reg[14]/NET0131 , \u0_L4_reg[15]/P0001 , \u0_L4_reg[16]/NET0131 , \u0_L4_reg[17]/NET0131 , \u0_L4_reg[18]/NET0131 , \u0_L4_reg[19]/NET0131 , \u0_L4_reg[1]/NET0131 , \u0_L4_reg[20]/NET0131 , \u0_L4_reg[21]/NET0131 , \u0_L4_reg[22]/NET0131 , \u0_L4_reg[23]/NET0131 , \u0_L4_reg[24]/NET0131 , \u0_L4_reg[25]/NET0131 , \u0_L4_reg[26]/NET0131 , \u0_L4_reg[27]/NET0131 , \u0_L4_reg[28]/NET0131 , \u0_L4_reg[29]/NET0131 , \u0_L4_reg[2]/NET0131 , \u0_L4_reg[30]/NET0131 , \u0_L4_reg[31]/NET0131 , \u0_L4_reg[32]/NET0131 , \u0_L4_reg[3]/NET0131 , \u0_L4_reg[4]/NET0131 , \u0_L4_reg[5]/NET0131 , \u0_L4_reg[6]/NET0131 , \u0_L4_reg[7]/NET0131 , \u0_L4_reg[8]/NET0131 , \u0_L4_reg[9]/NET0131 , \u0_L5_reg[10]/NET0131 , \u0_L5_reg[11]/NET0131 , \u0_L5_reg[12]/NET0131 , \u0_L5_reg[13]/NET0131 , \u0_L5_reg[14]/NET0131 , \u0_L5_reg[15]/P0001 , \u0_L5_reg[16]/NET0131 , \u0_L5_reg[17]/NET0131 , \u0_L5_reg[18]/NET0131 , \u0_L5_reg[19]/P0001 , \u0_L5_reg[1]/NET0131 , \u0_L5_reg[20]/NET0131 , \u0_L5_reg[21]/NET0131 , \u0_L5_reg[22]/NET0131 , \u0_L5_reg[23]/NET0131 , \u0_L5_reg[24]/NET0131 , \u0_L5_reg[25]/NET0131 , \u0_L5_reg[26]/NET0131 , \u0_L5_reg[27]/NET0131 , \u0_L5_reg[28]/NET0131 , \u0_L5_reg[29]/NET0131 , \u0_L5_reg[2]/NET0131 , \u0_L5_reg[30]/NET0131 , \u0_L5_reg[31]/NET0131 , \u0_L5_reg[32]/NET0131 , \u0_L5_reg[3]/NET0131 , \u0_L5_reg[4]/NET0131 , \u0_L5_reg[5]/NET0131 , \u0_L5_reg[6]/NET0131 , \u0_L5_reg[7]/NET0131 , \u0_L5_reg[8]/NET0131 , \u0_L5_reg[9]/NET0131 , \u0_L6_reg[10]/NET0131 , \u0_L6_reg[11]/NET0131 , \u0_L6_reg[12]/NET0131 , \u0_L6_reg[13]/NET0131 , \u0_L6_reg[14]/NET0131 , \u0_L6_reg[15]/P0001 , \u0_L6_reg[16]/NET0131 , \u0_L6_reg[17]/NET0131 , \u0_L6_reg[18]/NET0131 , \u0_L6_reg[19]/P0001 , \u0_L6_reg[1]/NET0131 , \u0_L6_reg[20]/NET0131 , \u0_L6_reg[21]/NET0131 , \u0_L6_reg[22]/NET0131 , \u0_L6_reg[23]/NET0131 , \u0_L6_reg[24]/NET0131 , \u0_L6_reg[25]/NET0131 , \u0_L6_reg[26]/NET0131 , \u0_L6_reg[27]/NET0131 , \u0_L6_reg[28]/NET0131 , \u0_L6_reg[29]/NET0131 , \u0_L6_reg[2]/NET0131 , \u0_L6_reg[30]/NET0131 , \u0_L6_reg[31]/NET0131 , \u0_L6_reg[32]/NET0131 , \u0_L6_reg[3]/NET0131 , \u0_L6_reg[4]/NET0131 , \u0_L6_reg[5]/NET0131 , \u0_L6_reg[6]/NET0131 , \u0_L6_reg[7]/NET0131 , \u0_L6_reg[8]/NET0131 , \u0_L6_reg[9]/NET0131 , \u0_L7_reg[10]/NET0131 , \u0_L7_reg[11]/NET0131 , \u0_L7_reg[12]/NET0131 , \u0_L7_reg[13]/NET0131 , \u0_L7_reg[14]/NET0131 , \u0_L7_reg[15]/P0001 , \u0_L7_reg[16]/NET0131 , \u0_L7_reg[17]/NET0131 , \u0_L7_reg[18]/NET0131 , \u0_L7_reg[19]/NET0131 , \u0_L7_reg[1]/NET0131 , \u0_L7_reg[20]/NET0131 , \u0_L7_reg[21]/NET0131 , \u0_L7_reg[22]/NET0131 , \u0_L7_reg[23]/NET0131 , \u0_L7_reg[24]/NET0131 , \u0_L7_reg[25]/NET0131 , \u0_L7_reg[26]/NET0131 , \u0_L7_reg[27]/NET0131 , \u0_L7_reg[28]/NET0131 , \u0_L7_reg[29]/NET0131 , \u0_L7_reg[2]/NET0131 , \u0_L7_reg[30]/NET0131 , \u0_L7_reg[31]/NET0131 , \u0_L7_reg[32]/NET0131 , \u0_L7_reg[3]/NET0131 , \u0_L7_reg[4]/NET0131 , \u0_L7_reg[5]/NET0131 , \u0_L7_reg[6]/NET0131 , \u0_L7_reg[7]/NET0131 , \u0_L7_reg[8]/NET0131 , \u0_L7_reg[9]/NET0131 , \u0_L8_reg[10]/NET0131 , \u0_L8_reg[11]/NET0131 , \u0_L8_reg[12]/NET0131 , \u0_L8_reg[13]/NET0131 , \u0_L8_reg[14]/NET0131 , \u0_L8_reg[15]/P0001 , \u0_L8_reg[16]/NET0131 , \u0_L8_reg[17]/NET0131 , \u0_L8_reg[18]/NET0131 , \u0_L8_reg[19]/NET0131 , \u0_L8_reg[1]/NET0131 , \u0_L8_reg[20]/NET0131 , \u0_L8_reg[21]/NET0131 , \u0_L8_reg[22]/NET0131 , \u0_L8_reg[23]/NET0131 , \u0_L8_reg[24]/NET0131 , \u0_L8_reg[25]/NET0131 , \u0_L8_reg[26]/NET0131 , \u0_L8_reg[27]/NET0131 , \u0_L8_reg[28]/NET0131 , \u0_L8_reg[29]/NET0131 , \u0_L8_reg[2]/NET0131 , \u0_L8_reg[30]/NET0131 , \u0_L8_reg[31]/NET0131 , \u0_L8_reg[32]/NET0131 , \u0_L8_reg[3]/NET0131 , \u0_L8_reg[4]/NET0131 , \u0_L8_reg[5]/NET0131 , \u0_L8_reg[6]/NET0131 , \u0_L8_reg[7]/NET0131 , \u0_L8_reg[8]/NET0131 , \u0_L8_reg[9]/NET0131 , \u0_L9_reg[10]/NET0131 , \u0_L9_reg[11]/NET0131 , \u0_L9_reg[12]/NET0131 , \u0_L9_reg[13]/NET0131 , \u0_L9_reg[14]/NET0131 , \u0_L9_reg[15]/P0001 , \u0_L9_reg[16]/NET0131 , \u0_L9_reg[17]/NET0131 , \u0_L9_reg[18]/NET0131 , \u0_L9_reg[19]/P0001 , \u0_L9_reg[1]/NET0131 , \u0_L9_reg[20]/NET0131 , \u0_L9_reg[21]/NET0131 , \u0_L9_reg[22]/NET0131 , \u0_L9_reg[23]/NET0131 , \u0_L9_reg[24]/NET0131 , \u0_L9_reg[25]/NET0131 , \u0_L9_reg[26]/NET0131 , \u0_L9_reg[27]/NET0131 , \u0_L9_reg[28]/NET0131 , \u0_L9_reg[29]/NET0131 , \u0_L9_reg[2]/NET0131 , \u0_L9_reg[30]/NET0131 , \u0_L9_reg[31]/NET0131 , \u0_L9_reg[32]/NET0131 , \u0_L9_reg[3]/NET0131 , \u0_L9_reg[4]/NET0131 , \u0_L9_reg[5]/NET0131 , \u0_L9_reg[6]/NET0131 , \u0_L9_reg[7]/NET0131 , \u0_L9_reg[8]/NET0131 , \u0_L9_reg[9]/NET0131 , \u0_R0_reg[10]/NET0131 , \u0_R0_reg[11]/NET0131 , \u0_R0_reg[12]/NET0131 , \u0_R0_reg[13]/NET0131 , \u0_R0_reg[14]/NET0131 , \u0_R0_reg[15]/NET0131 , \u0_R0_reg[16]/NET0131 , \u0_R0_reg[17]/NET0131 , \u0_R0_reg[18]/NET0131 , \u0_R0_reg[19]/NET0131 , \u0_R0_reg[1]/NET0131 , \u0_R0_reg[20]/NET0131 , \u0_R0_reg[21]/NET0131 , \u0_R0_reg[22]/NET0131 , \u0_R0_reg[23]/NET0131 , \u0_R0_reg[24]/NET0131 , \u0_R0_reg[25]/NET0131 , \u0_R0_reg[26]/NET0131 , \u0_R0_reg[27]/NET0131 , \u0_R0_reg[28]/NET0131 , \u0_R0_reg[29]/NET0131 , \u0_R0_reg[2]/NET0131 , \u0_R0_reg[30]/NET0131 , \u0_R0_reg[31]/NET0131 , \u0_R0_reg[32]/NET0131 , \u0_R0_reg[3]/NET0131 , \u0_R0_reg[4]/NET0131 , \u0_R0_reg[5]/NET0131 , \u0_R0_reg[6]/NET0131 , \u0_R0_reg[7]/NET0131 , \u0_R0_reg[8]/NET0131 , \u0_R0_reg[9]/NET0131 , \u0_R10_reg[10]/NET0131 , \u0_R10_reg[11]/NET0131 , \u0_R10_reg[12]/NET0131 , \u0_R10_reg[13]/NET0131 , \u0_R10_reg[14]/NET0131 , \u0_R10_reg[15]/NET0131 , \u0_R10_reg[16]/NET0131 , \u0_R10_reg[17]/NET0131 , \u0_R10_reg[18]/NET0131 , \u0_R10_reg[19]/NET0131 , \u0_R10_reg[1]/NET0131 , \u0_R10_reg[20]/NET0131 , \u0_R10_reg[21]/NET0131 , \u0_R10_reg[22]/NET0131 , \u0_R10_reg[23]/NET0131 , \u0_R10_reg[24]/NET0131 , \u0_R10_reg[25]/NET0131 , \u0_R10_reg[26]/NET0131 , \u0_R10_reg[27]/NET0131 , \u0_R10_reg[28]/NET0131 , \u0_R10_reg[29]/NET0131 , \u0_R10_reg[2]/NET0131 , \u0_R10_reg[30]/NET0131 , \u0_R10_reg[31]/P0001 , \u0_R10_reg[32]/NET0131 , \u0_R10_reg[3]/NET0131 , \u0_R10_reg[4]/NET0131 , \u0_R10_reg[5]/NET0131 , \u0_R10_reg[6]/NET0131 , \u0_R10_reg[7]/NET0131 , \u0_R10_reg[8]/NET0131 , \u0_R10_reg[9]/NET0131 , \u0_R11_reg[10]/NET0131 , \u0_R11_reg[11]/P0001 , \u0_R11_reg[12]/NET0131 , \u0_R11_reg[13]/NET0131 , \u0_R11_reg[14]/NET0131 , \u0_R11_reg[15]/NET0131 , \u0_R11_reg[16]/NET0131 , \u0_R11_reg[17]/NET0131 , \u0_R11_reg[18]/NET0131 , \u0_R11_reg[19]/NET0131 , \u0_R11_reg[1]/NET0131 , \u0_R11_reg[20]/NET0131 , \u0_R11_reg[21]/NET0131 , \u0_R11_reg[22]/NET0131 , \u0_R11_reg[23]/NET0131 , \u0_R11_reg[24]/NET0131 , \u0_R11_reg[25]/NET0131 , \u0_R11_reg[26]/NET0131 , \u0_R11_reg[27]/NET0131 , \u0_R11_reg[28]/NET0131 , \u0_R11_reg[29]/NET0131 , \u0_R11_reg[2]/NET0131 , \u0_R11_reg[30]/NET0131 , \u0_R11_reg[31]/P0001 , \u0_R11_reg[32]/NET0131 , \u0_R11_reg[3]/NET0131 , \u0_R11_reg[4]/NET0131 , \u0_R11_reg[5]/NET0131 , \u0_R11_reg[6]/NET0131 , \u0_R11_reg[7]/NET0131 , \u0_R11_reg[8]/NET0131 , \u0_R11_reg[9]/NET0131 , \u0_R12_reg[10]/NET0131 , \u0_R12_reg[11]/NET0131 , \u0_R12_reg[12]/NET0131 , \u0_R12_reg[13]/NET0131 , \u0_R12_reg[14]/NET0131 , \u0_R12_reg[15]/NET0131 , \u0_R12_reg[16]/NET0131 , \u0_R12_reg[17]/NET0131 , \u0_R12_reg[18]/NET0131 , \u0_R12_reg[19]/NET0131 , \u0_R12_reg[1]/NET0131 , \u0_R12_reg[20]/NET0131 , \u0_R12_reg[21]/NET0131 , \u0_R12_reg[22]/NET0131 , \u0_R12_reg[23]/NET0131 , \u0_R12_reg[24]/NET0131 , \u0_R12_reg[25]/NET0131 , \u0_R12_reg[26]/NET0131 , \u0_R12_reg[27]/NET0131 , \u0_R12_reg[28]/NET0131 , \u0_R12_reg[29]/NET0131 , \u0_R12_reg[2]/NET0131 , \u0_R12_reg[30]/NET0131 , \u0_R12_reg[31]/P0001 , \u0_R12_reg[32]/NET0131 , \u0_R12_reg[3]/NET0131 , \u0_R12_reg[4]/NET0131 , \u0_R12_reg[5]/NET0131 , \u0_R12_reg[6]/NET0131 , \u0_R12_reg[7]/NET0131 , \u0_R12_reg[8]/NET0131 , \u0_R12_reg[9]/NET0131 , \u0_R13_reg[10]/NET0131 , \u0_R13_reg[11]/NET0131 , \u0_R13_reg[12]/NET0131 , \u0_R13_reg[13]/NET0131 , \u0_R13_reg[14]/NET0131 , \u0_R13_reg[15]/NET0131 , \u0_R13_reg[16]/NET0131 , \u0_R13_reg[17]/NET0131 , \u0_R13_reg[18]/NET0131 , \u0_R13_reg[19]/NET0131 , \u0_R13_reg[1]/NET0131 , \u0_R13_reg[20]/NET0131 , \u0_R13_reg[21]/NET0131 , \u0_R13_reg[22]/P0001 , \u0_R13_reg[23]/NET0131 , \u0_R13_reg[24]/NET0131 , \u0_R13_reg[25]/NET0131 , \u0_R13_reg[26]/NET0131 , \u0_R13_reg[27]/P0001 , \u0_R13_reg[28]/NET0131 , \u0_R13_reg[29]/NET0131 , \u0_R13_reg[2]/NET0131 , \u0_R13_reg[30]/NET0131 , \u0_R13_reg[31]/NET0131 , \u0_R13_reg[32]/NET0131 , \u0_R13_reg[3]/NET0131 , \u0_R13_reg[4]/NET0131 , \u0_R13_reg[5]/NET0131 , \u0_R13_reg[6]/NET0131 , \u0_R13_reg[7]/NET0131 , \u0_R13_reg[8]/NET0131 , \u0_R13_reg[9]/NET0131 , \u0_R14_reg[10]/NET0131 , \u0_R14_reg[11]/P0001 , \u0_R14_reg[12]/NET0131 , \u0_R14_reg[13]/NET0131 , \u0_R14_reg[14]/NET0131 , \u0_R14_reg[15]/NET0131 , \u0_R14_reg[16]/NET0131 , \u0_R14_reg[17]/NET0131 , \u0_R14_reg[18]/NET0131 , \u0_R14_reg[19]/NET0131 , \u0_R14_reg[1]/NET0131 , \u0_R14_reg[20]/NET0131 , \u0_R14_reg[21]/NET0131 , \u0_R14_reg[22]/P0001 , \u0_R14_reg[23]/NET0131 , \u0_R14_reg[24]/NET0131 , \u0_R14_reg[25]/NET0131 , \u0_R14_reg[26]/P0001 , \u0_R14_reg[27]/P0001 , \u0_R14_reg[28]/NET0131 , \u0_R14_reg[29]/NET0131 , \u0_R14_reg[2]/NET0131 , \u0_R14_reg[30]/NET0131 , \u0_R14_reg[31]/P0001 , \u0_R14_reg[32]/NET0131 , \u0_R14_reg[3]/NET0131 , \u0_R14_reg[4]/NET0131 , \u0_R14_reg[5]/NET0131 , \u0_R14_reg[6]/NET0131 , \u0_R14_reg[7]/NET0131 , \u0_R14_reg[8]/NET0131 , \u0_R14_reg[9]/NET0131 , \u0_R1_reg[10]/NET0131 , \u0_R1_reg[11]/NET0131 , \u0_R1_reg[12]/NET0131 , \u0_R1_reg[13]/NET0131 , \u0_R1_reg[14]/NET0131 , \u0_R1_reg[15]/NET0131 , \u0_R1_reg[16]/NET0131 , \u0_R1_reg[17]/NET0131 , \u0_R1_reg[18]/NET0131 , \u0_R1_reg[19]/NET0131 , \u0_R1_reg[1]/NET0131 , \u0_R1_reg[20]/NET0131 , \u0_R1_reg[21]/NET0131 , \u0_R1_reg[22]/NET0131 , \u0_R1_reg[23]/NET0131 , \u0_R1_reg[24]/NET0131 , \u0_R1_reg[25]/NET0131 , \u0_R1_reg[26]/NET0131 , \u0_R1_reg[27]/NET0131 , \u0_R1_reg[28]/NET0131 , \u0_R1_reg[29]/NET0131 , \u0_R1_reg[2]/NET0131 , \u0_R1_reg[30]/NET0131 , \u0_R1_reg[31]/NET0131 , \u0_R1_reg[32]/NET0131 , \u0_R1_reg[3]/NET0131 , \u0_R1_reg[4]/NET0131 , \u0_R1_reg[5]/NET0131 , \u0_R1_reg[6]/NET0131 , \u0_R1_reg[7]/NET0131 , \u0_R1_reg[8]/NET0131 , \u0_R1_reg[9]/NET0131 , \u0_R2_reg[10]/NET0131 , \u0_R2_reg[11]/NET0131 , \u0_R2_reg[12]/NET0131 , \u0_R2_reg[13]/NET0131 , \u0_R2_reg[14]/NET0131 , \u0_R2_reg[15]/NET0131 , \u0_R2_reg[16]/NET0131 , \u0_R2_reg[17]/NET0131 , \u0_R2_reg[18]/NET0131 , \u0_R2_reg[19]/NET0131 , \u0_R2_reg[1]/NET0131 , \u0_R2_reg[20]/NET0131 , \u0_R2_reg[21]/NET0131 , \u0_R2_reg[22]/NET0131 , \u0_R2_reg[23]/NET0131 , \u0_R2_reg[24]/NET0131 , \u0_R2_reg[25]/NET0131 , \u0_R2_reg[26]/NET0131 , \u0_R2_reg[27]/NET0131 , \u0_R2_reg[28]/NET0131 , \u0_R2_reg[29]/NET0131 , \u0_R2_reg[2]/NET0131 , \u0_R2_reg[30]/NET0131 , \u0_R2_reg[31]/NET0131 , \u0_R2_reg[32]/NET0131 , \u0_R2_reg[3]/NET0131 , \u0_R2_reg[4]/NET0131 , \u0_R2_reg[5]/NET0131 , \u0_R2_reg[6]/NET0131 , \u0_R2_reg[7]/NET0131 , \u0_R2_reg[8]/NET0131 , \u0_R2_reg[9]/NET0131 , \u0_R3_reg[10]/NET0131 , \u0_R3_reg[11]/NET0131 , \u0_R3_reg[12]/NET0131 , \u0_R3_reg[13]/NET0131 , \u0_R3_reg[14]/NET0131 , \u0_R3_reg[15]/NET0131 , \u0_R3_reg[16]/NET0131 , \u0_R3_reg[17]/NET0131 , \u0_R3_reg[18]/NET0131 , \u0_R3_reg[19]/NET0131 , \u0_R3_reg[1]/NET0131 , \u0_R3_reg[20]/NET0131 , \u0_R3_reg[21]/NET0131 , \u0_R3_reg[22]/NET0131 , \u0_R3_reg[23]/NET0131 , \u0_R3_reg[24]/NET0131 , \u0_R3_reg[25]/NET0131 , \u0_R3_reg[26]/NET0131 , \u0_R3_reg[27]/NET0131 , \u0_R3_reg[28]/NET0131 , \u0_R3_reg[29]/NET0131 , \u0_R3_reg[2]/NET0131 , \u0_R3_reg[30]/NET0131 , \u0_R3_reg[31]/P0001 , \u0_R3_reg[32]/NET0131 , \u0_R3_reg[3]/NET0131 , \u0_R3_reg[4]/NET0131 , \u0_R3_reg[5]/NET0131 , \u0_R3_reg[6]/NET0131 , \u0_R3_reg[7]/NET0131 , \u0_R3_reg[8]/NET0131 , \u0_R3_reg[9]/NET0131 , \u0_R4_reg[10]/NET0131 , \u0_R4_reg[11]/NET0131 , \u0_R4_reg[12]/NET0131 , \u0_R4_reg[13]/NET0131 , \u0_R4_reg[14]/NET0131 , \u0_R4_reg[15]/NET0131 , \u0_R4_reg[16]/NET0131 , \u0_R4_reg[17]/NET0131 , \u0_R4_reg[18]/NET0131 , \u0_R4_reg[19]/NET0131 , \u0_R4_reg[1]/NET0131 , \u0_R4_reg[20]/NET0131 , \u0_R4_reg[21]/NET0131 , \u0_R4_reg[22]/NET0131 , \u0_R4_reg[23]/NET0131 , \u0_R4_reg[24]/NET0131 , \u0_R4_reg[25]/NET0131 , \u0_R4_reg[26]/NET0131 , \u0_R4_reg[27]/NET0131 , \u0_R4_reg[28]/NET0131 , \u0_R4_reg[29]/NET0131 , \u0_R4_reg[2]/NET0131 , \u0_R4_reg[30]/NET0131 , \u0_R4_reg[31]/P0001 , \u0_R4_reg[32]/NET0131 , \u0_R4_reg[3]/NET0131 , \u0_R4_reg[4]/NET0131 , \u0_R4_reg[5]/NET0131 , \u0_R4_reg[6]/NET0131 , \u0_R4_reg[7]/NET0131 , \u0_R4_reg[8]/NET0131 , \u0_R4_reg[9]/NET0131 , \u0_R5_reg[10]/NET0131 , \u0_R5_reg[11]/P0001 , \u0_R5_reg[12]/NET0131 , \u0_R5_reg[13]/NET0131 , \u0_R5_reg[14]/NET0131 , \u0_R5_reg[15]/NET0131 , \u0_R5_reg[16]/NET0131 , \u0_R5_reg[17]/NET0131 , \u0_R5_reg[18]/NET0131 , \u0_R5_reg[19]/NET0131 , \u0_R5_reg[1]/NET0131 , \u0_R5_reg[20]/NET0131 , \u0_R5_reg[21]/NET0131 , \u0_R5_reg[22]/NET0131 , \u0_R5_reg[23]/NET0131 , \u0_R5_reg[24]/NET0131 , \u0_R5_reg[25]/NET0131 , \u0_R5_reg[26]/NET0131 , \u0_R5_reg[27]/NET0131 , \u0_R5_reg[28]/NET0131 , \u0_R5_reg[29]/NET0131 , \u0_R5_reg[2]/NET0131 , \u0_R5_reg[30]/NET0131 , \u0_R5_reg[31]/P0001 , \u0_R5_reg[32]/NET0131 , \u0_R5_reg[3]/NET0131 , \u0_R5_reg[4]/NET0131 , \u0_R5_reg[5]/NET0131 , \u0_R5_reg[6]/NET0131 , \u0_R5_reg[7]/NET0131 , \u0_R5_reg[8]/NET0131 , \u0_R5_reg[9]/NET0131 , \u0_R6_reg[10]/NET0131 , \u0_R6_reg[11]/NET0131 , \u0_R6_reg[12]/NET0131 , \u0_R6_reg[13]/NET0131 , \u0_R6_reg[14]/NET0131 , \u0_R6_reg[15]/NET0131 , \u0_R6_reg[16]/NET0131 , \u0_R6_reg[17]/NET0131 , \u0_R6_reg[18]/NET0131 , \u0_R6_reg[19]/NET0131 , \u0_R6_reg[1]/NET0131 , \u0_R6_reg[20]/NET0131 , \u0_R6_reg[21]/NET0131 , \u0_R6_reg[22]/NET0131 , \u0_R6_reg[23]/NET0131 , \u0_R6_reg[24]/NET0131 , \u0_R6_reg[25]/NET0131 , \u0_R6_reg[26]/NET0131 , \u0_R6_reg[27]/NET0131 , \u0_R6_reg[28]/NET0131 , \u0_R6_reg[29]/NET0131 , \u0_R6_reg[2]/NET0131 , \u0_R6_reg[30]/NET0131 , \u0_R6_reg[31]/P0001 , \u0_R6_reg[32]/NET0131 , \u0_R6_reg[3]/NET0131 , \u0_R6_reg[4]/NET0131 , \u0_R6_reg[5]/NET0131 , \u0_R6_reg[6]/NET0131 , \u0_R6_reg[7]/NET0131 , \u0_R6_reg[8]/NET0131 , \u0_R6_reg[9]/NET0131 , \u0_R7_reg[10]/NET0131 , \u0_R7_reg[11]/P0001 , \u0_R7_reg[12]/NET0131 , \u0_R7_reg[13]/NET0131 , \u0_R7_reg[14]/NET0131 , \u0_R7_reg[15]/NET0131 , \u0_R7_reg[16]/NET0131 , \u0_R7_reg[17]/NET0131 , \u0_R7_reg[18]/NET0131 , \u0_R7_reg[19]/NET0131 , \u0_R7_reg[1]/NET0131 , \u0_R7_reg[20]/NET0131 , \u0_R7_reg[21]/NET0131 , \u0_R7_reg[22]/NET0131 , \u0_R7_reg[23]/NET0131 , \u0_R7_reg[24]/NET0131 , \u0_R7_reg[25]/NET0131 , \u0_R7_reg[26]/NET0131 , \u0_R7_reg[27]/NET0131 , \u0_R7_reg[28]/NET0131 , \u0_R7_reg[29]/NET0131 , \u0_R7_reg[2]/NET0131 , \u0_R7_reg[30]/NET0131 , \u0_R7_reg[31]/P0001 , \u0_R7_reg[32]/NET0131 , \u0_R7_reg[3]/NET0131 , \u0_R7_reg[4]/NET0131 , \u0_R7_reg[5]/NET0131 , \u0_R7_reg[6]/NET0131 , \u0_R7_reg[7]/NET0131 , \u0_R7_reg[8]/NET0131 , \u0_R7_reg[9]/NET0131 , \u0_R8_reg[10]/NET0131 , \u0_R8_reg[11]/NET0131 , \u0_R8_reg[12]/NET0131 , \u0_R8_reg[13]/NET0131 , \u0_R8_reg[14]/NET0131 , \u0_R8_reg[15]/NET0131 , \u0_R8_reg[16]/NET0131 , \u0_R8_reg[17]/NET0131 , \u0_R8_reg[18]/NET0131 , \u0_R8_reg[19]/NET0131 , \u0_R8_reg[1]/NET0131 , \u0_R8_reg[20]/NET0131 , \u0_R8_reg[21]/NET0131 , \u0_R8_reg[22]/NET0131 , \u0_R8_reg[23]/NET0131 , \u0_R8_reg[24]/NET0131 , \u0_R8_reg[25]/NET0131 , \u0_R8_reg[26]/NET0131 , \u0_R8_reg[27]/NET0131 , \u0_R8_reg[28]/NET0131 , \u0_R8_reg[29]/NET0131 , \u0_R8_reg[2]/NET0131 , \u0_R8_reg[30]/NET0131 , \u0_R8_reg[31]/P0001 , \u0_R8_reg[32]/NET0131 , \u0_R8_reg[3]/NET0131 , \u0_R8_reg[4]/NET0131 , \u0_R8_reg[5]/NET0131 , \u0_R8_reg[6]/NET0131 , \u0_R8_reg[7]/NET0131 , \u0_R8_reg[8]/NET0131 , \u0_R8_reg[9]/NET0131 , \u0_R9_reg[10]/NET0131 , \u0_R9_reg[11]/P0001 , \u0_R9_reg[12]/NET0131 , \u0_R9_reg[13]/NET0131 , \u0_R9_reg[14]/NET0131 , \u0_R9_reg[15]/NET0131 , \u0_R9_reg[16]/NET0131 , \u0_R9_reg[17]/NET0131 , \u0_R9_reg[18]/NET0131 , \u0_R9_reg[19]/NET0131 , \u0_R9_reg[1]/NET0131 , \u0_R9_reg[20]/NET0131 , \u0_R9_reg[21]/NET0131 , \u0_R9_reg[22]/NET0131 , \u0_R9_reg[23]/NET0131 , \u0_R9_reg[24]/NET0131 , \u0_R9_reg[25]/NET0131 , \u0_R9_reg[26]/NET0131 , \u0_R9_reg[27]/NET0131 , \u0_R9_reg[28]/NET0131 , \u0_R9_reg[29]/NET0131 , \u0_R9_reg[2]/NET0131 , \u0_R9_reg[30]/NET0131 , \u0_R9_reg[31]/P0001 , \u0_R9_reg[32]/NET0131 , \u0_R9_reg[3]/NET0131 , \u0_R9_reg[4]/NET0131 , \u0_R9_reg[5]/NET0131 , \u0_R9_reg[6]/NET0131 , \u0_R9_reg[7]/NET0131 , \u0_R9_reg[8]/NET0131 , \u0_R9_reg[9]/NET0131 , \u0_desIn_r_reg[0]/NET0131 , \u0_desIn_r_reg[10]/NET0131 , \u0_desIn_r_reg[11]/NET0131 , \u0_desIn_r_reg[12]/NET0131 , \u0_desIn_r_reg[13]/NET0131 , \u0_desIn_r_reg[14]/NET0131 , \u0_desIn_r_reg[15]/NET0131 , \u0_desIn_r_reg[16]/NET0131 , \u0_desIn_r_reg[17]/NET0131 , \u0_desIn_r_reg[18]/NET0131 , \u0_desIn_r_reg[19]/NET0131 , \u0_desIn_r_reg[1]/NET0131 , \u0_desIn_r_reg[20]/NET0131 , \u0_desIn_r_reg[21]/NET0131 , \u0_desIn_r_reg[22]/NET0131 , \u0_desIn_r_reg[23]/NET0131 , \u0_desIn_r_reg[24]/NET0131 , \u0_desIn_r_reg[25]/NET0131 , \u0_desIn_r_reg[26]/NET0131 , \u0_desIn_r_reg[27]/NET0131 , \u0_desIn_r_reg[28]/NET0131 , \u0_desIn_r_reg[29]/NET0131 , \u0_desIn_r_reg[2]/NET0131 , \u0_desIn_r_reg[30]/NET0131 , \u0_desIn_r_reg[31]/NET0131 , \u0_desIn_r_reg[32]/NET0131 , \u0_desIn_r_reg[33]/NET0131 , \u0_desIn_r_reg[34]/NET0131 , \u0_desIn_r_reg[35]/NET0131 , \u0_desIn_r_reg[36]/NET0131 , \u0_desIn_r_reg[37]/NET0131 , \u0_desIn_r_reg[38]/NET0131 , \u0_desIn_r_reg[39]/NET0131 , \u0_desIn_r_reg[3]/NET0131 , \u0_desIn_r_reg[40]/NET0131 , \u0_desIn_r_reg[41]/NET0131 , \u0_desIn_r_reg[42]/NET0131 , \u0_desIn_r_reg[43]/NET0131 , \u0_desIn_r_reg[44]/NET0131 , \u0_desIn_r_reg[45]/NET0131 , \u0_desIn_r_reg[46]/NET0131 , \u0_desIn_r_reg[47]/NET0131 , \u0_desIn_r_reg[48]/NET0131 , \u0_desIn_r_reg[49]/NET0131 , \u0_desIn_r_reg[4]/NET0131 , \u0_desIn_r_reg[50]/NET0131 , \u0_desIn_r_reg[51]/NET0131 , \u0_desIn_r_reg[52]/NET0131 , \u0_desIn_r_reg[53]/NET0131 , \u0_desIn_r_reg[54]/NET0131 , \u0_desIn_r_reg[55]/NET0131 , \u0_desIn_r_reg[56]/NET0131 , \u0_desIn_r_reg[57]/NET0131 , \u0_desIn_r_reg[58]/NET0131 , \u0_desIn_r_reg[59]/NET0131 , \u0_desIn_r_reg[5]/NET0131 , \u0_desIn_r_reg[60]/NET0131 , \u0_desIn_r_reg[61]/NET0131 , \u0_desIn_r_reg[62]/NET0131 , \u0_desIn_r_reg[63]/NET0131 , \u0_desIn_r_reg[6]/NET0131 , \u0_desIn_r_reg[7]/NET0131 , \u0_desIn_r_reg[8]/NET0131 , \u0_desIn_r_reg[9]/NET0131 , \u0_key_r_reg[0]/NET0131 , \u0_key_r_reg[10]/P0001 , \u0_key_r_reg[11]/NET0131 , \u0_key_r_reg[12]/NET0131 , \u0_key_r_reg[13]/NET0131 , \u0_key_r_reg[14]/NET0131 , \u0_key_r_reg[15]/NET0131 , \u0_key_r_reg[16]/NET0131 , \u0_key_r_reg[17]/NET0131 , \u0_key_r_reg[18]/NET0131 , \u0_key_r_reg[19]/NET0131 , \u0_key_r_reg[1]/NET0131 , \u0_key_r_reg[20]/NET0131 , \u0_key_r_reg[21]/NET0131 , \u0_key_r_reg[22]/NET0131 , \u0_key_r_reg[23]/NET0131 , \u0_key_r_reg[24]/NET0131 , \u0_key_r_reg[25]/NET0131 , \u0_key_r_reg[26]/NET0131 , \u0_key_r_reg[27]/NET0131 , \u0_key_r_reg[28]/NET0131 , \u0_key_r_reg[29]/NET0131 , \u0_key_r_reg[2]/NET0131 , \u0_key_r_reg[30]/NET0131 , \u0_key_r_reg[31]/NET0131 , \u0_key_r_reg[32]/NET0131 , \u0_key_r_reg[33]/NET0131 , \u0_key_r_reg[34]/NET0131 , \u0_key_r_reg[35]/P0001 , \u0_key_r_reg[36]/NET0131 , \u0_key_r_reg[37]/NET0131 , \u0_key_r_reg[38]/NET0131 , \u0_key_r_reg[39]/P0001 , \u0_key_r_reg[3]/NET0131 , \u0_key_r_reg[40]/NET0131 , \u0_key_r_reg[41]/NET0131 , \u0_key_r_reg[42]/P0001 , \u0_key_r_reg[43]/NET0131 , \u0_key_r_reg[44]/NET0131 , \u0_key_r_reg[45]/NET0131 , \u0_key_r_reg[46]/NET0131 , \u0_key_r_reg[47]/NET0131 , \u0_key_r_reg[48]/NET0131 , \u0_key_r_reg[49]/NET0131 , \u0_key_r_reg[4]/NET0131 , \u0_key_r_reg[50]/NET0131 , \u0_key_r_reg[51]/NET0131 , \u0_key_r_reg[52]/NET0131 , \u0_key_r_reg[53]/NET0131 , \u0_key_r_reg[54]/NET0131 , \u0_key_r_reg[55]/NET0131 , \u0_key_r_reg[5]/NET0131 , \u0_key_r_reg[6]/NET0131 , \u0_key_r_reg[7]/NET0131 , \u0_key_r_reg[8]/NET0131 , \u0_key_r_reg[9]/NET0131 , \u0_uk_K_r0_reg[0]/NET0131 , \u0_uk_K_r0_reg[10]/NET0131 , \u0_uk_K_r0_reg[11]/NET0131 , \u0_uk_K_r0_reg[12]/NET0131 , \u0_uk_K_r0_reg[13]/NET0131 , \u0_uk_K_r0_reg[14]/NET0131 , \u0_uk_K_r0_reg[15]/NET0131 , \u0_uk_K_r0_reg[16]/NET0131 , \u0_uk_K_r0_reg[17]/NET0131 , \u0_uk_K_r0_reg[18]/NET0131 , \u0_uk_K_r0_reg[19]/NET0131 , \u0_uk_K_r0_reg[20]/NET0131 , \u0_uk_K_r0_reg[21]/NET0131 , \u0_uk_K_r0_reg[22]/NET0131 , \u0_uk_K_r0_reg[23]/NET0131 , \u0_uk_K_r0_reg[24]/P0001 , \u0_uk_K_r0_reg[25]/P0001 , \u0_uk_K_r0_reg[26]/NET0131 , \u0_uk_K_r0_reg[27]/NET0131 , \u0_uk_K_r0_reg[28]/NET0131 , \u0_uk_K_r0_reg[29]/NET0131 , \u0_uk_K_r0_reg[2]/NET0131 , \u0_uk_K_r0_reg[30]/NET0131 , \u0_uk_K_r0_reg[31]/NET0131 , \u0_uk_K_r0_reg[32]/NET0131 , \u0_uk_K_r0_reg[33]/NET0131 , \u0_uk_K_r0_reg[34]/NET0131 , \u0_uk_K_r0_reg[35]/NET0131 , \u0_uk_K_r0_reg[36]/NET0131 , \u0_uk_K_r0_reg[37]/NET0131 , \u0_uk_K_r0_reg[38]/NET0131 , \u0_uk_K_r0_reg[39]/NET0131 , \u0_uk_K_r0_reg[3]/NET0131 , \u0_uk_K_r0_reg[40]/NET0131 , \u0_uk_K_r0_reg[41]/NET0131 , \u0_uk_K_r0_reg[42]/NET0131 , \u0_uk_K_r0_reg[43]/NET0131 , \u0_uk_K_r0_reg[44]/NET0131 , \u0_uk_K_r0_reg[45]/NET0131 , \u0_uk_K_r0_reg[46]/NET0131 , \u0_uk_K_r0_reg[47]/NET0131 , \u0_uk_K_r0_reg[48]/NET0131 , \u0_uk_K_r0_reg[49]/NET0131 , \u0_uk_K_r0_reg[4]/NET0131 , \u0_uk_K_r0_reg[50]/NET0131 , \u0_uk_K_r0_reg[51]/NET0131 , \u0_uk_K_r0_reg[52]/NET0131 , \u0_uk_K_r0_reg[54]/NET0131 , \u0_uk_K_r0_reg[55]/NET0131 , \u0_uk_K_r0_reg[5]/NET0131 , \u0_uk_K_r0_reg[6]/NET0131 , \u0_uk_K_r0_reg[7]/NET0131 , \u0_uk_K_r0_reg[8]/NET0131 , \u0_uk_K_r0_reg[9]/NET0131 , \u0_uk_K_r10_reg[0]/NET0131 , \u0_uk_K_r10_reg[10]/NET0131 , \u0_uk_K_r10_reg[11]/NET0131 , \u0_uk_K_r10_reg[12]/NET0131 , \u0_uk_K_r10_reg[14]/NET0131 , \u0_uk_K_r10_reg[15]/NET0131 , \u0_uk_K_r10_reg[16]/NET0131 , \u0_uk_K_r10_reg[17]/NET0131 , \u0_uk_K_r10_reg[18]/NET0131 , \u0_uk_K_r10_reg[19]/NET0131 , \u0_uk_K_r10_reg[1]/NET0131 , \u0_uk_K_r10_reg[20]/NET0131 , \u0_uk_K_r10_reg[21]/NET0131 , \u0_uk_K_r10_reg[22]/NET0131 , \u0_uk_K_r10_reg[23]/NET0131 , \u0_uk_K_r10_reg[24]/NET0131 , \u0_uk_K_r10_reg[25]/NET0131 , \u0_uk_K_r10_reg[26]/NET0131 , \u0_uk_K_r10_reg[27]/NET0131 , \u0_uk_K_r10_reg[28]/NET0131 , \u0_uk_K_r10_reg[29]/NET0131 , \u0_uk_K_r10_reg[2]/NET0131 , \u0_uk_K_r10_reg[30]/NET0131 , \u0_uk_K_r10_reg[31]/NET0131 , \u0_uk_K_r10_reg[32]/NET0131 , \u0_uk_K_r10_reg[33]/NET0131 , \u0_uk_K_r10_reg[34]/NET0131 , \u0_uk_K_r10_reg[35]/NET0131 , \u0_uk_K_r10_reg[36]/NET0131 , \u0_uk_K_r10_reg[37]/NET0131 , \u0_uk_K_r10_reg[38]/NET0131 , \u0_uk_K_r10_reg[39]/NET0131 , \u0_uk_K_r10_reg[3]/NET0131 , \u0_uk_K_r10_reg[40]/NET0131 , \u0_uk_K_r10_reg[41]/P0001 , \u0_uk_K_r10_reg[42]/NET0131 , \u0_uk_K_r10_reg[43]/NET0131 , \u0_uk_K_r10_reg[44]/NET0131 , \u0_uk_K_r10_reg[45]/P0001 , \u0_uk_K_r10_reg[46]/NET0131 , \u0_uk_K_r10_reg[47]/NET0131 , \u0_uk_K_r10_reg[48]/NET0131 , \u0_uk_K_r10_reg[49]/NET0131 , \u0_uk_K_r10_reg[4]/NET0131 , \u0_uk_K_r10_reg[50]/NET0131 , \u0_uk_K_r10_reg[51]/NET0131 , \u0_uk_K_r10_reg[52]/NET0131 , \u0_uk_K_r10_reg[53]/NET0131 , \u0_uk_K_r10_reg[54]/NET0131 , \u0_uk_K_r10_reg[55]/NET0131 , \u0_uk_K_r10_reg[5]/NET0131 , \u0_uk_K_r10_reg[6]/NET0131 , \u0_uk_K_r10_reg[7]/NET0131 , \u0_uk_K_r10_reg[8]/NET0131 , \u0_uk_K_r10_reg[9]/NET0131 , \u0_uk_K_r11_reg[0]/NET0131 , \u0_uk_K_r11_reg[10]/NET0131 , \u0_uk_K_r11_reg[11]/NET0131 , \u0_uk_K_r11_reg[12]/NET0131 , \u0_uk_K_r11_reg[13]/NET0131 , \u0_uk_K_r11_reg[14]/NET0131 , \u0_uk_K_r11_reg[15]/NET0131 , \u0_uk_K_r11_reg[16]/NET0131 , \u0_uk_K_r11_reg[17]/NET0131 , \u0_uk_K_r11_reg[18]/NET0131 , \u0_uk_K_r11_reg[19]/NET0131 , \u0_uk_K_r11_reg[1]/NET0131 , \u0_uk_K_r11_reg[20]/NET0131 , \u0_uk_K_r11_reg[21]/NET0131 , \u0_uk_K_r11_reg[22]/NET0131 , \u0_uk_K_r11_reg[23]/NET0131 , \u0_uk_K_r11_reg[24]/NET0131 , \u0_uk_K_r11_reg[25]/NET0131 , \u0_uk_K_r11_reg[26]/NET0131 , \u0_uk_K_r11_reg[27]/P0001 , \u0_uk_K_r11_reg[28]/NET0131 , \u0_uk_K_r11_reg[29]/NET0131 , \u0_uk_K_r11_reg[2]/NET0131 , \u0_uk_K_r11_reg[31]/NET0131 , \u0_uk_K_r11_reg[32]/NET0131 , \u0_uk_K_r11_reg[33]/NET0131 , \u0_uk_K_r11_reg[34]/NET0131 , \u0_uk_K_r11_reg[35]/NET0131 , \u0_uk_K_r11_reg[36]/NET0131 , \u0_uk_K_r11_reg[37]/NET0131 , \u0_uk_K_r11_reg[38]/NET0131 , \u0_uk_K_r11_reg[39]/NET0131 , \u0_uk_K_r11_reg[3]/NET0131 , \u0_uk_K_r11_reg[40]/NET0131 , \u0_uk_K_r11_reg[41]/NET0131 , \u0_uk_K_r11_reg[42]/NET0131 , \u0_uk_K_r11_reg[43]/NET0131 , \u0_uk_K_r11_reg[44]/NET0131 , \u0_uk_K_r11_reg[45]/NET0131 , \u0_uk_K_r11_reg[46]/NET0131 , \u0_uk_K_r11_reg[47]/NET0131 , \u0_uk_K_r11_reg[48]/NET0131 , \u0_uk_K_r11_reg[49]/NET0131 , \u0_uk_K_r11_reg[4]/NET0131 , \u0_uk_K_r11_reg[50]/NET0131 , \u0_uk_K_r11_reg[51]/NET0131 , \u0_uk_K_r11_reg[52]/NET0131 , \u0_uk_K_r11_reg[53]/P0001 , \u0_uk_K_r11_reg[54]/NET0131 , \u0_uk_K_r11_reg[55]/NET0131 , \u0_uk_K_r11_reg[5]/NET0131 , \u0_uk_K_r11_reg[6]/NET0131 , \u0_uk_K_r11_reg[7]/NET0131 , \u0_uk_K_r11_reg[8]/NET0131 , \u0_uk_K_r11_reg[9]/NET0131 , \u0_uk_K_r12_reg[0]/NET0131 , \u0_uk_K_r12_reg[10]/P0001 , \u0_uk_K_r12_reg[11]/NET0131 , \u0_uk_K_r12_reg[12]/NET0131 , \u0_uk_K_r12_reg[13]/NET0131 , \u0_uk_K_r12_reg[14]/NET0131 , \u0_uk_K_r12_reg[15]/NET0131 , \u0_uk_K_r12_reg[16]/NET0131 , \u0_uk_K_r12_reg[17]/NET0131 , \u0_uk_K_r12_reg[18]/NET0131 , \u0_uk_K_r12_reg[19]/NET0131 , \u0_uk_K_r12_reg[1]/NET0131 , \u0_uk_K_r12_reg[20]/NET0131 , \u0_uk_K_r12_reg[21]/NET0131 , \u0_uk_K_r12_reg[22]/NET0131 , \u0_uk_K_r12_reg[23]/NET0131 , \u0_uk_K_r12_reg[24]/NET0131 , \u0_uk_K_r12_reg[25]/NET0131 , \u0_uk_K_r12_reg[26]/NET0131 , \u0_uk_K_r12_reg[27]/NET0131 , \u0_uk_K_r12_reg[28]/NET0131 , \u0_uk_K_r12_reg[29]/NET0131 , \u0_uk_K_r12_reg[2]/NET0131 , \u0_uk_K_r12_reg[30]/NET0131 , \u0_uk_K_r12_reg[31]/NET0131 , \u0_uk_K_r12_reg[32]/NET0131 , \u0_uk_K_r12_reg[33]/NET0131 , \u0_uk_K_r12_reg[34]/NET0131 , \u0_uk_K_r12_reg[35]/NET0131 , \u0_uk_K_r12_reg[36]/NET0131 , \u0_uk_K_r12_reg[37]/NET0131 , \u0_uk_K_r12_reg[38]/NET0131 , \u0_uk_K_r12_reg[3]/NET0131 , \u0_uk_K_r12_reg[40]/NET0131 , \u0_uk_K_r12_reg[41]/NET0131 , \u0_uk_K_r12_reg[42]/NET0131 , \u0_uk_K_r12_reg[43]/NET0131 , \u0_uk_K_r12_reg[44]/P0001 , \u0_uk_K_r12_reg[45]/NET0131 , \u0_uk_K_r12_reg[46]/NET0131 , \u0_uk_K_r12_reg[47]/NET0131 , \u0_uk_K_r12_reg[48]/NET0131 , \u0_uk_K_r12_reg[49]/NET0131 , \u0_uk_K_r12_reg[4]/NET0131 , \u0_uk_K_r12_reg[50]/NET0131 , \u0_uk_K_r12_reg[51]/NET0131 , \u0_uk_K_r12_reg[52]/NET0131 , \u0_uk_K_r12_reg[53]/NET0131 , \u0_uk_K_r12_reg[54]/NET0131 , \u0_uk_K_r12_reg[55]/NET0131 , \u0_uk_K_r12_reg[5]/NET0131 , \u0_uk_K_r12_reg[6]/NET0131 , \u0_uk_K_r12_reg[7]/P0001 , \u0_uk_K_r12_reg[8]/NET0131 , \u0_uk_K_r12_reg[9]/NET0131 , \u0_uk_K_r13_reg[0]/NET0131 , \u0_uk_K_r13_reg[10]/NET0131 , \u0_uk_K_r13_reg[11]/NET0131 , \u0_uk_K_r13_reg[12]/NET0131 , \u0_uk_K_r13_reg[13]/NET0131 , \u0_uk_K_r13_reg[14]/NET0131 , \u0_uk_K_r13_reg[15]/NET0131 , \u0_uk_K_r13_reg[16]/NET0131 , \u0_uk_K_r13_reg[17]/NET0131 , \u0_uk_K_r13_reg[18]/NET0131 , \u0_uk_K_r13_reg[19]/NET0131 , \u0_uk_K_r13_reg[20]/NET0131 , \u0_uk_K_r13_reg[21]/NET0131 , \u0_uk_K_r13_reg[22]/NET0131 , \u0_uk_K_r13_reg[23]/NET0131 , \u0_uk_K_r13_reg[24]/NET0131 , \u0_uk_K_r13_reg[25]/P0001 , \u0_uk_K_r13_reg[26]/NET0131 , \u0_uk_K_r13_reg[27]/NET0131 , \u0_uk_K_r13_reg[28]/NET0131 , \u0_uk_K_r13_reg[29]/NET0131 , \u0_uk_K_r13_reg[2]/NET0131 , \u0_uk_K_r13_reg[30]/NET0131 , \u0_uk_K_r13_reg[31]/NET0131 , \u0_uk_K_r13_reg[32]/NET0131 , \u0_uk_K_r13_reg[33]/NET0131 , \u0_uk_K_r13_reg[34]/NET0131 , \u0_uk_K_r13_reg[35]/NET0131 , \u0_uk_K_r13_reg[36]/NET0131 , \u0_uk_K_r13_reg[37]/NET0131 , \u0_uk_K_r13_reg[38]/NET0131 , \u0_uk_K_r13_reg[39]/NET0131 , \u0_uk_K_r13_reg[3]/NET0131 , \u0_uk_K_r13_reg[40]/NET0131 , \u0_uk_K_r13_reg[41]/NET0131 , \u0_uk_K_r13_reg[42]/NET0131 , \u0_uk_K_r13_reg[43]/NET0131 , \u0_uk_K_r13_reg[44]/NET0131 , \u0_uk_K_r13_reg[45]/NET0131 , \u0_uk_K_r13_reg[46]/NET0131 , \u0_uk_K_r13_reg[47]/NET0131 , \u0_uk_K_r13_reg[48]/NET0131 , \u0_uk_K_r13_reg[49]/NET0131 , \u0_uk_K_r13_reg[4]/NET0131 , \u0_uk_K_r13_reg[50]/NET0131 , \u0_uk_K_r13_reg[51]/NET0131 , \u0_uk_K_r13_reg[52]/P0001 , \u0_uk_K_r13_reg[54]/NET0131 , \u0_uk_K_r13_reg[55]/NET0131 , \u0_uk_K_r13_reg[5]/NET0131 , \u0_uk_K_r13_reg[6]/NET0131 , \u0_uk_K_r13_reg[7]/NET0131 , \u0_uk_K_r13_reg[8]/NET0131 , \u0_uk_K_r13_reg[9]/NET0131 , \u0_uk_K_r14_reg[0]/NET0131 , \u0_uk_K_r14_reg[10]/P0001 , \u0_uk_K_r14_reg[11]/NET0131 , \u0_uk_K_r14_reg[12]/NET0131 , \u0_uk_K_r14_reg[13]/NET0131 , \u0_uk_K_r14_reg[14]/NET0131 , \u0_uk_K_r14_reg[15]/NET0131 , \u0_uk_K_r14_reg[16]/NET0131 , \u0_uk_K_r14_reg[17]/NET0131 , \u0_uk_K_r14_reg[18]/NET0131 , \u0_uk_K_r14_reg[19]/NET0131 , \u0_uk_K_r14_reg[1]/NET0131 , \u0_uk_K_r14_reg[20]/NET0131 , \u0_uk_K_r14_reg[21]/NET0131 , \u0_uk_K_r14_reg[22]/NET0131 , \u0_uk_K_r14_reg[23]/NET0131 , \u0_uk_K_r14_reg[24]/NET0131 , \u0_uk_K_r14_reg[25]/NET0131 , \u0_uk_K_r14_reg[26]/NET0131 , \u0_uk_K_r14_reg[27]/NET0131 , \u0_uk_K_r14_reg[28]/NET0131 , \u0_uk_K_r14_reg[29]/NET0131 , \u0_uk_K_r14_reg[2]/NET0131 , \u0_uk_K_r14_reg[30]/NET0131 , \u0_uk_K_r14_reg[31]/NET0131 , \u0_uk_K_r14_reg[32]/NET0131 , \u0_uk_K_r14_reg[33]/NET0131 , \u0_uk_K_r14_reg[34]/NET0131 , \u0_uk_K_r14_reg[35]/P0001 , \u0_uk_K_r14_reg[36]/NET0131 , \u0_uk_K_r14_reg[37]/NET0131 , \u0_uk_K_r14_reg[38]/NET0131 , \u0_uk_K_r14_reg[39]/P0001 , \u0_uk_K_r14_reg[3]/NET0131 , \u0_uk_K_r14_reg[40]/NET0131 , \u0_uk_K_r14_reg[41]/NET0131 , \u0_uk_K_r14_reg[42]/P0001 , \u0_uk_K_r14_reg[43]/NET0131 , \u0_uk_K_r14_reg[44]/NET0131 , \u0_uk_K_r14_reg[45]/NET0131 , \u0_uk_K_r14_reg[46]/NET0131 , \u0_uk_K_r14_reg[47]/NET0131 , \u0_uk_K_r14_reg[48]/NET0131 , \u0_uk_K_r14_reg[49]/NET0131 , \u0_uk_K_r14_reg[4]/NET0131 , \u0_uk_K_r14_reg[50]/NET0131 , \u0_uk_K_r14_reg[51]/NET0131 , \u0_uk_K_r14_reg[52]/NET0131 , \u0_uk_K_r14_reg[53]/NET0131 , \u0_uk_K_r14_reg[54]/NET0131 , \u0_uk_K_r14_reg[55]/NET0131 , \u0_uk_K_r14_reg[5]/NET0131 , \u0_uk_K_r14_reg[6]/NET0131 , \u0_uk_K_r14_reg[7]/NET0131 , \u0_uk_K_r14_reg[8]/NET0131 , \u0_uk_K_r14_reg[9]/NET0131 , \u0_uk_K_r1_reg[0]/NET0131 , \u0_uk_K_r1_reg[10]/P0001 , \u0_uk_K_r1_reg[11]/NET0131 , \u0_uk_K_r1_reg[12]/NET0131 , \u0_uk_K_r1_reg[13]/NET0131 , \u0_uk_K_r1_reg[14]/NET0131 , \u0_uk_K_r1_reg[15]/NET0131 , \u0_uk_K_r1_reg[16]/NET0131 , \u0_uk_K_r1_reg[17]/NET0131 , \u0_uk_K_r1_reg[18]/NET0131 , \u0_uk_K_r1_reg[19]/NET0131 , \u0_uk_K_r1_reg[1]/NET0131 , \u0_uk_K_r1_reg[20]/NET0131 , \u0_uk_K_r1_reg[21]/NET0131 , \u0_uk_K_r1_reg[22]/NET0131 , \u0_uk_K_r1_reg[23]/NET0131 , \u0_uk_K_r1_reg[24]/NET0131 , \u0_uk_K_r1_reg[25]/NET0131 , \u0_uk_K_r1_reg[26]/NET0131 , \u0_uk_K_r1_reg[27]/NET0131 , \u0_uk_K_r1_reg[28]/NET0131 , \u0_uk_K_r1_reg[29]/NET0131 , \u0_uk_K_r1_reg[2]/NET0131 , \u0_uk_K_r1_reg[30]/NET0131 , \u0_uk_K_r1_reg[31]/NET0131 , \u0_uk_K_r1_reg[32]/NET0131 , \u0_uk_K_r1_reg[33]/NET0131 , \u0_uk_K_r1_reg[34]/NET0131 , \u0_uk_K_r1_reg[35]/NET0131 , \u0_uk_K_r1_reg[36]/NET0131 , \u0_uk_K_r1_reg[37]/NET0131 , \u0_uk_K_r1_reg[38]/NET0131 , \u0_uk_K_r1_reg[3]/NET0131 , \u0_uk_K_r1_reg[40]/NET0131 , \u0_uk_K_r1_reg[41]/NET0131 , \u0_uk_K_r1_reg[42]/NET0131 , \u0_uk_K_r1_reg[43]/NET0131 , \u0_uk_K_r1_reg[44]/P0001 , \u0_uk_K_r1_reg[45]/NET0131 , \u0_uk_K_r1_reg[46]/NET0131 , \u0_uk_K_r1_reg[47]/NET0131 , \u0_uk_K_r1_reg[48]/NET0131 , \u0_uk_K_r1_reg[49]/NET0131 , \u0_uk_K_r1_reg[4]/NET0131 , \u0_uk_K_r1_reg[50]/NET0131 , \u0_uk_K_r1_reg[51]/NET0131 , \u0_uk_K_r1_reg[52]/NET0131 , \u0_uk_K_r1_reg[53]/NET0131 , \u0_uk_K_r1_reg[54]/NET0131 , \u0_uk_K_r1_reg[55]/NET0131 , \u0_uk_K_r1_reg[5]/NET0131 , \u0_uk_K_r1_reg[6]/NET0131 , \u0_uk_K_r1_reg[7]/P0001 , \u0_uk_K_r1_reg[8]/NET0131 , \u0_uk_K_r1_reg[9]/NET0131 , \u0_uk_K_r2_reg[0]/NET0131 , \u0_uk_K_r2_reg[10]/NET0131 , \u0_uk_K_r2_reg[11]/NET0131 , \u0_uk_K_r2_reg[12]/NET0131 , \u0_uk_K_r2_reg[13]/NET0131 , \u0_uk_K_r2_reg[14]/NET0131 , \u0_uk_K_r2_reg[15]/NET0131 , \u0_uk_K_r2_reg[16]/NET0131 , \u0_uk_K_r2_reg[17]/NET0131 , \u0_uk_K_r2_reg[18]/NET0131 , \u0_uk_K_r2_reg[19]/NET0131 , \u0_uk_K_r2_reg[1]/NET0131 , \u0_uk_K_r2_reg[20]/NET0131 , \u0_uk_K_r2_reg[21]/NET0131 , \u0_uk_K_r2_reg[22]/NET0131 , \u0_uk_K_r2_reg[23]/NET0131 , \u0_uk_K_r2_reg[24]/NET0131 , \u0_uk_K_r2_reg[25]/NET0131 , \u0_uk_K_r2_reg[26]/NET0131 , \u0_uk_K_r2_reg[27]/P0001 , \u0_uk_K_r2_reg[28]/NET0131 , \u0_uk_K_r2_reg[29]/NET0131 , \u0_uk_K_r2_reg[2]/NET0131 , \u0_uk_K_r2_reg[31]/NET0131 , \u0_uk_K_r2_reg[32]/NET0131 , \u0_uk_K_r2_reg[33]/NET0131 , \u0_uk_K_r2_reg[34]/NET0131 , \u0_uk_K_r2_reg[35]/NET0131 , \u0_uk_K_r2_reg[36]/NET0131 , \u0_uk_K_r2_reg[37]/NET0131 , \u0_uk_K_r2_reg[38]/NET0131 , \u0_uk_K_r2_reg[39]/NET0131 , \u0_uk_K_r2_reg[3]/NET0131 , \u0_uk_K_r2_reg[40]/NET0131 , \u0_uk_K_r2_reg[41]/NET0131 , \u0_uk_K_r2_reg[42]/NET0131 , \u0_uk_K_r2_reg[43]/NET0131 , \u0_uk_K_r2_reg[44]/NET0131 , \u0_uk_K_r2_reg[45]/NET0131 , \u0_uk_K_r2_reg[46]/NET0131 , \u0_uk_K_r2_reg[47]/NET0131 , \u0_uk_K_r2_reg[48]/NET0131 , \u0_uk_K_r2_reg[49]/NET0131 , \u0_uk_K_r2_reg[4]/NET0131 , \u0_uk_K_r2_reg[50]/NET0131 , \u0_uk_K_r2_reg[51]/NET0131 , \u0_uk_K_r2_reg[52]/NET0131 , \u0_uk_K_r2_reg[53]/P0001 , \u0_uk_K_r2_reg[54]/NET0131 , \u0_uk_K_r2_reg[55]/NET0131 , \u0_uk_K_r2_reg[5]/NET0131 , \u0_uk_K_r2_reg[6]/NET0131 , \u0_uk_K_r2_reg[7]/NET0131 , \u0_uk_K_r2_reg[8]/NET0131 , \u0_uk_K_r2_reg[9]/NET0131 , \u0_uk_K_r3_reg[0]/NET0131 , \u0_uk_K_r3_reg[10]/NET0131 , \u0_uk_K_r3_reg[11]/NET0131 , \u0_uk_K_r3_reg[12]/NET0131 , \u0_uk_K_r3_reg[14]/NET0131 , \u0_uk_K_r3_reg[15]/NET0131 , \u0_uk_K_r3_reg[16]/NET0131 , \u0_uk_K_r3_reg[17]/NET0131 , \u0_uk_K_r3_reg[18]/NET0131 , \u0_uk_K_r3_reg[19]/NET0131 , \u0_uk_K_r3_reg[1]/NET0131 , \u0_uk_K_r3_reg[20]/NET0131 , \u0_uk_K_r3_reg[21]/NET0131 , \u0_uk_K_r3_reg[22]/NET0131 , \u0_uk_K_r3_reg[23]/NET0131 , \u0_uk_K_r3_reg[24]/NET0131 , \u0_uk_K_r3_reg[25]/NET0131 , \u0_uk_K_r3_reg[26]/NET0131 , \u0_uk_K_r3_reg[27]/NET0131 , \u0_uk_K_r3_reg[28]/NET0131 , \u0_uk_K_r3_reg[29]/NET0131 , \u0_uk_K_r3_reg[2]/NET0131 , \u0_uk_K_r3_reg[30]/NET0131 , \u0_uk_K_r3_reg[31]/NET0131 , \u0_uk_K_r3_reg[32]/NET0131 , \u0_uk_K_r3_reg[33]/NET0131 , \u0_uk_K_r3_reg[34]/NET0131 , \u0_uk_K_r3_reg[35]/NET0131 , \u0_uk_K_r3_reg[36]/NET0131 , \u0_uk_K_r3_reg[37]/NET0131 , \u0_uk_K_r3_reg[38]/NET0131 , \u0_uk_K_r3_reg[39]/NET0131 , \u0_uk_K_r3_reg[3]/NET0131 , \u0_uk_K_r3_reg[40]/NET0131 , \u0_uk_K_r3_reg[41]/NET0131 , \u0_uk_K_r3_reg[42]/NET0131 , \u0_uk_K_r3_reg[43]/NET0131 , \u0_uk_K_r3_reg[44]/NET0131 , \u0_uk_K_r3_reg[45]/P0001 , \u0_uk_K_r3_reg[46]/NET0131 , \u0_uk_K_r3_reg[47]/NET0131 , \u0_uk_K_r3_reg[48]/NET0131 , \u0_uk_K_r3_reg[49]/NET0131 , \u0_uk_K_r3_reg[4]/NET0131 , \u0_uk_K_r3_reg[50]/NET0131 , \u0_uk_K_r3_reg[51]/NET0131 , \u0_uk_K_r3_reg[52]/NET0131 , \u0_uk_K_r3_reg[53]/NET0131 , \u0_uk_K_r3_reg[54]/NET0131 , \u0_uk_K_r3_reg[55]/NET0131 , \u0_uk_K_r3_reg[5]/NET0131 , \u0_uk_K_r3_reg[6]/NET0131 , \u0_uk_K_r3_reg[7]/NET0131 , \u0_uk_K_r3_reg[8]/NET0131 , \u0_uk_K_r3_reg[9]/NET0131 , \u0_uk_K_r4_reg[0]/P0001 , \u0_uk_K_r4_reg[10]/NET0131 , \u0_uk_K_r4_reg[11]/NET0131 , \u0_uk_K_r4_reg[12]/NET0131 , \u0_uk_K_r4_reg[13]/NET0131 , \u0_uk_K_r4_reg[14]/NET0131 , \u0_uk_K_r4_reg[15]/NET0131 , \u0_uk_K_r4_reg[16]/NET0131 , \u0_uk_K_r4_reg[17]/NET0131 , \u0_uk_K_r4_reg[18]/NET0131 , \u0_uk_K_r4_reg[19]/NET0131 , \u0_uk_K_r4_reg[1]/NET0131 , \u0_uk_K_r4_reg[20]/NET0131 , \u0_uk_K_r4_reg[21]/NET0131 , \u0_uk_K_r4_reg[22]/NET0131 , \u0_uk_K_r4_reg[23]/P0001 , \u0_uk_K_r4_reg[25]/NET0131 , \u0_uk_K_r4_reg[26]/NET0131 , \u0_uk_K_r4_reg[27]/P0001 , \u0_uk_K_r4_reg[28]/NET0131 , \u0_uk_K_r4_reg[29]/NET0131 , \u0_uk_K_r4_reg[30]/NET0131 , \u0_uk_K_r4_reg[31]/P0001 , \u0_uk_K_r4_reg[32]/NET0131 , \u0_uk_K_r4_reg[33]/NET0131 , \u0_uk_K_r4_reg[34]/NET0131 , \u0_uk_K_r4_reg[35]/NET0131 , \u0_uk_K_r4_reg[36]/NET0131 , \u0_uk_K_r4_reg[37]/NET0131 , \u0_uk_K_r4_reg[38]/NET0131 , \u0_uk_K_r4_reg[39]/NET0131 , \u0_uk_K_r4_reg[3]/NET0131 , \u0_uk_K_r4_reg[40]/NET0131 , \u0_uk_K_r4_reg[41]/NET0131 , \u0_uk_K_r4_reg[42]/NET0131 , \u0_uk_K_r4_reg[43]/NET0131 , \u0_uk_K_r4_reg[44]/NET0131 , \u0_uk_K_r4_reg[45]/NET0131 , \u0_uk_K_r4_reg[46]/NET0131 , \u0_uk_K_r4_reg[47]/NET0131 , \u0_uk_K_r4_reg[48]/NET0131 , \u0_uk_K_r4_reg[49]/NET0131 , \u0_uk_K_r4_reg[4]/NET0131 , \u0_uk_K_r4_reg[50]/NET0131 , \u0_uk_K_r4_reg[51]/NET0131 , \u0_uk_K_r4_reg[52]/NET0131 , \u0_uk_K_r4_reg[53]/NET0131 , \u0_uk_K_r4_reg[54]/NET0131 , \u0_uk_K_r4_reg[55]/NET0131 , \u0_uk_K_r4_reg[5]/NET0131 , \u0_uk_K_r4_reg[6]/NET0131 , \u0_uk_K_r4_reg[7]/NET0131 , \u0_uk_K_r4_reg[8]/NET0131 , \u0_uk_K_r4_reg[9]/NET0131 , \u0_uk_K_r5_reg[0]/NET0131 , \u0_uk_K_r5_reg[10]/NET0131 , \u0_uk_K_r5_reg[11]/NET0131 , \u0_uk_K_r5_reg[12]/NET0131 , \u0_uk_K_r5_reg[13]/P0001 , \u0_uk_K_r5_reg[14]/NET0131 , \u0_uk_K_r5_reg[15]/NET0131 , \u0_uk_K_r5_reg[16]/NET0131 , \u0_uk_K_r5_reg[17]/NET0131 , \u0_uk_K_r5_reg[18]/NET0131 , \u0_uk_K_r5_reg[19]/NET0131 , \u0_uk_K_r5_reg[1]/NET0131 , \u0_uk_K_r5_reg[20]/NET0131 , \u0_uk_K_r5_reg[21]/NET0131 , \u0_uk_K_r5_reg[22]/NET0131 , \u0_uk_K_r5_reg[23]/NET0131 , \u0_uk_K_r5_reg[24]/NET0131 , \u0_uk_K_r5_reg[25]/NET0131 , \u0_uk_K_r5_reg[26]/NET0131 , \u0_uk_K_r5_reg[27]/NET0131 , \u0_uk_K_r5_reg[28]/NET0131 , \u0_uk_K_r5_reg[29]/NET0131 , \u0_uk_K_r5_reg[2]/NET0131 , \u0_uk_K_r5_reg[30]/NET0131 , \u0_uk_K_r5_reg[31]/NET0131 , \u0_uk_K_r5_reg[32]/NET0131 , \u0_uk_K_r5_reg[33]/NET0131 , \u0_uk_K_r5_reg[34]/NET0131 , \u0_uk_K_r5_reg[35]/NET0131 , \u0_uk_K_r5_reg[36]/NET0131 , \u0_uk_K_r5_reg[37]/P0001 , \u0_uk_K_r5_reg[38]/NET0131 , \u0_uk_K_r5_reg[39]/NET0131 , \u0_uk_K_r5_reg[3]/NET0131 , \u0_uk_K_r5_reg[40]/NET0131 , \u0_uk_K_r5_reg[41]/NET0131 , \u0_uk_K_r5_reg[42]/NET0131 , \u0_uk_K_r5_reg[43]/NET0131 , \u0_uk_K_r5_reg[44]/NET0131 , \u0_uk_K_r5_reg[46]/NET0131 , \u0_uk_K_r5_reg[47]/NET0131 , \u0_uk_K_r5_reg[48]/NET0131 , \u0_uk_K_r5_reg[49]/NET0131 , \u0_uk_K_r5_reg[4]/NET0131 , \u0_uk_K_r5_reg[50]/NET0131 , \u0_uk_K_r5_reg[51]/NET0131 , \u0_uk_K_r5_reg[52]/NET0131 , \u0_uk_K_r5_reg[53]/NET0131 , \u0_uk_K_r5_reg[54]/NET0131 , \u0_uk_K_r5_reg[55]/NET0131 , \u0_uk_K_r5_reg[5]/NET0131 , \u0_uk_K_r5_reg[6]/NET0131 , \u0_uk_K_r5_reg[7]/NET0131 , \u0_uk_K_r5_reg[8]/NET0131 , \u0_uk_K_r5_reg[9]/NET0131 , \u0_uk_K_r6_reg[0]/NET0131 , \u0_uk_K_r6_reg[10]/NET0131 , \u0_uk_K_r6_reg[11]/NET0131 , \u0_uk_K_r6_reg[12]/NET0131 , \u0_uk_K_r6_reg[13]/NET0131 , \u0_uk_K_r6_reg[14]/NET0131 , \u0_uk_K_r6_reg[15]/NET0131 , \u0_uk_K_r6_reg[16]/NET0131 , \u0_uk_K_r6_reg[17]/NET0131 , \u0_uk_K_r6_reg[18]/NET0131 , \u0_uk_K_r6_reg[19]/NET0131 , \u0_uk_K_r6_reg[1]/NET0131 , \u0_uk_K_r6_reg[20]/NET0131 , \u0_uk_K_r6_reg[21]/NET0131 , \u0_uk_K_r6_reg[22]/NET0131 , \u0_uk_K_r6_reg[23]/P0001 , \u0_uk_K_r6_reg[24]/NET0131 , \u0_uk_K_r6_reg[25]/NET0131 , \u0_uk_K_r6_reg[26]/P0001 , \u0_uk_K_r6_reg[27]/NET0131 , \u0_uk_K_r6_reg[28]/NET0131 , \u0_uk_K_r6_reg[29]/NET0131 , \u0_uk_K_r6_reg[2]/NET0131 , \u0_uk_K_r6_reg[30]/P0001 , \u0_uk_K_r6_reg[31]/NET0131 , \u0_uk_K_r6_reg[32]/NET0131 , \u0_uk_K_r6_reg[33]/NET0131 , \u0_uk_K_r6_reg[34]/NET0131 , \u0_uk_K_r6_reg[35]/NET0131 , \u0_uk_K_r6_reg[36]/NET0131 , \u0_uk_K_r6_reg[37]/NET0131 , \u0_uk_K_r6_reg[38]/NET0131 , \u0_uk_K_r6_reg[39]/NET0131 , \u0_uk_K_r6_reg[3]/NET0131 , \u0_uk_K_r6_reg[40]/NET0131 , \u0_uk_K_r6_reg[41]/NET0131 , \u0_uk_K_r6_reg[42]/NET0131 , \u0_uk_K_r6_reg[43]/NET0131 , \u0_uk_K_r6_reg[44]/NET0131 , \u0_uk_K_r6_reg[45]/NET0131 , \u0_uk_K_r6_reg[46]/NET0131 , \u0_uk_K_r6_reg[47]/NET0131 , \u0_uk_K_r6_reg[48]/NET0131 , \u0_uk_K_r6_reg[49]/NET0131 , \u0_uk_K_r6_reg[4]/NET0131 , \u0_uk_K_r6_reg[50]/NET0131 , \u0_uk_K_r6_reg[51]/NET0131 , \u0_uk_K_r6_reg[52]/NET0131 , \u0_uk_K_r6_reg[53]/NET0131 , \u0_uk_K_r6_reg[54]/NET0131 , \u0_uk_K_r6_reg[55]/P0001 , \u0_uk_K_r6_reg[5]/NET0131 , \u0_uk_K_r6_reg[6]/NET0131 , \u0_uk_K_r6_reg[7]/NET0131 , \u0_uk_K_r6_reg[8]/NET0131 , \u0_uk_K_r6_reg[9]/NET0131 , \u0_uk_K_r7_reg[0]/NET0131 , \u0_uk_K_r7_reg[10]/NET0131 , \u0_uk_K_r7_reg[11]/NET0131 , \u0_uk_K_r7_reg[12]/NET0131 , \u0_uk_K_r7_reg[13]/NET0131 , \u0_uk_K_r7_reg[14]/NET0131 , \u0_uk_K_r7_reg[15]/NET0131 , \u0_uk_K_r7_reg[16]/NET0131 , \u0_uk_K_r7_reg[17]/NET0131 , \u0_uk_K_r7_reg[18]/NET0131 , \u0_uk_K_r7_reg[19]/NET0131 , \u0_uk_K_r7_reg[1]/NET0131 , \u0_uk_K_r7_reg[20]/NET0131 , \u0_uk_K_r7_reg[21]/NET0131 , \u0_uk_K_r7_reg[22]/NET0131 , \u0_uk_K_r7_reg[23]/P0001 , \u0_uk_K_r7_reg[24]/NET0131 , \u0_uk_K_r7_reg[25]/NET0131 , \u0_uk_K_r7_reg[26]/P0001 , \u0_uk_K_r7_reg[27]/NET0131 , \u0_uk_K_r7_reg[28]/NET0131 , \u0_uk_K_r7_reg[29]/NET0131 , \u0_uk_K_r7_reg[2]/NET0131 , \u0_uk_K_r7_reg[30]/P0001 , \u0_uk_K_r7_reg[31]/NET0131 , \u0_uk_K_r7_reg[32]/NET0131 , \u0_uk_K_r7_reg[33]/NET0131 , \u0_uk_K_r7_reg[34]/NET0131 , \u0_uk_K_r7_reg[35]/NET0131 , \u0_uk_K_r7_reg[36]/NET0131 , \u0_uk_K_r7_reg[37]/NET0131 , \u0_uk_K_r7_reg[38]/NET0131 , \u0_uk_K_r7_reg[39]/NET0131 , \u0_uk_K_r7_reg[3]/NET0131 , \u0_uk_K_r7_reg[40]/NET0131 , \u0_uk_K_r7_reg[41]/NET0131 , \u0_uk_K_r7_reg[42]/NET0131 , \u0_uk_K_r7_reg[43]/NET0131 , \u0_uk_K_r7_reg[44]/NET0131 , \u0_uk_K_r7_reg[45]/NET0131 , \u0_uk_K_r7_reg[46]/NET0131 , \u0_uk_K_r7_reg[47]/NET0131 , \u0_uk_K_r7_reg[48]/NET0131 , \u0_uk_K_r7_reg[49]/NET0131 , \u0_uk_K_r7_reg[4]/NET0131 , \u0_uk_K_r7_reg[50]/NET0131 , \u0_uk_K_r7_reg[51]/NET0131 , \u0_uk_K_r7_reg[52]/NET0131 , \u0_uk_K_r7_reg[53]/NET0131 , \u0_uk_K_r7_reg[54]/NET0131 , \u0_uk_K_r7_reg[55]/P0001 , \u0_uk_K_r7_reg[5]/NET0131 , \u0_uk_K_r7_reg[6]/NET0131 , \u0_uk_K_r7_reg[7]/NET0131 , \u0_uk_K_r7_reg[8]/NET0131 , \u0_uk_K_r7_reg[9]/NET0131 , \u0_uk_K_r8_reg[0]/NET0131 , \u0_uk_K_r8_reg[10]/NET0131 , \u0_uk_K_r8_reg[11]/NET0131 , \u0_uk_K_r8_reg[12]/NET0131 , \u0_uk_K_r8_reg[13]/P0001 , \u0_uk_K_r8_reg[14]/NET0131 , \u0_uk_K_r8_reg[15]/NET0131 , \u0_uk_K_r8_reg[16]/NET0131 , \u0_uk_K_r8_reg[17]/NET0131 , \u0_uk_K_r8_reg[18]/NET0131 , \u0_uk_K_r8_reg[19]/NET0131 , \u0_uk_K_r8_reg[1]/NET0131 , \u0_uk_K_r8_reg[20]/NET0131 , \u0_uk_K_r8_reg[21]/NET0131 , \u0_uk_K_r8_reg[22]/NET0131 , \u0_uk_K_r8_reg[23]/NET0131 , \u0_uk_K_r8_reg[24]/NET0131 , \u0_uk_K_r8_reg[25]/NET0131 , \u0_uk_K_r8_reg[26]/NET0131 , \u0_uk_K_r8_reg[27]/NET0131 , \u0_uk_K_r8_reg[28]/NET0131 , \u0_uk_K_r8_reg[29]/NET0131 , \u0_uk_K_r8_reg[2]/NET0131 , \u0_uk_K_r8_reg[30]/NET0131 , \u0_uk_K_r8_reg[31]/NET0131 , \u0_uk_K_r8_reg[32]/NET0131 , \u0_uk_K_r8_reg[33]/NET0131 , \u0_uk_K_r8_reg[34]/NET0131 , \u0_uk_K_r8_reg[35]/NET0131 , \u0_uk_K_r8_reg[36]/NET0131 , \u0_uk_K_r8_reg[37]/P0001 , \u0_uk_K_r8_reg[38]/NET0131 , \u0_uk_K_r8_reg[39]/NET0131 , \u0_uk_K_r8_reg[3]/NET0131 , \u0_uk_K_r8_reg[40]/NET0131 , \u0_uk_K_r8_reg[41]/NET0131 , \u0_uk_K_r8_reg[42]/NET0131 , \u0_uk_K_r8_reg[43]/NET0131 , \u0_uk_K_r8_reg[44]/NET0131 , \u0_uk_K_r8_reg[46]/NET0131 , \u0_uk_K_r8_reg[47]/NET0131 , \u0_uk_K_r8_reg[48]/NET0131 , \u0_uk_K_r8_reg[49]/NET0131 , \u0_uk_K_r8_reg[4]/NET0131 , \u0_uk_K_r8_reg[50]/NET0131 , \u0_uk_K_r8_reg[51]/NET0131 , \u0_uk_K_r8_reg[52]/NET0131 , \u0_uk_K_r8_reg[53]/NET0131 , \u0_uk_K_r8_reg[54]/NET0131 , \u0_uk_K_r8_reg[55]/NET0131 , \u0_uk_K_r8_reg[5]/NET0131 , \u0_uk_K_r8_reg[6]/NET0131 , \u0_uk_K_r8_reg[7]/NET0131 , \u0_uk_K_r8_reg[8]/NET0131 , \u0_uk_K_r8_reg[9]/P0001 , \u0_uk_K_r9_reg[0]/P0001 , \u0_uk_K_r9_reg[10]/NET0131 , \u0_uk_K_r9_reg[11]/NET0131 , \u0_uk_K_r9_reg[12]/NET0131 , \u0_uk_K_r9_reg[13]/NET0131 , \u0_uk_K_r9_reg[14]/NET0131 , \u0_uk_K_r9_reg[15]/NET0131 , \u0_uk_K_r9_reg[16]/NET0131 , \u0_uk_K_r9_reg[17]/NET0131 , \u0_uk_K_r9_reg[18]/NET0131 , \u0_uk_K_r9_reg[19]/NET0131 , \u0_uk_K_r9_reg[1]/NET0131 , \u0_uk_K_r9_reg[20]/NET0131 , \u0_uk_K_r9_reg[21]/NET0131 , \u0_uk_K_r9_reg[22]/NET0131 , \u0_uk_K_r9_reg[23]/P0001 , \u0_uk_K_r9_reg[25]/NET0131 , \u0_uk_K_r9_reg[26]/NET0131 , \u0_uk_K_r9_reg[27]/P0001 , \u0_uk_K_r9_reg[28]/NET0131 , \u0_uk_K_r9_reg[29]/NET0131 , \u0_uk_K_r9_reg[30]/NET0131 , \u0_uk_K_r9_reg[31]/P0001 , \u0_uk_K_r9_reg[32]/NET0131 , \u0_uk_K_r9_reg[33]/NET0131 , \u0_uk_K_r9_reg[34]/NET0131 , \u0_uk_K_r9_reg[35]/NET0131 , \u0_uk_K_r9_reg[36]/NET0131 , \u0_uk_K_r9_reg[37]/NET0131 , \u0_uk_K_r9_reg[38]/NET0131 , \u0_uk_K_r9_reg[39]/NET0131 , \u0_uk_K_r9_reg[3]/NET0131 , \u0_uk_K_r9_reg[40]/NET0131 , \u0_uk_K_r9_reg[41]/NET0131 , \u0_uk_K_r9_reg[42]/NET0131 , \u0_uk_K_r9_reg[43]/NET0131 , \u0_uk_K_r9_reg[44]/NET0131 , \u0_uk_K_r9_reg[45]/NET0131 , \u0_uk_K_r9_reg[46]/NET0131 , \u0_uk_K_r9_reg[47]/NET0131 , \u0_uk_K_r9_reg[48]/NET0131 , \u0_uk_K_r9_reg[49]/NET0131 , \u0_uk_K_r9_reg[4]/NET0131 , \u0_uk_K_r9_reg[50]/NET0131 , \u0_uk_K_r9_reg[51]/NET0131 , \u0_uk_K_r9_reg[52]/NET0131 , \u0_uk_K_r9_reg[53]/NET0131 , \u0_uk_K_r9_reg[54]/NET0131 , \u0_uk_K_r9_reg[55]/NET0131 , \u0_uk_K_r9_reg[5]/NET0131 , \u0_uk_K_r9_reg[6]/NET0131 , \u0_uk_K_r9_reg[7]/NET0131 , \u0_uk_K_r9_reg[8]/NET0131 , \u0_uk_K_r9_reg[9]/NET0131 , \u1_L0_reg[10]/NET0131 , \u1_L0_reg[11]/NET0131 , \u1_L0_reg[12]/NET0131 , \u1_L0_reg[13]/NET0131 , \u1_L0_reg[14]/NET0131 , \u1_L0_reg[15]/P0001 , \u1_L0_reg[16]/NET0131 , \u1_L0_reg[17]/NET0131 , \u1_L0_reg[18]/NET0131 , \u1_L0_reg[19]/NET0131 , \u1_L0_reg[1]/NET0131 , \u1_L0_reg[20]/NET0131 , \u1_L0_reg[21]/NET0131 , \u1_L0_reg[22]/NET0131 , \u1_L0_reg[23]/NET0131 , \u1_L0_reg[24]/NET0131 , \u1_L0_reg[25]/NET0131 , \u1_L0_reg[26]/NET0131 , \u1_L0_reg[27]/NET0131 , \u1_L0_reg[28]/NET0131 , \u1_L0_reg[29]/NET0131 , \u1_L0_reg[2]/NET0131 , \u1_L0_reg[30]/NET0131 , \u1_L0_reg[31]/NET0131 , \u1_L0_reg[32]/NET0131 , \u1_L0_reg[3]/NET0131 , \u1_L0_reg[4]/NET0131 , \u1_L0_reg[5]/NET0131 , \u1_L0_reg[6]/NET0131 , \u1_L0_reg[7]/NET0131 , \u1_L0_reg[8]/NET0131 , \u1_L0_reg[9]/NET0131 , \u1_L10_reg[10]/NET0131 , \u1_L10_reg[11]/NET0131 , \u1_L10_reg[12]/NET0131 , \u1_L10_reg[13]/NET0131 , \u1_L10_reg[14]/NET0131 , \u1_L10_reg[15]/P0001 , \u1_L10_reg[16]/NET0131 , \u1_L10_reg[17]/NET0131 , \u1_L10_reg[18]/P0001 , \u1_L10_reg[19]/P0001 , \u1_L10_reg[1]/NET0131 , \u1_L10_reg[20]/NET0131 , \u1_L10_reg[21]/NET0131 , \u1_L10_reg[22]/NET0131 , \u1_L10_reg[23]/NET0131 , \u1_L10_reg[24]/NET0131 , \u1_L10_reg[25]/NET0131 , \u1_L10_reg[26]/NET0131 , \u1_L10_reg[27]/NET0131 , \u1_L10_reg[28]/NET0131 , \u1_L10_reg[29]/NET0131 , \u1_L10_reg[2]/NET0131 , \u1_L10_reg[30]/NET0131 , \u1_L10_reg[31]/NET0131 , \u1_L10_reg[32]/NET0131 , \u1_L10_reg[3]/NET0131 , \u1_L10_reg[4]/NET0131 , \u1_L10_reg[5]/NET0131 , \u1_L10_reg[6]/NET0131 , \u1_L10_reg[7]/NET0131 , \u1_L10_reg[8]/NET0131 , \u1_L10_reg[9]/NET0131 , \u1_L11_reg[10]/NET0131 , \u1_L11_reg[11]/NET0131 , \u1_L11_reg[12]/NET0131 , \u1_L11_reg[13]/NET0131 , \u1_L11_reg[14]/NET0131 , \u1_L11_reg[15]/P0001 , \u1_L11_reg[16]/NET0131 , \u1_L11_reg[17]/NET0131 , \u1_L11_reg[18]/P0001 , \u1_L11_reg[19]/P0001 , \u1_L11_reg[1]/NET0131 , \u1_L11_reg[20]/NET0131 , \u1_L11_reg[21]/NET0131 , \u1_L11_reg[22]/NET0131 , \u1_L11_reg[23]/NET0131 , \u1_L11_reg[24]/NET0131 , \u1_L11_reg[25]/NET0131 , \u1_L11_reg[26]/NET0131 , \u1_L11_reg[27]/NET0131 , \u1_L11_reg[28]/NET0131 , \u1_L11_reg[29]/NET0131 , \u1_L11_reg[2]/NET0131 , \u1_L11_reg[30]/NET0131 , \u1_L11_reg[31]/NET0131 , \u1_L11_reg[32]/NET0131 , \u1_L11_reg[3]/NET0131 , \u1_L11_reg[4]/NET0131 , \u1_L11_reg[5]/NET0131 , \u1_L11_reg[6]/NET0131 , \u1_L11_reg[7]/NET0131 , \u1_L11_reg[8]/NET0131 , \u1_L11_reg[9]/NET0131 , \u1_L12_reg[10]/NET0131 , \u1_L12_reg[11]/NET0131 , \u1_L12_reg[12]/NET0131 , \u1_L12_reg[13]/NET0131 , \u1_L12_reg[14]/NET0131 , \u1_L12_reg[15]/P0001 , \u1_L12_reg[16]/NET0131 , \u1_L12_reg[17]/NET0131 , \u1_L12_reg[18]/P0001 , \u1_L12_reg[19]/NET0131 , \u1_L12_reg[1]/NET0131 , \u1_L12_reg[20]/NET0131 , \u1_L12_reg[21]/NET0131 , \u1_L12_reg[22]/NET0131 , \u1_L12_reg[23]/P0001 , \u1_L12_reg[24]/NET0131 , \u1_L12_reg[25]/NET0131 , \u1_L12_reg[26]/NET0131 , \u1_L12_reg[27]/NET0131 , \u1_L12_reg[28]/NET0131 , \u1_L12_reg[29]/NET0131 , \u1_L12_reg[2]/NET0131 , \u1_L12_reg[30]/NET0131 , \u1_L12_reg[31]/NET0131 , \u1_L12_reg[32]/NET0131 , \u1_L12_reg[3]/NET0131 , \u1_L12_reg[4]/NET0131 , \u1_L12_reg[5]/NET0131 , \u1_L12_reg[6]/NET0131 , \u1_L12_reg[7]/NET0131 , \u1_L12_reg[8]/NET0131 , \u1_L12_reg[9]/NET0131 , \u1_L13_reg[10]/NET0131 , \u1_L13_reg[11]/NET0131 , \u1_L13_reg[12]/NET0131 , \u1_L13_reg[13]/NET0131 , \u1_L13_reg[14]/NET0131 , \u1_L13_reg[15]/P0001 , \u1_L13_reg[16]/NET0131 , \u1_L13_reg[17]/NET0131 , \u1_L13_reg[18]/P0001 , \u1_L13_reg[19]/P0001 , \u1_L13_reg[1]/NET0131 , \u1_L13_reg[20]/NET0131 , \u1_L13_reg[21]/NET0131 , \u1_L13_reg[22]/NET0131 , \u1_L13_reg[23]/P0001 , \u1_L13_reg[24]/NET0131 , \u1_L13_reg[25]/NET0131 , \u1_L13_reg[26]/NET0131 , \u1_L13_reg[27]/NET0131 , \u1_L13_reg[28]/NET0131 , \u1_L13_reg[29]/NET0131 , \u1_L13_reg[2]/NET0131 , \u1_L13_reg[30]/NET0131 , \u1_L13_reg[31]/NET0131 , \u1_L13_reg[32]/NET0131 , \u1_L13_reg[3]/NET0131 , \u1_L13_reg[4]/NET0131 , \u1_L13_reg[5]/NET0131 , \u1_L13_reg[6]/NET0131 , \u1_L13_reg[7]/NET0131 , \u1_L13_reg[8]/NET0131 , \u1_L13_reg[9]/NET0131 , \u1_L14_reg[10]/P0001 , \u1_L14_reg[11]/P0001 , \u1_L14_reg[12]/P0001 , \u1_L14_reg[13]/P0001 , \u1_L14_reg[14]/P0001 , \u1_L14_reg[15]/P0001 , \u1_L14_reg[16]/P0001 , \u1_L14_reg[17]/P0001 , \u1_L14_reg[18]/P0001 , \u1_L14_reg[19]/P0001 , \u1_L14_reg[1]/P0001 , \u1_L14_reg[20]/P0001 , \u1_L14_reg[21]/P0001 , \u1_L14_reg[22]/P0001 , \u1_L14_reg[23]/P0001 , \u1_L14_reg[24]/P0001 , \u1_L14_reg[25]/P0001 , \u1_L14_reg[26]/P0001 , \u1_L14_reg[27]/P0001 , \u1_L14_reg[28]/P0001 , \u1_L14_reg[29]/P0001 , \u1_L14_reg[2]/P0001 , \u1_L14_reg[30]/P0001 , \u1_L14_reg[31]/P0001 , \u1_L14_reg[32]/P0001 , \u1_L14_reg[3]/P0001 , \u1_L14_reg[4]/P0001 , \u1_L14_reg[5]/P0001 , \u1_L14_reg[6]/P0001 , \u1_L14_reg[7]/P0001 , \u1_L14_reg[8]/P0001 , \u1_L14_reg[9]/P0001 , \u1_L1_reg[10]/NET0131 , \u1_L1_reg[11]/NET0131 , \u1_L1_reg[12]/NET0131 , \u1_L1_reg[13]/NET0131 , \u1_L1_reg[14]/NET0131 , \u1_L1_reg[15]/P0001 , \u1_L1_reg[16]/NET0131 , \u1_L1_reg[17]/NET0131 , \u1_L1_reg[18]/NET0131 , \u1_L1_reg[19]/P0001 , \u1_L1_reg[1]/NET0131 , \u1_L1_reg[20]/NET0131 , \u1_L1_reg[21]/NET0131 , \u1_L1_reg[22]/NET0131 , \u1_L1_reg[23]/NET0131 , \u1_L1_reg[24]/NET0131 , \u1_L1_reg[25]/NET0131 , \u1_L1_reg[26]/NET0131 , \u1_L1_reg[27]/NET0131 , \u1_L1_reg[28]/NET0131 , \u1_L1_reg[29]/NET0131 , \u1_L1_reg[2]/NET0131 , \u1_L1_reg[30]/NET0131 , \u1_L1_reg[31]/NET0131 , \u1_L1_reg[32]/NET0131 , \u1_L1_reg[3]/NET0131 , \u1_L1_reg[4]/NET0131 , \u1_L1_reg[5]/NET0131 , \u1_L1_reg[6]/NET0131 , \u1_L1_reg[7]/NET0131 , \u1_L1_reg[8]/NET0131 , \u1_L1_reg[9]/NET0131 , \u1_L2_reg[10]/NET0131 , \u1_L2_reg[11]/NET0131 , \u1_L2_reg[12]/NET0131 , \u1_L2_reg[13]/NET0131 , \u1_L2_reg[14]/NET0131 , \u1_L2_reg[15]/P0001 , \u1_L2_reg[16]/NET0131 , \u1_L2_reg[17]/NET0131 , \u1_L2_reg[18]/NET0131 , \u1_L2_reg[19]/NET0131 , \u1_L2_reg[1]/NET0131 , \u1_L2_reg[20]/NET0131 , \u1_L2_reg[21]/NET0131 , \u1_L2_reg[22]/NET0131 , \u1_L2_reg[23]/NET0131 , \u1_L2_reg[24]/NET0131 , \u1_L2_reg[25]/NET0131 , \u1_L2_reg[26]/NET0131 , \u1_L2_reg[27]/NET0131 , \u1_L2_reg[28]/NET0131 , \u1_L2_reg[29]/NET0131 , \u1_L2_reg[2]/NET0131 , \u1_L2_reg[30]/NET0131 , \u1_L2_reg[31]/NET0131 , \u1_L2_reg[32]/NET0131 , \u1_L2_reg[3]/NET0131 , \u1_L2_reg[4]/NET0131 , \u1_L2_reg[5]/NET0131 , \u1_L2_reg[6]/NET0131 , \u1_L2_reg[7]/NET0131 , \u1_L2_reg[8]/NET0131 , \u1_L2_reg[9]/NET0131 , \u1_L3_reg[10]/NET0131 , \u1_L3_reg[11]/NET0131 , \u1_L3_reg[12]/NET0131 , \u1_L3_reg[13]/NET0131 , \u1_L3_reg[14]/NET0131 , \u1_L3_reg[15]/P0001 , \u1_L3_reg[16]/NET0131 , \u1_L3_reg[17]/NET0131 , \u1_L3_reg[18]/NET0131 , \u1_L3_reg[19]/NET0131 , \u1_L3_reg[1]/NET0131 , \u1_L3_reg[20]/NET0131 , \u1_L3_reg[21]/NET0131 , \u1_L3_reg[22]/NET0131 , \u1_L3_reg[23]/NET0131 , \u1_L3_reg[24]/NET0131 , \u1_L3_reg[25]/NET0131 , \u1_L3_reg[26]/NET0131 , \u1_L3_reg[27]/NET0131 , \u1_L3_reg[28]/NET0131 , \u1_L3_reg[29]/NET0131 , \u1_L3_reg[2]/NET0131 , \u1_L3_reg[30]/NET0131 , \u1_L3_reg[31]/NET0131 , \u1_L3_reg[32]/NET0131 , \u1_L3_reg[3]/NET0131 , \u1_L3_reg[4]/NET0131 , \u1_L3_reg[5]/NET0131 , \u1_L3_reg[6]/NET0131 , \u1_L3_reg[7]/NET0131 , \u1_L3_reg[8]/NET0131 , \u1_L3_reg[9]/NET0131 , \u1_L4_reg[10]/NET0131 , \u1_L4_reg[11]/P0001 , \u1_L4_reg[12]/NET0131 , \u1_L4_reg[13]/NET0131 , \u1_L4_reg[14]/NET0131 , \u1_L4_reg[15]/P0001 , \u1_L4_reg[16]/NET0131 , \u1_L4_reg[17]/NET0131 , \u1_L4_reg[18]/NET0131 , \u1_L4_reg[19]/P0001 , \u1_L4_reg[1]/NET0131 , \u1_L4_reg[20]/NET0131 , \u1_L4_reg[21]/NET0131 , \u1_L4_reg[22]/NET0131 , \u1_L4_reg[23]/NET0131 , \u1_L4_reg[24]/NET0131 , \u1_L4_reg[25]/NET0131 , \u1_L4_reg[26]/NET0131 , \u1_L4_reg[27]/NET0131 , \u1_L4_reg[28]/NET0131 , \u1_L4_reg[29]/NET0131 , \u1_L4_reg[2]/NET0131 , \u1_L4_reg[30]/NET0131 , \u1_L4_reg[31]/NET0131 , \u1_L4_reg[32]/NET0131 , \u1_L4_reg[3]/NET0131 , \u1_L4_reg[4]/NET0131 , \u1_L4_reg[5]/NET0131 , \u1_L4_reg[6]/NET0131 , \u1_L4_reg[7]/NET0131 , \u1_L4_reg[8]/NET0131 , \u1_L4_reg[9]/NET0131 , \u1_L5_reg[10]/NET0131 , \u1_L5_reg[11]/NET0131 , \u1_L5_reg[12]/NET0131 , \u1_L5_reg[13]/NET0131 , \u1_L5_reg[14]/NET0131 , \u1_L5_reg[15]/P0001 , \u1_L5_reg[16]/NET0131 , \u1_L5_reg[17]/NET0131 , \u1_L5_reg[18]/NET0131 , \u1_L5_reg[19]/NET0131 , \u1_L5_reg[1]/NET0131 , \u1_L5_reg[20]/NET0131 , \u1_L5_reg[21]/NET0131 , \u1_L5_reg[22]/NET0131 , \u1_L5_reg[23]/NET0131 , \u1_L5_reg[24]/NET0131 , \u1_L5_reg[25]/NET0131 , \u1_L5_reg[26]/NET0131 , \u1_L5_reg[27]/NET0131 , \u1_L5_reg[28]/NET0131 , \u1_L5_reg[29]/NET0131 , \u1_L5_reg[2]/NET0131 , \u1_L5_reg[30]/NET0131 , \u1_L5_reg[31]/NET0131 , \u1_L5_reg[32]/NET0131 , \u1_L5_reg[3]/NET0131 , \u1_L5_reg[4]/NET0131 , \u1_L5_reg[5]/NET0131 , \u1_L5_reg[6]/NET0131 , \u1_L5_reg[7]/NET0131 , \u1_L5_reg[8]/NET0131 , \u1_L5_reg[9]/NET0131 , \u1_L6_reg[10]/NET0131 , \u1_L6_reg[11]/NET0131 , \u1_L6_reg[12]/NET0131 , \u1_L6_reg[13]/NET0131 , \u1_L6_reg[14]/NET0131 , \u1_L6_reg[15]/P0001 , \u1_L6_reg[16]/NET0131 , \u1_L6_reg[17]/NET0131 , \u1_L6_reg[18]/NET0131 , \u1_L6_reg[19]/NET0131 , \u1_L6_reg[1]/NET0131 , \u1_L6_reg[20]/NET0131 , \u1_L6_reg[21]/NET0131 , \u1_L6_reg[22]/NET0131 , \u1_L6_reg[23]/NET0131 , \u1_L6_reg[24]/NET0131 , \u1_L6_reg[25]/NET0131 , \u1_L6_reg[26]/NET0131 , \u1_L6_reg[27]/NET0131 , \u1_L6_reg[28]/NET0131 , \u1_L6_reg[29]/NET0131 , \u1_L6_reg[2]/NET0131 , \u1_L6_reg[30]/NET0131 , \u1_L6_reg[31]/NET0131 , \u1_L6_reg[32]/NET0131 , \u1_L6_reg[3]/NET0131 , \u1_L6_reg[4]/NET0131 , \u1_L6_reg[5]/NET0131 , \u1_L6_reg[6]/NET0131 , \u1_L6_reg[7]/NET0131 , \u1_L6_reg[8]/NET0131 , \u1_L6_reg[9]/NET0131 , \u1_L7_reg[10]/NET0131 , \u1_L7_reg[11]/NET0131 , \u1_L7_reg[12]/NET0131 , \u1_L7_reg[13]/NET0131 , \u1_L7_reg[14]/NET0131 , \u1_L7_reg[15]/P0001 , \u1_L7_reg[16]/NET0131 , \u1_L7_reg[17]/NET0131 , \u1_L7_reg[18]/NET0131 , \u1_L7_reg[19]/P0001 , \u1_L7_reg[1]/NET0131 , \u1_L7_reg[20]/NET0131 , \u1_L7_reg[21]/NET0131 , \u1_L7_reg[22]/NET0131 , \u1_L7_reg[23]/NET0131 , \u1_L7_reg[24]/NET0131 , \u1_L7_reg[25]/NET0131 , \u1_L7_reg[26]/NET0131 , \u1_L7_reg[27]/NET0131 , \u1_L7_reg[28]/NET0131 , \u1_L7_reg[29]/NET0131 , \u1_L7_reg[2]/NET0131 , \u1_L7_reg[30]/NET0131 , \u1_L7_reg[31]/NET0131 , \u1_L7_reg[32]/NET0131 , \u1_L7_reg[3]/NET0131 , \u1_L7_reg[4]/NET0131 , \u1_L7_reg[5]/NET0131 , \u1_L7_reg[6]/NET0131 , \u1_L7_reg[7]/NET0131 , \u1_L7_reg[8]/NET0131 , \u1_L7_reg[9]/NET0131 , \u1_L8_reg[10]/NET0131 , \u1_L8_reg[11]/NET0131 , \u1_L8_reg[12]/NET0131 , \u1_L8_reg[13]/NET0131 , \u1_L8_reg[14]/NET0131 , \u1_L8_reg[15]/P0001 , \u1_L8_reg[16]/NET0131 , \u1_L8_reg[17]/NET0131 , \u1_L8_reg[18]/NET0131 , \u1_L8_reg[19]/P0001 , \u1_L8_reg[1]/NET0131 , \u1_L8_reg[20]/NET0131 , \u1_L8_reg[21]/NET0131 , \u1_L8_reg[22]/NET0131 , \u1_L8_reg[23]/NET0131 , \u1_L8_reg[24]/NET0131 , \u1_L8_reg[25]/NET0131 , \u1_L8_reg[26]/NET0131 , \u1_L8_reg[27]/NET0131 , \u1_L8_reg[28]/NET0131 , \u1_L8_reg[29]/NET0131 , \u1_L8_reg[2]/NET0131 , \u1_L8_reg[30]/NET0131 , \u1_L8_reg[31]/NET0131 , \u1_L8_reg[32]/NET0131 , \u1_L8_reg[3]/NET0131 , \u1_L8_reg[4]/NET0131 , \u1_L8_reg[5]/NET0131 , \u1_L8_reg[6]/NET0131 , \u1_L8_reg[7]/NET0131 , \u1_L8_reg[8]/NET0131 , \u1_L8_reg[9]/NET0131 , \u1_L9_reg[10]/NET0131 , \u1_L9_reg[11]/NET0131 , \u1_L9_reg[12]/NET0131 , \u1_L9_reg[13]/NET0131 , \u1_L9_reg[14]/NET0131 , \u1_L9_reg[15]/P0001 , \u1_L9_reg[16]/NET0131 , \u1_L9_reg[17]/NET0131 , \u1_L9_reg[18]/P0001 , \u1_L9_reg[19]/NET0131 , \u1_L9_reg[1]/NET0131 , \u1_L9_reg[20]/NET0131 , \u1_L9_reg[21]/NET0131 , \u1_L9_reg[22]/NET0131 , \u1_L9_reg[23]/NET0131 , \u1_L9_reg[24]/NET0131 , \u1_L9_reg[25]/NET0131 , \u1_L9_reg[26]/NET0131 , \u1_L9_reg[27]/NET0131 , \u1_L9_reg[28]/NET0131 , \u1_L9_reg[29]/NET0131 , \u1_L9_reg[2]/NET0131 , \u1_L9_reg[30]/NET0131 , \u1_L9_reg[31]/NET0131 , \u1_L9_reg[32]/NET0131 , \u1_L9_reg[3]/NET0131 , \u1_L9_reg[4]/NET0131 , \u1_L9_reg[5]/NET0131 , \u1_L9_reg[6]/NET0131 , \u1_L9_reg[7]/NET0131 , \u1_L9_reg[8]/NET0131 , \u1_L9_reg[9]/NET0131 , \u1_R0_reg[10]/NET0131 , \u1_R0_reg[11]/NET0131 , \u1_R0_reg[12]/NET0131 , \u1_R0_reg[13]/NET0131 , \u1_R0_reg[14]/NET0131 , \u1_R0_reg[15]/NET0131 , \u1_R0_reg[16]/NET0131 , \u1_R0_reg[17]/NET0131 , \u1_R0_reg[18]/NET0131 , \u1_R0_reg[19]/NET0131 , \u1_R0_reg[1]/NET0131 , \u1_R0_reg[20]/NET0131 , \u1_R0_reg[21]/NET0131 , \u1_R0_reg[22]/NET0131 , \u1_R0_reg[23]/NET0131 , \u1_R0_reg[24]/NET0131 , \u1_R0_reg[25]/NET0131 , \u1_R0_reg[26]/NET0131 , \u1_R0_reg[27]/NET0131 , \u1_R0_reg[28]/NET0131 , \u1_R0_reg[29]/NET0131 , \u1_R0_reg[2]/NET0131 , \u1_R0_reg[30]/NET0131 , \u1_R0_reg[31]/P0001 , \u1_R0_reg[32]/NET0131 , \u1_R0_reg[3]/NET0131 , \u1_R0_reg[4]/NET0131 , \u1_R0_reg[5]/NET0131 , \u1_R0_reg[6]/NET0131 , \u1_R0_reg[7]/NET0131 , \u1_R0_reg[8]/NET0131 , \u1_R0_reg[9]/NET0131 , \u1_R10_reg[10]/NET0131 , \u1_R10_reg[11]/NET0131 , \u1_R10_reg[12]/NET0131 , \u1_R10_reg[13]/NET0131 , \u1_R10_reg[14]/NET0131 , \u1_R10_reg[15]/NET0131 , \u1_R10_reg[16]/NET0131 , \u1_R10_reg[17]/NET0131 , \u1_R10_reg[18]/NET0131 , \u1_R10_reg[19]/NET0131 , \u1_R10_reg[1]/NET0131 , \u1_R10_reg[20]/NET0131 , \u1_R10_reg[21]/NET0131 , \u1_R10_reg[22]/NET0131 , \u1_R10_reg[23]/NET0131 , \u1_R10_reg[24]/NET0131 , \u1_R10_reg[25]/NET0131 , \u1_R10_reg[26]/NET0131 , \u1_R10_reg[27]/NET0131 , \u1_R10_reg[28]/NET0131 , \u1_R10_reg[29]/NET0131 , \u1_R10_reg[2]/NET0131 , \u1_R10_reg[30]/NET0131 , \u1_R10_reg[31]/P0001 , \u1_R10_reg[32]/NET0131 , \u1_R10_reg[3]/NET0131 , \u1_R10_reg[4]/NET0131 , \u1_R10_reg[5]/NET0131 , \u1_R10_reg[6]/NET0131 , \u1_R10_reg[7]/NET0131 , \u1_R10_reg[8]/NET0131 , \u1_R10_reg[9]/NET0131 , \u1_R11_reg[10]/NET0131 , \u1_R11_reg[11]/NET0131 , \u1_R11_reg[12]/NET0131 , \u1_R11_reg[13]/NET0131 , \u1_R11_reg[14]/NET0131 , \u1_R11_reg[15]/NET0131 , \u1_R11_reg[16]/NET0131 , \u1_R11_reg[17]/NET0131 , \u1_R11_reg[18]/NET0131 , \u1_R11_reg[19]/NET0131 , \u1_R11_reg[1]/NET0131 , \u1_R11_reg[20]/NET0131 , \u1_R11_reg[21]/NET0131 , \u1_R11_reg[22]/NET0131 , \u1_R11_reg[23]/NET0131 , \u1_R11_reg[24]/NET0131 , \u1_R11_reg[25]/NET0131 , \u1_R11_reg[26]/NET0131 , \u1_R11_reg[27]/NET0131 , \u1_R11_reg[28]/NET0131 , \u1_R11_reg[29]/NET0131 , \u1_R11_reg[2]/NET0131 , \u1_R11_reg[30]/NET0131 , \u1_R11_reg[31]/NET0131 , \u1_R11_reg[32]/NET0131 , \u1_R11_reg[3]/NET0131 , \u1_R11_reg[4]/NET0131 , \u1_R11_reg[5]/NET0131 , \u1_R11_reg[6]/NET0131 , \u1_R11_reg[7]/NET0131 , \u1_R11_reg[8]/NET0131 , \u1_R11_reg[9]/NET0131 , \u1_R12_reg[10]/NET0131 , \u1_R12_reg[11]/NET0131 , \u1_R12_reg[12]/NET0131 , \u1_R12_reg[13]/NET0131 , \u1_R12_reg[14]/NET0131 , \u1_R12_reg[15]/NET0131 , \u1_R12_reg[16]/NET0131 , \u1_R12_reg[17]/NET0131 , \u1_R12_reg[18]/NET0131 , \u1_R12_reg[19]/NET0131 , \u1_R12_reg[1]/NET0131 , \u1_R12_reg[20]/NET0131 , \u1_R12_reg[21]/NET0131 , \u1_R12_reg[22]/NET0131 , \u1_R12_reg[23]/NET0131 , \u1_R12_reg[24]/NET0131 , \u1_R12_reg[25]/NET0131 , \u1_R12_reg[26]/NET0131 , \u1_R12_reg[27]/NET0131 , \u1_R12_reg[28]/NET0131 , \u1_R12_reg[29]/NET0131 , \u1_R12_reg[2]/NET0131 , \u1_R12_reg[30]/NET0131 , \u1_R12_reg[31]/NET0131 , \u1_R12_reg[32]/NET0131 , \u1_R12_reg[3]/NET0131 , \u1_R12_reg[4]/NET0131 , \u1_R12_reg[5]/NET0131 , \u1_R12_reg[6]/NET0131 , \u1_R12_reg[7]/NET0131 , \u1_R12_reg[8]/NET0131 , \u1_R12_reg[9]/NET0131 , \u1_R13_reg[10]/NET0131 , \u1_R13_reg[11]/P0001 , \u1_R13_reg[12]/NET0131 , \u1_R13_reg[13]/NET0131 , \u1_R13_reg[14]/NET0131 , \u1_R13_reg[15]/NET0131 , \u1_R13_reg[16]/NET0131 , \u1_R13_reg[17]/NET0131 , \u1_R13_reg[18]/NET0131 , \u1_R13_reg[19]/NET0131 , \u1_R13_reg[1]/NET0131 , \u1_R13_reg[20]/NET0131 , \u1_R13_reg[21]/NET0131 , \u1_R13_reg[22]/NET0131 , \u1_R13_reg[23]/P0001 , \u1_R13_reg[24]/NET0131 , \u1_R13_reg[25]/NET0131 , \u1_R13_reg[26]/NET0131 , \u1_R13_reg[27]/P0001 , \u1_R13_reg[28]/NET0131 , \u1_R13_reg[29]/NET0131 , \u1_R13_reg[2]/NET0131 , \u1_R13_reg[30]/NET0131 , \u1_R13_reg[31]/P0001 , \u1_R13_reg[32]/NET0131 , \u1_R13_reg[3]/NET0131 , \u1_R13_reg[4]/NET0131 , \u1_R13_reg[5]/NET0131 , \u1_R13_reg[6]/NET0131 , \u1_R13_reg[7]/NET0131 , \u1_R13_reg[8]/NET0131 , \u1_R13_reg[9]/NET0131 , \u1_R14_reg[10]/P0001 , \u1_R14_reg[11]/P0001 , \u1_R14_reg[12]/NET0131 , \u1_R14_reg[13]/NET0131 , \u1_R14_reg[14]/NET0131 , \u1_R14_reg[15]/NET0131 , \u1_R14_reg[16]/NET0131 , \u1_R14_reg[17]/NET0131 , \u1_R14_reg[18]/NET0131 , \u1_R14_reg[19]/P0001 , \u1_R14_reg[1]/NET0131 , \u1_R14_reg[20]/NET0131 , \u1_R14_reg[21]/NET0131 , \u1_R14_reg[22]/P0001 , \u1_R14_reg[23]/P0001 , \u1_R14_reg[24]/NET0131 , \u1_R14_reg[25]/NET0131 , \u1_R14_reg[26]/NET0131 , \u1_R14_reg[27]/P0001 , \u1_R14_reg[28]/NET0131 , \u1_R14_reg[29]/NET0131 , \u1_R14_reg[2]/NET0131 , \u1_R14_reg[30]/NET0131 , \u1_R14_reg[31]/P0001 , \u1_R14_reg[32]/NET0131 , \u1_R14_reg[3]/NET0131 , \u1_R14_reg[4]/NET0131 , \u1_R14_reg[5]/NET0131 , \u1_R14_reg[6]/NET0131 , \u1_R14_reg[7]/P0001 , \u1_R14_reg[8]/NET0131 , \u1_R14_reg[9]/NET0131 , \u1_R1_reg[10]/NET0131 , \u1_R1_reg[11]/NET0131 , \u1_R1_reg[12]/NET0131 , \u1_R1_reg[13]/NET0131 , \u1_R1_reg[14]/NET0131 , \u1_R1_reg[15]/NET0131 , \u1_R1_reg[16]/NET0131 , \u1_R1_reg[17]/NET0131 , \u1_R1_reg[18]/NET0131 , \u1_R1_reg[19]/NET0131 , \u1_R1_reg[1]/NET0131 , \u1_R1_reg[20]/NET0131 , \u1_R1_reg[21]/NET0131 , \u1_R1_reg[22]/NET0131 , \u1_R1_reg[23]/NET0131 , \u1_R1_reg[24]/NET0131 , \u1_R1_reg[25]/NET0131 , \u1_R1_reg[26]/NET0131 , \u1_R1_reg[27]/NET0131 , \u1_R1_reg[28]/NET0131 , \u1_R1_reg[29]/NET0131 , \u1_R1_reg[2]/NET0131 , \u1_R1_reg[30]/NET0131 , \u1_R1_reg[31]/P0001 , \u1_R1_reg[32]/NET0131 , \u1_R1_reg[3]/NET0131 , \u1_R1_reg[4]/NET0131 , \u1_R1_reg[5]/NET0131 , \u1_R1_reg[6]/NET0131 , \u1_R1_reg[7]/NET0131 , \u1_R1_reg[8]/NET0131 , \u1_R1_reg[9]/NET0131 , \u1_R2_reg[10]/NET0131 , \u1_R2_reg[11]/NET0131 , \u1_R2_reg[12]/NET0131 , \u1_R2_reg[13]/NET0131 , \u1_R2_reg[14]/NET0131 , \u1_R2_reg[15]/NET0131 , \u1_R2_reg[16]/NET0131 , \u1_R2_reg[17]/NET0131 , \u1_R2_reg[18]/NET0131 , \u1_R2_reg[19]/NET0131 , \u1_R2_reg[1]/NET0131 , \u1_R2_reg[20]/NET0131 , \u1_R2_reg[21]/NET0131 , \u1_R2_reg[22]/NET0131 , \u1_R2_reg[23]/NET0131 , \u1_R2_reg[24]/NET0131 , \u1_R2_reg[25]/NET0131 , \u1_R2_reg[26]/NET0131 , \u1_R2_reg[27]/NET0131 , \u1_R2_reg[28]/NET0131 , \u1_R2_reg[29]/NET0131 , \u1_R2_reg[2]/NET0131 , \u1_R2_reg[30]/NET0131 , \u1_R2_reg[31]/P0001 , \u1_R2_reg[32]/NET0131 , \u1_R2_reg[3]/NET0131 , \u1_R2_reg[4]/NET0131 , \u1_R2_reg[5]/NET0131 , \u1_R2_reg[6]/NET0131 , \u1_R2_reg[7]/NET0131 , \u1_R2_reg[8]/NET0131 , \u1_R2_reg[9]/NET0131 , \u1_R3_reg[10]/NET0131 , \u1_R3_reg[11]/NET0131 , \u1_R3_reg[12]/NET0131 , \u1_R3_reg[13]/NET0131 , \u1_R3_reg[14]/NET0131 , \u1_R3_reg[15]/NET0131 , \u1_R3_reg[16]/NET0131 , \u1_R3_reg[17]/NET0131 , \u1_R3_reg[18]/NET0131 , \u1_R3_reg[19]/NET0131 , \u1_R3_reg[1]/NET0131 , \u1_R3_reg[20]/NET0131 , \u1_R3_reg[21]/NET0131 , \u1_R3_reg[22]/NET0131 , \u1_R3_reg[23]/NET0131 , \u1_R3_reg[24]/NET0131 , \u1_R3_reg[25]/NET0131 , \u1_R3_reg[26]/NET0131 , \u1_R3_reg[27]/NET0131 , \u1_R3_reg[28]/NET0131 , \u1_R3_reg[29]/NET0131 , \u1_R3_reg[2]/NET0131 , \u1_R3_reg[30]/NET0131 , \u1_R3_reg[31]/P0001 , \u1_R3_reg[32]/NET0131 , \u1_R3_reg[3]/NET0131 , \u1_R3_reg[4]/NET0131 , \u1_R3_reg[5]/NET0131 , \u1_R3_reg[6]/NET0131 , \u1_R3_reg[7]/NET0131 , \u1_R3_reg[8]/NET0131 , \u1_R3_reg[9]/NET0131 , \u1_R4_reg[10]/NET0131 , \u1_R4_reg[11]/P0001 , \u1_R4_reg[12]/NET0131 , \u1_R4_reg[13]/NET0131 , \u1_R4_reg[14]/NET0131 , \u1_R4_reg[15]/NET0131 , \u1_R4_reg[16]/NET0131 , \u1_R4_reg[17]/NET0131 , \u1_R4_reg[18]/NET0131 , \u1_R4_reg[19]/NET0131 , \u1_R4_reg[1]/NET0131 , \u1_R4_reg[20]/NET0131 , \u1_R4_reg[21]/NET0131 , \u1_R4_reg[22]/NET0131 , \u1_R4_reg[23]/NET0131 , \u1_R4_reg[24]/NET0131 , \u1_R4_reg[25]/NET0131 , \u1_R4_reg[26]/NET0131 , \u1_R4_reg[27]/NET0131 , \u1_R4_reg[28]/NET0131 , \u1_R4_reg[29]/NET0131 , \u1_R4_reg[2]/NET0131 , \u1_R4_reg[30]/NET0131 , \u1_R4_reg[31]/P0001 , \u1_R4_reg[32]/NET0131 , \u1_R4_reg[3]/NET0131 , \u1_R4_reg[4]/NET0131 , \u1_R4_reg[5]/NET0131 , \u1_R4_reg[6]/NET0131 , \u1_R4_reg[7]/NET0131 , \u1_R4_reg[8]/NET0131 , \u1_R4_reg[9]/NET0131 , \u1_R5_reg[10]/NET0131 , \u1_R5_reg[11]/NET0131 , \u1_R5_reg[12]/NET0131 , \u1_R5_reg[13]/NET0131 , \u1_R5_reg[14]/NET0131 , \u1_R5_reg[15]/NET0131 , \u1_R5_reg[16]/NET0131 , \u1_R5_reg[17]/NET0131 , \u1_R5_reg[18]/NET0131 , \u1_R5_reg[19]/NET0131 , \u1_R5_reg[1]/NET0131 , \u1_R5_reg[20]/NET0131 , \u1_R5_reg[21]/NET0131 , \u1_R5_reg[22]/NET0131 , \u1_R5_reg[23]/NET0131 , \u1_R5_reg[24]/NET0131 , \u1_R5_reg[25]/NET0131 , \u1_R5_reg[26]/NET0131 , \u1_R5_reg[27]/NET0131 , \u1_R5_reg[28]/NET0131 , \u1_R5_reg[29]/NET0131 , \u1_R5_reg[2]/NET0131 , \u1_R5_reg[30]/NET0131 , \u1_R5_reg[31]/P0001 , \u1_R5_reg[32]/NET0131 , \u1_R5_reg[3]/NET0131 , \u1_R5_reg[4]/NET0131 , \u1_R5_reg[5]/NET0131 , \u1_R5_reg[6]/NET0131 , \u1_R5_reg[7]/NET0131 , \u1_R5_reg[8]/NET0131 , \u1_R5_reg[9]/NET0131 , \u1_R6_reg[10]/NET0131 , \u1_R6_reg[11]/NET0131 , \u1_R6_reg[12]/NET0131 , \u1_R6_reg[13]/NET0131 , \u1_R6_reg[14]/NET0131 , \u1_R6_reg[15]/NET0131 , \u1_R6_reg[16]/NET0131 , \u1_R6_reg[17]/NET0131 , \u1_R6_reg[18]/NET0131 , \u1_R6_reg[19]/NET0131 , \u1_R6_reg[1]/NET0131 , \u1_R6_reg[20]/NET0131 , \u1_R6_reg[21]/NET0131 , \u1_R6_reg[22]/NET0131 , \u1_R6_reg[23]/NET0131 , \u1_R6_reg[24]/NET0131 , \u1_R6_reg[25]/NET0131 , \u1_R6_reg[26]/NET0131 , \u1_R6_reg[27]/NET0131 , \u1_R6_reg[28]/NET0131 , \u1_R6_reg[29]/NET0131 , \u1_R6_reg[2]/NET0131 , \u1_R6_reg[30]/NET0131 , \u1_R6_reg[31]/P0001 , \u1_R6_reg[32]/NET0131 , \u1_R6_reg[3]/NET0131 , \u1_R6_reg[4]/NET0131 , \u1_R6_reg[5]/NET0131 , \u1_R6_reg[6]/NET0131 , \u1_R6_reg[7]/NET0131 , \u1_R6_reg[8]/NET0131 , \u1_R6_reg[9]/NET0131 , \u1_R7_reg[10]/NET0131 , \u1_R7_reg[11]/NET0131 , \u1_R7_reg[12]/NET0131 , \u1_R7_reg[13]/NET0131 , \u1_R7_reg[14]/NET0131 , \u1_R7_reg[15]/NET0131 , \u1_R7_reg[16]/NET0131 , \u1_R7_reg[17]/NET0131 , \u1_R7_reg[18]/NET0131 , \u1_R7_reg[19]/NET0131 , \u1_R7_reg[1]/NET0131 , \u1_R7_reg[20]/NET0131 , \u1_R7_reg[21]/NET0131 , \u1_R7_reg[22]/NET0131 , \u1_R7_reg[23]/NET0131 , \u1_R7_reg[24]/NET0131 , \u1_R7_reg[25]/NET0131 , \u1_R7_reg[26]/NET0131 , \u1_R7_reg[27]/NET0131 , \u1_R7_reg[28]/NET0131 , \u1_R7_reg[29]/NET0131 , \u1_R7_reg[2]/NET0131 , \u1_R7_reg[30]/NET0131 , \u1_R7_reg[31]/P0001 , \u1_R7_reg[32]/NET0131 , \u1_R7_reg[3]/NET0131 , \u1_R7_reg[4]/NET0131 , \u1_R7_reg[5]/NET0131 , \u1_R7_reg[6]/NET0131 , \u1_R7_reg[7]/NET0131 , \u1_R7_reg[8]/NET0131 , \u1_R7_reg[9]/NET0131 , \u1_R8_reg[10]/NET0131 , \u1_R8_reg[11]/NET0131 , \u1_R8_reg[12]/NET0131 , \u1_R8_reg[13]/NET0131 , \u1_R8_reg[14]/NET0131 , \u1_R8_reg[15]/NET0131 , \u1_R8_reg[16]/NET0131 , \u1_R8_reg[17]/NET0131 , \u1_R8_reg[18]/NET0131 , \u1_R8_reg[19]/NET0131 , \u1_R8_reg[1]/NET0131 , \u1_R8_reg[20]/NET0131 , \u1_R8_reg[21]/NET0131 , \u1_R8_reg[22]/NET0131 , \u1_R8_reg[23]/NET0131 , \u1_R8_reg[24]/NET0131 , \u1_R8_reg[25]/NET0131 , \u1_R8_reg[26]/NET0131 , \u1_R8_reg[27]/NET0131 , \u1_R8_reg[28]/NET0131 , \u1_R8_reg[29]/NET0131 , \u1_R8_reg[2]/NET0131 , \u1_R8_reg[30]/NET0131 , \u1_R8_reg[31]/P0001 , \u1_R8_reg[32]/NET0131 , \u1_R8_reg[3]/NET0131 , \u1_R8_reg[4]/NET0131 , \u1_R8_reg[5]/NET0131 , \u1_R8_reg[6]/NET0131 , \u1_R8_reg[7]/NET0131 , \u1_R8_reg[8]/NET0131 , \u1_R8_reg[9]/NET0131 , \u1_R9_reg[10]/NET0131 , \u1_R9_reg[11]/NET0131 , \u1_R9_reg[12]/NET0131 , \u1_R9_reg[13]/NET0131 , \u1_R9_reg[14]/NET0131 , \u1_R9_reg[15]/NET0131 , \u1_R9_reg[16]/NET0131 , \u1_R9_reg[17]/NET0131 , \u1_R9_reg[18]/NET0131 , \u1_R9_reg[19]/NET0131 , \u1_R9_reg[1]/NET0131 , \u1_R9_reg[20]/NET0131 , \u1_R9_reg[21]/NET0131 , \u1_R9_reg[22]/NET0131 , \u1_R9_reg[23]/NET0131 , \u1_R9_reg[24]/NET0131 , \u1_R9_reg[25]/NET0131 , \u1_R9_reg[26]/NET0131 , \u1_R9_reg[27]/NET0131 , \u1_R9_reg[28]/NET0131 , \u1_R9_reg[29]/NET0131 , \u1_R9_reg[2]/NET0131 , \u1_R9_reg[30]/NET0131 , \u1_R9_reg[31]/NET0131 , \u1_R9_reg[32]/NET0131 , \u1_R9_reg[3]/NET0131 , \u1_R9_reg[4]/NET0131 , \u1_R9_reg[5]/NET0131 , \u1_R9_reg[6]/NET0131 , \u1_R9_reg[7]/NET0131 , \u1_R9_reg[8]/NET0131 , \u1_R9_reg[9]/NET0131 , \u1_desIn_r_reg[0]/NET0131 , \u1_desIn_r_reg[10]/NET0131 , \u1_desIn_r_reg[11]/NET0131 , \u1_desIn_r_reg[12]/NET0131 , \u1_desIn_r_reg[13]/NET0131 , \u1_desIn_r_reg[14]/NET0131 , \u1_desIn_r_reg[15]/NET0131 , \u1_desIn_r_reg[16]/NET0131 , \u1_desIn_r_reg[17]/NET0131 , \u1_desIn_r_reg[18]/P0001 , \u1_desIn_r_reg[19]/NET0131 , \u1_desIn_r_reg[1]/NET0131 , \u1_desIn_r_reg[20]/NET0131 , \u1_desIn_r_reg[21]/NET0131 , \u1_desIn_r_reg[22]/NET0131 , \u1_desIn_r_reg[23]/NET0131 , \u1_desIn_r_reg[24]/NET0131 , \u1_desIn_r_reg[25]/NET0131 , \u1_desIn_r_reg[26]/NET0131 , \u1_desIn_r_reg[27]/NET0131 , \u1_desIn_r_reg[28]/NET0131 , \u1_desIn_r_reg[29]/NET0131 , \u1_desIn_r_reg[2]/NET0131 , \u1_desIn_r_reg[30]/NET0131 , \u1_desIn_r_reg[31]/NET0131 , \u1_desIn_r_reg[32]/NET0131 , \u1_desIn_r_reg[33]/NET0131 , \u1_desIn_r_reg[34]/NET0131 , \u1_desIn_r_reg[35]/NET0131 , \u1_desIn_r_reg[36]/NET0131 , \u1_desIn_r_reg[37]/NET0131 , \u1_desIn_r_reg[38]/NET0131 , \u1_desIn_r_reg[39]/NET0131 , \u1_desIn_r_reg[3]/NET0131 , \u1_desIn_r_reg[40]/NET0131 , \u1_desIn_r_reg[41]/NET0131 , \u1_desIn_r_reg[42]/NET0131 , \u1_desIn_r_reg[43]/NET0131 , \u1_desIn_r_reg[44]/NET0131 , \u1_desIn_r_reg[45]/NET0131 , \u1_desIn_r_reg[46]/NET0131 , \u1_desIn_r_reg[47]/NET0131 , \u1_desIn_r_reg[48]/NET0131 , \u1_desIn_r_reg[49]/NET0131 , \u1_desIn_r_reg[4]/NET0131 , \u1_desIn_r_reg[50]/NET0131 , \u1_desIn_r_reg[51]/NET0131 , \u1_desIn_r_reg[52]/P0001 , \u1_desIn_r_reg[53]/NET0131 , \u1_desIn_r_reg[54]/NET0131 , \u1_desIn_r_reg[55]/NET0131 , \u1_desIn_r_reg[56]/NET0131 , \u1_desIn_r_reg[57]/NET0131 , \u1_desIn_r_reg[58]/NET0131 , \u1_desIn_r_reg[59]/NET0131 , \u1_desIn_r_reg[5]/NET0131 , \u1_desIn_r_reg[60]/NET0131 , \u1_desIn_r_reg[61]/NET0131 , \u1_desIn_r_reg[62]/NET0131 , \u1_desIn_r_reg[63]/NET0131 , \u1_desIn_r_reg[6]/NET0131 , \u1_desIn_r_reg[7]/NET0131 , \u1_desIn_r_reg[8]/NET0131 , \u1_desIn_r_reg[9]/NET0131 , \u1_key_r_reg[0]/NET0131 , \u1_key_r_reg[10]/NET0131 , \u1_key_r_reg[11]/NET0131 , \u1_key_r_reg[12]/NET0131 , \u1_key_r_reg[13]/NET0131 , \u1_key_r_reg[14]/NET0131 , \u1_key_r_reg[15]/NET0131 , \u1_key_r_reg[16]/NET0131 , \u1_key_r_reg[17]/NET0131 , \u1_key_r_reg[18]/NET0131 , \u1_key_r_reg[19]/NET0131 , \u1_key_r_reg[1]/NET0131 , \u1_key_r_reg[20]/NET0131 , \u1_key_r_reg[21]/NET0131 , \u1_key_r_reg[22]/NET0131 , \u1_key_r_reg[23]/NET0131 , \u1_key_r_reg[24]/NET0131 , \u1_key_r_reg[25]/NET0131 , \u1_key_r_reg[26]/NET0131 , \u1_key_r_reg[27]/NET0131 , \u1_key_r_reg[28]/NET0131 , \u1_key_r_reg[29]/NET0131 , \u1_key_r_reg[2]/NET0131 , \u1_key_r_reg[30]/NET0131 , \u1_key_r_reg[31]/NET0131 , \u1_key_r_reg[32]/NET0131 , \u1_key_r_reg[33]/NET0131 , \u1_key_r_reg[34]/NET0131 , \u1_key_r_reg[35]/P0001 , \u1_key_r_reg[36]/NET0131 , \u1_key_r_reg[37]/NET0131 , \u1_key_r_reg[38]/NET0131 , \u1_key_r_reg[39]/P0001 , \u1_key_r_reg[3]/NET0131 , \u1_key_r_reg[40]/NET0131 , \u1_key_r_reg[41]/NET0131 , \u1_key_r_reg[42]/P0001 , \u1_key_r_reg[43]/NET0131 , \u1_key_r_reg[44]/NET0131 , \u1_key_r_reg[45]/NET0131 , \u1_key_r_reg[46]/NET0131 , \u1_key_r_reg[47]/NET0131 , \u1_key_r_reg[48]/NET0131 , \u1_key_r_reg[49]/NET0131 , \u1_key_r_reg[4]/NET0131 , \u1_key_r_reg[50]/NET0131 , \u1_key_r_reg[51]/NET0131 , \u1_key_r_reg[52]/NET0131 , \u1_key_r_reg[53]/NET0131 , \u1_key_r_reg[54]/NET0131 , \u1_key_r_reg[55]/NET0131 , \u1_key_r_reg[5]/NET0131 , \u1_key_r_reg[6]/NET0131 , \u1_key_r_reg[7]/NET0131 , \u1_key_r_reg[8]/NET0131 , \u1_key_r_reg[9]/NET0131 , \u1_uk_K_r0_reg[0]/NET0131 , \u1_uk_K_r0_reg[10]/NET0131 , \u1_uk_K_r0_reg[11]/NET0131 , \u1_uk_K_r0_reg[12]/NET0131 , \u1_uk_K_r0_reg[13]/NET0131 , \u1_uk_K_r0_reg[14]/NET0131 , \u1_uk_K_r0_reg[15]/NET0131 , \u1_uk_K_r0_reg[16]/NET0131 , \u1_uk_K_r0_reg[17]/NET0131 , \u1_uk_K_r0_reg[18]/NET0131 , \u1_uk_K_r0_reg[19]/NET0131 , \u1_uk_K_r0_reg[20]/NET0131 , \u1_uk_K_r0_reg[21]/NET0131 , \u1_uk_K_r0_reg[22]/NET0131 , \u1_uk_K_r0_reg[23]/NET0131 , \u1_uk_K_r0_reg[24]/NET0131 , \u1_uk_K_r0_reg[25]/P0001 , \u1_uk_K_r0_reg[26]/NET0131 , \u1_uk_K_r0_reg[27]/NET0131 , \u1_uk_K_r0_reg[28]/NET0131 , \u1_uk_K_r0_reg[29]/NET0131 , \u1_uk_K_r0_reg[2]/NET0131 , \u1_uk_K_r0_reg[30]/NET0131 , \u1_uk_K_r0_reg[31]/NET0131 , \u1_uk_K_r0_reg[32]/NET0131 , \u1_uk_K_r0_reg[33]/NET0131 , \u1_uk_K_r0_reg[34]/NET0131 , \u1_uk_K_r0_reg[35]/NET0131 , \u1_uk_K_r0_reg[36]/NET0131 , \u1_uk_K_r0_reg[37]/NET0131 , \u1_uk_K_r0_reg[38]/NET0131 , \u1_uk_K_r0_reg[39]/NET0131 , \u1_uk_K_r0_reg[3]/NET0131 , \u1_uk_K_r0_reg[40]/NET0131 , \u1_uk_K_r0_reg[41]/NET0131 , \u1_uk_K_r0_reg[42]/NET0131 , \u1_uk_K_r0_reg[43]/NET0131 , \u1_uk_K_r0_reg[44]/NET0131 , \u1_uk_K_r0_reg[45]/NET0131 , \u1_uk_K_r0_reg[46]/NET0131 , \u1_uk_K_r0_reg[47]/NET0131 , \u1_uk_K_r0_reg[48]/NET0131 , \u1_uk_K_r0_reg[49]/NET0131 , \u1_uk_K_r0_reg[4]/NET0131 , \u1_uk_K_r0_reg[50]/NET0131 , \u1_uk_K_r0_reg[51]/NET0131 , \u1_uk_K_r0_reg[52]/P0001 , \u1_uk_K_r0_reg[54]/NET0131 , \u1_uk_K_r0_reg[55]/NET0131 , \u1_uk_K_r0_reg[5]/NET0131 , \u1_uk_K_r0_reg[6]/NET0131 , \u1_uk_K_r0_reg[7]/NET0131 , \u1_uk_K_r0_reg[8]/NET0131 , \u1_uk_K_r0_reg[9]/NET0131 , \u1_uk_K_r10_reg[0]/NET0131 , \u1_uk_K_r10_reg[10]/NET0131 , \u1_uk_K_r10_reg[11]/NET0131 , \u1_uk_K_r10_reg[12]/NET0131 , \u1_uk_K_r10_reg[14]/NET0131 , \u1_uk_K_r10_reg[15]/NET0131 , \u1_uk_K_r10_reg[16]/NET0131 , \u1_uk_K_r10_reg[17]/NET0131 , \u1_uk_K_r10_reg[18]/NET0131 , \u1_uk_K_r10_reg[19]/NET0131 , \u1_uk_K_r10_reg[1]/NET0131 , \u1_uk_K_r10_reg[20]/NET0131 , \u1_uk_K_r10_reg[21]/NET0131 , \u1_uk_K_r10_reg[22]/NET0131 , \u1_uk_K_r10_reg[23]/NET0131 , \u1_uk_K_r10_reg[24]/NET0131 , \u1_uk_K_r10_reg[25]/NET0131 , \u1_uk_K_r10_reg[26]/NET0131 , \u1_uk_K_r10_reg[27]/NET0131 , \u1_uk_K_r10_reg[28]/NET0131 , \u1_uk_K_r10_reg[29]/NET0131 , \u1_uk_K_r10_reg[2]/NET0131 , \u1_uk_K_r10_reg[30]/NET0131 , \u1_uk_K_r10_reg[31]/NET0131 , \u1_uk_K_r10_reg[32]/NET0131 , \u1_uk_K_r10_reg[33]/NET0131 , \u1_uk_K_r10_reg[34]/NET0131 , \u1_uk_K_r10_reg[35]/NET0131 , \u1_uk_K_r10_reg[36]/NET0131 , \u1_uk_K_r10_reg[37]/NET0131 , \u1_uk_K_r10_reg[38]/NET0131 , \u1_uk_K_r10_reg[39]/NET0131 , \u1_uk_K_r10_reg[3]/NET0131 , \u1_uk_K_r10_reg[40]/NET0131 , \u1_uk_K_r10_reg[41]/P0001 , \u1_uk_K_r10_reg[42]/NET0131 , \u1_uk_K_r10_reg[43]/NET0131 , \u1_uk_K_r10_reg[44]/NET0131 , \u1_uk_K_r10_reg[45]/P0001 , \u1_uk_K_r10_reg[46]/NET0131 , \u1_uk_K_r10_reg[47]/NET0131 , \u1_uk_K_r10_reg[48]/NET0131 , \u1_uk_K_r10_reg[49]/NET0131 , \u1_uk_K_r10_reg[4]/NET0131 , \u1_uk_K_r10_reg[50]/NET0131 , \u1_uk_K_r10_reg[51]/NET0131 , \u1_uk_K_r10_reg[52]/NET0131 , \u1_uk_K_r10_reg[53]/NET0131 , \u1_uk_K_r10_reg[54]/NET0131 , \u1_uk_K_r10_reg[55]/NET0131 , \u1_uk_K_r10_reg[5]/NET0131 , \u1_uk_K_r10_reg[6]/NET0131 , \u1_uk_K_r10_reg[7]/NET0131 , \u1_uk_K_r10_reg[8]/NET0131 , \u1_uk_K_r10_reg[9]/NET0131 , \u1_uk_K_r11_reg[0]/NET0131 , \u1_uk_K_r11_reg[10]/NET0131 , \u1_uk_K_r11_reg[11]/NET0131 , \u1_uk_K_r11_reg[12]/NET0131 , \u1_uk_K_r11_reg[13]/NET0131 , \u1_uk_K_r11_reg[14]/NET0131 , \u1_uk_K_r11_reg[15]/NET0131 , \u1_uk_K_r11_reg[16]/NET0131 , \u1_uk_K_r11_reg[17]/NET0131 , \u1_uk_K_r11_reg[18]/NET0131 , \u1_uk_K_r11_reg[19]/NET0131 , \u1_uk_K_r11_reg[1]/NET0131 , \u1_uk_K_r11_reg[20]/NET0131 , \u1_uk_K_r11_reg[21]/NET0131 , \u1_uk_K_r11_reg[22]/NET0131 , \u1_uk_K_r11_reg[23]/NET0131 , \u1_uk_K_r11_reg[24]/NET0131 , \u1_uk_K_r11_reg[25]/NET0131 , \u1_uk_K_r11_reg[26]/NET0131 , \u1_uk_K_r11_reg[27]/P0001 , \u1_uk_K_r11_reg[28]/NET0131 , \u1_uk_K_r11_reg[29]/NET0131 , \u1_uk_K_r11_reg[2]/NET0131 , \u1_uk_K_r11_reg[31]/NET0131 , \u1_uk_K_r11_reg[32]/NET0131 , \u1_uk_K_r11_reg[33]/NET0131 , \u1_uk_K_r11_reg[34]/NET0131 , \u1_uk_K_r11_reg[35]/NET0131 , \u1_uk_K_r11_reg[36]/NET0131 , \u1_uk_K_r11_reg[37]/NET0131 , \u1_uk_K_r11_reg[38]/NET0131 , \u1_uk_K_r11_reg[39]/NET0131 , \u1_uk_K_r11_reg[3]/NET0131 , \u1_uk_K_r11_reg[40]/NET0131 , \u1_uk_K_r11_reg[41]/NET0131 , \u1_uk_K_r11_reg[42]/NET0131 , \u1_uk_K_r11_reg[43]/NET0131 , \u1_uk_K_r11_reg[44]/NET0131 , \u1_uk_K_r11_reg[45]/NET0131 , \u1_uk_K_r11_reg[46]/NET0131 , \u1_uk_K_r11_reg[47]/NET0131 , \u1_uk_K_r11_reg[48]/NET0131 , \u1_uk_K_r11_reg[49]/NET0131 , \u1_uk_K_r11_reg[4]/NET0131 , \u1_uk_K_r11_reg[50]/NET0131 , \u1_uk_K_r11_reg[51]/NET0131 , \u1_uk_K_r11_reg[52]/NET0131 , \u1_uk_K_r11_reg[53]/P0001 , \u1_uk_K_r11_reg[54]/NET0131 , \u1_uk_K_r11_reg[55]/NET0131 , \u1_uk_K_r11_reg[5]/NET0131 , \u1_uk_K_r11_reg[6]/NET0131 , \u1_uk_K_r11_reg[7]/NET0131 , \u1_uk_K_r11_reg[8]/NET0131 , \u1_uk_K_r11_reg[9]/NET0131 , \u1_uk_K_r12_reg[0]/NET0131 , \u1_uk_K_r12_reg[10]/P0001 , \u1_uk_K_r12_reg[11]/NET0131 , \u1_uk_K_r12_reg[12]/NET0131 , \u1_uk_K_r12_reg[13]/NET0131 , \u1_uk_K_r12_reg[14]/NET0131 , \u1_uk_K_r12_reg[15]/NET0131 , \u1_uk_K_r12_reg[16]/NET0131 , \u1_uk_K_r12_reg[17]/NET0131 , \u1_uk_K_r12_reg[18]/NET0131 , \u1_uk_K_r12_reg[19]/NET0131 , \u1_uk_K_r12_reg[1]/NET0131 , \u1_uk_K_r12_reg[20]/NET0131 , \u1_uk_K_r12_reg[21]/NET0131 , \u1_uk_K_r12_reg[22]/NET0131 , \u1_uk_K_r12_reg[23]/NET0131 , \u1_uk_K_r12_reg[24]/NET0131 , \u1_uk_K_r12_reg[25]/NET0131 , \u1_uk_K_r12_reg[26]/NET0131 , \u1_uk_K_r12_reg[27]/NET0131 , \u1_uk_K_r12_reg[28]/NET0131 , \u1_uk_K_r12_reg[29]/NET0131 , \u1_uk_K_r12_reg[2]/NET0131 , \u1_uk_K_r12_reg[30]/NET0131 , \u1_uk_K_r12_reg[31]/NET0131 , \u1_uk_K_r12_reg[32]/NET0131 , \u1_uk_K_r12_reg[33]/NET0131 , \u1_uk_K_r12_reg[34]/NET0131 , \u1_uk_K_r12_reg[35]/NET0131 , \u1_uk_K_r12_reg[36]/NET0131 , \u1_uk_K_r12_reg[37]/NET0131 , \u1_uk_K_r12_reg[38]/NET0131 , \u1_uk_K_r12_reg[3]/NET0131 , \u1_uk_K_r12_reg[40]/NET0131 , \u1_uk_K_r12_reg[41]/NET0131 , \u1_uk_K_r12_reg[42]/NET0131 , \u1_uk_K_r12_reg[43]/NET0131 , \u1_uk_K_r12_reg[44]/P0001 , \u1_uk_K_r12_reg[45]/NET0131 , \u1_uk_K_r12_reg[46]/NET0131 , \u1_uk_K_r12_reg[47]/NET0131 , \u1_uk_K_r12_reg[48]/NET0131 , \u1_uk_K_r12_reg[49]/NET0131 , \u1_uk_K_r12_reg[4]/NET0131 , \u1_uk_K_r12_reg[50]/NET0131 , \u1_uk_K_r12_reg[51]/NET0131 , \u1_uk_K_r12_reg[52]/NET0131 , \u1_uk_K_r12_reg[53]/NET0131 , \u1_uk_K_r12_reg[54]/NET0131 , \u1_uk_K_r12_reg[55]/NET0131 , \u1_uk_K_r12_reg[5]/NET0131 , \u1_uk_K_r12_reg[6]/NET0131 , \u1_uk_K_r12_reg[7]/P0001 , \u1_uk_K_r12_reg[8]/NET0131 , \u1_uk_K_r12_reg[9]/NET0131 , \u1_uk_K_r13_reg[0]/NET0131 , \u1_uk_K_r13_reg[10]/NET0131 , \u1_uk_K_r13_reg[11]/NET0131 , \u1_uk_K_r13_reg[12]/NET0131 , \u1_uk_K_r13_reg[13]/NET0131 , \u1_uk_K_r13_reg[14]/NET0131 , \u1_uk_K_r13_reg[15]/NET0131 , \u1_uk_K_r13_reg[16]/NET0131 , \u1_uk_K_r13_reg[17]/NET0131 , \u1_uk_K_r13_reg[18]/NET0131 , \u1_uk_K_r13_reg[19]/NET0131 , \u1_uk_K_r13_reg[20]/NET0131 , \u1_uk_K_r13_reg[21]/NET0131 , \u1_uk_K_r13_reg[22]/NET0131 , \u1_uk_K_r13_reg[23]/NET0131 , \u1_uk_K_r13_reg[24]/NET0131 , \u1_uk_K_r13_reg[25]/P0001 , \u1_uk_K_r13_reg[26]/NET0131 , \u1_uk_K_r13_reg[27]/NET0131 , \u1_uk_K_r13_reg[28]/NET0131 , \u1_uk_K_r13_reg[29]/NET0131 , \u1_uk_K_r13_reg[2]/NET0131 , \u1_uk_K_r13_reg[30]/NET0131 , \u1_uk_K_r13_reg[31]/NET0131 , \u1_uk_K_r13_reg[32]/NET0131 , \u1_uk_K_r13_reg[33]/NET0131 , \u1_uk_K_r13_reg[34]/NET0131 , \u1_uk_K_r13_reg[35]/NET0131 , \u1_uk_K_r13_reg[36]/NET0131 , \u1_uk_K_r13_reg[37]/NET0131 , \u1_uk_K_r13_reg[38]/NET0131 , \u1_uk_K_r13_reg[39]/NET0131 , \u1_uk_K_r13_reg[3]/NET0131 , \u1_uk_K_r13_reg[40]/NET0131 , \u1_uk_K_r13_reg[41]/NET0131 , \u1_uk_K_r13_reg[42]/NET0131 , \u1_uk_K_r13_reg[43]/NET0131 , \u1_uk_K_r13_reg[44]/NET0131 , \u1_uk_K_r13_reg[45]/NET0131 , \u1_uk_K_r13_reg[46]/NET0131 , \u1_uk_K_r13_reg[47]/NET0131 , \u1_uk_K_r13_reg[48]/NET0131 , \u1_uk_K_r13_reg[49]/NET0131 , \u1_uk_K_r13_reg[4]/NET0131 , \u1_uk_K_r13_reg[50]/NET0131 , \u1_uk_K_r13_reg[51]/NET0131 , \u1_uk_K_r13_reg[52]/P0001 , \u1_uk_K_r13_reg[54]/NET0131 , \u1_uk_K_r13_reg[55]/NET0131 , \u1_uk_K_r13_reg[5]/NET0131 , \u1_uk_K_r13_reg[6]/NET0131 , \u1_uk_K_r13_reg[7]/NET0131 , \u1_uk_K_r13_reg[8]/NET0131 , \u1_uk_K_r13_reg[9]/NET0131 , \u1_uk_K_r14_reg[0]/P0001 , \u1_uk_K_r14_reg[10]/P0001 , \u1_uk_K_r14_reg[11]/NET0131 , \u1_uk_K_r14_reg[12]/NET0131 , \u1_uk_K_r14_reg[13]/NET0131 , \u1_uk_K_r14_reg[14]/NET0131 , \u1_uk_K_r14_reg[15]/NET0131 , \u1_uk_K_r14_reg[16]/NET0131 , \u1_uk_K_r14_reg[17]/NET0131 , \u1_uk_K_r14_reg[18]/NET0131 , \u1_uk_K_r14_reg[19]/NET0131 , \u1_uk_K_r14_reg[1]/NET0131 , \u1_uk_K_r14_reg[20]/NET0131 , \u1_uk_K_r14_reg[21]/NET0131 , \u1_uk_K_r14_reg[22]/NET0131 , \u1_uk_K_r14_reg[23]/NET0131 , \u1_uk_K_r14_reg[24]/NET0131 , \u1_uk_K_r14_reg[25]/NET0131 , \u1_uk_K_r14_reg[26]/NET0131 , \u1_uk_K_r14_reg[27]/NET0131 , \u1_uk_K_r14_reg[28]/NET0131 , \u1_uk_K_r14_reg[29]/NET0131 , \u1_uk_K_r14_reg[2]/NET0131 , \u1_uk_K_r14_reg[30]/NET0131 , \u1_uk_K_r14_reg[31]/NET0131 , \u1_uk_K_r14_reg[32]/NET0131 , \u1_uk_K_r14_reg[33]/NET0131 , \u1_uk_K_r14_reg[34]/NET0131 , \u1_uk_K_r14_reg[35]/P0001 , \u1_uk_K_r14_reg[36]/NET0131 , \u1_uk_K_r14_reg[37]/NET0131 , \u1_uk_K_r14_reg[38]/NET0131 , \u1_uk_K_r14_reg[39]/P0001 , \u1_uk_K_r14_reg[3]/NET0131 , \u1_uk_K_r14_reg[40]/NET0131 , \u1_uk_K_r14_reg[41]/NET0131 , \u1_uk_K_r14_reg[42]/P0001 , \u1_uk_K_r14_reg[43]/NET0131 , \u1_uk_K_r14_reg[44]/NET0131 , \u1_uk_K_r14_reg[45]/NET0131 , \u1_uk_K_r14_reg[46]/NET0131 , \u1_uk_K_r14_reg[47]/NET0131 , \u1_uk_K_r14_reg[48]/NET0131 , \u1_uk_K_r14_reg[49]/NET0131 , \u1_uk_K_r14_reg[4]/NET0131 , \u1_uk_K_r14_reg[50]/NET0131 , \u1_uk_K_r14_reg[51]/NET0131 , \u1_uk_K_r14_reg[52]/NET0131 , \u1_uk_K_r14_reg[53]/NET0131 , \u1_uk_K_r14_reg[54]/NET0131 , \u1_uk_K_r14_reg[55]/NET0131 , \u1_uk_K_r14_reg[5]/NET0131 , \u1_uk_K_r14_reg[6]/NET0131 , \u1_uk_K_r14_reg[7]/NET0131 , \u1_uk_K_r14_reg[8]/P0001 , \u1_uk_K_r14_reg[9]/NET0131 , \u1_uk_K_r1_reg[0]/NET0131 , \u1_uk_K_r1_reg[10]/P0001 , \u1_uk_K_r1_reg[11]/NET0131 , \u1_uk_K_r1_reg[12]/NET0131 , \u1_uk_K_r1_reg[13]/NET0131 , \u1_uk_K_r1_reg[14]/NET0131 , \u1_uk_K_r1_reg[15]/NET0131 , \u1_uk_K_r1_reg[16]/NET0131 , \u1_uk_K_r1_reg[17]/NET0131 , \u1_uk_K_r1_reg[18]/NET0131 , \u1_uk_K_r1_reg[19]/NET0131 , \u1_uk_K_r1_reg[1]/NET0131 , \u1_uk_K_r1_reg[20]/NET0131 , \u1_uk_K_r1_reg[21]/NET0131 , \u1_uk_K_r1_reg[22]/NET0131 , \u1_uk_K_r1_reg[23]/NET0131 , \u1_uk_K_r1_reg[24]/NET0131 , \u1_uk_K_r1_reg[25]/NET0131 , \u1_uk_K_r1_reg[26]/NET0131 , \u1_uk_K_r1_reg[27]/NET0131 , \u1_uk_K_r1_reg[28]/NET0131 , \u1_uk_K_r1_reg[29]/NET0131 , \u1_uk_K_r1_reg[2]/NET0131 , \u1_uk_K_r1_reg[30]/NET0131 , \u1_uk_K_r1_reg[31]/NET0131 , \u1_uk_K_r1_reg[32]/NET0131 , \u1_uk_K_r1_reg[33]/NET0131 , \u1_uk_K_r1_reg[34]/NET0131 , \u1_uk_K_r1_reg[35]/NET0131 , \u1_uk_K_r1_reg[36]/NET0131 , \u1_uk_K_r1_reg[37]/NET0131 , \u1_uk_K_r1_reg[38]/NET0131 , \u1_uk_K_r1_reg[3]/NET0131 , \u1_uk_K_r1_reg[40]/NET0131 , \u1_uk_K_r1_reg[41]/NET0131 , \u1_uk_K_r1_reg[42]/NET0131 , \u1_uk_K_r1_reg[43]/NET0131 , \u1_uk_K_r1_reg[44]/P0001 , \u1_uk_K_r1_reg[45]/NET0131 , \u1_uk_K_r1_reg[46]/NET0131 , \u1_uk_K_r1_reg[47]/NET0131 , \u1_uk_K_r1_reg[48]/NET0131 , \u1_uk_K_r1_reg[49]/NET0131 , \u1_uk_K_r1_reg[4]/NET0131 , \u1_uk_K_r1_reg[50]/NET0131 , \u1_uk_K_r1_reg[51]/NET0131 , \u1_uk_K_r1_reg[52]/NET0131 , \u1_uk_K_r1_reg[53]/NET0131 , \u1_uk_K_r1_reg[54]/NET0131 , \u1_uk_K_r1_reg[55]/NET0131 , \u1_uk_K_r1_reg[5]/NET0131 , \u1_uk_K_r1_reg[6]/NET0131 , \u1_uk_K_r1_reg[7]/P0001 , \u1_uk_K_r1_reg[8]/NET0131 , \u1_uk_K_r1_reg[9]/NET0131 , \u1_uk_K_r2_reg[0]/NET0131 , \u1_uk_K_r2_reg[10]/NET0131 , \u1_uk_K_r2_reg[11]/NET0131 , \u1_uk_K_r2_reg[12]/NET0131 , \u1_uk_K_r2_reg[13]/NET0131 , \u1_uk_K_r2_reg[14]/NET0131 , \u1_uk_K_r2_reg[15]/NET0131 , \u1_uk_K_r2_reg[16]/NET0131 , \u1_uk_K_r2_reg[17]/NET0131 , \u1_uk_K_r2_reg[18]/NET0131 , \u1_uk_K_r2_reg[19]/NET0131 , \u1_uk_K_r2_reg[1]/NET0131 , \u1_uk_K_r2_reg[20]/NET0131 , \u1_uk_K_r2_reg[21]/NET0131 , \u1_uk_K_r2_reg[22]/NET0131 , \u1_uk_K_r2_reg[23]/NET0131 , \u1_uk_K_r2_reg[24]/NET0131 , \u1_uk_K_r2_reg[25]/NET0131 , \u1_uk_K_r2_reg[26]/NET0131 , \u1_uk_K_r2_reg[27]/NET0131 , \u1_uk_K_r2_reg[28]/NET0131 , \u1_uk_K_r2_reg[29]/NET0131 , \u1_uk_K_r2_reg[2]/NET0131 , \u1_uk_K_r2_reg[31]/NET0131 , \u1_uk_K_r2_reg[32]/NET0131 , \u1_uk_K_r2_reg[33]/NET0131 , \u1_uk_K_r2_reg[34]/NET0131 , \u1_uk_K_r2_reg[35]/NET0131 , \u1_uk_K_r2_reg[36]/NET0131 , \u1_uk_K_r2_reg[37]/NET0131 , \u1_uk_K_r2_reg[38]/NET0131 , \u1_uk_K_r2_reg[39]/NET0131 , \u1_uk_K_r2_reg[3]/NET0131 , \u1_uk_K_r2_reg[40]/NET0131 , \u1_uk_K_r2_reg[41]/NET0131 , \u1_uk_K_r2_reg[42]/NET0131 , \u1_uk_K_r2_reg[43]/NET0131 , \u1_uk_K_r2_reg[44]/NET0131 , \u1_uk_K_r2_reg[45]/NET0131 , \u1_uk_K_r2_reg[46]/NET0131 , \u1_uk_K_r2_reg[47]/NET0131 , \u1_uk_K_r2_reg[48]/NET0131 , \u1_uk_K_r2_reg[49]/NET0131 , \u1_uk_K_r2_reg[4]/NET0131 , \u1_uk_K_r2_reg[50]/NET0131 , \u1_uk_K_r2_reg[51]/NET0131 , \u1_uk_K_r2_reg[52]/NET0131 , \u1_uk_K_r2_reg[53]/P0001 , \u1_uk_K_r2_reg[54]/NET0131 , \u1_uk_K_r2_reg[55]/NET0131 , \u1_uk_K_r2_reg[5]/NET0131 , \u1_uk_K_r2_reg[6]/NET0131 , \u1_uk_K_r2_reg[7]/NET0131 , \u1_uk_K_r2_reg[8]/NET0131 , \u1_uk_K_r2_reg[9]/NET0131 , \u1_uk_K_r3_reg[0]/NET0131 , \u1_uk_K_r3_reg[10]/NET0131 , \u1_uk_K_r3_reg[11]/NET0131 , \u1_uk_K_r3_reg[12]/NET0131 , \u1_uk_K_r3_reg[14]/NET0131 , \u1_uk_K_r3_reg[15]/NET0131 , \u1_uk_K_r3_reg[16]/NET0131 , \u1_uk_K_r3_reg[17]/NET0131 , \u1_uk_K_r3_reg[18]/NET0131 , \u1_uk_K_r3_reg[19]/NET0131 , \u1_uk_K_r3_reg[1]/NET0131 , \u1_uk_K_r3_reg[20]/NET0131 , \u1_uk_K_r3_reg[21]/NET0131 , \u1_uk_K_r3_reg[22]/NET0131 , \u1_uk_K_r3_reg[23]/NET0131 , \u1_uk_K_r3_reg[24]/NET0131 , \u1_uk_K_r3_reg[25]/NET0131 , \u1_uk_K_r3_reg[26]/NET0131 , \u1_uk_K_r3_reg[27]/NET0131 , \u1_uk_K_r3_reg[28]/NET0131 , \u1_uk_K_r3_reg[29]/NET0131 , \u1_uk_K_r3_reg[2]/NET0131 , \u1_uk_K_r3_reg[30]/NET0131 , \u1_uk_K_r3_reg[31]/NET0131 , \u1_uk_K_r3_reg[32]/NET0131 , \u1_uk_K_r3_reg[33]/NET0131 , \u1_uk_K_r3_reg[34]/NET0131 , \u1_uk_K_r3_reg[35]/NET0131 , \u1_uk_K_r3_reg[36]/NET0131 , \u1_uk_K_r3_reg[37]/NET0131 , \u1_uk_K_r3_reg[38]/NET0131 , \u1_uk_K_r3_reg[39]/NET0131 , \u1_uk_K_r3_reg[3]/NET0131 , \u1_uk_K_r3_reg[40]/NET0131 , \u1_uk_K_r3_reg[41]/NET0131 , \u1_uk_K_r3_reg[42]/NET0131 , \u1_uk_K_r3_reg[43]/NET0131 , \u1_uk_K_r3_reg[44]/NET0131 , \u1_uk_K_r3_reg[45]/NET0131 , \u1_uk_K_r3_reg[46]/NET0131 , \u1_uk_K_r3_reg[47]/NET0131 , \u1_uk_K_r3_reg[48]/NET0131 , \u1_uk_K_r3_reg[49]/NET0131 , \u1_uk_K_r3_reg[4]/NET0131 , \u1_uk_K_r3_reg[50]/NET0131 , \u1_uk_K_r3_reg[51]/NET0131 , \u1_uk_K_r3_reg[52]/NET0131 , \u1_uk_K_r3_reg[53]/NET0131 , \u1_uk_K_r3_reg[54]/NET0131 , \u1_uk_K_r3_reg[55]/NET0131 , \u1_uk_K_r3_reg[5]/NET0131 , \u1_uk_K_r3_reg[6]/NET0131 , \u1_uk_K_r3_reg[7]/NET0131 , \u1_uk_K_r3_reg[8]/NET0131 , \u1_uk_K_r3_reg[9]/NET0131 , \u1_uk_K_r4_reg[0]/P0001 , \u1_uk_K_r4_reg[10]/NET0131 , \u1_uk_K_r4_reg[11]/NET0131 , \u1_uk_K_r4_reg[12]/NET0131 , \u1_uk_K_r4_reg[13]/NET0131 , \u1_uk_K_r4_reg[14]/NET0131 , \u1_uk_K_r4_reg[15]/NET0131 , \u1_uk_K_r4_reg[16]/NET0131 , \u1_uk_K_r4_reg[17]/NET0131 , \u1_uk_K_r4_reg[18]/NET0131 , \u1_uk_K_r4_reg[19]/NET0131 , \u1_uk_K_r4_reg[1]/NET0131 , \u1_uk_K_r4_reg[20]/NET0131 , \u1_uk_K_r4_reg[21]/NET0131 , \u1_uk_K_r4_reg[22]/NET0131 , \u1_uk_K_r4_reg[23]/P0001 , \u1_uk_K_r4_reg[25]/NET0131 , \u1_uk_K_r4_reg[26]/NET0131 , \u1_uk_K_r4_reg[27]/P0001 , \u1_uk_K_r4_reg[28]/NET0131 , \u1_uk_K_r4_reg[29]/NET0131 , \u1_uk_K_r4_reg[30]/NET0131 , \u1_uk_K_r4_reg[31]/P0001 , \u1_uk_K_r4_reg[32]/NET0131 , \u1_uk_K_r4_reg[33]/NET0131 , \u1_uk_K_r4_reg[34]/NET0131 , \u1_uk_K_r4_reg[35]/NET0131 , \u1_uk_K_r4_reg[36]/NET0131 , \u1_uk_K_r4_reg[37]/NET0131 , \u1_uk_K_r4_reg[38]/NET0131 , \u1_uk_K_r4_reg[39]/NET0131 , \u1_uk_K_r4_reg[3]/NET0131 , \u1_uk_K_r4_reg[40]/NET0131 , \u1_uk_K_r4_reg[41]/NET0131 , \u1_uk_K_r4_reg[42]/NET0131 , \u1_uk_K_r4_reg[43]/NET0131 , \u1_uk_K_r4_reg[44]/NET0131 , \u1_uk_K_r4_reg[45]/NET0131 , \u1_uk_K_r4_reg[46]/NET0131 , \u1_uk_K_r4_reg[47]/NET0131 , \u1_uk_K_r4_reg[48]/NET0131 , \u1_uk_K_r4_reg[49]/NET0131 , \u1_uk_K_r4_reg[4]/NET0131 , \u1_uk_K_r4_reg[50]/NET0131 , \u1_uk_K_r4_reg[51]/NET0131 , \u1_uk_K_r4_reg[52]/NET0131 , \u1_uk_K_r4_reg[53]/NET0131 , \u1_uk_K_r4_reg[54]/NET0131 , \u1_uk_K_r4_reg[55]/NET0131 , \u1_uk_K_r4_reg[5]/NET0131 , \u1_uk_K_r4_reg[6]/NET0131 , \u1_uk_K_r4_reg[7]/NET0131 , \u1_uk_K_r4_reg[8]/NET0131 , \u1_uk_K_r4_reg[9]/NET0131 , \u1_uk_K_r5_reg[0]/NET0131 , \u1_uk_K_r5_reg[10]/NET0131 , \u1_uk_K_r5_reg[11]/NET0131 , \u1_uk_K_r5_reg[12]/P0001 , \u1_uk_K_r5_reg[13]/P0001 , \u1_uk_K_r5_reg[14]/NET0131 , \u1_uk_K_r5_reg[15]/NET0131 , \u1_uk_K_r5_reg[16]/NET0131 , \u1_uk_K_r5_reg[17]/NET0131 , \u1_uk_K_r5_reg[18]/NET0131 , \u1_uk_K_r5_reg[19]/NET0131 , \u1_uk_K_r5_reg[1]/NET0131 , \u1_uk_K_r5_reg[20]/NET0131 , \u1_uk_K_r5_reg[21]/NET0131 , \u1_uk_K_r5_reg[22]/NET0131 , \u1_uk_K_r5_reg[23]/NET0131 , \u1_uk_K_r5_reg[24]/NET0131 , \u1_uk_K_r5_reg[25]/NET0131 , \u1_uk_K_r5_reg[26]/NET0131 , \u1_uk_K_r5_reg[27]/NET0131 , \u1_uk_K_r5_reg[28]/NET0131 , \u1_uk_K_r5_reg[29]/NET0131 , \u1_uk_K_r5_reg[2]/NET0131 , \u1_uk_K_r5_reg[30]/NET0131 , \u1_uk_K_r5_reg[31]/NET0131 , \u1_uk_K_r5_reg[32]/NET0131 , \u1_uk_K_r5_reg[33]/NET0131 , \u1_uk_K_r5_reg[34]/NET0131 , \u1_uk_K_r5_reg[35]/NET0131 , \u1_uk_K_r5_reg[36]/NET0131 , \u1_uk_K_r5_reg[37]/P0001 , \u1_uk_K_r5_reg[38]/NET0131 , \u1_uk_K_r5_reg[39]/NET0131 , \u1_uk_K_r5_reg[3]/NET0131 , \u1_uk_K_r5_reg[40]/NET0131 , \u1_uk_K_r5_reg[41]/NET0131 , \u1_uk_K_r5_reg[42]/NET0131 , \u1_uk_K_r5_reg[43]/NET0131 , \u1_uk_K_r5_reg[44]/NET0131 , \u1_uk_K_r5_reg[46]/NET0131 , \u1_uk_K_r5_reg[47]/NET0131 , \u1_uk_K_r5_reg[48]/NET0131 , \u1_uk_K_r5_reg[49]/NET0131 , \u1_uk_K_r5_reg[4]/NET0131 , \u1_uk_K_r5_reg[50]/NET0131 , \u1_uk_K_r5_reg[51]/NET0131 , \u1_uk_K_r5_reg[52]/NET0131 , \u1_uk_K_r5_reg[53]/NET0131 , \u1_uk_K_r5_reg[54]/NET0131 , \u1_uk_K_r5_reg[55]/NET0131 , \u1_uk_K_r5_reg[5]/NET0131 , \u1_uk_K_r5_reg[6]/NET0131 , \u1_uk_K_r5_reg[7]/NET0131 , \u1_uk_K_r5_reg[8]/NET0131 , \u1_uk_K_r5_reg[9]/NET0131 , \u1_uk_K_r6_reg[0]/NET0131 , \u1_uk_K_r6_reg[10]/NET0131 , \u1_uk_K_r6_reg[11]/NET0131 , \u1_uk_K_r6_reg[12]/NET0131 , \u1_uk_K_r6_reg[13]/NET0131 , \u1_uk_K_r6_reg[14]/NET0131 , \u1_uk_K_r6_reg[15]/NET0131 , \u1_uk_K_r6_reg[16]/NET0131 , \u1_uk_K_r6_reg[17]/NET0131 , \u1_uk_K_r6_reg[18]/NET0131 , \u1_uk_K_r6_reg[19]/NET0131 , \u1_uk_K_r6_reg[1]/NET0131 , \u1_uk_K_r6_reg[20]/NET0131 , \u1_uk_K_r6_reg[21]/NET0131 , \u1_uk_K_r6_reg[22]/NET0131 , \u1_uk_K_r6_reg[23]/P0001 , \u1_uk_K_r6_reg[24]/NET0131 , \u1_uk_K_r6_reg[25]/NET0131 , \u1_uk_K_r6_reg[26]/NET0131 , \u1_uk_K_r6_reg[27]/NET0131 , \u1_uk_K_r6_reg[28]/NET0131 , \u1_uk_K_r6_reg[29]/NET0131 , \u1_uk_K_r6_reg[2]/NET0131 , \u1_uk_K_r6_reg[30]/P0001 , \u1_uk_K_r6_reg[31]/NET0131 , \u1_uk_K_r6_reg[32]/NET0131 , \u1_uk_K_r6_reg[33]/NET0131 , \u1_uk_K_r6_reg[34]/NET0131 , \u1_uk_K_r6_reg[35]/NET0131 , \u1_uk_K_r6_reg[36]/NET0131 , \u1_uk_K_r6_reg[37]/NET0131 , \u1_uk_K_r6_reg[38]/NET0131 , \u1_uk_K_r6_reg[39]/NET0131 , \u1_uk_K_r6_reg[3]/NET0131 , \u1_uk_K_r6_reg[40]/NET0131 , \u1_uk_K_r6_reg[41]/NET0131 , \u1_uk_K_r6_reg[42]/NET0131 , \u1_uk_K_r6_reg[43]/NET0131 , \u1_uk_K_r6_reg[44]/NET0131 , \u1_uk_K_r6_reg[45]/NET0131 , \u1_uk_K_r6_reg[46]/NET0131 , \u1_uk_K_r6_reg[47]/NET0131 , \u1_uk_K_r6_reg[48]/NET0131 , \u1_uk_K_r6_reg[49]/NET0131 , \u1_uk_K_r6_reg[4]/NET0131 , \u1_uk_K_r6_reg[50]/NET0131 , \u1_uk_K_r6_reg[51]/NET0131 , \u1_uk_K_r6_reg[52]/NET0131 , \u1_uk_K_r6_reg[53]/NET0131 , \u1_uk_K_r6_reg[54]/NET0131 , \u1_uk_K_r6_reg[55]/P0001 , \u1_uk_K_r6_reg[5]/NET0131 , \u1_uk_K_r6_reg[6]/NET0131 , \u1_uk_K_r6_reg[7]/NET0131 , \u1_uk_K_r6_reg[8]/NET0131 , \u1_uk_K_r6_reg[9]/NET0131 , \u1_uk_K_r7_reg[0]/NET0131 , \u1_uk_K_r7_reg[10]/NET0131 , \u1_uk_K_r7_reg[11]/NET0131 , \u1_uk_K_r7_reg[12]/NET0131 , \u1_uk_K_r7_reg[13]/NET0131 , \u1_uk_K_r7_reg[14]/NET0131 , \u1_uk_K_r7_reg[15]/NET0131 , \u1_uk_K_r7_reg[16]/NET0131 , \u1_uk_K_r7_reg[17]/NET0131 , \u1_uk_K_r7_reg[18]/NET0131 , \u1_uk_K_r7_reg[19]/NET0131 , \u1_uk_K_r7_reg[1]/NET0131 , \u1_uk_K_r7_reg[20]/NET0131 , \u1_uk_K_r7_reg[21]/NET0131 , \u1_uk_K_r7_reg[22]/NET0131 , \u1_uk_K_r7_reg[23]/P0001 , \u1_uk_K_r7_reg[24]/NET0131 , \u1_uk_K_r7_reg[25]/NET0131 , \u1_uk_K_r7_reg[26]/P0001 , \u1_uk_K_r7_reg[27]/NET0131 , \u1_uk_K_r7_reg[28]/NET0131 , \u1_uk_K_r7_reg[29]/NET0131 , \u1_uk_K_r7_reg[2]/NET0131 , \u1_uk_K_r7_reg[30]/P0001 , \u1_uk_K_r7_reg[31]/NET0131 , \u1_uk_K_r7_reg[32]/NET0131 , \u1_uk_K_r7_reg[33]/NET0131 , \u1_uk_K_r7_reg[34]/NET0131 , \u1_uk_K_r7_reg[35]/NET0131 , \u1_uk_K_r7_reg[36]/NET0131 , \u1_uk_K_r7_reg[37]/NET0131 , \u1_uk_K_r7_reg[38]/NET0131 , \u1_uk_K_r7_reg[39]/NET0131 , \u1_uk_K_r7_reg[3]/NET0131 , \u1_uk_K_r7_reg[40]/NET0131 , \u1_uk_K_r7_reg[41]/NET0131 , \u1_uk_K_r7_reg[42]/NET0131 , \u1_uk_K_r7_reg[43]/NET0131 , \u1_uk_K_r7_reg[44]/NET0131 , \u1_uk_K_r7_reg[45]/NET0131 , \u1_uk_K_r7_reg[46]/NET0131 , \u1_uk_K_r7_reg[47]/NET0131 , \u1_uk_K_r7_reg[48]/NET0131 , \u1_uk_K_r7_reg[49]/NET0131 , \u1_uk_K_r7_reg[4]/NET0131 , \u1_uk_K_r7_reg[50]/NET0131 , \u1_uk_K_r7_reg[51]/NET0131 , \u1_uk_K_r7_reg[52]/NET0131 , \u1_uk_K_r7_reg[53]/NET0131 , \u1_uk_K_r7_reg[54]/NET0131 , \u1_uk_K_r7_reg[55]/P0001 , \u1_uk_K_r7_reg[5]/NET0131 , \u1_uk_K_r7_reg[6]/NET0131 , \u1_uk_K_r7_reg[7]/NET0131 , \u1_uk_K_r7_reg[8]/NET0131 , \u1_uk_K_r7_reg[9]/NET0131 , \u1_uk_K_r8_reg[0]/NET0131 , \u1_uk_K_r8_reg[10]/NET0131 , \u1_uk_K_r8_reg[11]/NET0131 , \u1_uk_K_r8_reg[12]/NET0131 , \u1_uk_K_r8_reg[13]/P0001 , \u1_uk_K_r8_reg[14]/NET0131 , \u1_uk_K_r8_reg[15]/NET0131 , \u1_uk_K_r8_reg[16]/NET0131 , \u1_uk_K_r8_reg[17]/NET0131 , \u1_uk_K_r8_reg[18]/NET0131 , \u1_uk_K_r8_reg[19]/NET0131 , \u1_uk_K_r8_reg[1]/NET0131 , \u1_uk_K_r8_reg[20]/NET0131 , \u1_uk_K_r8_reg[21]/NET0131 , \u1_uk_K_r8_reg[22]/NET0131 , \u1_uk_K_r8_reg[23]/NET0131 , \u1_uk_K_r8_reg[24]/NET0131 , \u1_uk_K_r8_reg[25]/NET0131 , \u1_uk_K_r8_reg[26]/NET0131 , \u1_uk_K_r8_reg[27]/NET0131 , \u1_uk_K_r8_reg[28]/NET0131 , \u1_uk_K_r8_reg[29]/NET0131 , \u1_uk_K_r8_reg[2]/NET0131 , \u1_uk_K_r8_reg[30]/NET0131 , \u1_uk_K_r8_reg[31]/NET0131 , \u1_uk_K_r8_reg[32]/NET0131 , \u1_uk_K_r8_reg[33]/NET0131 , \u1_uk_K_r8_reg[34]/NET0131 , \u1_uk_K_r8_reg[35]/NET0131 , \u1_uk_K_r8_reg[36]/NET0131 , \u1_uk_K_r8_reg[37]/P0001 , \u1_uk_K_r8_reg[38]/NET0131 , \u1_uk_K_r8_reg[39]/NET0131 , \u1_uk_K_r8_reg[3]/NET0131 , \u1_uk_K_r8_reg[40]/NET0131 , \u1_uk_K_r8_reg[41]/NET0131 , \u1_uk_K_r8_reg[42]/NET0131 , \u1_uk_K_r8_reg[43]/NET0131 , \u1_uk_K_r8_reg[44]/NET0131 , \u1_uk_K_r8_reg[46]/NET0131 , \u1_uk_K_r8_reg[47]/NET0131 , \u1_uk_K_r8_reg[48]/NET0131 , \u1_uk_K_r8_reg[49]/NET0131 , \u1_uk_K_r8_reg[4]/NET0131 , \u1_uk_K_r8_reg[50]/NET0131 , \u1_uk_K_r8_reg[51]/NET0131 , \u1_uk_K_r8_reg[52]/NET0131 , \u1_uk_K_r8_reg[53]/NET0131 , \u1_uk_K_r8_reg[54]/NET0131 , \u1_uk_K_r8_reg[55]/NET0131 , \u1_uk_K_r8_reg[5]/NET0131 , \u1_uk_K_r8_reg[6]/NET0131 , \u1_uk_K_r8_reg[7]/NET0131 , \u1_uk_K_r8_reg[8]/NET0131 , \u1_uk_K_r8_reg[9]/NET0131 , \u1_uk_K_r9_reg[0]/P0001 , \u1_uk_K_r9_reg[10]/NET0131 , \u1_uk_K_r9_reg[11]/NET0131 , \u1_uk_K_r9_reg[12]/NET0131 , \u1_uk_K_r9_reg[13]/NET0131 , \u1_uk_K_r9_reg[14]/NET0131 , \u1_uk_K_r9_reg[15]/NET0131 , \u1_uk_K_r9_reg[16]/NET0131 , \u1_uk_K_r9_reg[17]/NET0131 , \u1_uk_K_r9_reg[18]/NET0131 , \u1_uk_K_r9_reg[19]/NET0131 , \u1_uk_K_r9_reg[1]/NET0131 , \u1_uk_K_r9_reg[20]/NET0131 , \u1_uk_K_r9_reg[21]/NET0131 , \u1_uk_K_r9_reg[22]/NET0131 , \u1_uk_K_r9_reg[23]/NET0131 , \u1_uk_K_r9_reg[25]/NET0131 , \u1_uk_K_r9_reg[26]/NET0131 , \u1_uk_K_r9_reg[27]/P0001 , \u1_uk_K_r9_reg[28]/NET0131 , \u1_uk_K_r9_reg[29]/NET0131 , \u1_uk_K_r9_reg[30]/NET0131 , \u1_uk_K_r9_reg[31]/P0001 , \u1_uk_K_r9_reg[32]/NET0131 , \u1_uk_K_r9_reg[33]/NET0131 , \u1_uk_K_r9_reg[34]/NET0131 , \u1_uk_K_r9_reg[35]/NET0131 , \u1_uk_K_r9_reg[36]/NET0131 , \u1_uk_K_r9_reg[37]/NET0131 , \u1_uk_K_r9_reg[38]/NET0131 , \u1_uk_K_r9_reg[39]/NET0131 , \u1_uk_K_r9_reg[3]/NET0131 , \u1_uk_K_r9_reg[40]/NET0131 , \u1_uk_K_r9_reg[41]/NET0131 , \u1_uk_K_r9_reg[42]/NET0131 , \u1_uk_K_r9_reg[43]/NET0131 , \u1_uk_K_r9_reg[44]/NET0131 , \u1_uk_K_r9_reg[45]/NET0131 , \u1_uk_K_r9_reg[46]/NET0131 , \u1_uk_K_r9_reg[47]/NET0131 , \u1_uk_K_r9_reg[48]/NET0131 , \u1_uk_K_r9_reg[49]/NET0131 , \u1_uk_K_r9_reg[4]/NET0131 , \u1_uk_K_r9_reg[50]/NET0131 , \u1_uk_K_r9_reg[51]/NET0131 , \u1_uk_K_r9_reg[52]/NET0131 , \u1_uk_K_r9_reg[53]/NET0131 , \u1_uk_K_r9_reg[54]/NET0131 , \u1_uk_K_r9_reg[55]/NET0131 , \u1_uk_K_r9_reg[5]/NET0131 , \u1_uk_K_r9_reg[6]/NET0131 , \u1_uk_K_r9_reg[7]/NET0131 , \u1_uk_K_r9_reg[8]/NET0131 , \u1_uk_K_r9_reg[9]/NET0131 , \u2_L0_reg[10]/NET0131 , \u2_L0_reg[11]/NET0131 , \u2_L0_reg[12]/NET0131 , \u2_L0_reg[13]/NET0131 , \u2_L0_reg[14]/NET0131 , \u2_L0_reg[15]/NET0131 , \u2_L0_reg[16]/NET0131 , \u2_L0_reg[17]/NET0131 , \u2_L0_reg[18]/P0001 , \u2_L0_reg[19]/NET0131 , \u2_L0_reg[1]/NET0131 , \u2_L0_reg[20]/NET0131 , \u2_L0_reg[21]/NET0131 , \u2_L0_reg[22]/NET0131 , \u2_L0_reg[23]/NET0131 , \u2_L0_reg[24]/NET0131 , \u2_L0_reg[25]/NET0131 , \u2_L0_reg[26]/NET0131 , \u2_L0_reg[27]/NET0131 , \u2_L0_reg[28]/NET0131 , \u2_L0_reg[29]/NET0131 , \u2_L0_reg[2]/NET0131 , \u2_L0_reg[30]/NET0131 , \u2_L0_reg[31]/NET0131 , \u2_L0_reg[32]/NET0131 , \u2_L0_reg[3]/NET0131 , \u2_L0_reg[4]/NET0131 , \u2_L0_reg[5]/NET0131 , \u2_L0_reg[6]/NET0131 , \u2_L0_reg[7]/NET0131 , \u2_L0_reg[8]/NET0131 , \u2_L0_reg[9]/NET0131 , \u2_L10_reg[10]/NET0131 , \u2_L10_reg[11]/NET0131 , \u2_L10_reg[12]/NET0131 , \u2_L10_reg[13]/NET0131 , \u2_L10_reg[14]/NET0131 , \u2_L10_reg[15]/NET0131 , \u2_L10_reg[16]/NET0131 , \u2_L10_reg[17]/NET0131 , \u2_L10_reg[18]/P0001 , \u2_L10_reg[19]/NET0131 , \u2_L10_reg[1]/NET0131 , \u2_L10_reg[20]/NET0131 , \u2_L10_reg[21]/NET0131 , \u2_L10_reg[22]/NET0131 , \u2_L10_reg[23]/NET0131 , \u2_L10_reg[24]/NET0131 , \u2_L10_reg[25]/NET0131 , \u2_L10_reg[26]/NET0131 , \u2_L10_reg[27]/NET0131 , \u2_L10_reg[28]/NET0131 , \u2_L10_reg[29]/NET0131 , \u2_L10_reg[2]/NET0131 , \u2_L10_reg[30]/NET0131 , \u2_L10_reg[31]/NET0131 , \u2_L10_reg[32]/NET0131 , \u2_L10_reg[3]/NET0131 , \u2_L10_reg[4]/NET0131 , \u2_L10_reg[5]/NET0131 , \u2_L10_reg[6]/NET0131 , \u2_L10_reg[7]/NET0131 , \u2_L10_reg[8]/NET0131 , \u2_L10_reg[9]/NET0131 , \u2_L11_reg[10]/NET0131 , \u2_L11_reg[11]/NET0131 , \u2_L11_reg[12]/NET0131 , \u2_L11_reg[13]/NET0131 , \u2_L11_reg[14]/NET0131 , \u2_L11_reg[15]/NET0131 , \u2_L11_reg[16]/NET0131 , \u2_L11_reg[17]/NET0131 , \u2_L11_reg[18]/P0001 , \u2_L11_reg[19]/NET0131 , \u2_L11_reg[1]/NET0131 , \u2_L11_reg[20]/NET0131 , \u2_L11_reg[21]/NET0131 , \u2_L11_reg[22]/NET0131 , \u2_L11_reg[23]/NET0131 , \u2_L11_reg[24]/NET0131 , \u2_L11_reg[25]/NET0131 , \u2_L11_reg[26]/NET0131 , \u2_L11_reg[27]/NET0131 , \u2_L11_reg[28]/NET0131 , \u2_L11_reg[29]/NET0131 , \u2_L11_reg[2]/NET0131 , \u2_L11_reg[30]/NET0131 , \u2_L11_reg[31]/NET0131 , \u2_L11_reg[32]/NET0131 , \u2_L11_reg[3]/NET0131 , \u2_L11_reg[4]/NET0131 , \u2_L11_reg[5]/NET0131 , \u2_L11_reg[6]/NET0131 , \u2_L11_reg[7]/NET0131 , \u2_L11_reg[8]/NET0131 , \u2_L11_reg[9]/NET0131 , \u2_L12_reg[10]/NET0131 , \u2_L12_reg[11]/NET0131 , \u2_L12_reg[12]/NET0131 , \u2_L12_reg[13]/NET0131 , \u2_L12_reg[14]/NET0131 , \u2_L12_reg[15]/NET0131 , \u2_L12_reg[16]/NET0131 , \u2_L12_reg[17]/NET0131 , \u2_L12_reg[18]/P0001 , \u2_L12_reg[19]/NET0131 , \u2_L12_reg[1]/NET0131 , \u2_L12_reg[20]/NET0131 , \u2_L12_reg[21]/NET0131 , \u2_L12_reg[22]/NET0131 , \u2_L12_reg[23]/NET0131 , \u2_L12_reg[24]/NET0131 , \u2_L12_reg[25]/NET0131 , \u2_L12_reg[26]/NET0131 , \u2_L12_reg[27]/NET0131 , \u2_L12_reg[28]/NET0131 , \u2_L12_reg[29]/NET0131 , \u2_L12_reg[2]/NET0131 , \u2_L12_reg[30]/NET0131 , \u2_L12_reg[31]/NET0131 , \u2_L12_reg[32]/NET0131 , \u2_L12_reg[3]/NET0131 , \u2_L12_reg[4]/NET0131 , \u2_L12_reg[5]/NET0131 , \u2_L12_reg[6]/NET0131 , \u2_L12_reg[7]/NET0131 , \u2_L12_reg[8]/NET0131 , \u2_L12_reg[9]/NET0131 , \u2_L13_reg[10]/NET0131 , \u2_L13_reg[11]/NET0131 , \u2_L13_reg[12]/NET0131 , \u2_L13_reg[13]/NET0131 , \u2_L13_reg[14]/NET0131 , \u2_L13_reg[15]/NET0131 , \u2_L13_reg[16]/NET0131 , \u2_L13_reg[17]/NET0131 , \u2_L13_reg[18]/P0001 , \u2_L13_reg[19]/P0001 , \u2_L13_reg[1]/NET0131 , \u2_L13_reg[20]/NET0131 , \u2_L13_reg[21]/NET0131 , \u2_L13_reg[22]/NET0131 , \u2_L13_reg[23]/P0001 , \u2_L13_reg[24]/NET0131 , \u2_L13_reg[25]/NET0131 , \u2_L13_reg[26]/NET0131 , \u2_L13_reg[27]/NET0131 , \u2_L13_reg[28]/NET0131 , \u2_L13_reg[29]/NET0131 , \u2_L13_reg[2]/NET0131 , \u2_L13_reg[30]/NET0131 , \u2_L13_reg[31]/NET0131 , \u2_L13_reg[32]/NET0131 , \u2_L13_reg[3]/NET0131 , \u2_L13_reg[4]/NET0131 , \u2_L13_reg[5]/NET0131 , \u2_L13_reg[6]/NET0131 , \u2_L13_reg[7]/NET0131 , \u2_L13_reg[8]/NET0131 , \u2_L13_reg[9]/NET0131 , \u2_L14_reg[10]/P0001 , \u2_L14_reg[11]/P0001 , \u2_L14_reg[12]/P0001 , \u2_L14_reg[13]/P0001 , \u2_L14_reg[14]/P0001 , \u2_L14_reg[15]/P0001 , \u2_L14_reg[16]/P0001 , \u2_L14_reg[17]/P0001 , \u2_L14_reg[18]/P0001 , \u2_L14_reg[19]/P0001 , \u2_L14_reg[1]/P0001 , \u2_L14_reg[20]/P0001 , \u2_L14_reg[21]/P0001 , \u2_L14_reg[22]/P0001 , \u2_L14_reg[23]/P0001 , \u2_L14_reg[24]/P0001 , \u2_L14_reg[25]/P0001 , \u2_L14_reg[26]/P0001 , \u2_L14_reg[27]/P0001 , \u2_L14_reg[28]/P0001 , \u2_L14_reg[29]/P0001 , \u2_L14_reg[2]/P0001 , \u2_L14_reg[30]/P0001 , \u2_L14_reg[31]/P0001 , \u2_L14_reg[32]/P0001 , \u2_L14_reg[3]/P0001 , \u2_L14_reg[4]/P0001 , \u2_L14_reg[5]/P0001 , \u2_L14_reg[6]/P0001 , \u2_L14_reg[7]/P0001 , \u2_L14_reg[8]/P0001 , \u2_L14_reg[9]/P0001 , \u2_L1_reg[10]/NET0131 , \u2_L1_reg[11]/NET0131 , \u2_L1_reg[12]/NET0131 , \u2_L1_reg[13]/NET0131 , \u2_L1_reg[14]/NET0131 , \u2_L1_reg[15]/NET0131 , \u2_L1_reg[16]/NET0131 , \u2_L1_reg[17]/NET0131 , \u2_L1_reg[18]/P0001 , \u2_L1_reg[19]/NET0131 , \u2_L1_reg[1]/NET0131 , \u2_L1_reg[20]/NET0131 , \u2_L1_reg[21]/NET0131 , \u2_L1_reg[22]/NET0131 , \u2_L1_reg[23]/NET0131 , \u2_L1_reg[24]/NET0131 , \u2_L1_reg[25]/NET0131 , \u2_L1_reg[26]/NET0131 , \u2_L1_reg[27]/NET0131 , \u2_L1_reg[28]/NET0131 , \u2_L1_reg[29]/NET0131 , \u2_L1_reg[2]/NET0131 , \u2_L1_reg[30]/NET0131 , \u2_L1_reg[31]/NET0131 , \u2_L1_reg[32]/NET0131 , \u2_L1_reg[3]/NET0131 , \u2_L1_reg[4]/NET0131 , \u2_L1_reg[5]/NET0131 , \u2_L1_reg[6]/NET0131 , \u2_L1_reg[7]/NET0131 , \u2_L1_reg[8]/NET0131 , \u2_L1_reg[9]/NET0131 , \u2_L2_reg[10]/NET0131 , \u2_L2_reg[11]/NET0131 , \u2_L2_reg[12]/NET0131 , \u2_L2_reg[13]/NET0131 , \u2_L2_reg[14]/NET0131 , \u2_L2_reg[15]/NET0131 , \u2_L2_reg[16]/NET0131 , \u2_L2_reg[17]/NET0131 , \u2_L2_reg[18]/P0001 , \u2_L2_reg[19]/NET0131 , \u2_L2_reg[1]/NET0131 , \u2_L2_reg[20]/NET0131 , \u2_L2_reg[21]/NET0131 , \u2_L2_reg[22]/NET0131 , \u2_L2_reg[23]/NET0131 , \u2_L2_reg[24]/NET0131 , \u2_L2_reg[25]/NET0131 , \u2_L2_reg[26]/NET0131 , \u2_L2_reg[27]/NET0131 , \u2_L2_reg[28]/NET0131 , \u2_L2_reg[29]/NET0131 , \u2_L2_reg[2]/NET0131 , \u2_L2_reg[30]/NET0131 , \u2_L2_reg[31]/NET0131 , \u2_L2_reg[32]/NET0131 , \u2_L2_reg[3]/NET0131 , \u2_L2_reg[4]/NET0131 , \u2_L2_reg[5]/NET0131 , \u2_L2_reg[6]/NET0131 , \u2_L2_reg[7]/NET0131 , \u2_L2_reg[8]/NET0131 , \u2_L2_reg[9]/NET0131 , \u2_L3_reg[10]/NET0131 , \u2_L3_reg[11]/NET0131 , \u2_L3_reg[12]/NET0131 , \u2_L3_reg[13]/NET0131 , \u2_L3_reg[14]/NET0131 , \u2_L3_reg[15]/NET0131 , \u2_L3_reg[16]/NET0131 , \u2_L3_reg[17]/NET0131 , \u2_L3_reg[18]/P0001 , \u2_L3_reg[19]/NET0131 , \u2_L3_reg[1]/NET0131 , \u2_L3_reg[20]/NET0131 , \u2_L3_reg[21]/NET0131 , \u2_L3_reg[22]/NET0131 , \u2_L3_reg[23]/NET0131 , \u2_L3_reg[24]/NET0131 , \u2_L3_reg[25]/NET0131 , \u2_L3_reg[26]/NET0131 , \u2_L3_reg[27]/NET0131 , \u2_L3_reg[28]/NET0131 , \u2_L3_reg[29]/NET0131 , \u2_L3_reg[2]/NET0131 , \u2_L3_reg[30]/NET0131 , \u2_L3_reg[31]/NET0131 , \u2_L3_reg[32]/NET0131 , \u2_L3_reg[3]/NET0131 , \u2_L3_reg[4]/NET0131 , \u2_L3_reg[5]/NET0131 , \u2_L3_reg[6]/NET0131 , \u2_L3_reg[7]/NET0131 , \u2_L3_reg[8]/NET0131 , \u2_L3_reg[9]/NET0131 , \u2_L4_reg[10]/NET0131 , \u2_L4_reg[11]/NET0131 , \u2_L4_reg[12]/NET0131 , \u2_L4_reg[13]/NET0131 , \u2_L4_reg[14]/NET0131 , \u2_L4_reg[15]/NET0131 , \u2_L4_reg[16]/NET0131 , \u2_L4_reg[17]/NET0131 , \u2_L4_reg[18]/P0001 , \u2_L4_reg[19]/NET0131 , \u2_L4_reg[1]/NET0131 , \u2_L4_reg[20]/NET0131 , \u2_L4_reg[21]/NET0131 , \u2_L4_reg[22]/NET0131 , \u2_L4_reg[23]/NET0131 , \u2_L4_reg[24]/NET0131 , \u2_L4_reg[25]/NET0131 , \u2_L4_reg[26]/NET0131 , \u2_L4_reg[27]/NET0131 , \u2_L4_reg[28]/NET0131 , \u2_L4_reg[29]/NET0131 , \u2_L4_reg[2]/NET0131 , \u2_L4_reg[30]/NET0131 , \u2_L4_reg[31]/NET0131 , \u2_L4_reg[32]/NET0131 , \u2_L4_reg[3]/NET0131 , \u2_L4_reg[4]/NET0131 , \u2_L4_reg[5]/NET0131 , \u2_L4_reg[6]/NET0131 , \u2_L4_reg[7]/NET0131 , \u2_L4_reg[8]/NET0131 , \u2_L4_reg[9]/NET0131 , \u2_L5_reg[10]/NET0131 , \u2_L5_reg[11]/NET0131 , \u2_L5_reg[12]/NET0131 , \u2_L5_reg[13]/NET0131 , \u2_L5_reg[14]/NET0131 , \u2_L5_reg[15]/NET0131 , \u2_L5_reg[16]/NET0131 , \u2_L5_reg[17]/NET0131 , \u2_L5_reg[18]/NET0131 , \u2_L5_reg[19]/NET0131 , \u2_L5_reg[1]/NET0131 , \u2_L5_reg[20]/NET0131 , \u2_L5_reg[21]/NET0131 , \u2_L5_reg[22]/NET0131 , \u2_L5_reg[23]/NET0131 , \u2_L5_reg[24]/NET0131 , \u2_L5_reg[25]/NET0131 , \u2_L5_reg[26]/NET0131 , \u2_L5_reg[27]/NET0131 , \u2_L5_reg[28]/NET0131 , \u2_L5_reg[29]/NET0131 , \u2_L5_reg[2]/NET0131 , \u2_L5_reg[30]/NET0131 , \u2_L5_reg[31]/NET0131 , \u2_L5_reg[32]/NET0131 , \u2_L5_reg[3]/NET0131 , \u2_L5_reg[4]/NET0131 , \u2_L5_reg[5]/NET0131 , \u2_L5_reg[6]/NET0131 , \u2_L5_reg[7]/NET0131 , \u2_L5_reg[8]/NET0131 , \u2_L5_reg[9]/NET0131 , \u2_L6_reg[10]/NET0131 , \u2_L6_reg[11]/NET0131 , \u2_L6_reg[12]/NET0131 , \u2_L6_reg[13]/NET0131 , \u2_L6_reg[14]/NET0131 , \u2_L6_reg[15]/NET0131 , \u2_L6_reg[16]/NET0131 , \u2_L6_reg[17]/NET0131 , \u2_L6_reg[18]/P0001 , \u2_L6_reg[19]/NET0131 , \u2_L6_reg[1]/NET0131 , \u2_L6_reg[20]/NET0131 , \u2_L6_reg[21]/NET0131 , \u2_L6_reg[22]/NET0131 , \u2_L6_reg[23]/NET0131 , \u2_L6_reg[24]/NET0131 , \u2_L6_reg[25]/NET0131 , \u2_L6_reg[26]/NET0131 , \u2_L6_reg[27]/NET0131 , \u2_L6_reg[28]/NET0131 , \u2_L6_reg[29]/NET0131 , \u2_L6_reg[2]/NET0131 , \u2_L6_reg[30]/NET0131 , \u2_L6_reg[31]/NET0131 , \u2_L6_reg[32]/NET0131 , \u2_L6_reg[3]/NET0131 , \u2_L6_reg[4]/NET0131 , \u2_L6_reg[5]/NET0131 , \u2_L6_reg[6]/NET0131 , \u2_L6_reg[7]/NET0131 , \u2_L6_reg[8]/NET0131 , \u2_L6_reg[9]/NET0131 , \u2_L7_reg[10]/NET0131 , \u2_L7_reg[11]/NET0131 , \u2_L7_reg[12]/NET0131 , \u2_L7_reg[13]/NET0131 , \u2_L7_reg[14]/NET0131 , \u2_L7_reg[15]/NET0131 , \u2_L7_reg[16]/NET0131 , \u2_L7_reg[17]/NET0131 , \u2_L7_reg[18]/P0001 , \u2_L7_reg[19]/NET0131 , \u2_L7_reg[1]/NET0131 , \u2_L7_reg[20]/NET0131 , \u2_L7_reg[21]/NET0131 , \u2_L7_reg[22]/NET0131 , \u2_L7_reg[23]/NET0131 , \u2_L7_reg[24]/NET0131 , \u2_L7_reg[25]/NET0131 , \u2_L7_reg[26]/NET0131 , \u2_L7_reg[27]/NET0131 , \u2_L7_reg[28]/NET0131 , \u2_L7_reg[29]/NET0131 , \u2_L7_reg[2]/NET0131 , \u2_L7_reg[30]/NET0131 , \u2_L7_reg[31]/NET0131 , \u2_L7_reg[32]/NET0131 , \u2_L7_reg[3]/NET0131 , \u2_L7_reg[4]/NET0131 , \u2_L7_reg[5]/NET0131 , \u2_L7_reg[6]/NET0131 , \u2_L7_reg[7]/NET0131 , \u2_L7_reg[8]/NET0131 , \u2_L7_reg[9]/NET0131 , \u2_L8_reg[10]/NET0131 , \u2_L8_reg[11]/NET0131 , \u2_L8_reg[12]/NET0131 , \u2_L8_reg[13]/NET0131 , \u2_L8_reg[14]/NET0131 , \u2_L8_reg[15]/NET0131 , \u2_L8_reg[16]/NET0131 , \u2_L8_reg[17]/NET0131 , \u2_L8_reg[18]/P0001 , \u2_L8_reg[19]/NET0131 , \u2_L8_reg[1]/NET0131 , \u2_L8_reg[20]/NET0131 , \u2_L8_reg[21]/NET0131 , \u2_L8_reg[22]/NET0131 , \u2_L8_reg[23]/NET0131 , \u2_L8_reg[24]/NET0131 , \u2_L8_reg[25]/NET0131 , \u2_L8_reg[26]/NET0131 , \u2_L8_reg[27]/NET0131 , \u2_L8_reg[28]/NET0131 , \u2_L8_reg[29]/NET0131 , \u2_L8_reg[2]/NET0131 , \u2_L8_reg[30]/NET0131 , \u2_L8_reg[31]/NET0131 , \u2_L8_reg[32]/NET0131 , \u2_L8_reg[3]/NET0131 , \u2_L8_reg[4]/NET0131 , \u2_L8_reg[5]/NET0131 , \u2_L8_reg[6]/NET0131 , \u2_L8_reg[7]/NET0131 , \u2_L8_reg[8]/NET0131 , \u2_L8_reg[9]/NET0131 , \u2_L9_reg[10]/NET0131 , \u2_L9_reg[11]/NET0131 , \u2_L9_reg[12]/NET0131 , \u2_L9_reg[13]/NET0131 , \u2_L9_reg[14]/NET0131 , \u2_L9_reg[15]/NET0131 , \u2_L9_reg[16]/NET0131 , \u2_L9_reg[17]/NET0131 , \u2_L9_reg[18]/P0001 , \u2_L9_reg[19]/NET0131 , \u2_L9_reg[1]/NET0131 , \u2_L9_reg[20]/NET0131 , \u2_L9_reg[21]/NET0131 , \u2_L9_reg[22]/NET0131 , \u2_L9_reg[23]/NET0131 , \u2_L9_reg[24]/NET0131 , \u2_L9_reg[25]/NET0131 , \u2_L9_reg[26]/NET0131 , \u2_L9_reg[27]/NET0131 , \u2_L9_reg[28]/NET0131 , \u2_L9_reg[29]/NET0131 , \u2_L9_reg[2]/NET0131 , \u2_L9_reg[30]/NET0131 , \u2_L9_reg[31]/NET0131 , \u2_L9_reg[32]/NET0131 , \u2_L9_reg[3]/NET0131 , \u2_L9_reg[4]/NET0131 , \u2_L9_reg[5]/NET0131 , \u2_L9_reg[6]/NET0131 , \u2_L9_reg[7]/NET0131 , \u2_L9_reg[8]/NET0131 , \u2_L9_reg[9]/NET0131 , \u2_R0_reg[10]/NET0131 , \u2_R0_reg[11]/P0001 , \u2_R0_reg[12]/NET0131 , \u2_R0_reg[13]/NET0131 , \u2_R0_reg[14]/NET0131 , \u2_R0_reg[15]/NET0131 , \u2_R0_reg[16]/NET0131 , \u2_R0_reg[17]/NET0131 , \u2_R0_reg[18]/NET0131 , \u2_R0_reg[19]/NET0131 , \u2_R0_reg[1]/NET0131 , \u2_R0_reg[20]/NET0131 , \u2_R0_reg[21]/NET0131 , \u2_R0_reg[22]/NET0131 , \u2_R0_reg[23]/NET0131 , \u2_R0_reg[24]/NET0131 , \u2_R0_reg[25]/NET0131 , \u2_R0_reg[26]/NET0131 , \u2_R0_reg[27]/NET0131 , \u2_R0_reg[28]/NET0131 , \u2_R0_reg[29]/NET0131 , \u2_R0_reg[2]/NET0131 , \u2_R0_reg[30]/NET0131 , \u2_R0_reg[31]/P0001 , \u2_R0_reg[32]/NET0131 , \u2_R0_reg[3]/NET0131 , \u2_R0_reg[4]/NET0131 , \u2_R0_reg[5]/NET0131 , \u2_R0_reg[6]/NET0131 , \u2_R0_reg[7]/NET0131 , \u2_R0_reg[8]/NET0131 , \u2_R0_reg[9]/NET0131 , \u2_R10_reg[10]/NET0131 , \u2_R10_reg[11]/NET0131 , \u2_R10_reg[12]/NET0131 , \u2_R10_reg[13]/NET0131 , \u2_R10_reg[14]/NET0131 , \u2_R10_reg[15]/NET0131 , \u2_R10_reg[16]/NET0131 , \u2_R10_reg[17]/NET0131 , \u2_R10_reg[18]/NET0131 , \u2_R10_reg[19]/NET0131 , \u2_R10_reg[1]/NET0131 , \u2_R10_reg[20]/NET0131 , \u2_R10_reg[21]/NET0131 , \u2_R10_reg[22]/NET0131 , \u2_R10_reg[23]/NET0131 , \u2_R10_reg[24]/NET0131 , \u2_R10_reg[25]/NET0131 , \u2_R10_reg[26]/NET0131 , \u2_R10_reg[27]/NET0131 , \u2_R10_reg[28]/NET0131 , \u2_R10_reg[29]/NET0131 , \u2_R10_reg[2]/NET0131 , \u2_R10_reg[30]/NET0131 , \u2_R10_reg[31]/P0001 , \u2_R10_reg[32]/NET0131 , \u2_R10_reg[3]/NET0131 , \u2_R10_reg[4]/NET0131 , \u2_R10_reg[5]/NET0131 , \u2_R10_reg[6]/NET0131 , \u2_R10_reg[7]/NET0131 , \u2_R10_reg[8]/NET0131 , \u2_R10_reg[9]/NET0131 , \u2_R11_reg[10]/NET0131 , \u2_R11_reg[11]/NET0131 , \u2_R11_reg[12]/NET0131 , \u2_R11_reg[13]/NET0131 , \u2_R11_reg[14]/NET0131 , \u2_R11_reg[15]/NET0131 , \u2_R11_reg[16]/NET0131 , \u2_R11_reg[17]/NET0131 , \u2_R11_reg[18]/NET0131 , \u2_R11_reg[19]/NET0131 , \u2_R11_reg[1]/NET0131 , \u2_R11_reg[20]/NET0131 , \u2_R11_reg[21]/NET0131 , \u2_R11_reg[22]/NET0131 , \u2_R11_reg[23]/NET0131 , \u2_R11_reg[24]/NET0131 , \u2_R11_reg[25]/NET0131 , \u2_R11_reg[26]/NET0131 , \u2_R11_reg[27]/NET0131 , \u2_R11_reg[28]/NET0131 , \u2_R11_reg[29]/NET0131 , \u2_R11_reg[2]/NET0131 , \u2_R11_reg[30]/NET0131 , \u2_R11_reg[31]/P0001 , \u2_R11_reg[32]/NET0131 , \u2_R11_reg[3]/NET0131 , \u2_R11_reg[4]/NET0131 , \u2_R11_reg[5]/NET0131 , \u2_R11_reg[6]/NET0131 , \u2_R11_reg[7]/NET0131 , \u2_R11_reg[8]/NET0131 , \u2_R11_reg[9]/NET0131 , \u2_R12_reg[10]/NET0131 , \u2_R12_reg[11]/NET0131 , \u2_R12_reg[12]/NET0131 , \u2_R12_reg[13]/NET0131 , \u2_R12_reg[14]/NET0131 , \u2_R12_reg[15]/NET0131 , \u2_R12_reg[16]/NET0131 , \u2_R12_reg[17]/NET0131 , \u2_R12_reg[18]/NET0131 , \u2_R12_reg[19]/NET0131 , \u2_R12_reg[1]/NET0131 , \u2_R12_reg[20]/NET0131 , \u2_R12_reg[21]/NET0131 , \u2_R12_reg[22]/NET0131 , \u2_R12_reg[23]/NET0131 , \u2_R12_reg[24]/NET0131 , \u2_R12_reg[25]/NET0131 , \u2_R12_reg[26]/NET0131 , \u2_R12_reg[27]/NET0131 , \u2_R12_reg[28]/NET0131 , \u2_R12_reg[29]/NET0131 , \u2_R12_reg[2]/NET0131 , \u2_R12_reg[30]/NET0131 , \u2_R12_reg[31]/P0001 , \u2_R12_reg[32]/NET0131 , \u2_R12_reg[3]/NET0131 , \u2_R12_reg[4]/NET0131 , \u2_R12_reg[5]/NET0131 , \u2_R12_reg[6]/NET0131 , \u2_R12_reg[7]/NET0131 , \u2_R12_reg[8]/NET0131 , \u2_R12_reg[9]/NET0131 , \u2_R13_reg[10]/NET0131 , \u2_R13_reg[11]/NET0131 , \u2_R13_reg[12]/NET0131 , \u2_R13_reg[13]/NET0131 , \u2_R13_reg[14]/NET0131 , \u2_R13_reg[15]/NET0131 , \u2_R13_reg[16]/NET0131 , \u2_R13_reg[17]/NET0131 , \u2_R13_reg[18]/NET0131 , \u2_R13_reg[19]/NET0131 , \u2_R13_reg[1]/NET0131 , \u2_R13_reg[20]/NET0131 , \u2_R13_reg[21]/NET0131 , \u2_R13_reg[22]/NET0131 , \u2_R13_reg[23]/NET0131 , \u2_R13_reg[24]/NET0131 , \u2_R13_reg[25]/NET0131 , \u2_R13_reg[26]/NET0131 , \u2_R13_reg[27]/P0001 , \u2_R13_reg[28]/NET0131 , \u2_R13_reg[29]/NET0131 , \u2_R13_reg[2]/NET0131 , \u2_R13_reg[30]/NET0131 , \u2_R13_reg[31]/P0001 , \u2_R13_reg[32]/NET0131 , \u2_R13_reg[3]/NET0131 , \u2_R13_reg[4]/NET0131 , \u2_R13_reg[5]/NET0131 , \u2_R13_reg[6]/NET0131 , \u2_R13_reg[7]/NET0131 , \u2_R13_reg[8]/NET0131 , \u2_R13_reg[9]/NET0131 , \u2_R14_reg[10]/P0001 , \u2_R14_reg[11]/P0001 , \u2_R14_reg[12]/NET0131 , \u2_R14_reg[13]/NET0131 , \u2_R14_reg[14]/NET0131 , \u2_R14_reg[15]/NET0131 , \u2_R14_reg[16]/NET0131 , \u2_R14_reg[17]/NET0131 , \u2_R14_reg[18]/NET0131 , \u2_R14_reg[19]/P0001 , \u2_R14_reg[1]/NET0131 , \u2_R14_reg[20]/NET0131 , \u2_R14_reg[21]/NET0131 , \u2_R14_reg[22]/P0001 , \u2_R14_reg[23]/P0001 , \u2_R14_reg[24]/NET0131 , \u2_R14_reg[25]/NET0131 , \u2_R14_reg[26]/P0001 , \u2_R14_reg[27]/P0001 , \u2_R14_reg[28]/NET0131 , \u2_R14_reg[29]/NET0131 , \u2_R14_reg[2]/NET0131 , \u2_R14_reg[30]/NET0131 , \u2_R14_reg[31]/P0001 , \u2_R14_reg[32]/NET0131 , \u2_R14_reg[3]/NET0131 , \u2_R14_reg[4]/NET0131 , \u2_R14_reg[5]/NET0131 , \u2_R14_reg[6]/NET0131 , \u2_R14_reg[7]/P0001 , \u2_R14_reg[8]/NET0131 , \u2_R14_reg[9]/NET0131 , \u2_R1_reg[10]/NET0131 , \u2_R1_reg[11]/P0001 , \u2_R1_reg[12]/NET0131 , \u2_R1_reg[13]/NET0131 , \u2_R1_reg[14]/NET0131 , \u2_R1_reg[15]/NET0131 , \u2_R1_reg[16]/NET0131 , \u2_R1_reg[17]/NET0131 , \u2_R1_reg[18]/NET0131 , \u2_R1_reg[19]/NET0131 , \u2_R1_reg[1]/NET0131 , \u2_R1_reg[20]/NET0131 , \u2_R1_reg[21]/NET0131 , \u2_R1_reg[22]/NET0131 , \u2_R1_reg[23]/NET0131 , \u2_R1_reg[24]/NET0131 , \u2_R1_reg[25]/NET0131 , \u2_R1_reg[26]/NET0131 , \u2_R1_reg[27]/NET0131 , \u2_R1_reg[28]/NET0131 , \u2_R1_reg[29]/NET0131 , \u2_R1_reg[2]/NET0131 , \u2_R1_reg[30]/NET0131 , \u2_R1_reg[31]/P0001 , \u2_R1_reg[32]/NET0131 , \u2_R1_reg[3]/NET0131 , \u2_R1_reg[4]/NET0131 , \u2_R1_reg[5]/NET0131 , \u2_R1_reg[6]/NET0131 , \u2_R1_reg[7]/NET0131 , \u2_R1_reg[8]/NET0131 , \u2_R1_reg[9]/NET0131 , \u2_R2_reg[10]/NET0131 , \u2_R2_reg[11]/NET0131 , \u2_R2_reg[12]/NET0131 , \u2_R2_reg[13]/NET0131 , \u2_R2_reg[14]/NET0131 , \u2_R2_reg[15]/NET0131 , \u2_R2_reg[16]/NET0131 , \u2_R2_reg[17]/NET0131 , \u2_R2_reg[18]/NET0131 , \u2_R2_reg[19]/NET0131 , \u2_R2_reg[1]/NET0131 , \u2_R2_reg[20]/NET0131 , \u2_R2_reg[21]/NET0131 , \u2_R2_reg[22]/NET0131 , \u2_R2_reg[23]/NET0131 , \u2_R2_reg[24]/NET0131 , \u2_R2_reg[25]/NET0131 , \u2_R2_reg[26]/NET0131 , \u2_R2_reg[27]/NET0131 , \u2_R2_reg[28]/NET0131 , \u2_R2_reg[29]/NET0131 , \u2_R2_reg[2]/NET0131 , \u2_R2_reg[30]/NET0131 , \u2_R2_reg[31]/P0001 , \u2_R2_reg[32]/NET0131 , \u2_R2_reg[3]/NET0131 , \u2_R2_reg[4]/NET0131 , \u2_R2_reg[5]/NET0131 , \u2_R2_reg[6]/NET0131 , \u2_R2_reg[7]/NET0131 , \u2_R2_reg[8]/NET0131 , \u2_R2_reg[9]/NET0131 , \u2_R3_reg[10]/NET0131 , \u2_R3_reg[11]/P0001 , \u2_R3_reg[12]/NET0131 , \u2_R3_reg[13]/NET0131 , \u2_R3_reg[14]/NET0131 , \u2_R3_reg[15]/NET0131 , \u2_R3_reg[16]/NET0131 , \u2_R3_reg[17]/NET0131 , \u2_R3_reg[18]/NET0131 , \u2_R3_reg[19]/NET0131 , \u2_R3_reg[1]/NET0131 , \u2_R3_reg[20]/NET0131 , \u2_R3_reg[21]/NET0131 , \u2_R3_reg[22]/NET0131 , \u2_R3_reg[23]/NET0131 , \u2_R3_reg[24]/NET0131 , \u2_R3_reg[25]/NET0131 , \u2_R3_reg[26]/NET0131 , \u2_R3_reg[27]/NET0131 , \u2_R3_reg[28]/NET0131 , \u2_R3_reg[29]/NET0131 , \u2_R3_reg[2]/NET0131 , \u2_R3_reg[30]/NET0131 , \u2_R3_reg[31]/P0001 , \u2_R3_reg[32]/NET0131 , \u2_R3_reg[3]/NET0131 , \u2_R3_reg[4]/NET0131 , \u2_R3_reg[5]/NET0131 , \u2_R3_reg[6]/NET0131 , \u2_R3_reg[7]/NET0131 , \u2_R3_reg[8]/NET0131 , \u2_R3_reg[9]/NET0131 , \u2_R4_reg[10]/NET0131 , \u2_R4_reg[11]/NET0131 , \u2_R4_reg[12]/NET0131 , \u2_R4_reg[13]/NET0131 , \u2_R4_reg[14]/NET0131 , \u2_R4_reg[15]/NET0131 , \u2_R4_reg[16]/NET0131 , \u2_R4_reg[17]/NET0131 , \u2_R4_reg[18]/NET0131 , \u2_R4_reg[19]/NET0131 , \u2_R4_reg[1]/NET0131 , \u2_R4_reg[20]/NET0131 , \u2_R4_reg[21]/NET0131 , \u2_R4_reg[22]/NET0131 , \u2_R4_reg[23]/NET0131 , \u2_R4_reg[24]/NET0131 , \u2_R4_reg[25]/NET0131 , \u2_R4_reg[26]/NET0131 , \u2_R4_reg[27]/NET0131 , \u2_R4_reg[28]/NET0131 , \u2_R4_reg[29]/NET0131 , \u2_R4_reg[2]/NET0131 , \u2_R4_reg[30]/NET0131 , \u2_R4_reg[31]/P0001 , \u2_R4_reg[32]/NET0131 , \u2_R4_reg[3]/NET0131 , \u2_R4_reg[4]/NET0131 , \u2_R4_reg[5]/NET0131 , \u2_R4_reg[6]/NET0131 , \u2_R4_reg[7]/NET0131 , \u2_R4_reg[8]/NET0131 , \u2_R4_reg[9]/NET0131 , \u2_R5_reg[10]/NET0131 , \u2_R5_reg[11]/NET0131 , \u2_R5_reg[12]/NET0131 , \u2_R5_reg[13]/NET0131 , \u2_R5_reg[14]/NET0131 , \u2_R5_reg[15]/NET0131 , \u2_R5_reg[16]/NET0131 , \u2_R5_reg[17]/NET0131 , \u2_R5_reg[18]/NET0131 , \u2_R5_reg[19]/NET0131 , \u2_R5_reg[1]/NET0131 , \u2_R5_reg[20]/NET0131 , \u2_R5_reg[21]/NET0131 , \u2_R5_reg[22]/NET0131 , \u2_R5_reg[23]/NET0131 , \u2_R5_reg[24]/NET0131 , \u2_R5_reg[25]/NET0131 , \u2_R5_reg[26]/NET0131 , \u2_R5_reg[27]/NET0131 , \u2_R5_reg[28]/NET0131 , \u2_R5_reg[29]/NET0131 , \u2_R5_reg[2]/NET0131 , \u2_R5_reg[30]/NET0131 , \u2_R5_reg[31]/P0001 , \u2_R5_reg[32]/NET0131 , \u2_R5_reg[3]/NET0131 , \u2_R5_reg[4]/NET0131 , \u2_R5_reg[5]/NET0131 , \u2_R5_reg[6]/NET0131 , \u2_R5_reg[7]/NET0131 , \u2_R5_reg[8]/NET0131 , \u2_R5_reg[9]/NET0131 , \u2_R6_reg[10]/NET0131 , \u2_R6_reg[11]/NET0131 , \u2_R6_reg[12]/NET0131 , \u2_R6_reg[13]/NET0131 , \u2_R6_reg[14]/NET0131 , \u2_R6_reg[15]/NET0131 , \u2_R6_reg[16]/NET0131 , \u2_R6_reg[17]/NET0131 , \u2_R6_reg[18]/NET0131 , \u2_R6_reg[19]/NET0131 , \u2_R6_reg[1]/NET0131 , \u2_R6_reg[20]/NET0131 , \u2_R6_reg[21]/NET0131 , \u2_R6_reg[22]/NET0131 , \u2_R6_reg[23]/NET0131 , \u2_R6_reg[24]/NET0131 , \u2_R6_reg[25]/NET0131 , \u2_R6_reg[26]/NET0131 , \u2_R6_reg[27]/NET0131 , \u2_R6_reg[28]/NET0131 , \u2_R6_reg[29]/NET0131 , \u2_R6_reg[2]/NET0131 , \u2_R6_reg[30]/NET0131 , \u2_R6_reg[31]/P0001 , \u2_R6_reg[32]/NET0131 , \u2_R6_reg[3]/NET0131 , \u2_R6_reg[4]/NET0131 , \u2_R6_reg[5]/NET0131 , \u2_R6_reg[6]/NET0131 , \u2_R6_reg[7]/NET0131 , \u2_R6_reg[8]/NET0131 , \u2_R6_reg[9]/NET0131 , \u2_R7_reg[10]/NET0131 , \u2_R7_reg[11]/NET0131 , \u2_R7_reg[12]/NET0131 , \u2_R7_reg[13]/NET0131 , \u2_R7_reg[14]/NET0131 , \u2_R7_reg[15]/NET0131 , \u2_R7_reg[16]/NET0131 , \u2_R7_reg[17]/NET0131 , \u2_R7_reg[18]/NET0131 , \u2_R7_reg[19]/NET0131 , \u2_R7_reg[1]/NET0131 , \u2_R7_reg[20]/NET0131 , \u2_R7_reg[21]/NET0131 , \u2_R7_reg[22]/NET0131 , \u2_R7_reg[23]/NET0131 , \u2_R7_reg[24]/NET0131 , \u2_R7_reg[25]/NET0131 , \u2_R7_reg[26]/NET0131 , \u2_R7_reg[27]/NET0131 , \u2_R7_reg[28]/NET0131 , \u2_R7_reg[29]/NET0131 , \u2_R7_reg[2]/NET0131 , \u2_R7_reg[30]/NET0131 , \u2_R7_reg[31]/P0001 , \u2_R7_reg[32]/NET0131 , \u2_R7_reg[3]/NET0131 , \u2_R7_reg[4]/NET0131 , \u2_R7_reg[5]/NET0131 , \u2_R7_reg[6]/NET0131 , \u2_R7_reg[7]/NET0131 , \u2_R7_reg[8]/NET0131 , \u2_R7_reg[9]/NET0131 , \u2_R8_reg[10]/NET0131 , \u2_R8_reg[11]/NET0131 , \u2_R8_reg[12]/NET0131 , \u2_R8_reg[13]/NET0131 , \u2_R8_reg[14]/NET0131 , \u2_R8_reg[15]/NET0131 , \u2_R8_reg[16]/NET0131 , \u2_R8_reg[17]/NET0131 , \u2_R8_reg[18]/NET0131 , \u2_R8_reg[19]/NET0131 , \u2_R8_reg[1]/NET0131 , \u2_R8_reg[20]/NET0131 , \u2_R8_reg[21]/NET0131 , \u2_R8_reg[22]/NET0131 , \u2_R8_reg[23]/NET0131 , \u2_R8_reg[24]/NET0131 , \u2_R8_reg[25]/NET0131 , \u2_R8_reg[26]/NET0131 , \u2_R8_reg[27]/NET0131 , \u2_R8_reg[28]/NET0131 , \u2_R8_reg[29]/NET0131 , \u2_R8_reg[2]/NET0131 , \u2_R8_reg[30]/NET0131 , \u2_R8_reg[31]/P0001 , \u2_R8_reg[32]/NET0131 , \u2_R8_reg[3]/NET0131 , \u2_R8_reg[4]/NET0131 , \u2_R8_reg[5]/NET0131 , \u2_R8_reg[6]/NET0131 , \u2_R8_reg[7]/NET0131 , \u2_R8_reg[8]/NET0131 , \u2_R8_reg[9]/NET0131 , \u2_R9_reg[10]/NET0131 , \u2_R9_reg[11]/NET0131 , \u2_R9_reg[12]/NET0131 , \u2_R9_reg[13]/NET0131 , \u2_R9_reg[14]/NET0131 , \u2_R9_reg[15]/NET0131 , \u2_R9_reg[16]/NET0131 , \u2_R9_reg[17]/NET0131 , \u2_R9_reg[18]/NET0131 , \u2_R9_reg[19]/NET0131 , \u2_R9_reg[1]/NET0131 , \u2_R9_reg[20]/NET0131 , \u2_R9_reg[21]/NET0131 , \u2_R9_reg[22]/NET0131 , \u2_R9_reg[23]/NET0131 , \u2_R9_reg[24]/NET0131 , \u2_R9_reg[25]/NET0131 , \u2_R9_reg[26]/NET0131 , \u2_R9_reg[27]/NET0131 , \u2_R9_reg[28]/NET0131 , \u2_R9_reg[29]/NET0131 , \u2_R9_reg[2]/NET0131 , \u2_R9_reg[30]/NET0131 , \u2_R9_reg[31]/P0001 , \u2_R9_reg[32]/NET0131 , \u2_R9_reg[3]/NET0131 , \u2_R9_reg[4]/NET0131 , \u2_R9_reg[5]/NET0131 , \u2_R9_reg[6]/NET0131 , \u2_R9_reg[7]/NET0131 , \u2_R9_reg[8]/NET0131 , \u2_R9_reg[9]/NET0131 , \u2_desIn_r_reg[0]/NET0131 , \u2_desIn_r_reg[10]/P0001 , \u2_desIn_r_reg[11]/NET0131 , \u2_desIn_r_reg[12]/NET0131 , \u2_desIn_r_reg[13]/NET0131 , \u2_desIn_r_reg[14]/NET0131 , \u2_desIn_r_reg[15]/NET0131 , \u2_desIn_r_reg[16]/NET0131 , \u2_desIn_r_reg[17]/NET0131 , \u2_desIn_r_reg[18]/NET0131 , \u2_desIn_r_reg[19]/NET0131 , \u2_desIn_r_reg[1]/NET0131 , \u2_desIn_r_reg[20]/NET0131 , \u2_desIn_r_reg[21]/NET0131 , \u2_desIn_r_reg[22]/NET0131 , \u2_desIn_r_reg[23]/NET0131 , \u2_desIn_r_reg[24]/NET0131 , \u2_desIn_r_reg[25]/NET0131 , \u2_desIn_r_reg[26]/NET0131 , \u2_desIn_r_reg[27]/NET0131 , \u2_desIn_r_reg[28]/NET0131 , \u2_desIn_r_reg[29]/NET0131 , \u2_desIn_r_reg[2]/NET0131 , \u2_desIn_r_reg[30]/NET0131 , \u2_desIn_r_reg[31]/NET0131 , \u2_desIn_r_reg[32]/NET0131 , \u2_desIn_r_reg[33]/NET0131 , \u2_desIn_r_reg[34]/NET0131 , \u2_desIn_r_reg[35]/NET0131 , \u2_desIn_r_reg[36]/NET0131 , \u2_desIn_r_reg[37]/NET0131 , \u2_desIn_r_reg[38]/NET0131 , \u2_desIn_r_reg[39]/NET0131 , \u2_desIn_r_reg[3]/NET0131 , \u2_desIn_r_reg[40]/NET0131 , \u2_desIn_r_reg[41]/NET0131 , \u2_desIn_r_reg[42]/NET0131 , \u2_desIn_r_reg[43]/NET0131 , \u2_desIn_r_reg[44]/NET0131 , \u2_desIn_r_reg[45]/NET0131 , \u2_desIn_r_reg[46]/NET0131 , \u2_desIn_r_reg[47]/NET0131 , \u2_desIn_r_reg[48]/NET0131 , \u2_desIn_r_reg[49]/NET0131 , \u2_desIn_r_reg[4]/NET0131 , \u2_desIn_r_reg[50]/NET0131 , \u2_desIn_r_reg[51]/NET0131 , \u2_desIn_r_reg[52]/NET0131 , \u2_desIn_r_reg[53]/NET0131 , \u2_desIn_r_reg[54]/NET0131 , \u2_desIn_r_reg[55]/NET0131 , \u2_desIn_r_reg[56]/NET0131 , \u2_desIn_r_reg[57]/NET0131 , \u2_desIn_r_reg[58]/NET0131 , \u2_desIn_r_reg[59]/NET0131 , \u2_desIn_r_reg[5]/NET0131 , \u2_desIn_r_reg[60]/NET0131 , \u2_desIn_r_reg[61]/NET0131 , \u2_desIn_r_reg[62]/NET0131 , \u2_desIn_r_reg[63]/NET0131 , \u2_desIn_r_reg[6]/NET0131 , \u2_desIn_r_reg[7]/NET0131 , \u2_desIn_r_reg[8]/NET0131 , \u2_desIn_r_reg[9]/NET0131 , \u2_key_r_reg[0]/NET0131 , \u2_key_r_reg[10]/NET0131 , \u2_key_r_reg[11]/NET0131 , \u2_key_r_reg[12]/NET0131 , \u2_key_r_reg[13]/NET0131 , \u2_key_r_reg[14]/NET0131 , \u2_key_r_reg[15]/NET0131 , \u2_key_r_reg[16]/NET0131 , \u2_key_r_reg[17]/NET0131 , \u2_key_r_reg[18]/NET0131 , \u2_key_r_reg[19]/NET0131 , \u2_key_r_reg[1]/NET0131 , \u2_key_r_reg[20]/NET0131 , \u2_key_r_reg[21]/NET0131 , \u2_key_r_reg[22]/NET0131 , \u2_key_r_reg[23]/NET0131 , \u2_key_r_reg[24]/NET0131 , \u2_key_r_reg[25]/NET0131 , \u2_key_r_reg[26]/NET0131 , \u2_key_r_reg[27]/NET0131 , \u2_key_r_reg[28]/NET0131 , \u2_key_r_reg[29]/NET0131 , \u2_key_r_reg[2]/NET0131 , \u2_key_r_reg[30]/NET0131 , \u2_key_r_reg[31]/NET0131 , \u2_key_r_reg[32]/NET0131 , \u2_key_r_reg[33]/NET0131 , \u2_key_r_reg[34]/NET0131 , \u2_key_r_reg[35]/P0001 , \u2_key_r_reg[36]/NET0131 , \u2_key_r_reg[37]/NET0131 , \u2_key_r_reg[38]/NET0131 , \u2_key_r_reg[39]/P0001 , \u2_key_r_reg[3]/NET0131 , \u2_key_r_reg[40]/NET0131 , \u2_key_r_reg[41]/NET0131 , \u2_key_r_reg[42]/P0001 , \u2_key_r_reg[43]/NET0131 , \u2_key_r_reg[44]/NET0131 , \u2_key_r_reg[45]/NET0131 , \u2_key_r_reg[46]/NET0131 , \u2_key_r_reg[47]/NET0131 , \u2_key_r_reg[48]/NET0131 , \u2_key_r_reg[49]/NET0131 , \u2_key_r_reg[4]/NET0131 , \u2_key_r_reg[50]/NET0131 , \u2_key_r_reg[51]/NET0131 , \u2_key_r_reg[52]/NET0131 , \u2_key_r_reg[53]/NET0131 , \u2_key_r_reg[54]/NET0131 , \u2_key_r_reg[55]/NET0131 , \u2_key_r_reg[5]/NET0131 , \u2_key_r_reg[6]/NET0131 , \u2_key_r_reg[7]/NET0131 , \u2_key_r_reg[8]/NET0131 , \u2_key_r_reg[9]/NET0131 , \u2_uk_K_r0_reg[0]/NET0131 , \u2_uk_K_r0_reg[10]/NET0131 , \u2_uk_K_r0_reg[11]/NET0131 , \u2_uk_K_r0_reg[12]/NET0131 , \u2_uk_K_r0_reg[13]/NET0131 , \u2_uk_K_r0_reg[14]/NET0131 , \u2_uk_K_r0_reg[15]/NET0131 , \u2_uk_K_r0_reg[16]/NET0131 , \u2_uk_K_r0_reg[17]/NET0131 , \u2_uk_K_r0_reg[18]/NET0131 , \u2_uk_K_r0_reg[19]/NET0131 , \u2_uk_K_r0_reg[20]/NET0131 , \u2_uk_K_r0_reg[21]/NET0131 , \u2_uk_K_r0_reg[22]/NET0131 , \u2_uk_K_r0_reg[23]/NET0131 , \u2_uk_K_r0_reg[24]/P0001 , \u2_uk_K_r0_reg[25]/P0001 , \u2_uk_K_r0_reg[26]/NET0131 , \u2_uk_K_r0_reg[27]/NET0131 , \u2_uk_K_r0_reg[28]/NET0131 , \u2_uk_K_r0_reg[29]/NET0131 , \u2_uk_K_r0_reg[2]/NET0131 , \u2_uk_K_r0_reg[30]/NET0131 , \u2_uk_K_r0_reg[31]/NET0131 , \u2_uk_K_r0_reg[32]/NET0131 , \u2_uk_K_r0_reg[33]/NET0131 , \u2_uk_K_r0_reg[34]/NET0131 , \u2_uk_K_r0_reg[35]/NET0131 , \u2_uk_K_r0_reg[36]/NET0131 , \u2_uk_K_r0_reg[37]/NET0131 , \u2_uk_K_r0_reg[38]/NET0131 , \u2_uk_K_r0_reg[39]/NET0131 , \u2_uk_K_r0_reg[3]/NET0131 , \u2_uk_K_r0_reg[40]/NET0131 , \u2_uk_K_r0_reg[41]/NET0131 , \u2_uk_K_r0_reg[42]/NET0131 , \u2_uk_K_r0_reg[43]/NET0131 , \u2_uk_K_r0_reg[44]/NET0131 , \u2_uk_K_r0_reg[45]/NET0131 , \u2_uk_K_r0_reg[46]/NET0131 , \u2_uk_K_r0_reg[47]/NET0131 , \u2_uk_K_r0_reg[48]/NET0131 , \u2_uk_K_r0_reg[49]/NET0131 , \u2_uk_K_r0_reg[4]/NET0131 , \u2_uk_K_r0_reg[50]/NET0131 , \u2_uk_K_r0_reg[51]/NET0131 , \u2_uk_K_r0_reg[52]/P0001 , \u2_uk_K_r0_reg[54]/NET0131 , \u2_uk_K_r0_reg[55]/NET0131 , \u2_uk_K_r0_reg[5]/NET0131 , \u2_uk_K_r0_reg[6]/NET0131 , \u2_uk_K_r0_reg[7]/NET0131 , \u2_uk_K_r0_reg[8]/NET0131 , \u2_uk_K_r0_reg[9]/NET0131 , \u2_uk_K_r10_reg[0]/NET0131 , \u2_uk_K_r10_reg[10]/NET0131 , \u2_uk_K_r10_reg[11]/NET0131 , \u2_uk_K_r10_reg[12]/NET0131 , \u2_uk_K_r10_reg[14]/NET0131 , \u2_uk_K_r10_reg[15]/NET0131 , \u2_uk_K_r10_reg[16]/NET0131 , \u2_uk_K_r10_reg[17]/NET0131 , \u2_uk_K_r10_reg[18]/NET0131 , \u2_uk_K_r10_reg[19]/NET0131 , \u2_uk_K_r10_reg[1]/NET0131 , \u2_uk_K_r10_reg[20]/NET0131 , \u2_uk_K_r10_reg[21]/NET0131 , \u2_uk_K_r10_reg[22]/NET0131 , \u2_uk_K_r10_reg[23]/NET0131 , \u2_uk_K_r10_reg[24]/NET0131 , \u2_uk_K_r10_reg[25]/NET0131 , \u2_uk_K_r10_reg[26]/NET0131 , \u2_uk_K_r10_reg[27]/NET0131 , \u2_uk_K_r10_reg[28]/NET0131 , \u2_uk_K_r10_reg[29]/NET0131 , \u2_uk_K_r10_reg[2]/NET0131 , \u2_uk_K_r10_reg[30]/NET0131 , \u2_uk_K_r10_reg[31]/NET0131 , \u2_uk_K_r10_reg[32]/NET0131 , \u2_uk_K_r10_reg[33]/NET0131 , \u2_uk_K_r10_reg[34]/NET0131 , \u2_uk_K_r10_reg[35]/NET0131 , \u2_uk_K_r10_reg[36]/NET0131 , \u2_uk_K_r10_reg[37]/NET0131 , \u2_uk_K_r10_reg[38]/NET0131 , \u2_uk_K_r10_reg[39]/NET0131 , \u2_uk_K_r10_reg[3]/NET0131 , \u2_uk_K_r10_reg[40]/NET0131 , \u2_uk_K_r10_reg[41]/NET0131 , \u2_uk_K_r10_reg[42]/NET0131 , \u2_uk_K_r10_reg[43]/NET0131 , \u2_uk_K_r10_reg[44]/NET0131 , \u2_uk_K_r10_reg[45]/P0001 , \u2_uk_K_r10_reg[46]/NET0131 , \u2_uk_K_r10_reg[47]/NET0131 , \u2_uk_K_r10_reg[48]/NET0131 , \u2_uk_K_r10_reg[49]/NET0131 , \u2_uk_K_r10_reg[4]/NET0131 , \u2_uk_K_r10_reg[50]/NET0131 , \u2_uk_K_r10_reg[51]/NET0131 , \u2_uk_K_r10_reg[52]/NET0131 , \u2_uk_K_r10_reg[53]/NET0131 , \u2_uk_K_r10_reg[54]/NET0131 , \u2_uk_K_r10_reg[55]/NET0131 , \u2_uk_K_r10_reg[5]/NET0131 , \u2_uk_K_r10_reg[6]/NET0131 , \u2_uk_K_r10_reg[7]/NET0131 , \u2_uk_K_r10_reg[8]/NET0131 , \u2_uk_K_r10_reg[9]/NET0131 , \u2_uk_K_r11_reg[0]/NET0131 , \u2_uk_K_r11_reg[10]/NET0131 , \u2_uk_K_r11_reg[11]/NET0131 , \u2_uk_K_r11_reg[12]/NET0131 , \u2_uk_K_r11_reg[13]/NET0131 , \u2_uk_K_r11_reg[14]/NET0131 , \u2_uk_K_r11_reg[15]/NET0131 , \u2_uk_K_r11_reg[16]/NET0131 , \u2_uk_K_r11_reg[17]/NET0131 , \u2_uk_K_r11_reg[18]/NET0131 , \u2_uk_K_r11_reg[19]/NET0131 , \u2_uk_K_r11_reg[1]/NET0131 , \u2_uk_K_r11_reg[20]/NET0131 , \u2_uk_K_r11_reg[21]/NET0131 , \u2_uk_K_r11_reg[22]/NET0131 , \u2_uk_K_r11_reg[23]/NET0131 , \u2_uk_K_r11_reg[24]/NET0131 , \u2_uk_K_r11_reg[25]/NET0131 , \u2_uk_K_r11_reg[26]/NET0131 , \u2_uk_K_r11_reg[27]/NET0131 , \u2_uk_K_r11_reg[28]/NET0131 , \u2_uk_K_r11_reg[29]/NET0131 , \u2_uk_K_r11_reg[2]/NET0131 , \u2_uk_K_r11_reg[31]/NET0131 , \u2_uk_K_r11_reg[32]/NET0131 , \u2_uk_K_r11_reg[33]/NET0131 , \u2_uk_K_r11_reg[34]/NET0131 , \u2_uk_K_r11_reg[35]/NET0131 , \u2_uk_K_r11_reg[36]/NET0131 , \u2_uk_K_r11_reg[37]/NET0131 , \u2_uk_K_r11_reg[38]/NET0131 , \u2_uk_K_r11_reg[39]/NET0131 , \u2_uk_K_r11_reg[3]/NET0131 , \u2_uk_K_r11_reg[40]/NET0131 , \u2_uk_K_r11_reg[41]/NET0131 , \u2_uk_K_r11_reg[42]/NET0131 , \u2_uk_K_r11_reg[43]/NET0131 , \u2_uk_K_r11_reg[44]/NET0131 , \u2_uk_K_r11_reg[45]/NET0131 , \u2_uk_K_r11_reg[46]/NET0131 , \u2_uk_K_r11_reg[47]/NET0131 , \u2_uk_K_r11_reg[48]/NET0131 , \u2_uk_K_r11_reg[49]/NET0131 , \u2_uk_K_r11_reg[4]/NET0131 , \u2_uk_K_r11_reg[50]/NET0131 , \u2_uk_K_r11_reg[51]/NET0131 , \u2_uk_K_r11_reg[52]/NET0131 , \u2_uk_K_r11_reg[53]/P0001 , \u2_uk_K_r11_reg[54]/NET0131 , \u2_uk_K_r11_reg[55]/NET0131 , \u2_uk_K_r11_reg[5]/NET0131 , \u2_uk_K_r11_reg[6]/NET0131 , \u2_uk_K_r11_reg[7]/NET0131 , \u2_uk_K_r11_reg[8]/NET0131 , \u2_uk_K_r11_reg[9]/NET0131 , \u2_uk_K_r12_reg[0]/NET0131 , \u2_uk_K_r12_reg[10]/P0001 , \u2_uk_K_r12_reg[11]/NET0131 , \u2_uk_K_r12_reg[12]/NET0131 , \u2_uk_K_r12_reg[13]/NET0131 , \u2_uk_K_r12_reg[14]/NET0131 , \u2_uk_K_r12_reg[15]/NET0131 , \u2_uk_K_r12_reg[16]/NET0131 , \u2_uk_K_r12_reg[17]/NET0131 , \u2_uk_K_r12_reg[18]/NET0131 , \u2_uk_K_r12_reg[19]/NET0131 , \u2_uk_K_r12_reg[1]/NET0131 , \u2_uk_K_r12_reg[20]/NET0131 , \u2_uk_K_r12_reg[21]/NET0131 , \u2_uk_K_r12_reg[22]/NET0131 , \u2_uk_K_r12_reg[23]/NET0131 , \u2_uk_K_r12_reg[24]/NET0131 , \u2_uk_K_r12_reg[25]/NET0131 , \u2_uk_K_r12_reg[26]/NET0131 , \u2_uk_K_r12_reg[27]/NET0131 , \u2_uk_K_r12_reg[28]/NET0131 , \u2_uk_K_r12_reg[29]/NET0131 , \u2_uk_K_r12_reg[2]/NET0131 , \u2_uk_K_r12_reg[30]/NET0131 , \u2_uk_K_r12_reg[31]/NET0131 , \u2_uk_K_r12_reg[32]/NET0131 , \u2_uk_K_r12_reg[33]/NET0131 , \u2_uk_K_r12_reg[34]/NET0131 , \u2_uk_K_r12_reg[35]/NET0131 , \u2_uk_K_r12_reg[36]/NET0131 , \u2_uk_K_r12_reg[37]/NET0131 , \u2_uk_K_r12_reg[38]/NET0131 , \u2_uk_K_r12_reg[3]/NET0131 , \u2_uk_K_r12_reg[40]/NET0131 , \u2_uk_K_r12_reg[41]/NET0131 , \u2_uk_K_r12_reg[42]/NET0131 , \u2_uk_K_r12_reg[43]/NET0131 , \u2_uk_K_r12_reg[44]/P0001 , \u2_uk_K_r12_reg[45]/NET0131 , \u2_uk_K_r12_reg[46]/NET0131 , \u2_uk_K_r12_reg[47]/NET0131 , \u2_uk_K_r12_reg[48]/NET0131 , \u2_uk_K_r12_reg[49]/NET0131 , \u2_uk_K_r12_reg[4]/NET0131 , \u2_uk_K_r12_reg[50]/NET0131 , \u2_uk_K_r12_reg[51]/NET0131 , \u2_uk_K_r12_reg[52]/NET0131 , \u2_uk_K_r12_reg[53]/NET0131 , \u2_uk_K_r12_reg[54]/NET0131 , \u2_uk_K_r12_reg[55]/NET0131 , \u2_uk_K_r12_reg[5]/NET0131 , \u2_uk_K_r12_reg[6]/NET0131 , \u2_uk_K_r12_reg[7]/P0001 , \u2_uk_K_r12_reg[8]/NET0131 , \u2_uk_K_r12_reg[9]/NET0131 , \u2_uk_K_r13_reg[0]/NET0131 , \u2_uk_K_r13_reg[10]/NET0131 , \u2_uk_K_r13_reg[11]/NET0131 , \u2_uk_K_r13_reg[12]/NET0131 , \u2_uk_K_r13_reg[13]/NET0131 , \u2_uk_K_r13_reg[14]/NET0131 , \u2_uk_K_r13_reg[15]/NET0131 , \u2_uk_K_r13_reg[16]/NET0131 , \u2_uk_K_r13_reg[17]/NET0131 , \u2_uk_K_r13_reg[18]/NET0131 , \u2_uk_K_r13_reg[19]/NET0131 , \u2_uk_K_r13_reg[20]/NET0131 , \u2_uk_K_r13_reg[21]/NET0131 , \u2_uk_K_r13_reg[22]/NET0131 , \u2_uk_K_r13_reg[23]/NET0131 , \u2_uk_K_r13_reg[24]/NET0131 , \u2_uk_K_r13_reg[25]/P0001 , \u2_uk_K_r13_reg[26]/NET0131 , \u2_uk_K_r13_reg[27]/NET0131 , \u2_uk_K_r13_reg[28]/NET0131 , \u2_uk_K_r13_reg[29]/NET0131 , \u2_uk_K_r13_reg[2]/NET0131 , \u2_uk_K_r13_reg[30]/NET0131 , \u2_uk_K_r13_reg[31]/NET0131 , \u2_uk_K_r13_reg[32]/NET0131 , \u2_uk_K_r13_reg[33]/NET0131 , \u2_uk_K_r13_reg[34]/NET0131 , \u2_uk_K_r13_reg[35]/NET0131 , \u2_uk_K_r13_reg[36]/NET0131 , \u2_uk_K_r13_reg[37]/NET0131 , \u2_uk_K_r13_reg[38]/NET0131 , \u2_uk_K_r13_reg[39]/NET0131 , \u2_uk_K_r13_reg[3]/NET0131 , \u2_uk_K_r13_reg[40]/NET0131 , \u2_uk_K_r13_reg[41]/NET0131 , \u2_uk_K_r13_reg[42]/NET0131 , \u2_uk_K_r13_reg[43]/NET0131 , \u2_uk_K_r13_reg[44]/NET0131 , \u2_uk_K_r13_reg[45]/NET0131 , \u2_uk_K_r13_reg[46]/NET0131 , \u2_uk_K_r13_reg[47]/NET0131 , \u2_uk_K_r13_reg[48]/NET0131 , \u2_uk_K_r13_reg[49]/NET0131 , \u2_uk_K_r13_reg[4]/NET0131 , \u2_uk_K_r13_reg[50]/NET0131 , \u2_uk_K_r13_reg[51]/NET0131 , \u2_uk_K_r13_reg[52]/NET0131 , \u2_uk_K_r13_reg[54]/NET0131 , \u2_uk_K_r13_reg[55]/NET0131 , \u2_uk_K_r13_reg[5]/NET0131 , \u2_uk_K_r13_reg[6]/NET0131 , \u2_uk_K_r13_reg[7]/NET0131 , \u2_uk_K_r13_reg[8]/NET0131 , \u2_uk_K_r13_reg[9]/NET0131 , \u2_uk_K_r14_reg[0]/NET0131 , \u2_uk_K_r14_reg[10]/P0001 , \u2_uk_K_r14_reg[11]/NET0131 , \u2_uk_K_r14_reg[12]/NET0131 , \u2_uk_K_r14_reg[13]/NET0131 , \u2_uk_K_r14_reg[14]/NET0131 , \u2_uk_K_r14_reg[15]/NET0131 , \u2_uk_K_r14_reg[16]/NET0131 , \u2_uk_K_r14_reg[17]/NET0131 , \u2_uk_K_r14_reg[18]/NET0131 , \u2_uk_K_r14_reg[19]/NET0131 , \u2_uk_K_r14_reg[1]/NET0131 , \u2_uk_K_r14_reg[20]/NET0131 , \u2_uk_K_r14_reg[21]/NET0131 , \u2_uk_K_r14_reg[22]/NET0131 , \u2_uk_K_r14_reg[23]/NET0131 , \u2_uk_K_r14_reg[24]/NET0131 , \u2_uk_K_r14_reg[25]/NET0131 , \u2_uk_K_r14_reg[26]/NET0131 , \u2_uk_K_r14_reg[27]/NET0131 , \u2_uk_K_r14_reg[28]/NET0131 , \u2_uk_K_r14_reg[29]/NET0131 , \u2_uk_K_r14_reg[2]/NET0131 , \u2_uk_K_r14_reg[30]/NET0131 , \u2_uk_K_r14_reg[31]/NET0131 , \u2_uk_K_r14_reg[32]/NET0131 , \u2_uk_K_r14_reg[33]/NET0131 , \u2_uk_K_r14_reg[34]/NET0131 , \u2_uk_K_r14_reg[35]/P0001 , \u2_uk_K_r14_reg[36]/NET0131 , \u2_uk_K_r14_reg[37]/NET0131 , \u2_uk_K_r14_reg[38]/NET0131 , \u2_uk_K_r14_reg[39]/P0001 , \u2_uk_K_r14_reg[3]/NET0131 , \u2_uk_K_r14_reg[40]/NET0131 , \u2_uk_K_r14_reg[41]/NET0131 , \u2_uk_K_r14_reg[42]/P0001 , \u2_uk_K_r14_reg[43]/NET0131 , \u2_uk_K_r14_reg[44]/NET0131 , \u2_uk_K_r14_reg[45]/NET0131 , \u2_uk_K_r14_reg[46]/NET0131 , \u2_uk_K_r14_reg[47]/NET0131 , \u2_uk_K_r14_reg[48]/NET0131 , \u2_uk_K_r14_reg[49]/P0001 , \u2_uk_K_r14_reg[4]/NET0131 , \u2_uk_K_r14_reg[50]/NET0131 , \u2_uk_K_r14_reg[51]/NET0131 , \u2_uk_K_r14_reg[52]/NET0131 , \u2_uk_K_r14_reg[53]/NET0131 , \u2_uk_K_r14_reg[54]/NET0131 , \u2_uk_K_r14_reg[55]/NET0131 , \u2_uk_K_r14_reg[5]/NET0131 , \u2_uk_K_r14_reg[6]/NET0131 , \u2_uk_K_r14_reg[7]/NET0131 , \u2_uk_K_r14_reg[8]/NET0131 , \u2_uk_K_r14_reg[9]/NET0131 , \u2_uk_K_r1_reg[0]/NET0131 , \u2_uk_K_r1_reg[10]/P0001 , \u2_uk_K_r1_reg[11]/NET0131 , \u2_uk_K_r1_reg[12]/NET0131 , \u2_uk_K_r1_reg[13]/NET0131 , \u2_uk_K_r1_reg[14]/NET0131 , \u2_uk_K_r1_reg[15]/NET0131 , \u2_uk_K_r1_reg[16]/NET0131 , \u2_uk_K_r1_reg[17]/NET0131 , \u2_uk_K_r1_reg[18]/NET0131 , \u2_uk_K_r1_reg[19]/NET0131 , \u2_uk_K_r1_reg[1]/NET0131 , \u2_uk_K_r1_reg[20]/NET0131 , \u2_uk_K_r1_reg[21]/NET0131 , \u2_uk_K_r1_reg[22]/NET0131 , \u2_uk_K_r1_reg[23]/NET0131 , \u2_uk_K_r1_reg[24]/NET0131 , \u2_uk_K_r1_reg[25]/NET0131 , \u2_uk_K_r1_reg[26]/NET0131 , \u2_uk_K_r1_reg[27]/NET0131 , \u2_uk_K_r1_reg[28]/NET0131 , \u2_uk_K_r1_reg[29]/NET0131 , \u2_uk_K_r1_reg[2]/NET0131 , \u2_uk_K_r1_reg[30]/NET0131 , \u2_uk_K_r1_reg[31]/NET0131 , \u2_uk_K_r1_reg[32]/NET0131 , \u2_uk_K_r1_reg[33]/NET0131 , \u2_uk_K_r1_reg[34]/NET0131 , \u2_uk_K_r1_reg[35]/NET0131 , \u2_uk_K_r1_reg[36]/NET0131 , \u2_uk_K_r1_reg[37]/NET0131 , \u2_uk_K_r1_reg[38]/NET0131 , \u2_uk_K_r1_reg[3]/NET0131 , \u2_uk_K_r1_reg[40]/NET0131 , \u2_uk_K_r1_reg[41]/NET0131 , \u2_uk_K_r1_reg[42]/NET0131 , \u2_uk_K_r1_reg[43]/NET0131 , \u2_uk_K_r1_reg[44]/P0001 , \u2_uk_K_r1_reg[45]/NET0131 , \u2_uk_K_r1_reg[46]/NET0131 , \u2_uk_K_r1_reg[47]/NET0131 , \u2_uk_K_r1_reg[48]/NET0131 , \u2_uk_K_r1_reg[49]/NET0131 , \u2_uk_K_r1_reg[4]/NET0131 , \u2_uk_K_r1_reg[50]/NET0131 , \u2_uk_K_r1_reg[51]/NET0131 , \u2_uk_K_r1_reg[52]/NET0131 , \u2_uk_K_r1_reg[53]/NET0131 , \u2_uk_K_r1_reg[54]/NET0131 , \u2_uk_K_r1_reg[55]/NET0131 , \u2_uk_K_r1_reg[5]/NET0131 , \u2_uk_K_r1_reg[6]/NET0131 , \u2_uk_K_r1_reg[7]/P0001 , \u2_uk_K_r1_reg[8]/NET0131 , \u2_uk_K_r1_reg[9]/NET0131 , \u2_uk_K_r2_reg[0]/NET0131 , \u2_uk_K_r2_reg[10]/NET0131 , \u2_uk_K_r2_reg[11]/NET0131 , \u2_uk_K_r2_reg[12]/NET0131 , \u2_uk_K_r2_reg[13]/NET0131 , \u2_uk_K_r2_reg[14]/NET0131 , \u2_uk_K_r2_reg[15]/NET0131 , \u2_uk_K_r2_reg[16]/NET0131 , \u2_uk_K_r2_reg[17]/NET0131 , \u2_uk_K_r2_reg[18]/NET0131 , \u2_uk_K_r2_reg[19]/NET0131 , \u2_uk_K_r2_reg[1]/NET0131 , \u2_uk_K_r2_reg[20]/NET0131 , \u2_uk_K_r2_reg[21]/NET0131 , \u2_uk_K_r2_reg[22]/NET0131 , \u2_uk_K_r2_reg[23]/NET0131 , \u2_uk_K_r2_reg[24]/NET0131 , \u2_uk_K_r2_reg[25]/NET0131 , \u2_uk_K_r2_reg[26]/NET0131 , \u2_uk_K_r2_reg[27]/NET0131 , \u2_uk_K_r2_reg[28]/NET0131 , \u2_uk_K_r2_reg[29]/NET0131 , \u2_uk_K_r2_reg[2]/NET0131 , \u2_uk_K_r2_reg[31]/NET0131 , \u2_uk_K_r2_reg[32]/NET0131 , \u2_uk_K_r2_reg[33]/NET0131 , \u2_uk_K_r2_reg[34]/NET0131 , \u2_uk_K_r2_reg[35]/NET0131 , \u2_uk_K_r2_reg[36]/NET0131 , \u2_uk_K_r2_reg[37]/NET0131 , \u2_uk_K_r2_reg[38]/NET0131 , \u2_uk_K_r2_reg[39]/NET0131 , \u2_uk_K_r2_reg[3]/NET0131 , \u2_uk_K_r2_reg[40]/NET0131 , \u2_uk_K_r2_reg[41]/NET0131 , \u2_uk_K_r2_reg[42]/NET0131 , \u2_uk_K_r2_reg[43]/NET0131 , \u2_uk_K_r2_reg[44]/NET0131 , \u2_uk_K_r2_reg[45]/NET0131 , \u2_uk_K_r2_reg[46]/NET0131 , \u2_uk_K_r2_reg[47]/NET0131 , \u2_uk_K_r2_reg[48]/NET0131 , \u2_uk_K_r2_reg[49]/NET0131 , \u2_uk_K_r2_reg[4]/NET0131 , \u2_uk_K_r2_reg[50]/NET0131 , \u2_uk_K_r2_reg[51]/NET0131 , \u2_uk_K_r2_reg[52]/NET0131 , \u2_uk_K_r2_reg[53]/P0001 , \u2_uk_K_r2_reg[54]/NET0131 , \u2_uk_K_r2_reg[55]/NET0131 , \u2_uk_K_r2_reg[5]/NET0131 , \u2_uk_K_r2_reg[6]/NET0131 , \u2_uk_K_r2_reg[7]/NET0131 , \u2_uk_K_r2_reg[8]/NET0131 , \u2_uk_K_r2_reg[9]/NET0131 , \u2_uk_K_r3_reg[0]/NET0131 , \u2_uk_K_r3_reg[10]/NET0131 , \u2_uk_K_r3_reg[11]/NET0131 , \u2_uk_K_r3_reg[12]/NET0131 , \u2_uk_K_r3_reg[14]/NET0131 , \u2_uk_K_r3_reg[15]/NET0131 , \u2_uk_K_r3_reg[16]/NET0131 , \u2_uk_K_r3_reg[17]/NET0131 , \u2_uk_K_r3_reg[18]/NET0131 , \u2_uk_K_r3_reg[19]/NET0131 , \u2_uk_K_r3_reg[1]/NET0131 , \u2_uk_K_r3_reg[20]/NET0131 , \u2_uk_K_r3_reg[21]/NET0131 , \u2_uk_K_r3_reg[22]/NET0131 , \u2_uk_K_r3_reg[23]/NET0131 , \u2_uk_K_r3_reg[24]/NET0131 , \u2_uk_K_r3_reg[25]/NET0131 , \u2_uk_K_r3_reg[26]/NET0131 , \u2_uk_K_r3_reg[27]/NET0131 , \u2_uk_K_r3_reg[28]/NET0131 , \u2_uk_K_r3_reg[29]/NET0131 , \u2_uk_K_r3_reg[2]/NET0131 , \u2_uk_K_r3_reg[30]/NET0131 , \u2_uk_K_r3_reg[31]/NET0131 , \u2_uk_K_r3_reg[32]/NET0131 , \u2_uk_K_r3_reg[33]/NET0131 , \u2_uk_K_r3_reg[34]/NET0131 , \u2_uk_K_r3_reg[35]/NET0131 , \u2_uk_K_r3_reg[36]/NET0131 , \u2_uk_K_r3_reg[37]/NET0131 , \u2_uk_K_r3_reg[38]/NET0131 , \u2_uk_K_r3_reg[39]/NET0131 , \u2_uk_K_r3_reg[3]/NET0131 , \u2_uk_K_r3_reg[40]/NET0131 , \u2_uk_K_r3_reg[41]/NET0131 , \u2_uk_K_r3_reg[42]/NET0131 , \u2_uk_K_r3_reg[43]/NET0131 , \u2_uk_K_r3_reg[44]/NET0131 , \u2_uk_K_r3_reg[45]/P0001 , \u2_uk_K_r3_reg[46]/NET0131 , \u2_uk_K_r3_reg[47]/NET0131 , \u2_uk_K_r3_reg[48]/NET0131 , \u2_uk_K_r3_reg[49]/NET0131 , \u2_uk_K_r3_reg[4]/NET0131 , \u2_uk_K_r3_reg[50]/NET0131 , \u2_uk_K_r3_reg[51]/NET0131 , \u2_uk_K_r3_reg[52]/NET0131 , \u2_uk_K_r3_reg[53]/NET0131 , \u2_uk_K_r3_reg[54]/NET0131 , \u2_uk_K_r3_reg[55]/NET0131 , \u2_uk_K_r3_reg[5]/NET0131 , \u2_uk_K_r3_reg[6]/NET0131 , \u2_uk_K_r3_reg[7]/NET0131 , \u2_uk_K_r3_reg[8]/NET0131 , \u2_uk_K_r3_reg[9]/NET0131 , \u2_uk_K_r4_reg[0]/P0001 , \u2_uk_K_r4_reg[10]/NET0131 , \u2_uk_K_r4_reg[11]/NET0131 , \u2_uk_K_r4_reg[12]/NET0131 , \u2_uk_K_r4_reg[13]/NET0131 , \u2_uk_K_r4_reg[14]/NET0131 , \u2_uk_K_r4_reg[15]/NET0131 , \u2_uk_K_r4_reg[16]/NET0131 , \u2_uk_K_r4_reg[17]/NET0131 , \u2_uk_K_r4_reg[18]/NET0131 , \u2_uk_K_r4_reg[19]/NET0131 , \u2_uk_K_r4_reg[1]/NET0131 , \u2_uk_K_r4_reg[20]/NET0131 , \u2_uk_K_r4_reg[21]/NET0131 , \u2_uk_K_r4_reg[22]/NET0131 , \u2_uk_K_r4_reg[23]/NET0131 , \u2_uk_K_r4_reg[25]/NET0131 , \u2_uk_K_r4_reg[26]/NET0131 , \u2_uk_K_r4_reg[27]/P0001 , \u2_uk_K_r4_reg[28]/NET0131 , \u2_uk_K_r4_reg[29]/NET0131 , \u2_uk_K_r4_reg[30]/NET0131 , \u2_uk_K_r4_reg[31]/P0001 , \u2_uk_K_r4_reg[32]/NET0131 , \u2_uk_K_r4_reg[33]/NET0131 , \u2_uk_K_r4_reg[34]/NET0131 , \u2_uk_K_r4_reg[35]/NET0131 , \u2_uk_K_r4_reg[36]/NET0131 , \u2_uk_K_r4_reg[37]/NET0131 , \u2_uk_K_r4_reg[38]/NET0131 , \u2_uk_K_r4_reg[39]/NET0131 , \u2_uk_K_r4_reg[3]/NET0131 , \u2_uk_K_r4_reg[40]/NET0131 , \u2_uk_K_r4_reg[41]/NET0131 , \u2_uk_K_r4_reg[42]/NET0131 , \u2_uk_K_r4_reg[43]/NET0131 , \u2_uk_K_r4_reg[44]/NET0131 , \u2_uk_K_r4_reg[45]/NET0131 , \u2_uk_K_r4_reg[46]/NET0131 , \u2_uk_K_r4_reg[47]/NET0131 , \u2_uk_K_r4_reg[48]/NET0131 , \u2_uk_K_r4_reg[49]/NET0131 , \u2_uk_K_r4_reg[4]/NET0131 , \u2_uk_K_r4_reg[50]/NET0131 , \u2_uk_K_r4_reg[51]/NET0131 , \u2_uk_K_r4_reg[52]/NET0131 , \u2_uk_K_r4_reg[53]/NET0131 , \u2_uk_K_r4_reg[54]/NET0131 , \u2_uk_K_r4_reg[55]/NET0131 , \u2_uk_K_r4_reg[5]/NET0131 , \u2_uk_K_r4_reg[6]/NET0131 , \u2_uk_K_r4_reg[7]/NET0131 , \u2_uk_K_r4_reg[8]/NET0131 , \u2_uk_K_r4_reg[9]/NET0131 , \u2_uk_K_r5_reg[0]/NET0131 , \u2_uk_K_r5_reg[10]/NET0131 , \u2_uk_K_r5_reg[11]/NET0131 , \u2_uk_K_r5_reg[12]/NET0131 , \u2_uk_K_r5_reg[13]/P0001 , \u2_uk_K_r5_reg[14]/NET0131 , \u2_uk_K_r5_reg[15]/NET0131 , \u2_uk_K_r5_reg[16]/NET0131 , \u2_uk_K_r5_reg[17]/NET0131 , \u2_uk_K_r5_reg[18]/NET0131 , \u2_uk_K_r5_reg[19]/NET0131 , \u2_uk_K_r5_reg[1]/NET0131 , \u2_uk_K_r5_reg[20]/NET0131 , \u2_uk_K_r5_reg[21]/NET0131 , \u2_uk_K_r5_reg[22]/NET0131 , \u2_uk_K_r5_reg[23]/NET0131 , \u2_uk_K_r5_reg[24]/NET0131 , \u2_uk_K_r5_reg[25]/NET0131 , \u2_uk_K_r5_reg[26]/NET0131 , \u2_uk_K_r5_reg[27]/NET0131 , \u2_uk_K_r5_reg[28]/NET0131 , \u2_uk_K_r5_reg[29]/NET0131 , \u2_uk_K_r5_reg[2]/NET0131 , \u2_uk_K_r5_reg[30]/NET0131 , \u2_uk_K_r5_reg[31]/NET0131 , \u2_uk_K_r5_reg[32]/NET0131 , \u2_uk_K_r5_reg[33]/NET0131 , \u2_uk_K_r5_reg[34]/NET0131 , \u2_uk_K_r5_reg[35]/NET0131 , \u2_uk_K_r5_reg[36]/NET0131 , \u2_uk_K_r5_reg[37]/P0001 , \u2_uk_K_r5_reg[38]/NET0131 , \u2_uk_K_r5_reg[39]/NET0131 , \u2_uk_K_r5_reg[3]/NET0131 , \u2_uk_K_r5_reg[40]/NET0131 , \u2_uk_K_r5_reg[41]/NET0131 , \u2_uk_K_r5_reg[42]/NET0131 , \u2_uk_K_r5_reg[43]/NET0131 , \u2_uk_K_r5_reg[44]/NET0131 , \u2_uk_K_r5_reg[46]/NET0131 , \u2_uk_K_r5_reg[47]/NET0131 , \u2_uk_K_r5_reg[48]/NET0131 , \u2_uk_K_r5_reg[49]/NET0131 , \u2_uk_K_r5_reg[4]/NET0131 , \u2_uk_K_r5_reg[50]/NET0131 , \u2_uk_K_r5_reg[51]/NET0131 , \u2_uk_K_r5_reg[52]/NET0131 , \u2_uk_K_r5_reg[53]/NET0131 , \u2_uk_K_r5_reg[54]/NET0131 , \u2_uk_K_r5_reg[55]/NET0131 , \u2_uk_K_r5_reg[5]/NET0131 , \u2_uk_K_r5_reg[6]/NET0131 , \u2_uk_K_r5_reg[7]/NET0131 , \u2_uk_K_r5_reg[8]/NET0131 , \u2_uk_K_r5_reg[9]/P0001 , \u2_uk_K_r6_reg[0]/NET0131 , \u2_uk_K_r6_reg[10]/NET0131 , \u2_uk_K_r6_reg[11]/NET0131 , \u2_uk_K_r6_reg[12]/NET0131 , \u2_uk_K_r6_reg[13]/NET0131 , \u2_uk_K_r6_reg[14]/NET0131 , \u2_uk_K_r6_reg[15]/NET0131 , \u2_uk_K_r6_reg[16]/NET0131 , \u2_uk_K_r6_reg[17]/NET0131 , \u2_uk_K_r6_reg[18]/NET0131 , \u2_uk_K_r6_reg[19]/NET0131 , \u2_uk_K_r6_reg[1]/NET0131 , \u2_uk_K_r6_reg[20]/NET0131 , \u2_uk_K_r6_reg[21]/NET0131 , \u2_uk_K_r6_reg[22]/NET0131 , \u2_uk_K_r6_reg[23]/P0001 , \u2_uk_K_r6_reg[24]/NET0131 , \u2_uk_K_r6_reg[25]/NET0131 , \u2_uk_K_r6_reg[26]/NET0131 , \u2_uk_K_r6_reg[27]/NET0131 , \u2_uk_K_r6_reg[28]/NET0131 , \u2_uk_K_r6_reg[29]/NET0131 , \u2_uk_K_r6_reg[2]/NET0131 , \u2_uk_K_r6_reg[30]/P0001 , \u2_uk_K_r6_reg[31]/NET0131 , \u2_uk_K_r6_reg[32]/NET0131 , \u2_uk_K_r6_reg[33]/NET0131 , \u2_uk_K_r6_reg[34]/NET0131 , \u2_uk_K_r6_reg[35]/NET0131 , \u2_uk_K_r6_reg[36]/NET0131 , \u2_uk_K_r6_reg[37]/NET0131 , \u2_uk_K_r6_reg[38]/NET0131 , \u2_uk_K_r6_reg[39]/NET0131 , \u2_uk_K_r6_reg[3]/NET0131 , \u2_uk_K_r6_reg[40]/NET0131 , \u2_uk_K_r6_reg[41]/NET0131 , \u2_uk_K_r6_reg[42]/NET0131 , \u2_uk_K_r6_reg[43]/NET0131 , \u2_uk_K_r6_reg[44]/NET0131 , \u2_uk_K_r6_reg[45]/NET0131 , \u2_uk_K_r6_reg[46]/NET0131 , \u2_uk_K_r6_reg[47]/NET0131 , \u2_uk_K_r6_reg[48]/NET0131 , \u2_uk_K_r6_reg[49]/NET0131 , \u2_uk_K_r6_reg[4]/NET0131 , \u2_uk_K_r6_reg[50]/NET0131 , \u2_uk_K_r6_reg[51]/NET0131 , \u2_uk_K_r6_reg[52]/NET0131 , \u2_uk_K_r6_reg[53]/NET0131 , \u2_uk_K_r6_reg[54]/NET0131 , \u2_uk_K_r6_reg[55]/P0001 , \u2_uk_K_r6_reg[5]/NET0131 , \u2_uk_K_r6_reg[6]/NET0131 , \u2_uk_K_r6_reg[7]/NET0131 , \u2_uk_K_r6_reg[8]/NET0131 , \u2_uk_K_r6_reg[9]/NET0131 , \u2_uk_K_r7_reg[0]/NET0131 , \u2_uk_K_r7_reg[10]/NET0131 , \u2_uk_K_r7_reg[11]/NET0131 , \u2_uk_K_r7_reg[12]/NET0131 , \u2_uk_K_r7_reg[13]/NET0131 , \u2_uk_K_r7_reg[14]/NET0131 , \u2_uk_K_r7_reg[15]/NET0131 , \u2_uk_K_r7_reg[16]/NET0131 , \u2_uk_K_r7_reg[17]/NET0131 , \u2_uk_K_r7_reg[18]/NET0131 , \u2_uk_K_r7_reg[19]/NET0131 , \u2_uk_K_r7_reg[1]/NET0131 , \u2_uk_K_r7_reg[20]/NET0131 , \u2_uk_K_r7_reg[21]/NET0131 , \u2_uk_K_r7_reg[22]/NET0131 , \u2_uk_K_r7_reg[23]/P0001 , \u2_uk_K_r7_reg[24]/NET0131 , \u2_uk_K_r7_reg[25]/NET0131 , \u2_uk_K_r7_reg[26]/NET0131 , \u2_uk_K_r7_reg[27]/NET0131 , \u2_uk_K_r7_reg[28]/NET0131 , \u2_uk_K_r7_reg[29]/NET0131 , \u2_uk_K_r7_reg[2]/NET0131 , \u2_uk_K_r7_reg[30]/P0001 , \u2_uk_K_r7_reg[31]/NET0131 , \u2_uk_K_r7_reg[32]/NET0131 , \u2_uk_K_r7_reg[33]/NET0131 , \u2_uk_K_r7_reg[34]/NET0131 , \u2_uk_K_r7_reg[35]/NET0131 , \u2_uk_K_r7_reg[36]/NET0131 , \u2_uk_K_r7_reg[37]/NET0131 , \u2_uk_K_r7_reg[38]/NET0131 , \u2_uk_K_r7_reg[39]/NET0131 , \u2_uk_K_r7_reg[3]/NET0131 , \u2_uk_K_r7_reg[40]/NET0131 , \u2_uk_K_r7_reg[41]/NET0131 , \u2_uk_K_r7_reg[42]/NET0131 , \u2_uk_K_r7_reg[43]/NET0131 , \u2_uk_K_r7_reg[44]/NET0131 , \u2_uk_K_r7_reg[45]/NET0131 , \u2_uk_K_r7_reg[46]/NET0131 , \u2_uk_K_r7_reg[47]/NET0131 , \u2_uk_K_r7_reg[48]/NET0131 , \u2_uk_K_r7_reg[49]/NET0131 , \u2_uk_K_r7_reg[4]/NET0131 , \u2_uk_K_r7_reg[50]/NET0131 , \u2_uk_K_r7_reg[51]/NET0131 , \u2_uk_K_r7_reg[52]/NET0131 , \u2_uk_K_r7_reg[53]/NET0131 , \u2_uk_K_r7_reg[54]/NET0131 , \u2_uk_K_r7_reg[55]/P0001 , \u2_uk_K_r7_reg[5]/NET0131 , \u2_uk_K_r7_reg[6]/NET0131 , \u2_uk_K_r7_reg[7]/NET0131 , \u2_uk_K_r7_reg[8]/NET0131 , \u2_uk_K_r7_reg[9]/NET0131 , \u2_uk_K_r8_reg[0]/NET0131 , \u2_uk_K_r8_reg[10]/NET0131 , \u2_uk_K_r8_reg[11]/NET0131 , \u2_uk_K_r8_reg[12]/NET0131 , \u2_uk_K_r8_reg[13]/P0001 , \u2_uk_K_r8_reg[14]/NET0131 , \u2_uk_K_r8_reg[15]/NET0131 , \u2_uk_K_r8_reg[16]/NET0131 , \u2_uk_K_r8_reg[17]/NET0131 , \u2_uk_K_r8_reg[18]/NET0131 , \u2_uk_K_r8_reg[19]/NET0131 , \u2_uk_K_r8_reg[1]/NET0131 , \u2_uk_K_r8_reg[20]/NET0131 , \u2_uk_K_r8_reg[21]/NET0131 , \u2_uk_K_r8_reg[22]/NET0131 , \u2_uk_K_r8_reg[23]/NET0131 , \u2_uk_K_r8_reg[24]/NET0131 , \u2_uk_K_r8_reg[25]/NET0131 , \u2_uk_K_r8_reg[26]/NET0131 , \u2_uk_K_r8_reg[27]/NET0131 , \u2_uk_K_r8_reg[28]/NET0131 , \u2_uk_K_r8_reg[29]/NET0131 , \u2_uk_K_r8_reg[2]/NET0131 , \u2_uk_K_r8_reg[30]/NET0131 , \u2_uk_K_r8_reg[31]/NET0131 , \u2_uk_K_r8_reg[32]/NET0131 , \u2_uk_K_r8_reg[33]/NET0131 , \u2_uk_K_r8_reg[34]/NET0131 , \u2_uk_K_r8_reg[35]/NET0131 , \u2_uk_K_r8_reg[36]/NET0131 , \u2_uk_K_r8_reg[37]/P0001 , \u2_uk_K_r8_reg[38]/NET0131 , \u2_uk_K_r8_reg[39]/NET0131 , \u2_uk_K_r8_reg[3]/NET0131 , \u2_uk_K_r8_reg[40]/NET0131 , \u2_uk_K_r8_reg[41]/NET0131 , \u2_uk_K_r8_reg[42]/NET0131 , \u2_uk_K_r8_reg[43]/NET0131 , \u2_uk_K_r8_reg[44]/NET0131 , \u2_uk_K_r8_reg[46]/NET0131 , \u2_uk_K_r8_reg[47]/NET0131 , \u2_uk_K_r8_reg[48]/NET0131 , \u2_uk_K_r8_reg[49]/NET0131 , \u2_uk_K_r8_reg[4]/NET0131 , \u2_uk_K_r8_reg[50]/NET0131 , \u2_uk_K_r8_reg[51]/NET0131 , \u2_uk_K_r8_reg[52]/NET0131 , \u2_uk_K_r8_reg[53]/NET0131 , \u2_uk_K_r8_reg[54]/NET0131 , \u2_uk_K_r8_reg[55]/NET0131 , \u2_uk_K_r8_reg[5]/NET0131 , \u2_uk_K_r8_reg[6]/NET0131 , \u2_uk_K_r8_reg[7]/NET0131 , \u2_uk_K_r8_reg[8]/NET0131 , \u2_uk_K_r8_reg[9]/NET0131 , \u2_uk_K_r9_reg[0]/P0001 , \u2_uk_K_r9_reg[10]/NET0131 , \u2_uk_K_r9_reg[11]/NET0131 , \u2_uk_K_r9_reg[12]/NET0131 , \u2_uk_K_r9_reg[13]/NET0131 , \u2_uk_K_r9_reg[14]/NET0131 , \u2_uk_K_r9_reg[15]/NET0131 , \u2_uk_K_r9_reg[16]/NET0131 , \u2_uk_K_r9_reg[17]/NET0131 , \u2_uk_K_r9_reg[18]/NET0131 , \u2_uk_K_r9_reg[19]/NET0131 , \u2_uk_K_r9_reg[1]/NET0131 , \u2_uk_K_r9_reg[20]/NET0131 , \u2_uk_K_r9_reg[21]/NET0131 , \u2_uk_K_r9_reg[22]/NET0131 , \u2_uk_K_r9_reg[23]/NET0131 , \u2_uk_K_r9_reg[25]/NET0131 , \u2_uk_K_r9_reg[26]/NET0131 , \u2_uk_K_r9_reg[27]/NET0131 , \u2_uk_K_r9_reg[28]/NET0131 , \u2_uk_K_r9_reg[29]/NET0131 , \u2_uk_K_r9_reg[30]/NET0131 , \u2_uk_K_r9_reg[31]/P0001 , \u2_uk_K_r9_reg[32]/NET0131 , \u2_uk_K_r9_reg[33]/NET0131 , \u2_uk_K_r9_reg[34]/NET0131 , \u2_uk_K_r9_reg[35]/NET0131 , \u2_uk_K_r9_reg[36]/NET0131 , \u2_uk_K_r9_reg[37]/NET0131 , \u2_uk_K_r9_reg[38]/NET0131 , \u2_uk_K_r9_reg[39]/NET0131 , \u2_uk_K_r9_reg[3]/NET0131 , \u2_uk_K_r9_reg[40]/NET0131 , \u2_uk_K_r9_reg[41]/NET0131 , \u2_uk_K_r9_reg[42]/NET0131 , \u2_uk_K_r9_reg[43]/NET0131 , \u2_uk_K_r9_reg[44]/NET0131 , \u2_uk_K_r9_reg[45]/NET0131 , \u2_uk_K_r9_reg[46]/NET0131 , \u2_uk_K_r9_reg[47]/NET0131 , \u2_uk_K_r9_reg[48]/NET0131 , \u2_uk_K_r9_reg[49]/NET0131 , \u2_uk_K_r9_reg[4]/NET0131 , \u2_uk_K_r9_reg[50]/NET0131 , \u2_uk_K_r9_reg[51]/NET0131 , \u2_uk_K_r9_reg[52]/NET0131 , \u2_uk_K_r9_reg[53]/NET0131 , \u2_uk_K_r9_reg[54]/NET0131 , \u2_uk_K_r9_reg[55]/NET0131 , \u2_uk_K_r9_reg[5]/NET0131 , \u2_uk_K_r9_reg[6]/NET0131 , \u2_uk_K_r9_reg[7]/NET0131 , \u2_uk_K_r9_reg[8]/NET0131 , \u2_uk_K_r9_reg[9]/NET0131 , \_al_n0 , \_al_n1 , \g16/_0_ , \g191647/_3_ , \g191648/_3_ , \g191819/_3_ , \g191821/_0_ , \g191940/_3_ , \g191941/_0_ , \g191942/_0_ , \g191944/_0_ , \g191945/_0_ , \g191946/_0_ , \g191947/_3_ , \g191948/_0_ , \g191949/_0_ , \g191950/_0_ , \g191951/_3_ , \g191952/_0_ , \g192015/_3_ , \g192016/_3_ , \g192017/_3_ , \g192018/_3_ , \g192019/_3_ , \g192020/_0_ , \g192021/_3_ , \g192022/_0_ , \g192047/_0_ , \g192048/_0_ , \g192049/_0_ , \g192050/_0_ , \g192051/_0_ , \g192081/_0_ , \g193428/_3_ , \g193720/_0_ , \g193721/_0_ , \g193877/_0_ , \g193878/_0_ , \g193879/_0_ , \g193880/_3_ , \g193881/_0_ , \g193882/_0_ , \g193998/_0_ , \g193999/_0_ , \g194000/_3_ , \g194001/_0_ , \g194002/_0_ , \g194003/_0_ , \g194004/_0_ , \g194005/_0_ , \g194006/_0_ , \g194007/_0_ , \g194008/_0_ , \g194009/_0_ , \g194010/_0_ , \g194055/_3_ , \g194056/_3_ , \g194057/_0_ , \g194058/_0_ , \g194059/_0_ , \g194060/_0_ , \g194090/_0_ , \g194091/_0_ , \g194092/_0_ , \g194093/_0_ , \g195671/_0_ , \g195672/_3_ , \g195868/_0_ , \g195869/_0_ , \g195870/_0_ , \g196010/_0_ , \g196011/_0_ , \g196012/_0_ , \g196013/_0_ , \g196014/_0_ , \g196015/_0_ , \g196016/_0_ , \g196017/_0_ , \g196018/_0_ , \g196019/_3_ , \g196020/_0_ , \g196021/_0_ , \g196022/_0_ , \g196096/_3_ , \g196097/_0_ , \g196098/_0_ , \g196099/_0_ , \g196100/_3_ , \g196101/_0_ , \g196102/_0_ , \g196103/_0_ , \g196136/_0_ , \g196137/_0_ , \g196138/_0_ , \g196139/_0_ , \g196140/_0_ , \g196170/_0_ , \g197520/_3_ , \g197821/_0_ , \g197923/_0_ , \g197996/_0_ , \g197997/_3_ , \g197998/_0_ , \g197999/_0_ , \g198000/_0_ , \g198071/_0_ , \g198123/_0_ , \g198124/_0_ , \g198125/_0_ , \g198126/_0_ , \g198127/_0_ , \g198128/_0_ , \g198129/_0_ , \g198130/_0_ , \g198131/_0_ , \g198132/_0_ , \g198133/_0_ , \g198134/_3_ , \g198135/_0_ , \g198182/_0_ , \g198183/_3_ , \g198184/_0_ , \g198185/_0_ , \g198186/_0_ , \g198187/_0_ , \g198219/_0_ , \g198220/_0_ , \g198221/_0_ , \g198222/_0_ , \g199794/_0_ , \g199795/_3_ , \g200006/_0_ , \g200007/_0_ , \g200008/_0_ , \g200139/_0_ , \g200140/_0_ , \g200141/_0_ , \g200142/_0_ , \g200143/_0_ , \g200144/_0_ , \g200145/_0_ , \g200146/_0_ , \g200147/_0_ , \g200148/_0_ , \g200149/_0_ , \g200150/_3_ , \g200151/_0_ , \g200228/_3_ , \g200229/_0_ , \g200230/_0_ , \g200231/_0_ , \g200232/_3_ , \g200233/_0_ , \g200234/_0_ , \g200235/_0_ , \g200268/_0_ , \g200269/_0_ , \g200270/_0_ , \g200271/_0_ , \g200272/_0_ , \g200299/_0_ , \g201655/_3_ , \g201960/_0_ , \g201961/_0_ , \g202131/_0_ , \g202132/_0_ , \g202133/_3_ , \g202134/_0_ , \g202135/_0_ , \g202136/_0_ , \g202257/_0_ , \g202258/_0_ , \g202259/_3_ , \g202260/_0_ , \g202261/_0_ , \g202262/_0_ , \g202263/_0_ , \g202264/_0_ , \g202265/_0_ , \g202266/_0_ , \g202267/_0_ , \g202268/_0_ , \g202269/_0_ , \g202317/_0_ , \g202318/_3_ , \g202319/_0_ , \g202320/_0_ , \g202321/_0_ , \g202322/_0_ , \g202354/_0_ , \g202355/_0_ , \g202356/_0_ , \g202357/_0_ , \g203927/_0_ , \g203928/_3_ , \g204142/_0_ , \g204143/_0_ , \g204144/_0_ , \g204275/_0_ , \g204276/_0_ , \g204277/_0_ , \g204278/_0_ , \g204279/_0_ , \g204280/_0_ , \g204281/_0_ , \g204282/_0_ , \g204283/_0_ , \g204284/_0_ , \g204285/_0_ , \g204286/_3_ , \g204287/_0_ , \g204363/_3_ , \g204364/_0_ , \g204365/_0_ , \g204366/_0_ , \g204367/_3_ , \g204368/_0_ , \g204369/_0_ , \g204370/_0_ , \g204403/_0_ , \g204404/_0_ , \g204405/_0_ , \g204406/_0_ , \g204407/_0_ , \g204434/_0_ , \g205833/_3_ , \g206103/_0_ , \g206104/_0_ , \g206266/_0_ , \g206267/_0_ , \g206268/_0_ , \g206269/_3_ , \g206270/_0_ , \g206271/_0_ , \g206387/_0_ , \g206388/_0_ , \g206389/_3_ , \g206390/_0_ , \g206391/_0_ , \g206392/_0_ , \g206393/_0_ , \g206394/_0_ , \g206395/_0_ , \g206396/_0_ , \g206397/_0_ , \g206398/_0_ , \g206399/_0_ , \g206446/_0_ , \g206447/_3_ , \g206448/_0_ , \g206449/_0_ , \g206450/_0_ , \g206451/_0_ , \g206483/_0_ , \g206484/_0_ , \g206485/_0_ , \g206486/_0_ , \g208069/_0_ , \g208070/_3_ , \g208253/_0_ , \g208254/_0_ , \g208255/_0_ , \g208406/_0_ , \g208407/_0_ , \g208408/_0_ , \g208409/_0_ , \g208410/_0_ , \g208411/_0_ , \g208412/_0_ , \g208413/_0_ , \g208414/_0_ , \g208415/_3_ , \g208416/_0_ , \g208417/_0_ , \g208418/_0_ , \g208493/_3_ , \g208494/_0_ , \g208495/_0_ , \g208496/_0_ , \g208497/_3_ , \g208498/_0_ , \g208499/_0_ , \g208500/_0_ , \g208533/_0_ , \g208534/_0_ , \g208535/_0_ , \g208536/_0_ , \g208537/_0_ , \g208564/_0_ , \g209938/_3_ , \g210205/_0_ , \g210206/_0_ , \g210380/_0_ , \g210381/_0_ , \g210382/_0_ , \g210383/_3_ , \g210384/_0_ , \g210385/_0_ , \g210499/_0_ , \g210500/_0_ , \g210501/_3_ , \g210502/_0_ , \g210503/_0_ , \g210504/_0_ , \g210505/_0_ , \g210506/_0_ , \g210507/_0_ , \g210508/_0_ , \g210509/_0_ , \g210510/_0_ , \g210511/_0_ , \g210558/_0_ , \g210559/_3_ , \g210560/_0_ , \g210561/_0_ , \g210562/_0_ , \g210563/_0_ , \g210595/_0_ , \g210596/_0_ , \g210597/_0_ , \g210598/_0_ , \g212159/_0_ , \g212160/_3_ , \g212384/_0_ , \g212385/_0_ , \g212386/_0_ , \g212536/_0_ , \g212537/_0_ , \g212538/_0_ , \g212539/_0_ , \g212540/_0_ , \g212541/_0_ , \g212542/_0_ , \g212543/_0_ , \g212544/_0_ , \g212545/_0_ , \g212546/_3_ , \g212547/_0_ , \g212623/_3_ , \g212624/_0_ , \g212625/_0_ , \g212626/_0_ , \g212627/_0_ , \g212628/_3_ , \g212629/_0_ , \g212630/_0_ , \g212631/_0_ , \g212667/_0_ , \g212668/_0_ , \g212669/_0_ , \g212670/_0_ , \g212671/_0_ , \g212699/_0_ , \g214033/_3_ , \g214309/_3_ , \g214310/_0_ , \g214494/_0_ , \g214495/_0_ , \g214496/_0_ , \g214497/_3_ , \g214632/_0_ , \g214633/_0_ , \g214634/_3_ , \g214635/_0_ , \g214636/_0_ , \g214637/_0_ , \g214638/_0_ , \g214639/_0_ , \g214640/_0_ , \g214641/_0_ , \g214642/_0_ , \g214643/_0_ , \g214691/_0_ , \g214692/_0_ , \g214693/_3_ , \g214694/_0_ , \g214695/_0_ , \g214696/_0_ , \g214697/_0_ , \g214729/_0_ , \g214730/_0_ , \g214731/_0_ , \g214732/_0_ , \g214733/_0_ , \g216157/_0_ , \g216158/_3_ , \g216492/_0_ , \g216493/_0_ , \g216671/_0_ , \g216672/_0_ , \g216673/_0_ , \g216674/_0_ , \g216675/_0_ , \g216676/_3_ , \g216677/_0_ , \g216735/_0_ , \g216736/_3_ , \g216737/_0_ , \g216738/_0_ , \g216739/_0_ , \g216740/_0_ , \g216741/_0_ , \g216742/_0_ , \g216743/_0_ , \g216744/_0_ , \g216745/_0_ , \g216746/_3_ , \g216747/_0_ , \g216748/_0_ , \g216749/_0_ , \g216788/_0_ , \g216789/_0_ , \g216790/_0_ , \g216791/_0_ , \g216792/_0_ , \g216829/_0_ , \g218407/_3_ , \g218408/_0_ , \g218423/_3_ , \g218601/_0_ , \g218602/_0_ , \g218603/_0_ , \g218604/_0_ , \g218724/_0_ , \g218725/_0_ , \g218726/_0_ , \g218727/_0_ , \g218728/_0_ , \g218729/_0_ , \g218730/_0_ , \g218731/_0_ , \g218732/_0_ , \g218733/_0_ , \g218734/_0_ , \g218735/_3_ , \g218736/_0_ , \g218808/_3_ , \g218809/_0_ , \g218810/_0_ , \g218811/_3_ , \g218812/_0_ , \g218813/_0_ , \g218814/_0_ , \g218846/_0_ , \g218847/_0_ , \g218848/_0_ , \g218849/_0_ , \g218877/_0_ , \g22/_0_ , \g220545/_0_ , \g220546/_3_ , \g220725/_3_ , \g220726/_0_ , \g220793/_0_ , \g220794/_0_ , \g220795/_0_ , \g220796/_0_ , \g220797/_0_ , \g220798/_0_ , \g220799/_0_ , \g220800/_0_ , \g220801/_0_ , \g220802/_0_ , \g220803/_0_ , \g220804/_3_ , \g220805/_0_ , \g220806/_0_ , \g220807/_0_ , \g220872/_3_ , \g220873/_0_ , \g220874/_3_ , \g220875/_0_ , \g220876/_0_ , \g220877/_0_ , \g220921/_0_ , \g220922/_0_ , \g220923/_0_ , \g220924/_0_ , \g220925/_0_ , \g220926/_0_ , \g220969/_0_ , \g221011/_3_ , \g221039/_3_ , \g221086/_3_ , \g221131/_0_ , \g224010/_3_ , \g224368/_3_ , \g224369/_3_ , \g224532/_0_ , \g224533/_0_ , \g224534/_0_ , \g224535/_3_ , \g224536/_0_ , \g224537/_0_ , \g224640/_3_ , \g224641/_0_ , \g224642/_0_ , \g224643/_3_ , \g224644/_0_ , \g224645/_0_ , \g224646/_3_ , \g224647/_0_ , \g224648/_3_ , \g224649/_0_ , \g224650/_0_ , \g224651/_0_ , \g224652/_0_ , \g224690/_0_ , \g224691/_3_ , \g224692/_3_ , \g224693/_0_ , \g224694/_0_ , \g224695/_3_ , \g224723/_0_ , \g224724/_0_ , \g224725/_0_ , \g224726/_0_ , \g226372/_0_ , \g226373/_3_ , \g226549/_3_ , \g226550/_0_ , \g226616/_0_ , \g226635/_0_ , \g226636/_0_ , \g226637/_0_ , \g226638/_0_ , \g226639/_0_ , \g226640/_0_ , \g226641/_3_ , \g226642/_0_ , \g226643/_0_ , \g226644/_0_ , \g226645/_0_ , \g226646/_0_ , \g226692/_3_ , \g226693/_0_ , \g226694/_3_ , \g226695/_3_ , \g226696/_3_ , \g226697/_0_ , \g226698/_0_ , \g226699/_0_ , \g226728/_0_ , \g226729/_0_ , \g226730/_0_ , \g226731/_0_ , \g226732/_0_ , \g226759/_0_ , \g228250/_0_ , \g228396/_0_ , \g228397/_0_ , \g228566/_0_ , \g228567/_0_ , \g228568/_0_ , \g228609/_0_ , \g228610/_3_ , \g228688/_0_ , \g228689/_0_ , \g228690/_3_ , \g228691/_0_ , \g228692/_0_ , \g228693/_0_ , \g228694/_0_ , \g228695/_0_ , \g228696/_0_ , \g228697/_0_ , \g228698/_0_ , \g228699/_0_ , \g228700/_0_ , \g228748/_0_ , \g228749/_3_ , \g228750/_0_ , \g228751/_0_ , \g228752/_0_ , \g228753/_0_ , \g228784/_0_ , \g228785/_0_ , \g228786/_0_ , \g228787/_3_ , \g230339/_0_ , \g230340/_0_ , \g230546/_0_ , \g230580/_0_ , \g230679/_0_ , \g230680/_0_ , \g230681/_0_ , \g230682/_0_ , \g230683/_0_ , \g230684/_0_ , \g230685/_0_ , \g230686/_0_ , \g230687/_0_ , \g230688/_0_ , \g230689/_3_ , \g230690/_0_ , \g230710/_0_ , \g230766/_0_ , \g230767/_0_ , \g230768/_0_ , \g230769/_3_ , \g230770/_0_ , \g230771/_0_ , \g230772/_0_ , \g230773/_3_ , \g230810/_0_ , \g230811/_0_ , \g230812/_0_ , \g230813/_0_ , \g230814/_0_ , \g230840/_3_ , \g232196/_3_ , \g232469/_0_ , \g232470/_0_ , \g232633/_0_ , \g232635/_3_ , \g232636/_0_ , \g232637/_0_ , \g232691/_0_ , \g232747/_0_ , \g232748/_0_ , \g232749/_3_ , \g232750/_0_ , \g232751/_0_ , \g232752/_0_ , \g232753/_0_ , \g232754/_0_ , \g232755/_0_ , \g232756/_0_ , \g232757/_0_ , \g232758/_0_ , \g232759/_0_ , \g232804/_0_ , \g232805/_0_ , \g232806/_0_ , \g232807/_0_ , \g232808/_3_ , \g232809/_0_ , \g232841/_0_ , \g232842/_3_ , \g232843/_0_ , \g232844/_0_ , \g234520/_0_ , \g234687/_0_ , \g234688/_0_ , \g234689/_0_ , \g234764/_0_ , \g234765/_0_ , \g234766/_0_ , \g234767/_3_ , \g234768/_0_ , \g234769/_0_ , \g234770/_0_ , \g234771/_0_ , \g234772/_0_ , \g234773/_0_ , \g234774/_3_ , \g234775/_0_ , \g234776/_0_ , \g234824/_3_ , \g234825/_0_ , \g234826/_0_ , \g234827/_0_ , \g234828/_3_ , \g234829/_0_ , \g234830/_0_ , \g234831/_0_ , \g234867/_0_ , \g234868/_0_ , \g234869/_0_ , \g234870/_0_ , \g234896/_0_ , \g236294/_3_ , \g236541/_0_ , \g236542/_0_ , \g236724/_0_ , \g236725/_0_ , \g236726/_0_ , \g236727/_3_ , \g236728/_0_ , \g236729/_0_ , \g236821/_0_ , \g236822/_3_ , \g236823/_0_ , \g236824/_3_ , \g236825/_0_ , \g236826/_0_ , \g236827/_0_ , \g236828/_0_ , \g236829/_0_ , \g236830/_0_ , \g236831/_0_ , \g236832/_0_ , \g236877/_0_ , \g236878/_3_ , \g236879/_0_ , \g236880/_0_ , \g236881/_0_ , \g236882/_0_ , \g236914/_0_ , \g236915/_0_ , \g236916/_0_ , \g236917/_0_ , \g238530/_0_ , \g238531/_3_ , \g238723/_0_ , \g238724/_0_ , \g238725/_0_ , \g238840/_0_ , \g238841/_0_ , \g238842/_0_ , \g238843/_3_ , \g238844/_0_ , \g238845/_0_ , \g238846/_0_ , \g238847/_0_ , \g238848/_0_ , \g238849/_0_ , \g238850/_0_ , \g238851/_3_ , \g238852/_0_ , \g238924/_0_ , \g238925/_0_ , \g238926/_0_ , \g238927/_3_ , \g238928/_0_ , \g238929/_0_ , \g238930/_0_ , \g238965/_0_ , \g238966/_0_ , \g238967/_0_ , \g238968/_0_ , \g238969/_0_ , \g238996/_0_ , \g240353/_3_ , \g240640/_0_ , \g240641/_0_ , \g240813/_0_ , \g240814/_0_ , \g240815/_3_ , \g240816/_0_ , \g240817/_0_ , \g240818/_0_ , \g240925/_0_ , \g240926/_0_ , \g240927/_3_ , \g240928/_0_ , \g240929/_3_ , \g240930/_0_ , \g240931/_0_ , \g240932/_0_ , \g240933/_0_ , \g240934/_0_ , \g240935/_0_ , \g240936/_0_ , \g240937/_0_ , \g240984/_0_ , \g240985/_3_ , \g240986/_0_ , \g240987/_0_ , \g240988/_0_ , \g240989/_0_ , \g241021/_0_ , \g241022/_0_ , \g241023/_0_ , \g241024/_0_ , \g242616/_0_ , \g242617/_3_ , \g242815/_0_ , \g242816/_0_ , \g242817/_0_ , \g242955/_0_ , \g242956/_0_ , \g242957/_0_ , \g242958/_3_ , \g242959/_0_ , \g242960/_0_ , \g242961/_0_ , \g242962/_0_ , \g242963/_3_ , \g242964/_0_ , \g242965/_0_ , \g242966/_0_ , \g242967/_0_ , \g243037/_3_ , \g243038/_0_ , \g243039/_0_ , \g243040/_0_ , \g243041/_3_ , \g243042/_0_ , \g243043/_0_ , \g243044/_0_ , \g243078/_0_ , \g243079/_0_ , \g243080/_0_ , \g243081/_0_ , \g243082/_0_ , \g243109/_0_ , \g244465/_3_ , \g244753/_3_ , \g244754/_0_ , \g244924/_0_ , \g244925/_0_ , \g244926/_3_ , \g244927/_0_ , \g244928/_0_ , \g245035/_0_ , \g245036/_0_ , \g245037/_0_ , \g245038/_3_ , \g245039/_3_ , \g245040/_0_ , \g245041/_0_ , \g245043/_0_ , \g245045/_0_ , \g245046/_0_ , \g245047/_0_ , \g245092/_0_ , \g245093/_3_ , \g245094/_0_ , \g245095/_0_ , \g245096/_0_ , \g245097/_0_ , \g245129/_0_ , \g245130/_0_ , \g245131/_0_ , \g245132/_0_ , \g246715/_0_ , \g246716/_3_ , \g246911/_0_ , \g246912/_0_ , \g246913/_0_ , \g247057/_0_ , \g247058/_0_ , \g247059/_0_ , \g247060/_0_ , \g247061/_0_ , \g247062/_3_ , \g247063/_0_ , \g247064/_0_ , \g247065/_0_ , \g247066/_0_ , \g247067/_3_ , \g247068/_0_ , \g247069/_0_ , \g247137/_3_ , \g247138/_0_ , \g247139/_0_ , \g247140/_0_ , \g247141/_3_ , \g247142/_0_ , \g247143/_0_ , \g247144/_0_ , \g247179/_0_ , \g247180/_0_ , \g247181/_0_ , \g247182/_0_ , \g247183/_0_ , \g247210/_0_ , \g248581/_3_ , \g248828/_0_ , \g248829/_0_ , \g249033/_0_ , \g249035/_0_ , \g249036/_3_ , \g249037/_0_ , \g249038/_0_ , \g249147/_0_ , \g249148/_0_ , \g249149/_3_ , \g249150/_0_ , \g249152/_0_ , \g249153/_0_ , \g249155/_0_ , \g249156/_0_ , \g249157/_0_ , \g249200/_3_ , \g249201/_0_ , \g249202/_0_ , \g249203/_3_ , \g249204/_0_ , \g249205/_0_ , \g249206/_0_ , \g249207/_0_ , \g249239/_0_ , \g249240/_0_ , \g249241/_0_ , \g249242/_0_ , \g250815/_0_ , \g251006/_0_ , \g251007/_0_ , \g251008/_0_ , \g251009/_3_ , \g251160/_0_ , \g251161/_0_ , \g251162/_0_ , \g251163/_3_ , \g251164/_0_ , \g251165/_0_ , \g251166/_0_ , \g251167/_0_ , \g251168/_0_ , \g251169/_0_ , \g251170/_3_ , \g251171/_0_ , \g251245/_3_ , \g251246/_0_ , \g251247/_0_ , \g251248/_0_ , \g251249/_3_ , \g251250/_0_ , \g251251/_0_ , \g251252/_0_ , \g251286/_0_ , \g251287/_0_ , \g251288/_0_ , \g251289/_0_ , \g251290/_0_ , \g251291/_0_ , \g251318/_0_ , \g252698/_3_ , \g252942/_0_ , \g252943/_0_ , \g253118/_0_ , \g253119/_0_ , \g253120/_0_ , \g253121/_0_ , \g253122/_3_ , \g253123/_0_ , \g253236/_0_ , \g253237/_3_ , \g253238/_3_ , \g253239/_0_ , \g253240/_0_ , \g253241/_0_ , \g253242/_0_ , \g253243/_0_ , \g253244/_0_ , \g253245/_0_ , \g253246/_0_ , \g253247/_0_ , \g253248/_0_ , \g253306/_0_ , \g253307/_3_ , \g253308/_0_ , \g253309/_0_ , \g253310/_0_ , \g253311/_0_ , \g253356/_0_ , \g253357/_0_ , \g253358/_0_ , \g253359/_0_ , \g253436/_3_ , \g253437/_0_ , \g253438/_0_ , \g253469/_3_ , \g253470/_3_ , \g253471/_3_ , \g253521/_0_ , \g253522/_0_ , \g253523/_0_ , \g253524/_3_ , \g256730/_3_ , \g256731/_3_ , \g256927/_0_ , \g256928/_0_ , \g256929/_3_ , \g257049/_0_ , \g257050/_0_ , \g257051/_3_ , \g257052/_0_ , \g257053/_0_ , \g257054/_0_ , \g257055/_3_ , \g257056/_0_ , \g257057/_0_ , \g257058/_3_ , \g257059/_0_ , \g257060/_0_ , \g257082/_0_ , \g257125/_3_ , \g257126/_0_ , \g257127/_0_ , \g257128/_3_ , \g257129/_3_ , \g257130/_0_ , \g257131/_0_ , \g257132/_0_ , \g257163/_0_ , \g257164/_0_ , \g257165/_0_ , \g257166/_0_ , \g257167/_0_ , \g257194/_0_ , \g258552/_0_ , \g258850/_0_ , \g258851/_3_ , \g258993/_0_ , \g258994/_0_ , \g258995/_0_ , \g258996/_0_ , \g259026/_3_ , \g259027/_0_ , \g259105/_0_ , \g259106/_0_ , \g259107/_3_ , \g259108/_0_ , \g259109/_3_ , \g259110/_0_ , \g259111/_0_ , \g259112/_0_ , \g259113/_0_ , \g259114/_0_ , \g259115/_0_ , \g259116/_0_ , \g259117/_0_ , \g259163/_3_ , \g259164/_3_ , \g259165/_0_ , \g259166/_0_ , \g259167/_0_ , \g259168/_0_ , \g259197/_0_ , \g259198/_0_ , \g259199/_0_ , \g259200/_0_ , \g260774/_0_ , \g260792/_3_ , \g260991/_0_ , \g261013/_0_ , \g261070/_0_ , \g261125/_0_ , \g261126/_0_ , \g261128/_0_ , \g261129/_0_ , \g261130/_0_ , \g261131/_0_ , \g261132/_0_ , \g261133/_0_ , \g261134/_3_ , \g261135/_0_ , \g261136/_0_ , \g261158/_3_ , \g261206/_0_ , \g261207/_0_ , \g261208/_0_ , \g261209/_0_ , \g261210/_3_ , \g261211/_0_ , \g261212/_3_ , \g261213/_0_ , \g261248/_0_ , \g261249/_0_ , \g261250/_0_ , \g261251/_0_ , \g261252/_0_ , \g261279/_0_ , \g262658/_3_ , \g262949/_0_ , \g263008/_3_ , \g263092/_0_ , \g263093/_0_ , \g263099/_0_ , \g263100/_0_ , \g263101/_0_ , \g263159/_3_ , \g263204/_3_ , \g263205/_0_ , \g263206/_0_ , \g263208/_0_ , \g263209/_0_ , \g263210/_0_ , \g263211/_0_ , \g263212/_0_ , \g263213/_0_ , \g263214/_0_ , \g263215/_3_ , \g263216/_0_ , \g263260/_0_ , \g263261/_0_ , \g263262/_3_ , \g263263/_0_ , \g263264/_0_ , \g263265/_0_ , \g263297/_0_ , \g263298/_0_ , \g263299/_0_ , \g263300/_0_ , \g264930/_0_ , \g264946/_3_ , \g265143/_0_ , \g265144/_0_ , \g265152/_0_ , \g265222/_0_ , \g265223/_0_ , \g265224/_0_ , \g265225/_0_ , \g265226/_0_ , \g265227/_3_ , \g265228/_0_ , \g265229/_0_ , \g265230/_0_ , \g265231/_0_ , \g265232/_0_ , \g265233/_3_ , \g265234/_0_ , \g265306/_0_ , \g265307/_0_ , \g265308/_3_ , \g265309/_3_ , \g265310/_0_ , \g265311/_0_ , \g265312/_0_ , \g265313/_0_ , \g265348/_0_ , \g265349/_0_ , \g265350/_0_ , \g265351/_0_ , \g265379/_0_ , \g266965/_3_ , \g267049/_3_ , \g267050/_0_ , \g267215/_0_ , \g267216/_0_ , \g267263/_0_ , \g267264/_3_ , \g267265/_0_ , \g267266/_0_ , \g267314/_3_ , \g267315/_0_ , \g267316/_0_ , \g267317/_0_ , \g267318/_0_ , \g267319/_0_ , \g267320/_3_ , \g267321/_0_ , \g267322/_0_ , \g267324/_0_ , \g267325/_0_ , \g267326/_0_ , \g267372/_0_ , \g267373/_3_ , \g267374/_0_ , \g267375/_0_ , \g267376/_0_ , \g267377/_0_ , \g267409/_0_ , \g267410/_0_ , \g267411/_0_ , \g267412/_0_ , \g269004/_0_ , \g269099/_3_ , \g269202/_0_ , \g269226/_0_ , \g269333/_3_ , \g269334/_0_ , \g269335/_0_ , \g269355/_0_ , \g269356/_0_ , \g269357/_3_ , \g269358/_0_ , \g269359/_0_ , \g269360/_0_ , \g269361/_0_ , \g269362/_0_ , \g269363/_0_ , \g269364/_0_ , \g269414/_0_ , \g269415/_0_ , \g269416/_0_ , \g269417/_0_ , \g269418/_3_ , \g269419/_0_ , \g269420/_3_ , \g269421/_0_ , \g269456/_0_ , \g269457/_0_ , \g269458/_0_ , \g269459/_0_ , \g269460/_0_ , \g269487/_0_ , \g271006/_3_ , \g271186/_3_ , \g271187/_0_ , \g271299/_0_ , \g271300/_0_ , \g271301/_3_ , \g271302/_0_ , \g271303/_0_ , \g271352/_0_ , \g271410/_0_ , \g271411/_0_ , \g271412/_0_ , \g271413/_0_ , \g271414/_0_ , \g271415/_0_ , \g271416/_0_ , \g271417/_3_ , \g271418/_3_ , \g271419/_0_ , \g271420/_0_ , \g271421/_0_ , \g271422/_0_ , \g271468/_3_ , \g271469/_0_ , \g271470/_0_ , \g271471/_0_ , \g271472/_0_ , \g271473/_0_ , \g271505/_0_ , \g271506/_0_ , \g271507/_0_ , \g271508/_0_ , \g273135/_0_ , \g273136/_3_ , \g273362/_0_ , \g273373/_0_ , \g273374/_0_ , \g273431/_0_ , \g273432/_0_ , \g273433/_3_ , \g273434/_0_ , \g273435/_0_ , \g273436/_0_ , \g273437/_3_ , \g273438/_0_ , \g273439/_0_ , \g273441/_0_ , \g273442/_0_ , \g273443/_0_ , \g273515/_3_ , \g273516/_0_ , \g273517/_0_ , \g273518/_3_ , \g273519/_0_ , \g273520/_0_ , \g273521/_0_ , \g273522/_0_ , \g273557/_0_ , \g273558/_0_ , \g273559/_0_ , \g273560/_0_ , \g273561/_0_ , \g273588/_0_ , \g274960/_3_ , \g275266/_3_ , \g275327/_0_ , \g275396/_0_ , \g275397/_3_ , \g275398/_0_ , \g275455/_0_ , \g275456/_0_ , \g275463/_0_ , \g275510/_3_ , \g275511/_0_ , \g275512/_0_ , \g275513/_0_ , \g275514/_3_ , \g275515/_0_ , \g275516/_0_ , \g275517/_0_ , \g275518/_0_ , \g275519/_0_ , \g275520/_0_ , \g275521/_0_ , \g275522/_0_ , \g275568/_0_ , \g275569/_0_ , \g275570/_0_ , \g275571/_0_ , \g275572/_3_ , \g275573/_0_ , \g275605/_0_ , \g275606/_0_ , \g275607/_0_ , \g275608/_0_ , \g277189/_0_ , \g277294/_3_ , \g277367/_0_ , \g277456/_0_ , \g277457/_0_ , \g277512/_0_ , \g277513/_0_ , \g277514/_3_ , \g277515/_0_ , \g277516/_0_ , \g277517/_3_ , \g277518/_0_ , \g277519/_0_ , \g277520/_0_ , \g277521/_0_ , \g277594/_0_ , \g277595/_0_ , \g277596/_3_ , \g277597/_0_ , \g277598/_0_ , \g277599/_0_ , \g277600/_0_ , \g277601/_3_ , \g277635/_0_ , \g277636/_0_ , \g277637/_0_ , \g277638/_0_ , \g277639/_0_ , \g277666/_0_ , \g279090/_3_ , \g279330/_0_ , \g279331/_0_ , \g279493/_3_ , \g279494/_0_ , \g279495/_0_ , \g279502/_0_ , \g279503/_0_ , \g279504/_0_ , \g279590/_0_ , \g279591/_0_ , \g279592/_0_ , \g279593/_0_ , \g279594/_3_ , \g279595/_3_ , \g279596/_0_ , \g279597/_0_ , \g279598/_0_ , \g279599/_0_ , \g279600/_0_ , \g279601/_0_ , \g279602/_0_ , \g279649/_0_ , \g279650/_0_ , \g279651/_0_ , \g279652/_0_ , \g279653/_0_ , \g279654/_3_ , \g279686/_0_ , \g279687/_0_ , \g279688/_0_ , \g279689/_0_ , \g281329/_0_ , \g281394/_0_ , \g281483/_0_ , \g281498/_0_ , \g281532/_0_ , \g281616/_0_ , \g281617/_0_ , \g281618/_0_ , \g281619/_0_ , \g281620/_0_ , \g281621/_0_ , \g281622/_0_ , \g281623/_3_ , \g281624/_0_ , \g281642/_0_ , \g281643/_0_ , \g281644/_3_ , \g281645/_0_ , \g281696/_0_ , \g281697/_3_ , \g281698/_0_ , \g281699/_0_ , \g281700/_0_ , \g281701/_0_ , \g281702/_3_ , \g281703/_0_ , \g281799/_0_ , \g281800/_0_ , \g281801/_0_ , \g281802/_0_ , \g281803/_0_ , \g281965/_0_ , \g287377/_0_ , \g287867/_0_ , \g287899/_0_ , \g288304/_0_ , \g288334/_0_ , \g288350/_0_ , \g288351/_0_ , \g288352/_3_ , \g288353/_0_ , \g288668/_0_ , \g288669/_0_ , \g288670/_0_ , \g288671/_0_ , \g288673/_0_ , \g288674/_3_ , \g288675/_0_ , \g288676/_0_ , \g288677/_0_ , \g288678/_0_ , \g288679/_0_ , \g288680/_3_ , \g288889/_0_ , \g288890/_0_ , \g288891/_0_ , \g288892/_0_ , \g288893/_3_ , \g288894/_0_ , \g288895/_0_ , \g288984/_0_ , \g288985/_0_ , \g288986/_0_ , \g294974/_0_ , \g295054/_0_ , \g295601/_0_ , \g295607/_0_ , \g296036/_0_ , \g296037/_0_ , \g296038/_0_ , \g296039/_0_ , \g296040/_0_ , \g296041/_0_ , \g296042/_0_ , \g296043/_3_ , \g296044/_0_ , \g296045/_0_ , \g296046/_0_ , \g296047/_0_ , \g296048/_0_ , \g296049/_3_ , \g296522/_3_ , \g296523/_3_ , \g296524/_0_ , \g296525/_0_ , \g296526/_0_ , \g296527/_0_ , \g296528/_3_ , \g296529/_0_ , \g296530/_0_ , \g296531/_0_ , \g297026/_0_ , \g297027/_0_ , \g305620/_3_ , \g305621/_3_ , \g305622/_3_ , \g305623/_3_ , \g305624/_3_ , \g305625/_3_ , \g305626/_3_ , \g305627/_3_ , \g305628/_3_ , \g305629/_3_ , \g305630/_3_ , \g305631/_3_ , \g305632/_3_ , \g305633/_3_ , \g305634/_3_ , \g305635/_3_ , \g305636/_3_ , \g305637/_3_ , \g305638/_3_ , \g305639/_3_ , \g305640/_3_ , \g305641/_3_ , \g305642/_3_ , \g305643/_3_ , \g305644/_3_ , \g305645/_3_ , \g305646/_3_ , \g305647/_3_ , \g305648/_3_ , \g305649/_3_ , \g305650/_3_ , \g305651/_3_ , \g305652/_3_ , \g305653/_3_ , \g305654/_3_ , \g305655/_3_ , \g305656/_3_ , \g305657/_3_ , \g305658/_3_ , \g305659/_3_ , \g305660/_3_ , \g305661/_3_ , \g305662/_3_ , \g305663/_3_ , \g305664/_3_ , \g305665/_3_ , \g305666/_3_ , \g305667/_3_ , \g305668/_3_ , \g305669/_3_ , \g305670/_3_ , \g305671/_3_ , \g305672/_3_ , \g305673/_3_ , \g305674/_3_ , \g305675/_3_ , \g305676/_3_ , \g305677/_3_ , \g305678/_3_ , \g305679/_3_ , \g305680/_3_ , \g305681/_3_ , \g305682/_3_ , \g305683/_3_ , \g305684/_3_ , \g305685/_3_ , \g305686/_3_ , \g305687/_3_ , \g305688/_3_ , \g305689/_3_ , \g305690/_3_ , \g305691/_3_ , \g305692/_3_ , \g305693/_3_ , \g305694/_3_ , \g305695/_3_ , \g305696/_3_ , \g305697/_3_ , \g305698/_3_ , \g305699/_3_ , \g305700/_3_ , \g305701/_3_ , \g305702/_3_ , \g305703/_3_ , \g305704/_3_ , \g305705/_3_ , \g305706/_3_ , \g305707/_3_ , \g305708/_3_ , \g305709/_3_ , \g305710/_3_ , \g305711/_3_ , \g305712/_3_ , \g305713/_3_ , \g305714/_3_ , \g305715/_3_ , \g305716/_3_ , \g305717/_3_ , \g305718/_3_ , \g305719/_3_ , \g305720/_3_ , \g305721/_3_ , \g305722/_3_ , \g305723/_3_ , \g305724/_3_ , \g305725/_3_ , \g305726/_3_ , \g305727/_3_ , \g305728/_3_ , \g305729/_3_ , \g305730/_3_ , \g305731/_3_ , \g321371/_0_ , \g321424/_0_ , \g321474/_3_ , \g321637/_3_ , \g321688/_0_ , \g321712/_0_ , \g321772/_3_ , \g321832/_0_ , \g321999/_0_ , \g322013/_3_ , \g322109/_0_ , \g322184/_0_ , \g322250/_0_ , \g322274/_0_ , \g322293/_3_ , \g322437/_0_ , \g322537/_3_ , \g322584/_0_ , \g322830/_0_ , \g322871/_0_ , \g322882/_0_ , \g322933/_0_ , \g323004/_0_ , \g323104/_0_ , \g323125/_0_ , \g323138/_3_ , \g323273/_0_ , \u0_desOut_reg[0]/_05_ , \u0_desOut_reg[12]/_05_ , \u0_desOut_reg[14]/_05_ , \u0_desOut_reg[18]/_05_ , \u0_desOut_reg[20]/_05_ , \u0_desOut_reg[24]/_05_ , \u0_desOut_reg[26]/_05_ , \u0_desOut_reg[28]/_05_ , \u0_desOut_reg[2]/_05_ , \u0_desOut_reg[30]/_05_ , \u0_desOut_reg[32]/_05_ , \u0_desOut_reg[34]/_05_ , \u0_desOut_reg[36]/_05_ , \u0_desOut_reg[42]/_05_ , \u0_desOut_reg[44]/_05_ , \u0_desOut_reg[46]/_05_ , \u0_desOut_reg[48]/_05_ , \u0_desOut_reg[54]/_05_ , \u0_desOut_reg[56]/_05_ , \u0_desOut_reg[62]/_05_ , \u0_desOut_reg[6]/_05_ , \u0_desOut_reg[8]/_05_ , \u1_desOut_reg[0]/_05_ , \u1_desOut_reg[12]/_05_ , \u1_desOut_reg[14]/_05_ , \u1_desOut_reg[16]/_05_ , \u1_desOut_reg[18]/_05_ , \u1_desOut_reg[20]/_05_ , \u1_desOut_reg[22]/_05_ , \u1_desOut_reg[24]/_05_ , \u1_desOut_reg[26]/_05_ , \u1_desOut_reg[28]/_05_ , \u1_desOut_reg[2]/_05_ , \u1_desOut_reg[30]/_05_ , \u1_desOut_reg[32]/_05_ , \u1_desOut_reg[34]/_05_ , \u1_desOut_reg[36]/_05_ , \u1_desOut_reg[38]/_05_ , \u1_desOut_reg[42]/_05_ , \u1_desOut_reg[44]/_05_ , \u1_desOut_reg[46]/_05_ , \u1_desOut_reg[48]/_05_ , \u1_desOut_reg[4]/_05_ , \u1_desOut_reg[54]/_05_ , \u1_desOut_reg[56]/_05_ , \u1_desOut_reg[58]/_05_ , \u1_desOut_reg[60]/_05_ , \u1_desOut_reg[62]/_05_ , \u1_desOut_reg[6]/_05_ , \u1_desOut_reg[8]/_05_ , \u2_desOut_reg[0]/_05_ , \u2_desOut_reg[10]/_05_ , \u2_desOut_reg[12]/_05_ , \u2_desOut_reg[14]/_05_ , \u2_desOut_reg[16]/_05_ , \u2_desOut_reg[18]/_05_ , \u2_desOut_reg[20]/_05_ , \u2_desOut_reg[22]/_05_ , \u2_desOut_reg[24]/_05_ , \u2_desOut_reg[26]/_05_ , \u2_desOut_reg[28]/_05_ , \u2_desOut_reg[2]/_05_ , \u2_desOut_reg[30]/_05_ , \u2_desOut_reg[32]/_05_ , \u2_desOut_reg[34]/_05_ , \u2_desOut_reg[36]/_05_ , \u2_desOut_reg[38]/_05_ , \u2_desOut_reg[40]/_05_ , \u2_desOut_reg[42]/_05_ , \u2_desOut_reg[44]/_05_ , \u2_desOut_reg[46]/_05_ , \u2_desOut_reg[48]/_05_ , \u2_desOut_reg[4]/_05_ , \u2_desOut_reg[50]/_05_ , \u2_desOut_reg[52]/_05_ , \u2_desOut_reg[54]/_05_ , \u2_desOut_reg[56]/_05_ , \u2_desOut_reg[58]/_05_ , \u2_desOut_reg[60]/_05_ , \u2_desOut_reg[62]/_05_ , \u2_desOut_reg[6]/_05_ , \u2_desOut_reg[8]/_05_ );
	input decrypt_pad ;
	input \key1[0]_pad  ;
	input \key1[10]_pad  ;
	input \key1[11]_pad  ;
	input \key1[12]_pad  ;
	input \key1[13]_pad  ;
	input \key1[14]_pad  ;
	input \key1[15]_pad  ;
	input \key1[16]_pad  ;
	input \key1[17]_pad  ;
	input \key1[18]_pad  ;
	input \key1[19]_pad  ;
	input \key1[1]_pad  ;
	input \key1[20]_pad  ;
	input \key1[21]_pad  ;
	input \key1[22]_pad  ;
	input \key1[23]_pad  ;
	input \key1[24]_pad  ;
	input \key1[25]_pad  ;
	input \key1[26]_pad  ;
	input \key1[27]_pad  ;
	input \key1[28]_pad  ;
	input \key1[29]_pad  ;
	input \key1[2]_pad  ;
	input \key1[30]_pad  ;
	input \key1[31]_pad  ;
	input \key1[32]_pad  ;
	input \key1[33]_pad  ;
	input \key1[34]_pad  ;
	input \key1[35]_pad  ;
	input \key1[36]_pad  ;
	input \key1[37]_pad  ;
	input \key1[38]_pad  ;
	input \key1[39]_pad  ;
	input \key1[3]_pad  ;
	input \key1[40]_pad  ;
	input \key1[41]_pad  ;
	input \key1[42]_pad  ;
	input \key1[43]_pad  ;
	input \key1[44]_pad  ;
	input \key1[45]_pad  ;
	input \key1[46]_pad  ;
	input \key1[47]_pad  ;
	input \key1[48]_pad  ;
	input \key1[49]_pad  ;
	input \key1[4]_pad  ;
	input \key1[50]_pad  ;
	input \key1[51]_pad  ;
	input \key1[52]_pad  ;
	input \key1[53]_pad  ;
	input \key1[54]_pad  ;
	input \key1[55]_pad  ;
	input \key1[5]_pad  ;
	input \key1[6]_pad  ;
	input \key1[7]_pad  ;
	input \key1[8]_pad  ;
	input \key1[9]_pad  ;
	input \key3[0]_pad  ;
	input \key3[10]_pad  ;
	input \key3[11]_pad  ;
	input \key3[12]_pad  ;
	input \key3[13]_pad  ;
	input \key3[14]_pad  ;
	input \key3[15]_pad  ;
	input \key3[16]_pad  ;
	input \key3[17]_pad  ;
	input \key3[18]_pad  ;
	input \key3[19]_pad  ;
	input \key3[1]_pad  ;
	input \key3[20]_pad  ;
	input \key3[21]_pad  ;
	input \key3[22]_pad  ;
	input \key3[23]_pad  ;
	input \key3[24]_pad  ;
	input \key3[25]_pad  ;
	input \key3[26]_pad  ;
	input \key3[27]_pad  ;
	input \key3[28]_pad  ;
	input \key3[29]_pad  ;
	input \key3[2]_pad  ;
	input \key3[30]_pad  ;
	input \key3[31]_pad  ;
	input \key3[32]_pad  ;
	input \key3[33]_pad  ;
	input \key3[34]_pad  ;
	input \key3[35]_pad  ;
	input \key3[36]_pad  ;
	input \key3[37]_pad  ;
	input \key3[38]_pad  ;
	input \key3[39]_pad  ;
	input \key3[3]_pad  ;
	input \key3[40]_pad  ;
	input \key3[41]_pad  ;
	input \key3[42]_pad  ;
	input \key3[43]_pad  ;
	input \key3[44]_pad  ;
	input \key3[45]_pad  ;
	input \key3[46]_pad  ;
	input \key3[47]_pad  ;
	input \key3[48]_pad  ;
	input \key3[49]_pad  ;
	input \key3[4]_pad  ;
	input \key3[50]_pad  ;
	input \key3[51]_pad  ;
	input \key3[52]_pad  ;
	input \key3[53]_pad  ;
	input \key3[54]_pad  ;
	input \key3[55]_pad  ;
	input \key3[5]_pad  ;
	input \key3[6]_pad  ;
	input \key3[7]_pad  ;
	input \key3[8]_pad  ;
	input \key3[9]_pad  ;
	input \u0_L0_reg[10]/NET0131  ;
	input \u0_L0_reg[11]/NET0131  ;
	input \u0_L0_reg[12]/NET0131  ;
	input \u0_L0_reg[13]/NET0131  ;
	input \u0_L0_reg[14]/NET0131  ;
	input \u0_L0_reg[15]/P0001  ;
	input \u0_L0_reg[16]/NET0131  ;
	input \u0_L0_reg[17]/NET0131  ;
	input \u0_L0_reg[18]/NET0131  ;
	input \u0_L0_reg[19]/P0001  ;
	input \u0_L0_reg[1]/NET0131  ;
	input \u0_L0_reg[20]/NET0131  ;
	input \u0_L0_reg[21]/NET0131  ;
	input \u0_L0_reg[22]/NET0131  ;
	input \u0_L0_reg[23]/NET0131  ;
	input \u0_L0_reg[24]/NET0131  ;
	input \u0_L0_reg[25]/NET0131  ;
	input \u0_L0_reg[26]/NET0131  ;
	input \u0_L0_reg[27]/NET0131  ;
	input \u0_L0_reg[28]/NET0131  ;
	input \u0_L0_reg[29]/NET0131  ;
	input \u0_L0_reg[2]/NET0131  ;
	input \u0_L0_reg[30]/P0001  ;
	input \u0_L0_reg[31]/NET0131  ;
	input \u0_L0_reg[32]/NET0131  ;
	input \u0_L0_reg[3]/NET0131  ;
	input \u0_L0_reg[4]/NET0131  ;
	input \u0_L0_reg[5]/NET0131  ;
	input \u0_L0_reg[6]/NET0131  ;
	input \u0_L0_reg[7]/NET0131  ;
	input \u0_L0_reg[8]/NET0131  ;
	input \u0_L0_reg[9]/NET0131  ;
	input \u0_L10_reg[10]/NET0131  ;
	input \u0_L10_reg[11]/NET0131  ;
	input \u0_L10_reg[12]/NET0131  ;
	input \u0_L10_reg[13]/NET0131  ;
	input \u0_L10_reg[14]/NET0131  ;
	input \u0_L10_reg[15]/P0001  ;
	input \u0_L10_reg[16]/NET0131  ;
	input \u0_L10_reg[17]/NET0131  ;
	input \u0_L10_reg[18]/NET0131  ;
	input \u0_L10_reg[19]/NET0131  ;
	input \u0_L10_reg[1]/NET0131  ;
	input \u0_L10_reg[20]/NET0131  ;
	input \u0_L10_reg[21]/NET0131  ;
	input \u0_L10_reg[22]/NET0131  ;
	input \u0_L10_reg[23]/NET0131  ;
	input \u0_L10_reg[24]/NET0131  ;
	input \u0_L10_reg[25]/NET0131  ;
	input \u0_L10_reg[26]/NET0131  ;
	input \u0_L10_reg[27]/NET0131  ;
	input \u0_L10_reg[28]/NET0131  ;
	input \u0_L10_reg[29]/NET0131  ;
	input \u0_L10_reg[2]/NET0131  ;
	input \u0_L10_reg[30]/NET0131  ;
	input \u0_L10_reg[31]/NET0131  ;
	input \u0_L10_reg[32]/NET0131  ;
	input \u0_L10_reg[3]/NET0131  ;
	input \u0_L10_reg[4]/NET0131  ;
	input \u0_L10_reg[5]/NET0131  ;
	input \u0_L10_reg[6]/NET0131  ;
	input \u0_L10_reg[7]/NET0131  ;
	input \u0_L10_reg[8]/NET0131  ;
	input \u0_L10_reg[9]/NET0131  ;
	input \u0_L11_reg[10]/NET0131  ;
	input \u0_L11_reg[11]/P0001  ;
	input \u0_L11_reg[12]/NET0131  ;
	input \u0_L11_reg[13]/NET0131  ;
	input \u0_L11_reg[14]/NET0131  ;
	input \u0_L11_reg[15]/P0001  ;
	input \u0_L11_reg[16]/NET0131  ;
	input \u0_L11_reg[17]/NET0131  ;
	input \u0_L11_reg[18]/NET0131  ;
	input \u0_L11_reg[19]/NET0131  ;
	input \u0_L11_reg[1]/NET0131  ;
	input \u0_L11_reg[20]/NET0131  ;
	input \u0_L11_reg[21]/NET0131  ;
	input \u0_L11_reg[22]/NET0131  ;
	input \u0_L11_reg[23]/NET0131  ;
	input \u0_L11_reg[24]/NET0131  ;
	input \u0_L11_reg[25]/NET0131  ;
	input \u0_L11_reg[26]/NET0131  ;
	input \u0_L11_reg[27]/NET0131  ;
	input \u0_L11_reg[28]/NET0131  ;
	input \u0_L11_reg[29]/NET0131  ;
	input \u0_L11_reg[2]/NET0131  ;
	input \u0_L11_reg[30]/NET0131  ;
	input \u0_L11_reg[31]/NET0131  ;
	input \u0_L11_reg[32]/NET0131  ;
	input \u0_L11_reg[3]/NET0131  ;
	input \u0_L11_reg[4]/NET0131  ;
	input \u0_L11_reg[5]/NET0131  ;
	input \u0_L11_reg[6]/NET0131  ;
	input \u0_L11_reg[7]/NET0131  ;
	input \u0_L11_reg[8]/NET0131  ;
	input \u0_L11_reg[9]/NET0131  ;
	input \u0_L12_reg[10]/NET0131  ;
	input \u0_L12_reg[11]/NET0131  ;
	input \u0_L12_reg[12]/NET0131  ;
	input \u0_L12_reg[13]/NET0131  ;
	input \u0_L12_reg[14]/NET0131  ;
	input \u0_L12_reg[15]/P0001  ;
	input \u0_L12_reg[16]/NET0131  ;
	input \u0_L12_reg[17]/NET0131  ;
	input \u0_L12_reg[18]/NET0131  ;
	input \u0_L12_reg[19]/P0001  ;
	input \u0_L12_reg[1]/NET0131  ;
	input \u0_L12_reg[20]/NET0131  ;
	input \u0_L12_reg[21]/NET0131  ;
	input \u0_L12_reg[22]/NET0131  ;
	input \u0_L12_reg[23]/NET0131  ;
	input \u0_L12_reg[24]/NET0131  ;
	input \u0_L12_reg[25]/NET0131  ;
	input \u0_L12_reg[26]/NET0131  ;
	input \u0_L12_reg[27]/NET0131  ;
	input \u0_L12_reg[28]/NET0131  ;
	input \u0_L12_reg[29]/NET0131  ;
	input \u0_L12_reg[2]/NET0131  ;
	input \u0_L12_reg[30]/NET0131  ;
	input \u0_L12_reg[31]/NET0131  ;
	input \u0_L12_reg[32]/NET0131  ;
	input \u0_L12_reg[3]/NET0131  ;
	input \u0_L12_reg[4]/NET0131  ;
	input \u0_L12_reg[5]/NET0131  ;
	input \u0_L12_reg[6]/NET0131  ;
	input \u0_L12_reg[7]/NET0131  ;
	input \u0_L12_reg[8]/NET0131  ;
	input \u0_L12_reg[9]/NET0131  ;
	input \u0_L13_reg[10]/NET0131  ;
	input \u0_L13_reg[11]/NET0131  ;
	input \u0_L13_reg[12]/NET0131  ;
	input \u0_L13_reg[13]/NET0131  ;
	input \u0_L13_reg[14]/NET0131  ;
	input \u0_L13_reg[15]/P0001  ;
	input \u0_L13_reg[16]/NET0131  ;
	input \u0_L13_reg[17]/NET0131  ;
	input \u0_L13_reg[18]/NET0131  ;
	input \u0_L13_reg[19]/NET0131  ;
	input \u0_L13_reg[1]/NET0131  ;
	input \u0_L13_reg[20]/NET0131  ;
	input \u0_L13_reg[21]/NET0131  ;
	input \u0_L13_reg[22]/NET0131  ;
	input \u0_L13_reg[23]/NET0131  ;
	input \u0_L13_reg[24]/NET0131  ;
	input \u0_L13_reg[25]/NET0131  ;
	input \u0_L13_reg[26]/NET0131  ;
	input \u0_L13_reg[27]/NET0131  ;
	input \u0_L13_reg[28]/NET0131  ;
	input \u0_L13_reg[29]/NET0131  ;
	input \u0_L13_reg[2]/NET0131  ;
	input \u0_L13_reg[30]/NET0131  ;
	input \u0_L13_reg[31]/NET0131  ;
	input \u0_L13_reg[32]/NET0131  ;
	input \u0_L13_reg[3]/NET0131  ;
	input \u0_L13_reg[4]/NET0131  ;
	input \u0_L13_reg[5]/NET0131  ;
	input \u0_L13_reg[6]/NET0131  ;
	input \u0_L13_reg[7]/NET0131  ;
	input \u0_L13_reg[8]/NET0131  ;
	input \u0_L13_reg[9]/NET0131  ;
	input \u0_L14_reg[10]/P0001  ;
	input \u0_L14_reg[11]/P0001  ;
	input \u0_L14_reg[12]/P0001  ;
	input \u0_L14_reg[13]/P0001  ;
	input \u0_L14_reg[14]/P0001  ;
	input \u0_L14_reg[15]/P0001  ;
	input \u0_L14_reg[16]/P0001  ;
	input \u0_L14_reg[17]/P0001  ;
	input \u0_L14_reg[18]/P0001  ;
	input \u0_L14_reg[19]/P0001  ;
	input \u0_L14_reg[1]/P0001  ;
	input \u0_L14_reg[20]/P0001  ;
	input \u0_L14_reg[21]/P0001  ;
	input \u0_L14_reg[22]/P0001  ;
	input \u0_L14_reg[23]/P0001  ;
	input \u0_L14_reg[24]/P0001  ;
	input \u0_L14_reg[25]/P0001  ;
	input \u0_L14_reg[26]/P0001  ;
	input \u0_L14_reg[27]/P0001  ;
	input \u0_L14_reg[28]/P0001  ;
	input \u0_L14_reg[29]/P0001  ;
	input \u0_L14_reg[2]/P0001  ;
	input \u0_L14_reg[30]/P0001  ;
	input \u0_L14_reg[31]/P0001  ;
	input \u0_L14_reg[32]/P0001  ;
	input \u0_L14_reg[3]/P0001  ;
	input \u0_L14_reg[4]/P0001  ;
	input \u0_L14_reg[5]/P0001  ;
	input \u0_L14_reg[6]/P0001  ;
	input \u0_L14_reg[7]/P0001  ;
	input \u0_L14_reg[8]/P0001  ;
	input \u0_L14_reg[9]/P0001  ;
	input \u0_L1_reg[10]/NET0131  ;
	input \u0_L1_reg[11]/NET0131  ;
	input \u0_L1_reg[12]/NET0131  ;
	input \u0_L1_reg[13]/NET0131  ;
	input \u0_L1_reg[14]/NET0131  ;
	input \u0_L1_reg[15]/P0001  ;
	input \u0_L1_reg[16]/NET0131  ;
	input \u0_L1_reg[17]/NET0131  ;
	input \u0_L1_reg[18]/NET0131  ;
	input \u0_L1_reg[19]/NET0131  ;
	input \u0_L1_reg[1]/NET0131  ;
	input \u0_L1_reg[20]/NET0131  ;
	input \u0_L1_reg[21]/NET0131  ;
	input \u0_L1_reg[22]/NET0131  ;
	input \u0_L1_reg[23]/NET0131  ;
	input \u0_L1_reg[24]/NET0131  ;
	input \u0_L1_reg[25]/NET0131  ;
	input \u0_L1_reg[26]/NET0131  ;
	input \u0_L1_reg[27]/NET0131  ;
	input \u0_L1_reg[28]/NET0131  ;
	input \u0_L1_reg[29]/NET0131  ;
	input \u0_L1_reg[2]/NET0131  ;
	input \u0_L1_reg[30]/NET0131  ;
	input \u0_L1_reg[31]/NET0131  ;
	input \u0_L1_reg[32]/NET0131  ;
	input \u0_L1_reg[3]/NET0131  ;
	input \u0_L1_reg[4]/NET0131  ;
	input \u0_L1_reg[5]/NET0131  ;
	input \u0_L1_reg[6]/NET0131  ;
	input \u0_L1_reg[7]/NET0131  ;
	input \u0_L1_reg[8]/NET0131  ;
	input \u0_L1_reg[9]/NET0131  ;
	input \u0_L2_reg[10]/NET0131  ;
	input \u0_L2_reg[11]/NET0131  ;
	input \u0_L2_reg[12]/NET0131  ;
	input \u0_L2_reg[13]/NET0131  ;
	input \u0_L2_reg[14]/NET0131  ;
	input \u0_L2_reg[15]/P0001  ;
	input \u0_L2_reg[16]/NET0131  ;
	input \u0_L2_reg[17]/NET0131  ;
	input \u0_L2_reg[18]/NET0131  ;
	input \u0_L2_reg[19]/P0001  ;
	input \u0_L2_reg[1]/NET0131  ;
	input \u0_L2_reg[20]/NET0131  ;
	input \u0_L2_reg[21]/NET0131  ;
	input \u0_L2_reg[22]/NET0131  ;
	input \u0_L2_reg[23]/NET0131  ;
	input \u0_L2_reg[24]/NET0131  ;
	input \u0_L2_reg[25]/NET0131  ;
	input \u0_L2_reg[26]/NET0131  ;
	input \u0_L2_reg[27]/NET0131  ;
	input \u0_L2_reg[28]/NET0131  ;
	input \u0_L2_reg[29]/NET0131  ;
	input \u0_L2_reg[2]/NET0131  ;
	input \u0_L2_reg[30]/NET0131  ;
	input \u0_L2_reg[31]/NET0131  ;
	input \u0_L2_reg[32]/NET0131  ;
	input \u0_L2_reg[3]/NET0131  ;
	input \u0_L2_reg[4]/NET0131  ;
	input \u0_L2_reg[5]/NET0131  ;
	input \u0_L2_reg[6]/NET0131  ;
	input \u0_L2_reg[7]/NET0131  ;
	input \u0_L2_reg[8]/NET0131  ;
	input \u0_L2_reg[9]/NET0131  ;
	input \u0_L3_reg[10]/NET0131  ;
	input \u0_L3_reg[11]/NET0131  ;
	input \u0_L3_reg[12]/NET0131  ;
	input \u0_L3_reg[13]/NET0131  ;
	input \u0_L3_reg[14]/NET0131  ;
	input \u0_L3_reg[15]/P0001  ;
	input \u0_L3_reg[16]/NET0131  ;
	input \u0_L3_reg[17]/NET0131  ;
	input \u0_L3_reg[18]/NET0131  ;
	input \u0_L3_reg[19]/P0001  ;
	input \u0_L3_reg[1]/NET0131  ;
	input \u0_L3_reg[20]/NET0131  ;
	input \u0_L3_reg[21]/NET0131  ;
	input \u0_L3_reg[22]/NET0131  ;
	input \u0_L3_reg[23]/NET0131  ;
	input \u0_L3_reg[24]/NET0131  ;
	input \u0_L3_reg[25]/NET0131  ;
	input \u0_L3_reg[26]/NET0131  ;
	input \u0_L3_reg[27]/NET0131  ;
	input \u0_L3_reg[28]/NET0131  ;
	input \u0_L3_reg[29]/NET0131  ;
	input \u0_L3_reg[2]/NET0131  ;
	input \u0_L3_reg[30]/NET0131  ;
	input \u0_L3_reg[31]/NET0131  ;
	input \u0_L3_reg[32]/NET0131  ;
	input \u0_L3_reg[3]/NET0131  ;
	input \u0_L3_reg[4]/NET0131  ;
	input \u0_L3_reg[5]/NET0131  ;
	input \u0_L3_reg[6]/NET0131  ;
	input \u0_L3_reg[7]/NET0131  ;
	input \u0_L3_reg[8]/NET0131  ;
	input \u0_L3_reg[9]/NET0131  ;
	input \u0_L4_reg[10]/NET0131  ;
	input \u0_L4_reg[11]/NET0131  ;
	input \u0_L4_reg[12]/NET0131  ;
	input \u0_L4_reg[13]/NET0131  ;
	input \u0_L4_reg[14]/NET0131  ;
	input \u0_L4_reg[15]/P0001  ;
	input \u0_L4_reg[16]/NET0131  ;
	input \u0_L4_reg[17]/NET0131  ;
	input \u0_L4_reg[18]/NET0131  ;
	input \u0_L4_reg[19]/NET0131  ;
	input \u0_L4_reg[1]/NET0131  ;
	input \u0_L4_reg[20]/NET0131  ;
	input \u0_L4_reg[21]/NET0131  ;
	input \u0_L4_reg[22]/NET0131  ;
	input \u0_L4_reg[23]/NET0131  ;
	input \u0_L4_reg[24]/NET0131  ;
	input \u0_L4_reg[25]/NET0131  ;
	input \u0_L4_reg[26]/NET0131  ;
	input \u0_L4_reg[27]/NET0131  ;
	input \u0_L4_reg[28]/NET0131  ;
	input \u0_L4_reg[29]/NET0131  ;
	input \u0_L4_reg[2]/NET0131  ;
	input \u0_L4_reg[30]/NET0131  ;
	input \u0_L4_reg[31]/NET0131  ;
	input \u0_L4_reg[32]/NET0131  ;
	input \u0_L4_reg[3]/NET0131  ;
	input \u0_L4_reg[4]/NET0131  ;
	input \u0_L4_reg[5]/NET0131  ;
	input \u0_L4_reg[6]/NET0131  ;
	input \u0_L4_reg[7]/NET0131  ;
	input \u0_L4_reg[8]/NET0131  ;
	input \u0_L4_reg[9]/NET0131  ;
	input \u0_L5_reg[10]/NET0131  ;
	input \u0_L5_reg[11]/NET0131  ;
	input \u0_L5_reg[12]/NET0131  ;
	input \u0_L5_reg[13]/NET0131  ;
	input \u0_L5_reg[14]/NET0131  ;
	input \u0_L5_reg[15]/P0001  ;
	input \u0_L5_reg[16]/NET0131  ;
	input \u0_L5_reg[17]/NET0131  ;
	input \u0_L5_reg[18]/NET0131  ;
	input \u0_L5_reg[19]/P0001  ;
	input \u0_L5_reg[1]/NET0131  ;
	input \u0_L5_reg[20]/NET0131  ;
	input \u0_L5_reg[21]/NET0131  ;
	input \u0_L5_reg[22]/NET0131  ;
	input \u0_L5_reg[23]/NET0131  ;
	input \u0_L5_reg[24]/NET0131  ;
	input \u0_L5_reg[25]/NET0131  ;
	input \u0_L5_reg[26]/NET0131  ;
	input \u0_L5_reg[27]/NET0131  ;
	input \u0_L5_reg[28]/NET0131  ;
	input \u0_L5_reg[29]/NET0131  ;
	input \u0_L5_reg[2]/NET0131  ;
	input \u0_L5_reg[30]/NET0131  ;
	input \u0_L5_reg[31]/NET0131  ;
	input \u0_L5_reg[32]/NET0131  ;
	input \u0_L5_reg[3]/NET0131  ;
	input \u0_L5_reg[4]/NET0131  ;
	input \u0_L5_reg[5]/NET0131  ;
	input \u0_L5_reg[6]/NET0131  ;
	input \u0_L5_reg[7]/NET0131  ;
	input \u0_L5_reg[8]/NET0131  ;
	input \u0_L5_reg[9]/NET0131  ;
	input \u0_L6_reg[10]/NET0131  ;
	input \u0_L6_reg[11]/NET0131  ;
	input \u0_L6_reg[12]/NET0131  ;
	input \u0_L6_reg[13]/NET0131  ;
	input \u0_L6_reg[14]/NET0131  ;
	input \u0_L6_reg[15]/P0001  ;
	input \u0_L6_reg[16]/NET0131  ;
	input \u0_L6_reg[17]/NET0131  ;
	input \u0_L6_reg[18]/NET0131  ;
	input \u0_L6_reg[19]/P0001  ;
	input \u0_L6_reg[1]/NET0131  ;
	input \u0_L6_reg[20]/NET0131  ;
	input \u0_L6_reg[21]/NET0131  ;
	input \u0_L6_reg[22]/NET0131  ;
	input \u0_L6_reg[23]/NET0131  ;
	input \u0_L6_reg[24]/NET0131  ;
	input \u0_L6_reg[25]/NET0131  ;
	input \u0_L6_reg[26]/NET0131  ;
	input \u0_L6_reg[27]/NET0131  ;
	input \u0_L6_reg[28]/NET0131  ;
	input \u0_L6_reg[29]/NET0131  ;
	input \u0_L6_reg[2]/NET0131  ;
	input \u0_L6_reg[30]/NET0131  ;
	input \u0_L6_reg[31]/NET0131  ;
	input \u0_L6_reg[32]/NET0131  ;
	input \u0_L6_reg[3]/NET0131  ;
	input \u0_L6_reg[4]/NET0131  ;
	input \u0_L6_reg[5]/NET0131  ;
	input \u0_L6_reg[6]/NET0131  ;
	input \u0_L6_reg[7]/NET0131  ;
	input \u0_L6_reg[8]/NET0131  ;
	input \u0_L6_reg[9]/NET0131  ;
	input \u0_L7_reg[10]/NET0131  ;
	input \u0_L7_reg[11]/NET0131  ;
	input \u0_L7_reg[12]/NET0131  ;
	input \u0_L7_reg[13]/NET0131  ;
	input \u0_L7_reg[14]/NET0131  ;
	input \u0_L7_reg[15]/P0001  ;
	input \u0_L7_reg[16]/NET0131  ;
	input \u0_L7_reg[17]/NET0131  ;
	input \u0_L7_reg[18]/NET0131  ;
	input \u0_L7_reg[19]/NET0131  ;
	input \u0_L7_reg[1]/NET0131  ;
	input \u0_L7_reg[20]/NET0131  ;
	input \u0_L7_reg[21]/NET0131  ;
	input \u0_L7_reg[22]/NET0131  ;
	input \u0_L7_reg[23]/NET0131  ;
	input \u0_L7_reg[24]/NET0131  ;
	input \u0_L7_reg[25]/NET0131  ;
	input \u0_L7_reg[26]/NET0131  ;
	input \u0_L7_reg[27]/NET0131  ;
	input \u0_L7_reg[28]/NET0131  ;
	input \u0_L7_reg[29]/NET0131  ;
	input \u0_L7_reg[2]/NET0131  ;
	input \u0_L7_reg[30]/NET0131  ;
	input \u0_L7_reg[31]/NET0131  ;
	input \u0_L7_reg[32]/NET0131  ;
	input \u0_L7_reg[3]/NET0131  ;
	input \u0_L7_reg[4]/NET0131  ;
	input \u0_L7_reg[5]/NET0131  ;
	input \u0_L7_reg[6]/NET0131  ;
	input \u0_L7_reg[7]/NET0131  ;
	input \u0_L7_reg[8]/NET0131  ;
	input \u0_L7_reg[9]/NET0131  ;
	input \u0_L8_reg[10]/NET0131  ;
	input \u0_L8_reg[11]/NET0131  ;
	input \u0_L8_reg[12]/NET0131  ;
	input \u0_L8_reg[13]/NET0131  ;
	input \u0_L8_reg[14]/NET0131  ;
	input \u0_L8_reg[15]/P0001  ;
	input \u0_L8_reg[16]/NET0131  ;
	input \u0_L8_reg[17]/NET0131  ;
	input \u0_L8_reg[18]/NET0131  ;
	input \u0_L8_reg[19]/NET0131  ;
	input \u0_L8_reg[1]/NET0131  ;
	input \u0_L8_reg[20]/NET0131  ;
	input \u0_L8_reg[21]/NET0131  ;
	input \u0_L8_reg[22]/NET0131  ;
	input \u0_L8_reg[23]/NET0131  ;
	input \u0_L8_reg[24]/NET0131  ;
	input \u0_L8_reg[25]/NET0131  ;
	input \u0_L8_reg[26]/NET0131  ;
	input \u0_L8_reg[27]/NET0131  ;
	input \u0_L8_reg[28]/NET0131  ;
	input \u0_L8_reg[29]/NET0131  ;
	input \u0_L8_reg[2]/NET0131  ;
	input \u0_L8_reg[30]/NET0131  ;
	input \u0_L8_reg[31]/NET0131  ;
	input \u0_L8_reg[32]/NET0131  ;
	input \u0_L8_reg[3]/NET0131  ;
	input \u0_L8_reg[4]/NET0131  ;
	input \u0_L8_reg[5]/NET0131  ;
	input \u0_L8_reg[6]/NET0131  ;
	input \u0_L8_reg[7]/NET0131  ;
	input \u0_L8_reg[8]/NET0131  ;
	input \u0_L8_reg[9]/NET0131  ;
	input \u0_L9_reg[10]/NET0131  ;
	input \u0_L9_reg[11]/NET0131  ;
	input \u0_L9_reg[12]/NET0131  ;
	input \u0_L9_reg[13]/NET0131  ;
	input \u0_L9_reg[14]/NET0131  ;
	input \u0_L9_reg[15]/P0001  ;
	input \u0_L9_reg[16]/NET0131  ;
	input \u0_L9_reg[17]/NET0131  ;
	input \u0_L9_reg[18]/NET0131  ;
	input \u0_L9_reg[19]/P0001  ;
	input \u0_L9_reg[1]/NET0131  ;
	input \u0_L9_reg[20]/NET0131  ;
	input \u0_L9_reg[21]/NET0131  ;
	input \u0_L9_reg[22]/NET0131  ;
	input \u0_L9_reg[23]/NET0131  ;
	input \u0_L9_reg[24]/NET0131  ;
	input \u0_L9_reg[25]/NET0131  ;
	input \u0_L9_reg[26]/NET0131  ;
	input \u0_L9_reg[27]/NET0131  ;
	input \u0_L9_reg[28]/NET0131  ;
	input \u0_L9_reg[29]/NET0131  ;
	input \u0_L9_reg[2]/NET0131  ;
	input \u0_L9_reg[30]/NET0131  ;
	input \u0_L9_reg[31]/NET0131  ;
	input \u0_L9_reg[32]/NET0131  ;
	input \u0_L9_reg[3]/NET0131  ;
	input \u0_L9_reg[4]/NET0131  ;
	input \u0_L9_reg[5]/NET0131  ;
	input \u0_L9_reg[6]/NET0131  ;
	input \u0_L9_reg[7]/NET0131  ;
	input \u0_L9_reg[8]/NET0131  ;
	input \u0_L9_reg[9]/NET0131  ;
	input \u0_R0_reg[10]/NET0131  ;
	input \u0_R0_reg[11]/NET0131  ;
	input \u0_R0_reg[12]/NET0131  ;
	input \u0_R0_reg[13]/NET0131  ;
	input \u0_R0_reg[14]/NET0131  ;
	input \u0_R0_reg[15]/NET0131  ;
	input \u0_R0_reg[16]/NET0131  ;
	input \u0_R0_reg[17]/NET0131  ;
	input \u0_R0_reg[18]/NET0131  ;
	input \u0_R0_reg[19]/NET0131  ;
	input \u0_R0_reg[1]/NET0131  ;
	input \u0_R0_reg[20]/NET0131  ;
	input \u0_R0_reg[21]/NET0131  ;
	input \u0_R0_reg[22]/NET0131  ;
	input \u0_R0_reg[23]/NET0131  ;
	input \u0_R0_reg[24]/NET0131  ;
	input \u0_R0_reg[25]/NET0131  ;
	input \u0_R0_reg[26]/NET0131  ;
	input \u0_R0_reg[27]/NET0131  ;
	input \u0_R0_reg[28]/NET0131  ;
	input \u0_R0_reg[29]/NET0131  ;
	input \u0_R0_reg[2]/NET0131  ;
	input \u0_R0_reg[30]/NET0131  ;
	input \u0_R0_reg[31]/NET0131  ;
	input \u0_R0_reg[32]/NET0131  ;
	input \u0_R0_reg[3]/NET0131  ;
	input \u0_R0_reg[4]/NET0131  ;
	input \u0_R0_reg[5]/NET0131  ;
	input \u0_R0_reg[6]/NET0131  ;
	input \u0_R0_reg[7]/NET0131  ;
	input \u0_R0_reg[8]/NET0131  ;
	input \u0_R0_reg[9]/NET0131  ;
	input \u0_R10_reg[10]/NET0131  ;
	input \u0_R10_reg[11]/NET0131  ;
	input \u0_R10_reg[12]/NET0131  ;
	input \u0_R10_reg[13]/NET0131  ;
	input \u0_R10_reg[14]/NET0131  ;
	input \u0_R10_reg[15]/NET0131  ;
	input \u0_R10_reg[16]/NET0131  ;
	input \u0_R10_reg[17]/NET0131  ;
	input \u0_R10_reg[18]/NET0131  ;
	input \u0_R10_reg[19]/NET0131  ;
	input \u0_R10_reg[1]/NET0131  ;
	input \u0_R10_reg[20]/NET0131  ;
	input \u0_R10_reg[21]/NET0131  ;
	input \u0_R10_reg[22]/NET0131  ;
	input \u0_R10_reg[23]/NET0131  ;
	input \u0_R10_reg[24]/NET0131  ;
	input \u0_R10_reg[25]/NET0131  ;
	input \u0_R10_reg[26]/NET0131  ;
	input \u0_R10_reg[27]/NET0131  ;
	input \u0_R10_reg[28]/NET0131  ;
	input \u0_R10_reg[29]/NET0131  ;
	input \u0_R10_reg[2]/NET0131  ;
	input \u0_R10_reg[30]/NET0131  ;
	input \u0_R10_reg[31]/P0001  ;
	input \u0_R10_reg[32]/NET0131  ;
	input \u0_R10_reg[3]/NET0131  ;
	input \u0_R10_reg[4]/NET0131  ;
	input \u0_R10_reg[5]/NET0131  ;
	input \u0_R10_reg[6]/NET0131  ;
	input \u0_R10_reg[7]/NET0131  ;
	input \u0_R10_reg[8]/NET0131  ;
	input \u0_R10_reg[9]/NET0131  ;
	input \u0_R11_reg[10]/NET0131  ;
	input \u0_R11_reg[11]/P0001  ;
	input \u0_R11_reg[12]/NET0131  ;
	input \u0_R11_reg[13]/NET0131  ;
	input \u0_R11_reg[14]/NET0131  ;
	input \u0_R11_reg[15]/NET0131  ;
	input \u0_R11_reg[16]/NET0131  ;
	input \u0_R11_reg[17]/NET0131  ;
	input \u0_R11_reg[18]/NET0131  ;
	input \u0_R11_reg[19]/NET0131  ;
	input \u0_R11_reg[1]/NET0131  ;
	input \u0_R11_reg[20]/NET0131  ;
	input \u0_R11_reg[21]/NET0131  ;
	input \u0_R11_reg[22]/NET0131  ;
	input \u0_R11_reg[23]/NET0131  ;
	input \u0_R11_reg[24]/NET0131  ;
	input \u0_R11_reg[25]/NET0131  ;
	input \u0_R11_reg[26]/NET0131  ;
	input \u0_R11_reg[27]/NET0131  ;
	input \u0_R11_reg[28]/NET0131  ;
	input \u0_R11_reg[29]/NET0131  ;
	input \u0_R11_reg[2]/NET0131  ;
	input \u0_R11_reg[30]/NET0131  ;
	input \u0_R11_reg[31]/P0001  ;
	input \u0_R11_reg[32]/NET0131  ;
	input \u0_R11_reg[3]/NET0131  ;
	input \u0_R11_reg[4]/NET0131  ;
	input \u0_R11_reg[5]/NET0131  ;
	input \u0_R11_reg[6]/NET0131  ;
	input \u0_R11_reg[7]/NET0131  ;
	input \u0_R11_reg[8]/NET0131  ;
	input \u0_R11_reg[9]/NET0131  ;
	input \u0_R12_reg[10]/NET0131  ;
	input \u0_R12_reg[11]/NET0131  ;
	input \u0_R12_reg[12]/NET0131  ;
	input \u0_R12_reg[13]/NET0131  ;
	input \u0_R12_reg[14]/NET0131  ;
	input \u0_R12_reg[15]/NET0131  ;
	input \u0_R12_reg[16]/NET0131  ;
	input \u0_R12_reg[17]/NET0131  ;
	input \u0_R12_reg[18]/NET0131  ;
	input \u0_R12_reg[19]/NET0131  ;
	input \u0_R12_reg[1]/NET0131  ;
	input \u0_R12_reg[20]/NET0131  ;
	input \u0_R12_reg[21]/NET0131  ;
	input \u0_R12_reg[22]/NET0131  ;
	input \u0_R12_reg[23]/NET0131  ;
	input \u0_R12_reg[24]/NET0131  ;
	input \u0_R12_reg[25]/NET0131  ;
	input \u0_R12_reg[26]/NET0131  ;
	input \u0_R12_reg[27]/NET0131  ;
	input \u0_R12_reg[28]/NET0131  ;
	input \u0_R12_reg[29]/NET0131  ;
	input \u0_R12_reg[2]/NET0131  ;
	input \u0_R12_reg[30]/NET0131  ;
	input \u0_R12_reg[31]/P0001  ;
	input \u0_R12_reg[32]/NET0131  ;
	input \u0_R12_reg[3]/NET0131  ;
	input \u0_R12_reg[4]/NET0131  ;
	input \u0_R12_reg[5]/NET0131  ;
	input \u0_R12_reg[6]/NET0131  ;
	input \u0_R12_reg[7]/NET0131  ;
	input \u0_R12_reg[8]/NET0131  ;
	input \u0_R12_reg[9]/NET0131  ;
	input \u0_R13_reg[10]/NET0131  ;
	input \u0_R13_reg[11]/NET0131  ;
	input \u0_R13_reg[12]/NET0131  ;
	input \u0_R13_reg[13]/NET0131  ;
	input \u0_R13_reg[14]/NET0131  ;
	input \u0_R13_reg[15]/NET0131  ;
	input \u0_R13_reg[16]/NET0131  ;
	input \u0_R13_reg[17]/NET0131  ;
	input \u0_R13_reg[18]/NET0131  ;
	input \u0_R13_reg[19]/NET0131  ;
	input \u0_R13_reg[1]/NET0131  ;
	input \u0_R13_reg[20]/NET0131  ;
	input \u0_R13_reg[21]/NET0131  ;
	input \u0_R13_reg[22]/P0001  ;
	input \u0_R13_reg[23]/NET0131  ;
	input \u0_R13_reg[24]/NET0131  ;
	input \u0_R13_reg[25]/NET0131  ;
	input \u0_R13_reg[26]/NET0131  ;
	input \u0_R13_reg[27]/P0001  ;
	input \u0_R13_reg[28]/NET0131  ;
	input \u0_R13_reg[29]/NET0131  ;
	input \u0_R13_reg[2]/NET0131  ;
	input \u0_R13_reg[30]/NET0131  ;
	input \u0_R13_reg[31]/NET0131  ;
	input \u0_R13_reg[32]/NET0131  ;
	input \u0_R13_reg[3]/NET0131  ;
	input \u0_R13_reg[4]/NET0131  ;
	input \u0_R13_reg[5]/NET0131  ;
	input \u0_R13_reg[6]/NET0131  ;
	input \u0_R13_reg[7]/NET0131  ;
	input \u0_R13_reg[8]/NET0131  ;
	input \u0_R13_reg[9]/NET0131  ;
	input \u0_R14_reg[10]/NET0131  ;
	input \u0_R14_reg[11]/P0001  ;
	input \u0_R14_reg[12]/NET0131  ;
	input \u0_R14_reg[13]/NET0131  ;
	input \u0_R14_reg[14]/NET0131  ;
	input \u0_R14_reg[15]/NET0131  ;
	input \u0_R14_reg[16]/NET0131  ;
	input \u0_R14_reg[17]/NET0131  ;
	input \u0_R14_reg[18]/NET0131  ;
	input \u0_R14_reg[19]/NET0131  ;
	input \u0_R14_reg[1]/NET0131  ;
	input \u0_R14_reg[20]/NET0131  ;
	input \u0_R14_reg[21]/NET0131  ;
	input \u0_R14_reg[22]/P0001  ;
	input \u0_R14_reg[23]/NET0131  ;
	input \u0_R14_reg[24]/NET0131  ;
	input \u0_R14_reg[25]/NET0131  ;
	input \u0_R14_reg[26]/P0001  ;
	input \u0_R14_reg[27]/P0001  ;
	input \u0_R14_reg[28]/NET0131  ;
	input \u0_R14_reg[29]/NET0131  ;
	input \u0_R14_reg[2]/NET0131  ;
	input \u0_R14_reg[30]/NET0131  ;
	input \u0_R14_reg[31]/P0001  ;
	input \u0_R14_reg[32]/NET0131  ;
	input \u0_R14_reg[3]/NET0131  ;
	input \u0_R14_reg[4]/NET0131  ;
	input \u0_R14_reg[5]/NET0131  ;
	input \u0_R14_reg[6]/NET0131  ;
	input \u0_R14_reg[7]/NET0131  ;
	input \u0_R14_reg[8]/NET0131  ;
	input \u0_R14_reg[9]/NET0131  ;
	input \u0_R1_reg[10]/NET0131  ;
	input \u0_R1_reg[11]/NET0131  ;
	input \u0_R1_reg[12]/NET0131  ;
	input \u0_R1_reg[13]/NET0131  ;
	input \u0_R1_reg[14]/NET0131  ;
	input \u0_R1_reg[15]/NET0131  ;
	input \u0_R1_reg[16]/NET0131  ;
	input \u0_R1_reg[17]/NET0131  ;
	input \u0_R1_reg[18]/NET0131  ;
	input \u0_R1_reg[19]/NET0131  ;
	input \u0_R1_reg[1]/NET0131  ;
	input \u0_R1_reg[20]/NET0131  ;
	input \u0_R1_reg[21]/NET0131  ;
	input \u0_R1_reg[22]/NET0131  ;
	input \u0_R1_reg[23]/NET0131  ;
	input \u0_R1_reg[24]/NET0131  ;
	input \u0_R1_reg[25]/NET0131  ;
	input \u0_R1_reg[26]/NET0131  ;
	input \u0_R1_reg[27]/NET0131  ;
	input \u0_R1_reg[28]/NET0131  ;
	input \u0_R1_reg[29]/NET0131  ;
	input \u0_R1_reg[2]/NET0131  ;
	input \u0_R1_reg[30]/NET0131  ;
	input \u0_R1_reg[31]/NET0131  ;
	input \u0_R1_reg[32]/NET0131  ;
	input \u0_R1_reg[3]/NET0131  ;
	input \u0_R1_reg[4]/NET0131  ;
	input \u0_R1_reg[5]/NET0131  ;
	input \u0_R1_reg[6]/NET0131  ;
	input \u0_R1_reg[7]/NET0131  ;
	input \u0_R1_reg[8]/NET0131  ;
	input \u0_R1_reg[9]/NET0131  ;
	input \u0_R2_reg[10]/NET0131  ;
	input \u0_R2_reg[11]/NET0131  ;
	input \u0_R2_reg[12]/NET0131  ;
	input \u0_R2_reg[13]/NET0131  ;
	input \u0_R2_reg[14]/NET0131  ;
	input \u0_R2_reg[15]/NET0131  ;
	input \u0_R2_reg[16]/NET0131  ;
	input \u0_R2_reg[17]/NET0131  ;
	input \u0_R2_reg[18]/NET0131  ;
	input \u0_R2_reg[19]/NET0131  ;
	input \u0_R2_reg[1]/NET0131  ;
	input \u0_R2_reg[20]/NET0131  ;
	input \u0_R2_reg[21]/NET0131  ;
	input \u0_R2_reg[22]/NET0131  ;
	input \u0_R2_reg[23]/NET0131  ;
	input \u0_R2_reg[24]/NET0131  ;
	input \u0_R2_reg[25]/NET0131  ;
	input \u0_R2_reg[26]/NET0131  ;
	input \u0_R2_reg[27]/NET0131  ;
	input \u0_R2_reg[28]/NET0131  ;
	input \u0_R2_reg[29]/NET0131  ;
	input \u0_R2_reg[2]/NET0131  ;
	input \u0_R2_reg[30]/NET0131  ;
	input \u0_R2_reg[31]/NET0131  ;
	input \u0_R2_reg[32]/NET0131  ;
	input \u0_R2_reg[3]/NET0131  ;
	input \u0_R2_reg[4]/NET0131  ;
	input \u0_R2_reg[5]/NET0131  ;
	input \u0_R2_reg[6]/NET0131  ;
	input \u0_R2_reg[7]/NET0131  ;
	input \u0_R2_reg[8]/NET0131  ;
	input \u0_R2_reg[9]/NET0131  ;
	input \u0_R3_reg[10]/NET0131  ;
	input \u0_R3_reg[11]/NET0131  ;
	input \u0_R3_reg[12]/NET0131  ;
	input \u0_R3_reg[13]/NET0131  ;
	input \u0_R3_reg[14]/NET0131  ;
	input \u0_R3_reg[15]/NET0131  ;
	input \u0_R3_reg[16]/NET0131  ;
	input \u0_R3_reg[17]/NET0131  ;
	input \u0_R3_reg[18]/NET0131  ;
	input \u0_R3_reg[19]/NET0131  ;
	input \u0_R3_reg[1]/NET0131  ;
	input \u0_R3_reg[20]/NET0131  ;
	input \u0_R3_reg[21]/NET0131  ;
	input \u0_R3_reg[22]/NET0131  ;
	input \u0_R3_reg[23]/NET0131  ;
	input \u0_R3_reg[24]/NET0131  ;
	input \u0_R3_reg[25]/NET0131  ;
	input \u0_R3_reg[26]/NET0131  ;
	input \u0_R3_reg[27]/NET0131  ;
	input \u0_R3_reg[28]/NET0131  ;
	input \u0_R3_reg[29]/NET0131  ;
	input \u0_R3_reg[2]/NET0131  ;
	input \u0_R3_reg[30]/NET0131  ;
	input \u0_R3_reg[31]/P0001  ;
	input \u0_R3_reg[32]/NET0131  ;
	input \u0_R3_reg[3]/NET0131  ;
	input \u0_R3_reg[4]/NET0131  ;
	input \u0_R3_reg[5]/NET0131  ;
	input \u0_R3_reg[6]/NET0131  ;
	input \u0_R3_reg[7]/NET0131  ;
	input \u0_R3_reg[8]/NET0131  ;
	input \u0_R3_reg[9]/NET0131  ;
	input \u0_R4_reg[10]/NET0131  ;
	input \u0_R4_reg[11]/NET0131  ;
	input \u0_R4_reg[12]/NET0131  ;
	input \u0_R4_reg[13]/NET0131  ;
	input \u0_R4_reg[14]/NET0131  ;
	input \u0_R4_reg[15]/NET0131  ;
	input \u0_R4_reg[16]/NET0131  ;
	input \u0_R4_reg[17]/NET0131  ;
	input \u0_R4_reg[18]/NET0131  ;
	input \u0_R4_reg[19]/NET0131  ;
	input \u0_R4_reg[1]/NET0131  ;
	input \u0_R4_reg[20]/NET0131  ;
	input \u0_R4_reg[21]/NET0131  ;
	input \u0_R4_reg[22]/NET0131  ;
	input \u0_R4_reg[23]/NET0131  ;
	input \u0_R4_reg[24]/NET0131  ;
	input \u0_R4_reg[25]/NET0131  ;
	input \u0_R4_reg[26]/NET0131  ;
	input \u0_R4_reg[27]/NET0131  ;
	input \u0_R4_reg[28]/NET0131  ;
	input \u0_R4_reg[29]/NET0131  ;
	input \u0_R4_reg[2]/NET0131  ;
	input \u0_R4_reg[30]/NET0131  ;
	input \u0_R4_reg[31]/P0001  ;
	input \u0_R4_reg[32]/NET0131  ;
	input \u0_R4_reg[3]/NET0131  ;
	input \u0_R4_reg[4]/NET0131  ;
	input \u0_R4_reg[5]/NET0131  ;
	input \u0_R4_reg[6]/NET0131  ;
	input \u0_R4_reg[7]/NET0131  ;
	input \u0_R4_reg[8]/NET0131  ;
	input \u0_R4_reg[9]/NET0131  ;
	input \u0_R5_reg[10]/NET0131  ;
	input \u0_R5_reg[11]/P0001  ;
	input \u0_R5_reg[12]/NET0131  ;
	input \u0_R5_reg[13]/NET0131  ;
	input \u0_R5_reg[14]/NET0131  ;
	input \u0_R5_reg[15]/NET0131  ;
	input \u0_R5_reg[16]/NET0131  ;
	input \u0_R5_reg[17]/NET0131  ;
	input \u0_R5_reg[18]/NET0131  ;
	input \u0_R5_reg[19]/NET0131  ;
	input \u0_R5_reg[1]/NET0131  ;
	input \u0_R5_reg[20]/NET0131  ;
	input \u0_R5_reg[21]/NET0131  ;
	input \u0_R5_reg[22]/NET0131  ;
	input \u0_R5_reg[23]/NET0131  ;
	input \u0_R5_reg[24]/NET0131  ;
	input \u0_R5_reg[25]/NET0131  ;
	input \u0_R5_reg[26]/NET0131  ;
	input \u0_R5_reg[27]/NET0131  ;
	input \u0_R5_reg[28]/NET0131  ;
	input \u0_R5_reg[29]/NET0131  ;
	input \u0_R5_reg[2]/NET0131  ;
	input \u0_R5_reg[30]/NET0131  ;
	input \u0_R5_reg[31]/P0001  ;
	input \u0_R5_reg[32]/NET0131  ;
	input \u0_R5_reg[3]/NET0131  ;
	input \u0_R5_reg[4]/NET0131  ;
	input \u0_R5_reg[5]/NET0131  ;
	input \u0_R5_reg[6]/NET0131  ;
	input \u0_R5_reg[7]/NET0131  ;
	input \u0_R5_reg[8]/NET0131  ;
	input \u0_R5_reg[9]/NET0131  ;
	input \u0_R6_reg[10]/NET0131  ;
	input \u0_R6_reg[11]/NET0131  ;
	input \u0_R6_reg[12]/NET0131  ;
	input \u0_R6_reg[13]/NET0131  ;
	input \u0_R6_reg[14]/NET0131  ;
	input \u0_R6_reg[15]/NET0131  ;
	input \u0_R6_reg[16]/NET0131  ;
	input \u0_R6_reg[17]/NET0131  ;
	input \u0_R6_reg[18]/NET0131  ;
	input \u0_R6_reg[19]/NET0131  ;
	input \u0_R6_reg[1]/NET0131  ;
	input \u0_R6_reg[20]/NET0131  ;
	input \u0_R6_reg[21]/NET0131  ;
	input \u0_R6_reg[22]/NET0131  ;
	input \u0_R6_reg[23]/NET0131  ;
	input \u0_R6_reg[24]/NET0131  ;
	input \u0_R6_reg[25]/NET0131  ;
	input \u0_R6_reg[26]/NET0131  ;
	input \u0_R6_reg[27]/NET0131  ;
	input \u0_R6_reg[28]/NET0131  ;
	input \u0_R6_reg[29]/NET0131  ;
	input \u0_R6_reg[2]/NET0131  ;
	input \u0_R6_reg[30]/NET0131  ;
	input \u0_R6_reg[31]/P0001  ;
	input \u0_R6_reg[32]/NET0131  ;
	input \u0_R6_reg[3]/NET0131  ;
	input \u0_R6_reg[4]/NET0131  ;
	input \u0_R6_reg[5]/NET0131  ;
	input \u0_R6_reg[6]/NET0131  ;
	input \u0_R6_reg[7]/NET0131  ;
	input \u0_R6_reg[8]/NET0131  ;
	input \u0_R6_reg[9]/NET0131  ;
	input \u0_R7_reg[10]/NET0131  ;
	input \u0_R7_reg[11]/P0001  ;
	input \u0_R7_reg[12]/NET0131  ;
	input \u0_R7_reg[13]/NET0131  ;
	input \u0_R7_reg[14]/NET0131  ;
	input \u0_R7_reg[15]/NET0131  ;
	input \u0_R7_reg[16]/NET0131  ;
	input \u0_R7_reg[17]/NET0131  ;
	input \u0_R7_reg[18]/NET0131  ;
	input \u0_R7_reg[19]/NET0131  ;
	input \u0_R7_reg[1]/NET0131  ;
	input \u0_R7_reg[20]/NET0131  ;
	input \u0_R7_reg[21]/NET0131  ;
	input \u0_R7_reg[22]/NET0131  ;
	input \u0_R7_reg[23]/NET0131  ;
	input \u0_R7_reg[24]/NET0131  ;
	input \u0_R7_reg[25]/NET0131  ;
	input \u0_R7_reg[26]/NET0131  ;
	input \u0_R7_reg[27]/NET0131  ;
	input \u0_R7_reg[28]/NET0131  ;
	input \u0_R7_reg[29]/NET0131  ;
	input \u0_R7_reg[2]/NET0131  ;
	input \u0_R7_reg[30]/NET0131  ;
	input \u0_R7_reg[31]/P0001  ;
	input \u0_R7_reg[32]/NET0131  ;
	input \u0_R7_reg[3]/NET0131  ;
	input \u0_R7_reg[4]/NET0131  ;
	input \u0_R7_reg[5]/NET0131  ;
	input \u0_R7_reg[6]/NET0131  ;
	input \u0_R7_reg[7]/NET0131  ;
	input \u0_R7_reg[8]/NET0131  ;
	input \u0_R7_reg[9]/NET0131  ;
	input \u0_R8_reg[10]/NET0131  ;
	input \u0_R8_reg[11]/NET0131  ;
	input \u0_R8_reg[12]/NET0131  ;
	input \u0_R8_reg[13]/NET0131  ;
	input \u0_R8_reg[14]/NET0131  ;
	input \u0_R8_reg[15]/NET0131  ;
	input \u0_R8_reg[16]/NET0131  ;
	input \u0_R8_reg[17]/NET0131  ;
	input \u0_R8_reg[18]/NET0131  ;
	input \u0_R8_reg[19]/NET0131  ;
	input \u0_R8_reg[1]/NET0131  ;
	input \u0_R8_reg[20]/NET0131  ;
	input \u0_R8_reg[21]/NET0131  ;
	input \u0_R8_reg[22]/NET0131  ;
	input \u0_R8_reg[23]/NET0131  ;
	input \u0_R8_reg[24]/NET0131  ;
	input \u0_R8_reg[25]/NET0131  ;
	input \u0_R8_reg[26]/NET0131  ;
	input \u0_R8_reg[27]/NET0131  ;
	input \u0_R8_reg[28]/NET0131  ;
	input \u0_R8_reg[29]/NET0131  ;
	input \u0_R8_reg[2]/NET0131  ;
	input \u0_R8_reg[30]/NET0131  ;
	input \u0_R8_reg[31]/P0001  ;
	input \u0_R8_reg[32]/NET0131  ;
	input \u0_R8_reg[3]/NET0131  ;
	input \u0_R8_reg[4]/NET0131  ;
	input \u0_R8_reg[5]/NET0131  ;
	input \u0_R8_reg[6]/NET0131  ;
	input \u0_R8_reg[7]/NET0131  ;
	input \u0_R8_reg[8]/NET0131  ;
	input \u0_R8_reg[9]/NET0131  ;
	input \u0_R9_reg[10]/NET0131  ;
	input \u0_R9_reg[11]/P0001  ;
	input \u0_R9_reg[12]/NET0131  ;
	input \u0_R9_reg[13]/NET0131  ;
	input \u0_R9_reg[14]/NET0131  ;
	input \u0_R9_reg[15]/NET0131  ;
	input \u0_R9_reg[16]/NET0131  ;
	input \u0_R9_reg[17]/NET0131  ;
	input \u0_R9_reg[18]/NET0131  ;
	input \u0_R9_reg[19]/NET0131  ;
	input \u0_R9_reg[1]/NET0131  ;
	input \u0_R9_reg[20]/NET0131  ;
	input \u0_R9_reg[21]/NET0131  ;
	input \u0_R9_reg[22]/NET0131  ;
	input \u0_R9_reg[23]/NET0131  ;
	input \u0_R9_reg[24]/NET0131  ;
	input \u0_R9_reg[25]/NET0131  ;
	input \u0_R9_reg[26]/NET0131  ;
	input \u0_R9_reg[27]/NET0131  ;
	input \u0_R9_reg[28]/NET0131  ;
	input \u0_R9_reg[29]/NET0131  ;
	input \u0_R9_reg[2]/NET0131  ;
	input \u0_R9_reg[30]/NET0131  ;
	input \u0_R9_reg[31]/P0001  ;
	input \u0_R9_reg[32]/NET0131  ;
	input \u0_R9_reg[3]/NET0131  ;
	input \u0_R9_reg[4]/NET0131  ;
	input \u0_R9_reg[5]/NET0131  ;
	input \u0_R9_reg[6]/NET0131  ;
	input \u0_R9_reg[7]/NET0131  ;
	input \u0_R9_reg[8]/NET0131  ;
	input \u0_R9_reg[9]/NET0131  ;
	input \u0_desIn_r_reg[0]/NET0131  ;
	input \u0_desIn_r_reg[10]/NET0131  ;
	input \u0_desIn_r_reg[11]/NET0131  ;
	input \u0_desIn_r_reg[12]/NET0131  ;
	input \u0_desIn_r_reg[13]/NET0131  ;
	input \u0_desIn_r_reg[14]/NET0131  ;
	input \u0_desIn_r_reg[15]/NET0131  ;
	input \u0_desIn_r_reg[16]/NET0131  ;
	input \u0_desIn_r_reg[17]/NET0131  ;
	input \u0_desIn_r_reg[18]/NET0131  ;
	input \u0_desIn_r_reg[19]/NET0131  ;
	input \u0_desIn_r_reg[1]/NET0131  ;
	input \u0_desIn_r_reg[20]/NET0131  ;
	input \u0_desIn_r_reg[21]/NET0131  ;
	input \u0_desIn_r_reg[22]/NET0131  ;
	input \u0_desIn_r_reg[23]/NET0131  ;
	input \u0_desIn_r_reg[24]/NET0131  ;
	input \u0_desIn_r_reg[25]/NET0131  ;
	input \u0_desIn_r_reg[26]/NET0131  ;
	input \u0_desIn_r_reg[27]/NET0131  ;
	input \u0_desIn_r_reg[28]/NET0131  ;
	input \u0_desIn_r_reg[29]/NET0131  ;
	input \u0_desIn_r_reg[2]/NET0131  ;
	input \u0_desIn_r_reg[30]/NET0131  ;
	input \u0_desIn_r_reg[31]/NET0131  ;
	input \u0_desIn_r_reg[32]/NET0131  ;
	input \u0_desIn_r_reg[33]/NET0131  ;
	input \u0_desIn_r_reg[34]/NET0131  ;
	input \u0_desIn_r_reg[35]/NET0131  ;
	input \u0_desIn_r_reg[36]/NET0131  ;
	input \u0_desIn_r_reg[37]/NET0131  ;
	input \u0_desIn_r_reg[38]/NET0131  ;
	input \u0_desIn_r_reg[39]/NET0131  ;
	input \u0_desIn_r_reg[3]/NET0131  ;
	input \u0_desIn_r_reg[40]/NET0131  ;
	input \u0_desIn_r_reg[41]/NET0131  ;
	input \u0_desIn_r_reg[42]/NET0131  ;
	input \u0_desIn_r_reg[43]/NET0131  ;
	input \u0_desIn_r_reg[44]/NET0131  ;
	input \u0_desIn_r_reg[45]/NET0131  ;
	input \u0_desIn_r_reg[46]/NET0131  ;
	input \u0_desIn_r_reg[47]/NET0131  ;
	input \u0_desIn_r_reg[48]/NET0131  ;
	input \u0_desIn_r_reg[49]/NET0131  ;
	input \u0_desIn_r_reg[4]/NET0131  ;
	input \u0_desIn_r_reg[50]/NET0131  ;
	input \u0_desIn_r_reg[51]/NET0131  ;
	input \u0_desIn_r_reg[52]/NET0131  ;
	input \u0_desIn_r_reg[53]/NET0131  ;
	input \u0_desIn_r_reg[54]/NET0131  ;
	input \u0_desIn_r_reg[55]/NET0131  ;
	input \u0_desIn_r_reg[56]/NET0131  ;
	input \u0_desIn_r_reg[57]/NET0131  ;
	input \u0_desIn_r_reg[58]/NET0131  ;
	input \u0_desIn_r_reg[59]/NET0131  ;
	input \u0_desIn_r_reg[5]/NET0131  ;
	input \u0_desIn_r_reg[60]/NET0131  ;
	input \u0_desIn_r_reg[61]/NET0131  ;
	input \u0_desIn_r_reg[62]/NET0131  ;
	input \u0_desIn_r_reg[63]/NET0131  ;
	input \u0_desIn_r_reg[6]/NET0131  ;
	input \u0_desIn_r_reg[7]/NET0131  ;
	input \u0_desIn_r_reg[8]/NET0131  ;
	input \u0_desIn_r_reg[9]/NET0131  ;
	input \u0_key_r_reg[0]/NET0131  ;
	input \u0_key_r_reg[10]/P0001  ;
	input \u0_key_r_reg[11]/NET0131  ;
	input \u0_key_r_reg[12]/NET0131  ;
	input \u0_key_r_reg[13]/NET0131  ;
	input \u0_key_r_reg[14]/NET0131  ;
	input \u0_key_r_reg[15]/NET0131  ;
	input \u0_key_r_reg[16]/NET0131  ;
	input \u0_key_r_reg[17]/NET0131  ;
	input \u0_key_r_reg[18]/NET0131  ;
	input \u0_key_r_reg[19]/NET0131  ;
	input \u0_key_r_reg[1]/NET0131  ;
	input \u0_key_r_reg[20]/NET0131  ;
	input \u0_key_r_reg[21]/NET0131  ;
	input \u0_key_r_reg[22]/NET0131  ;
	input \u0_key_r_reg[23]/NET0131  ;
	input \u0_key_r_reg[24]/NET0131  ;
	input \u0_key_r_reg[25]/NET0131  ;
	input \u0_key_r_reg[26]/NET0131  ;
	input \u0_key_r_reg[27]/NET0131  ;
	input \u0_key_r_reg[28]/NET0131  ;
	input \u0_key_r_reg[29]/NET0131  ;
	input \u0_key_r_reg[2]/NET0131  ;
	input \u0_key_r_reg[30]/NET0131  ;
	input \u0_key_r_reg[31]/NET0131  ;
	input \u0_key_r_reg[32]/NET0131  ;
	input \u0_key_r_reg[33]/NET0131  ;
	input \u0_key_r_reg[34]/NET0131  ;
	input \u0_key_r_reg[35]/P0001  ;
	input \u0_key_r_reg[36]/NET0131  ;
	input \u0_key_r_reg[37]/NET0131  ;
	input \u0_key_r_reg[38]/NET0131  ;
	input \u0_key_r_reg[39]/P0001  ;
	input \u0_key_r_reg[3]/NET0131  ;
	input \u0_key_r_reg[40]/NET0131  ;
	input \u0_key_r_reg[41]/NET0131  ;
	input \u0_key_r_reg[42]/P0001  ;
	input \u0_key_r_reg[43]/NET0131  ;
	input \u0_key_r_reg[44]/NET0131  ;
	input \u0_key_r_reg[45]/NET0131  ;
	input \u0_key_r_reg[46]/NET0131  ;
	input \u0_key_r_reg[47]/NET0131  ;
	input \u0_key_r_reg[48]/NET0131  ;
	input \u0_key_r_reg[49]/NET0131  ;
	input \u0_key_r_reg[4]/NET0131  ;
	input \u0_key_r_reg[50]/NET0131  ;
	input \u0_key_r_reg[51]/NET0131  ;
	input \u0_key_r_reg[52]/NET0131  ;
	input \u0_key_r_reg[53]/NET0131  ;
	input \u0_key_r_reg[54]/NET0131  ;
	input \u0_key_r_reg[55]/NET0131  ;
	input \u0_key_r_reg[5]/NET0131  ;
	input \u0_key_r_reg[6]/NET0131  ;
	input \u0_key_r_reg[7]/NET0131  ;
	input \u0_key_r_reg[8]/NET0131  ;
	input \u0_key_r_reg[9]/NET0131  ;
	input \u0_uk_K_r0_reg[0]/NET0131  ;
	input \u0_uk_K_r0_reg[10]/NET0131  ;
	input \u0_uk_K_r0_reg[11]/NET0131  ;
	input \u0_uk_K_r0_reg[12]/NET0131  ;
	input \u0_uk_K_r0_reg[13]/NET0131  ;
	input \u0_uk_K_r0_reg[14]/NET0131  ;
	input \u0_uk_K_r0_reg[15]/NET0131  ;
	input \u0_uk_K_r0_reg[16]/NET0131  ;
	input \u0_uk_K_r0_reg[17]/NET0131  ;
	input \u0_uk_K_r0_reg[18]/NET0131  ;
	input \u0_uk_K_r0_reg[19]/NET0131  ;
	input \u0_uk_K_r0_reg[20]/NET0131  ;
	input \u0_uk_K_r0_reg[21]/NET0131  ;
	input \u0_uk_K_r0_reg[22]/NET0131  ;
	input \u0_uk_K_r0_reg[23]/NET0131  ;
	input \u0_uk_K_r0_reg[24]/P0001  ;
	input \u0_uk_K_r0_reg[25]/P0001  ;
	input \u0_uk_K_r0_reg[26]/NET0131  ;
	input \u0_uk_K_r0_reg[27]/NET0131  ;
	input \u0_uk_K_r0_reg[28]/NET0131  ;
	input \u0_uk_K_r0_reg[29]/NET0131  ;
	input \u0_uk_K_r0_reg[2]/NET0131  ;
	input \u0_uk_K_r0_reg[30]/NET0131  ;
	input \u0_uk_K_r0_reg[31]/NET0131  ;
	input \u0_uk_K_r0_reg[32]/NET0131  ;
	input \u0_uk_K_r0_reg[33]/NET0131  ;
	input \u0_uk_K_r0_reg[34]/NET0131  ;
	input \u0_uk_K_r0_reg[35]/NET0131  ;
	input \u0_uk_K_r0_reg[36]/NET0131  ;
	input \u0_uk_K_r0_reg[37]/NET0131  ;
	input \u0_uk_K_r0_reg[38]/NET0131  ;
	input \u0_uk_K_r0_reg[39]/NET0131  ;
	input \u0_uk_K_r0_reg[3]/NET0131  ;
	input \u0_uk_K_r0_reg[40]/NET0131  ;
	input \u0_uk_K_r0_reg[41]/NET0131  ;
	input \u0_uk_K_r0_reg[42]/NET0131  ;
	input \u0_uk_K_r0_reg[43]/NET0131  ;
	input \u0_uk_K_r0_reg[44]/NET0131  ;
	input \u0_uk_K_r0_reg[45]/NET0131  ;
	input \u0_uk_K_r0_reg[46]/NET0131  ;
	input \u0_uk_K_r0_reg[47]/NET0131  ;
	input \u0_uk_K_r0_reg[48]/NET0131  ;
	input \u0_uk_K_r0_reg[49]/NET0131  ;
	input \u0_uk_K_r0_reg[4]/NET0131  ;
	input \u0_uk_K_r0_reg[50]/NET0131  ;
	input \u0_uk_K_r0_reg[51]/NET0131  ;
	input \u0_uk_K_r0_reg[52]/NET0131  ;
	input \u0_uk_K_r0_reg[54]/NET0131  ;
	input \u0_uk_K_r0_reg[55]/NET0131  ;
	input \u0_uk_K_r0_reg[5]/NET0131  ;
	input \u0_uk_K_r0_reg[6]/NET0131  ;
	input \u0_uk_K_r0_reg[7]/NET0131  ;
	input \u0_uk_K_r0_reg[8]/NET0131  ;
	input \u0_uk_K_r0_reg[9]/NET0131  ;
	input \u0_uk_K_r10_reg[0]/NET0131  ;
	input \u0_uk_K_r10_reg[10]/NET0131  ;
	input \u0_uk_K_r10_reg[11]/NET0131  ;
	input \u0_uk_K_r10_reg[12]/NET0131  ;
	input \u0_uk_K_r10_reg[14]/NET0131  ;
	input \u0_uk_K_r10_reg[15]/NET0131  ;
	input \u0_uk_K_r10_reg[16]/NET0131  ;
	input \u0_uk_K_r10_reg[17]/NET0131  ;
	input \u0_uk_K_r10_reg[18]/NET0131  ;
	input \u0_uk_K_r10_reg[19]/NET0131  ;
	input \u0_uk_K_r10_reg[1]/NET0131  ;
	input \u0_uk_K_r10_reg[20]/NET0131  ;
	input \u0_uk_K_r10_reg[21]/NET0131  ;
	input \u0_uk_K_r10_reg[22]/NET0131  ;
	input \u0_uk_K_r10_reg[23]/NET0131  ;
	input \u0_uk_K_r10_reg[24]/NET0131  ;
	input \u0_uk_K_r10_reg[25]/NET0131  ;
	input \u0_uk_K_r10_reg[26]/NET0131  ;
	input \u0_uk_K_r10_reg[27]/NET0131  ;
	input \u0_uk_K_r10_reg[28]/NET0131  ;
	input \u0_uk_K_r10_reg[29]/NET0131  ;
	input \u0_uk_K_r10_reg[2]/NET0131  ;
	input \u0_uk_K_r10_reg[30]/NET0131  ;
	input \u0_uk_K_r10_reg[31]/NET0131  ;
	input \u0_uk_K_r10_reg[32]/NET0131  ;
	input \u0_uk_K_r10_reg[33]/NET0131  ;
	input \u0_uk_K_r10_reg[34]/NET0131  ;
	input \u0_uk_K_r10_reg[35]/NET0131  ;
	input \u0_uk_K_r10_reg[36]/NET0131  ;
	input \u0_uk_K_r10_reg[37]/NET0131  ;
	input \u0_uk_K_r10_reg[38]/NET0131  ;
	input \u0_uk_K_r10_reg[39]/NET0131  ;
	input \u0_uk_K_r10_reg[3]/NET0131  ;
	input \u0_uk_K_r10_reg[40]/NET0131  ;
	input \u0_uk_K_r10_reg[41]/P0001  ;
	input \u0_uk_K_r10_reg[42]/NET0131  ;
	input \u0_uk_K_r10_reg[43]/NET0131  ;
	input \u0_uk_K_r10_reg[44]/NET0131  ;
	input \u0_uk_K_r10_reg[45]/P0001  ;
	input \u0_uk_K_r10_reg[46]/NET0131  ;
	input \u0_uk_K_r10_reg[47]/NET0131  ;
	input \u0_uk_K_r10_reg[48]/NET0131  ;
	input \u0_uk_K_r10_reg[49]/NET0131  ;
	input \u0_uk_K_r10_reg[4]/NET0131  ;
	input \u0_uk_K_r10_reg[50]/NET0131  ;
	input \u0_uk_K_r10_reg[51]/NET0131  ;
	input \u0_uk_K_r10_reg[52]/NET0131  ;
	input \u0_uk_K_r10_reg[53]/NET0131  ;
	input \u0_uk_K_r10_reg[54]/NET0131  ;
	input \u0_uk_K_r10_reg[55]/NET0131  ;
	input \u0_uk_K_r10_reg[5]/NET0131  ;
	input \u0_uk_K_r10_reg[6]/NET0131  ;
	input \u0_uk_K_r10_reg[7]/NET0131  ;
	input \u0_uk_K_r10_reg[8]/NET0131  ;
	input \u0_uk_K_r10_reg[9]/NET0131  ;
	input \u0_uk_K_r11_reg[0]/NET0131  ;
	input \u0_uk_K_r11_reg[10]/NET0131  ;
	input \u0_uk_K_r11_reg[11]/NET0131  ;
	input \u0_uk_K_r11_reg[12]/NET0131  ;
	input \u0_uk_K_r11_reg[13]/NET0131  ;
	input \u0_uk_K_r11_reg[14]/NET0131  ;
	input \u0_uk_K_r11_reg[15]/NET0131  ;
	input \u0_uk_K_r11_reg[16]/NET0131  ;
	input \u0_uk_K_r11_reg[17]/NET0131  ;
	input \u0_uk_K_r11_reg[18]/NET0131  ;
	input \u0_uk_K_r11_reg[19]/NET0131  ;
	input \u0_uk_K_r11_reg[1]/NET0131  ;
	input \u0_uk_K_r11_reg[20]/NET0131  ;
	input \u0_uk_K_r11_reg[21]/NET0131  ;
	input \u0_uk_K_r11_reg[22]/NET0131  ;
	input \u0_uk_K_r11_reg[23]/NET0131  ;
	input \u0_uk_K_r11_reg[24]/NET0131  ;
	input \u0_uk_K_r11_reg[25]/NET0131  ;
	input \u0_uk_K_r11_reg[26]/NET0131  ;
	input \u0_uk_K_r11_reg[27]/P0001  ;
	input \u0_uk_K_r11_reg[28]/NET0131  ;
	input \u0_uk_K_r11_reg[29]/NET0131  ;
	input \u0_uk_K_r11_reg[2]/NET0131  ;
	input \u0_uk_K_r11_reg[31]/NET0131  ;
	input \u0_uk_K_r11_reg[32]/NET0131  ;
	input \u0_uk_K_r11_reg[33]/NET0131  ;
	input \u0_uk_K_r11_reg[34]/NET0131  ;
	input \u0_uk_K_r11_reg[35]/NET0131  ;
	input \u0_uk_K_r11_reg[36]/NET0131  ;
	input \u0_uk_K_r11_reg[37]/NET0131  ;
	input \u0_uk_K_r11_reg[38]/NET0131  ;
	input \u0_uk_K_r11_reg[39]/NET0131  ;
	input \u0_uk_K_r11_reg[3]/NET0131  ;
	input \u0_uk_K_r11_reg[40]/NET0131  ;
	input \u0_uk_K_r11_reg[41]/NET0131  ;
	input \u0_uk_K_r11_reg[42]/NET0131  ;
	input \u0_uk_K_r11_reg[43]/NET0131  ;
	input \u0_uk_K_r11_reg[44]/NET0131  ;
	input \u0_uk_K_r11_reg[45]/NET0131  ;
	input \u0_uk_K_r11_reg[46]/NET0131  ;
	input \u0_uk_K_r11_reg[47]/NET0131  ;
	input \u0_uk_K_r11_reg[48]/NET0131  ;
	input \u0_uk_K_r11_reg[49]/NET0131  ;
	input \u0_uk_K_r11_reg[4]/NET0131  ;
	input \u0_uk_K_r11_reg[50]/NET0131  ;
	input \u0_uk_K_r11_reg[51]/NET0131  ;
	input \u0_uk_K_r11_reg[52]/NET0131  ;
	input \u0_uk_K_r11_reg[53]/P0001  ;
	input \u0_uk_K_r11_reg[54]/NET0131  ;
	input \u0_uk_K_r11_reg[55]/NET0131  ;
	input \u0_uk_K_r11_reg[5]/NET0131  ;
	input \u0_uk_K_r11_reg[6]/NET0131  ;
	input \u0_uk_K_r11_reg[7]/NET0131  ;
	input \u0_uk_K_r11_reg[8]/NET0131  ;
	input \u0_uk_K_r11_reg[9]/NET0131  ;
	input \u0_uk_K_r12_reg[0]/NET0131  ;
	input \u0_uk_K_r12_reg[10]/P0001  ;
	input \u0_uk_K_r12_reg[11]/NET0131  ;
	input \u0_uk_K_r12_reg[12]/NET0131  ;
	input \u0_uk_K_r12_reg[13]/NET0131  ;
	input \u0_uk_K_r12_reg[14]/NET0131  ;
	input \u0_uk_K_r12_reg[15]/NET0131  ;
	input \u0_uk_K_r12_reg[16]/NET0131  ;
	input \u0_uk_K_r12_reg[17]/NET0131  ;
	input \u0_uk_K_r12_reg[18]/NET0131  ;
	input \u0_uk_K_r12_reg[19]/NET0131  ;
	input \u0_uk_K_r12_reg[1]/NET0131  ;
	input \u0_uk_K_r12_reg[20]/NET0131  ;
	input \u0_uk_K_r12_reg[21]/NET0131  ;
	input \u0_uk_K_r12_reg[22]/NET0131  ;
	input \u0_uk_K_r12_reg[23]/NET0131  ;
	input \u0_uk_K_r12_reg[24]/NET0131  ;
	input \u0_uk_K_r12_reg[25]/NET0131  ;
	input \u0_uk_K_r12_reg[26]/NET0131  ;
	input \u0_uk_K_r12_reg[27]/NET0131  ;
	input \u0_uk_K_r12_reg[28]/NET0131  ;
	input \u0_uk_K_r12_reg[29]/NET0131  ;
	input \u0_uk_K_r12_reg[2]/NET0131  ;
	input \u0_uk_K_r12_reg[30]/NET0131  ;
	input \u0_uk_K_r12_reg[31]/NET0131  ;
	input \u0_uk_K_r12_reg[32]/NET0131  ;
	input \u0_uk_K_r12_reg[33]/NET0131  ;
	input \u0_uk_K_r12_reg[34]/NET0131  ;
	input \u0_uk_K_r12_reg[35]/NET0131  ;
	input \u0_uk_K_r12_reg[36]/NET0131  ;
	input \u0_uk_K_r12_reg[37]/NET0131  ;
	input \u0_uk_K_r12_reg[38]/NET0131  ;
	input \u0_uk_K_r12_reg[3]/NET0131  ;
	input \u0_uk_K_r12_reg[40]/NET0131  ;
	input \u0_uk_K_r12_reg[41]/NET0131  ;
	input \u0_uk_K_r12_reg[42]/NET0131  ;
	input \u0_uk_K_r12_reg[43]/NET0131  ;
	input \u0_uk_K_r12_reg[44]/P0001  ;
	input \u0_uk_K_r12_reg[45]/NET0131  ;
	input \u0_uk_K_r12_reg[46]/NET0131  ;
	input \u0_uk_K_r12_reg[47]/NET0131  ;
	input \u0_uk_K_r12_reg[48]/NET0131  ;
	input \u0_uk_K_r12_reg[49]/NET0131  ;
	input \u0_uk_K_r12_reg[4]/NET0131  ;
	input \u0_uk_K_r12_reg[50]/NET0131  ;
	input \u0_uk_K_r12_reg[51]/NET0131  ;
	input \u0_uk_K_r12_reg[52]/NET0131  ;
	input \u0_uk_K_r12_reg[53]/NET0131  ;
	input \u0_uk_K_r12_reg[54]/NET0131  ;
	input \u0_uk_K_r12_reg[55]/NET0131  ;
	input \u0_uk_K_r12_reg[5]/NET0131  ;
	input \u0_uk_K_r12_reg[6]/NET0131  ;
	input \u0_uk_K_r12_reg[7]/P0001  ;
	input \u0_uk_K_r12_reg[8]/NET0131  ;
	input \u0_uk_K_r12_reg[9]/NET0131  ;
	input \u0_uk_K_r13_reg[0]/NET0131  ;
	input \u0_uk_K_r13_reg[10]/NET0131  ;
	input \u0_uk_K_r13_reg[11]/NET0131  ;
	input \u0_uk_K_r13_reg[12]/NET0131  ;
	input \u0_uk_K_r13_reg[13]/NET0131  ;
	input \u0_uk_K_r13_reg[14]/NET0131  ;
	input \u0_uk_K_r13_reg[15]/NET0131  ;
	input \u0_uk_K_r13_reg[16]/NET0131  ;
	input \u0_uk_K_r13_reg[17]/NET0131  ;
	input \u0_uk_K_r13_reg[18]/NET0131  ;
	input \u0_uk_K_r13_reg[19]/NET0131  ;
	input \u0_uk_K_r13_reg[20]/NET0131  ;
	input \u0_uk_K_r13_reg[21]/NET0131  ;
	input \u0_uk_K_r13_reg[22]/NET0131  ;
	input \u0_uk_K_r13_reg[23]/NET0131  ;
	input \u0_uk_K_r13_reg[24]/NET0131  ;
	input \u0_uk_K_r13_reg[25]/P0001  ;
	input \u0_uk_K_r13_reg[26]/NET0131  ;
	input \u0_uk_K_r13_reg[27]/NET0131  ;
	input \u0_uk_K_r13_reg[28]/NET0131  ;
	input \u0_uk_K_r13_reg[29]/NET0131  ;
	input \u0_uk_K_r13_reg[2]/NET0131  ;
	input \u0_uk_K_r13_reg[30]/NET0131  ;
	input \u0_uk_K_r13_reg[31]/NET0131  ;
	input \u0_uk_K_r13_reg[32]/NET0131  ;
	input \u0_uk_K_r13_reg[33]/NET0131  ;
	input \u0_uk_K_r13_reg[34]/NET0131  ;
	input \u0_uk_K_r13_reg[35]/NET0131  ;
	input \u0_uk_K_r13_reg[36]/NET0131  ;
	input \u0_uk_K_r13_reg[37]/NET0131  ;
	input \u0_uk_K_r13_reg[38]/NET0131  ;
	input \u0_uk_K_r13_reg[39]/NET0131  ;
	input \u0_uk_K_r13_reg[3]/NET0131  ;
	input \u0_uk_K_r13_reg[40]/NET0131  ;
	input \u0_uk_K_r13_reg[41]/NET0131  ;
	input \u0_uk_K_r13_reg[42]/NET0131  ;
	input \u0_uk_K_r13_reg[43]/NET0131  ;
	input \u0_uk_K_r13_reg[44]/NET0131  ;
	input \u0_uk_K_r13_reg[45]/NET0131  ;
	input \u0_uk_K_r13_reg[46]/NET0131  ;
	input \u0_uk_K_r13_reg[47]/NET0131  ;
	input \u0_uk_K_r13_reg[48]/NET0131  ;
	input \u0_uk_K_r13_reg[49]/NET0131  ;
	input \u0_uk_K_r13_reg[4]/NET0131  ;
	input \u0_uk_K_r13_reg[50]/NET0131  ;
	input \u0_uk_K_r13_reg[51]/NET0131  ;
	input \u0_uk_K_r13_reg[52]/P0001  ;
	input \u0_uk_K_r13_reg[54]/NET0131  ;
	input \u0_uk_K_r13_reg[55]/NET0131  ;
	input \u0_uk_K_r13_reg[5]/NET0131  ;
	input \u0_uk_K_r13_reg[6]/NET0131  ;
	input \u0_uk_K_r13_reg[7]/NET0131  ;
	input \u0_uk_K_r13_reg[8]/NET0131  ;
	input \u0_uk_K_r13_reg[9]/NET0131  ;
	input \u0_uk_K_r14_reg[0]/NET0131  ;
	input \u0_uk_K_r14_reg[10]/P0001  ;
	input \u0_uk_K_r14_reg[11]/NET0131  ;
	input \u0_uk_K_r14_reg[12]/NET0131  ;
	input \u0_uk_K_r14_reg[13]/NET0131  ;
	input \u0_uk_K_r14_reg[14]/NET0131  ;
	input \u0_uk_K_r14_reg[15]/NET0131  ;
	input \u0_uk_K_r14_reg[16]/NET0131  ;
	input \u0_uk_K_r14_reg[17]/NET0131  ;
	input \u0_uk_K_r14_reg[18]/NET0131  ;
	input \u0_uk_K_r14_reg[19]/NET0131  ;
	input \u0_uk_K_r14_reg[1]/NET0131  ;
	input \u0_uk_K_r14_reg[20]/NET0131  ;
	input \u0_uk_K_r14_reg[21]/NET0131  ;
	input \u0_uk_K_r14_reg[22]/NET0131  ;
	input \u0_uk_K_r14_reg[23]/NET0131  ;
	input \u0_uk_K_r14_reg[24]/NET0131  ;
	input \u0_uk_K_r14_reg[25]/NET0131  ;
	input \u0_uk_K_r14_reg[26]/NET0131  ;
	input \u0_uk_K_r14_reg[27]/NET0131  ;
	input \u0_uk_K_r14_reg[28]/NET0131  ;
	input \u0_uk_K_r14_reg[29]/NET0131  ;
	input \u0_uk_K_r14_reg[2]/NET0131  ;
	input \u0_uk_K_r14_reg[30]/NET0131  ;
	input \u0_uk_K_r14_reg[31]/NET0131  ;
	input \u0_uk_K_r14_reg[32]/NET0131  ;
	input \u0_uk_K_r14_reg[33]/NET0131  ;
	input \u0_uk_K_r14_reg[34]/NET0131  ;
	input \u0_uk_K_r14_reg[35]/P0001  ;
	input \u0_uk_K_r14_reg[36]/NET0131  ;
	input \u0_uk_K_r14_reg[37]/NET0131  ;
	input \u0_uk_K_r14_reg[38]/NET0131  ;
	input \u0_uk_K_r14_reg[39]/P0001  ;
	input \u0_uk_K_r14_reg[3]/NET0131  ;
	input \u0_uk_K_r14_reg[40]/NET0131  ;
	input \u0_uk_K_r14_reg[41]/NET0131  ;
	input \u0_uk_K_r14_reg[42]/P0001  ;
	input \u0_uk_K_r14_reg[43]/NET0131  ;
	input \u0_uk_K_r14_reg[44]/NET0131  ;
	input \u0_uk_K_r14_reg[45]/NET0131  ;
	input \u0_uk_K_r14_reg[46]/NET0131  ;
	input \u0_uk_K_r14_reg[47]/NET0131  ;
	input \u0_uk_K_r14_reg[48]/NET0131  ;
	input \u0_uk_K_r14_reg[49]/NET0131  ;
	input \u0_uk_K_r14_reg[4]/NET0131  ;
	input \u0_uk_K_r14_reg[50]/NET0131  ;
	input \u0_uk_K_r14_reg[51]/NET0131  ;
	input \u0_uk_K_r14_reg[52]/NET0131  ;
	input \u0_uk_K_r14_reg[53]/NET0131  ;
	input \u0_uk_K_r14_reg[54]/NET0131  ;
	input \u0_uk_K_r14_reg[55]/NET0131  ;
	input \u0_uk_K_r14_reg[5]/NET0131  ;
	input \u0_uk_K_r14_reg[6]/NET0131  ;
	input \u0_uk_K_r14_reg[7]/NET0131  ;
	input \u0_uk_K_r14_reg[8]/NET0131  ;
	input \u0_uk_K_r14_reg[9]/NET0131  ;
	input \u0_uk_K_r1_reg[0]/NET0131  ;
	input \u0_uk_K_r1_reg[10]/P0001  ;
	input \u0_uk_K_r1_reg[11]/NET0131  ;
	input \u0_uk_K_r1_reg[12]/NET0131  ;
	input \u0_uk_K_r1_reg[13]/NET0131  ;
	input \u0_uk_K_r1_reg[14]/NET0131  ;
	input \u0_uk_K_r1_reg[15]/NET0131  ;
	input \u0_uk_K_r1_reg[16]/NET0131  ;
	input \u0_uk_K_r1_reg[17]/NET0131  ;
	input \u0_uk_K_r1_reg[18]/NET0131  ;
	input \u0_uk_K_r1_reg[19]/NET0131  ;
	input \u0_uk_K_r1_reg[1]/NET0131  ;
	input \u0_uk_K_r1_reg[20]/NET0131  ;
	input \u0_uk_K_r1_reg[21]/NET0131  ;
	input \u0_uk_K_r1_reg[22]/NET0131  ;
	input \u0_uk_K_r1_reg[23]/NET0131  ;
	input \u0_uk_K_r1_reg[24]/NET0131  ;
	input \u0_uk_K_r1_reg[25]/NET0131  ;
	input \u0_uk_K_r1_reg[26]/NET0131  ;
	input \u0_uk_K_r1_reg[27]/NET0131  ;
	input \u0_uk_K_r1_reg[28]/NET0131  ;
	input \u0_uk_K_r1_reg[29]/NET0131  ;
	input \u0_uk_K_r1_reg[2]/NET0131  ;
	input \u0_uk_K_r1_reg[30]/NET0131  ;
	input \u0_uk_K_r1_reg[31]/NET0131  ;
	input \u0_uk_K_r1_reg[32]/NET0131  ;
	input \u0_uk_K_r1_reg[33]/NET0131  ;
	input \u0_uk_K_r1_reg[34]/NET0131  ;
	input \u0_uk_K_r1_reg[35]/NET0131  ;
	input \u0_uk_K_r1_reg[36]/NET0131  ;
	input \u0_uk_K_r1_reg[37]/NET0131  ;
	input \u0_uk_K_r1_reg[38]/NET0131  ;
	input \u0_uk_K_r1_reg[3]/NET0131  ;
	input \u0_uk_K_r1_reg[40]/NET0131  ;
	input \u0_uk_K_r1_reg[41]/NET0131  ;
	input \u0_uk_K_r1_reg[42]/NET0131  ;
	input \u0_uk_K_r1_reg[43]/NET0131  ;
	input \u0_uk_K_r1_reg[44]/P0001  ;
	input \u0_uk_K_r1_reg[45]/NET0131  ;
	input \u0_uk_K_r1_reg[46]/NET0131  ;
	input \u0_uk_K_r1_reg[47]/NET0131  ;
	input \u0_uk_K_r1_reg[48]/NET0131  ;
	input \u0_uk_K_r1_reg[49]/NET0131  ;
	input \u0_uk_K_r1_reg[4]/NET0131  ;
	input \u0_uk_K_r1_reg[50]/NET0131  ;
	input \u0_uk_K_r1_reg[51]/NET0131  ;
	input \u0_uk_K_r1_reg[52]/NET0131  ;
	input \u0_uk_K_r1_reg[53]/NET0131  ;
	input \u0_uk_K_r1_reg[54]/NET0131  ;
	input \u0_uk_K_r1_reg[55]/NET0131  ;
	input \u0_uk_K_r1_reg[5]/NET0131  ;
	input \u0_uk_K_r1_reg[6]/NET0131  ;
	input \u0_uk_K_r1_reg[7]/P0001  ;
	input \u0_uk_K_r1_reg[8]/NET0131  ;
	input \u0_uk_K_r1_reg[9]/NET0131  ;
	input \u0_uk_K_r2_reg[0]/NET0131  ;
	input \u0_uk_K_r2_reg[10]/NET0131  ;
	input \u0_uk_K_r2_reg[11]/NET0131  ;
	input \u0_uk_K_r2_reg[12]/NET0131  ;
	input \u0_uk_K_r2_reg[13]/NET0131  ;
	input \u0_uk_K_r2_reg[14]/NET0131  ;
	input \u0_uk_K_r2_reg[15]/NET0131  ;
	input \u0_uk_K_r2_reg[16]/NET0131  ;
	input \u0_uk_K_r2_reg[17]/NET0131  ;
	input \u0_uk_K_r2_reg[18]/NET0131  ;
	input \u0_uk_K_r2_reg[19]/NET0131  ;
	input \u0_uk_K_r2_reg[1]/NET0131  ;
	input \u0_uk_K_r2_reg[20]/NET0131  ;
	input \u0_uk_K_r2_reg[21]/NET0131  ;
	input \u0_uk_K_r2_reg[22]/NET0131  ;
	input \u0_uk_K_r2_reg[23]/NET0131  ;
	input \u0_uk_K_r2_reg[24]/NET0131  ;
	input \u0_uk_K_r2_reg[25]/NET0131  ;
	input \u0_uk_K_r2_reg[26]/NET0131  ;
	input \u0_uk_K_r2_reg[27]/P0001  ;
	input \u0_uk_K_r2_reg[28]/NET0131  ;
	input \u0_uk_K_r2_reg[29]/NET0131  ;
	input \u0_uk_K_r2_reg[2]/NET0131  ;
	input \u0_uk_K_r2_reg[31]/NET0131  ;
	input \u0_uk_K_r2_reg[32]/NET0131  ;
	input \u0_uk_K_r2_reg[33]/NET0131  ;
	input \u0_uk_K_r2_reg[34]/NET0131  ;
	input \u0_uk_K_r2_reg[35]/NET0131  ;
	input \u0_uk_K_r2_reg[36]/NET0131  ;
	input \u0_uk_K_r2_reg[37]/NET0131  ;
	input \u0_uk_K_r2_reg[38]/NET0131  ;
	input \u0_uk_K_r2_reg[39]/NET0131  ;
	input \u0_uk_K_r2_reg[3]/NET0131  ;
	input \u0_uk_K_r2_reg[40]/NET0131  ;
	input \u0_uk_K_r2_reg[41]/NET0131  ;
	input \u0_uk_K_r2_reg[42]/NET0131  ;
	input \u0_uk_K_r2_reg[43]/NET0131  ;
	input \u0_uk_K_r2_reg[44]/NET0131  ;
	input \u0_uk_K_r2_reg[45]/NET0131  ;
	input \u0_uk_K_r2_reg[46]/NET0131  ;
	input \u0_uk_K_r2_reg[47]/NET0131  ;
	input \u0_uk_K_r2_reg[48]/NET0131  ;
	input \u0_uk_K_r2_reg[49]/NET0131  ;
	input \u0_uk_K_r2_reg[4]/NET0131  ;
	input \u0_uk_K_r2_reg[50]/NET0131  ;
	input \u0_uk_K_r2_reg[51]/NET0131  ;
	input \u0_uk_K_r2_reg[52]/NET0131  ;
	input \u0_uk_K_r2_reg[53]/P0001  ;
	input \u0_uk_K_r2_reg[54]/NET0131  ;
	input \u0_uk_K_r2_reg[55]/NET0131  ;
	input \u0_uk_K_r2_reg[5]/NET0131  ;
	input \u0_uk_K_r2_reg[6]/NET0131  ;
	input \u0_uk_K_r2_reg[7]/NET0131  ;
	input \u0_uk_K_r2_reg[8]/NET0131  ;
	input \u0_uk_K_r2_reg[9]/NET0131  ;
	input \u0_uk_K_r3_reg[0]/NET0131  ;
	input \u0_uk_K_r3_reg[10]/NET0131  ;
	input \u0_uk_K_r3_reg[11]/NET0131  ;
	input \u0_uk_K_r3_reg[12]/NET0131  ;
	input \u0_uk_K_r3_reg[14]/NET0131  ;
	input \u0_uk_K_r3_reg[15]/NET0131  ;
	input \u0_uk_K_r3_reg[16]/NET0131  ;
	input \u0_uk_K_r3_reg[17]/NET0131  ;
	input \u0_uk_K_r3_reg[18]/NET0131  ;
	input \u0_uk_K_r3_reg[19]/NET0131  ;
	input \u0_uk_K_r3_reg[1]/NET0131  ;
	input \u0_uk_K_r3_reg[20]/NET0131  ;
	input \u0_uk_K_r3_reg[21]/NET0131  ;
	input \u0_uk_K_r3_reg[22]/NET0131  ;
	input \u0_uk_K_r3_reg[23]/NET0131  ;
	input \u0_uk_K_r3_reg[24]/NET0131  ;
	input \u0_uk_K_r3_reg[25]/NET0131  ;
	input \u0_uk_K_r3_reg[26]/NET0131  ;
	input \u0_uk_K_r3_reg[27]/NET0131  ;
	input \u0_uk_K_r3_reg[28]/NET0131  ;
	input \u0_uk_K_r3_reg[29]/NET0131  ;
	input \u0_uk_K_r3_reg[2]/NET0131  ;
	input \u0_uk_K_r3_reg[30]/NET0131  ;
	input \u0_uk_K_r3_reg[31]/NET0131  ;
	input \u0_uk_K_r3_reg[32]/NET0131  ;
	input \u0_uk_K_r3_reg[33]/NET0131  ;
	input \u0_uk_K_r3_reg[34]/NET0131  ;
	input \u0_uk_K_r3_reg[35]/NET0131  ;
	input \u0_uk_K_r3_reg[36]/NET0131  ;
	input \u0_uk_K_r3_reg[37]/NET0131  ;
	input \u0_uk_K_r3_reg[38]/NET0131  ;
	input \u0_uk_K_r3_reg[39]/NET0131  ;
	input \u0_uk_K_r3_reg[3]/NET0131  ;
	input \u0_uk_K_r3_reg[40]/NET0131  ;
	input \u0_uk_K_r3_reg[41]/NET0131  ;
	input \u0_uk_K_r3_reg[42]/NET0131  ;
	input \u0_uk_K_r3_reg[43]/NET0131  ;
	input \u0_uk_K_r3_reg[44]/NET0131  ;
	input \u0_uk_K_r3_reg[45]/P0001  ;
	input \u0_uk_K_r3_reg[46]/NET0131  ;
	input \u0_uk_K_r3_reg[47]/NET0131  ;
	input \u0_uk_K_r3_reg[48]/NET0131  ;
	input \u0_uk_K_r3_reg[49]/NET0131  ;
	input \u0_uk_K_r3_reg[4]/NET0131  ;
	input \u0_uk_K_r3_reg[50]/NET0131  ;
	input \u0_uk_K_r3_reg[51]/NET0131  ;
	input \u0_uk_K_r3_reg[52]/NET0131  ;
	input \u0_uk_K_r3_reg[53]/NET0131  ;
	input \u0_uk_K_r3_reg[54]/NET0131  ;
	input \u0_uk_K_r3_reg[55]/NET0131  ;
	input \u0_uk_K_r3_reg[5]/NET0131  ;
	input \u0_uk_K_r3_reg[6]/NET0131  ;
	input \u0_uk_K_r3_reg[7]/NET0131  ;
	input \u0_uk_K_r3_reg[8]/NET0131  ;
	input \u0_uk_K_r3_reg[9]/NET0131  ;
	input \u0_uk_K_r4_reg[0]/P0001  ;
	input \u0_uk_K_r4_reg[10]/NET0131  ;
	input \u0_uk_K_r4_reg[11]/NET0131  ;
	input \u0_uk_K_r4_reg[12]/NET0131  ;
	input \u0_uk_K_r4_reg[13]/NET0131  ;
	input \u0_uk_K_r4_reg[14]/NET0131  ;
	input \u0_uk_K_r4_reg[15]/NET0131  ;
	input \u0_uk_K_r4_reg[16]/NET0131  ;
	input \u0_uk_K_r4_reg[17]/NET0131  ;
	input \u0_uk_K_r4_reg[18]/NET0131  ;
	input \u0_uk_K_r4_reg[19]/NET0131  ;
	input \u0_uk_K_r4_reg[1]/NET0131  ;
	input \u0_uk_K_r4_reg[20]/NET0131  ;
	input \u0_uk_K_r4_reg[21]/NET0131  ;
	input \u0_uk_K_r4_reg[22]/NET0131  ;
	input \u0_uk_K_r4_reg[23]/P0001  ;
	input \u0_uk_K_r4_reg[25]/NET0131  ;
	input \u0_uk_K_r4_reg[26]/NET0131  ;
	input \u0_uk_K_r4_reg[27]/P0001  ;
	input \u0_uk_K_r4_reg[28]/NET0131  ;
	input \u0_uk_K_r4_reg[29]/NET0131  ;
	input \u0_uk_K_r4_reg[30]/NET0131  ;
	input \u0_uk_K_r4_reg[31]/P0001  ;
	input \u0_uk_K_r4_reg[32]/NET0131  ;
	input \u0_uk_K_r4_reg[33]/NET0131  ;
	input \u0_uk_K_r4_reg[34]/NET0131  ;
	input \u0_uk_K_r4_reg[35]/NET0131  ;
	input \u0_uk_K_r4_reg[36]/NET0131  ;
	input \u0_uk_K_r4_reg[37]/NET0131  ;
	input \u0_uk_K_r4_reg[38]/NET0131  ;
	input \u0_uk_K_r4_reg[39]/NET0131  ;
	input \u0_uk_K_r4_reg[3]/NET0131  ;
	input \u0_uk_K_r4_reg[40]/NET0131  ;
	input \u0_uk_K_r4_reg[41]/NET0131  ;
	input \u0_uk_K_r4_reg[42]/NET0131  ;
	input \u0_uk_K_r4_reg[43]/NET0131  ;
	input \u0_uk_K_r4_reg[44]/NET0131  ;
	input \u0_uk_K_r4_reg[45]/NET0131  ;
	input \u0_uk_K_r4_reg[46]/NET0131  ;
	input \u0_uk_K_r4_reg[47]/NET0131  ;
	input \u0_uk_K_r4_reg[48]/NET0131  ;
	input \u0_uk_K_r4_reg[49]/NET0131  ;
	input \u0_uk_K_r4_reg[4]/NET0131  ;
	input \u0_uk_K_r4_reg[50]/NET0131  ;
	input \u0_uk_K_r4_reg[51]/NET0131  ;
	input \u0_uk_K_r4_reg[52]/NET0131  ;
	input \u0_uk_K_r4_reg[53]/NET0131  ;
	input \u0_uk_K_r4_reg[54]/NET0131  ;
	input \u0_uk_K_r4_reg[55]/NET0131  ;
	input \u0_uk_K_r4_reg[5]/NET0131  ;
	input \u0_uk_K_r4_reg[6]/NET0131  ;
	input \u0_uk_K_r4_reg[7]/NET0131  ;
	input \u0_uk_K_r4_reg[8]/NET0131  ;
	input \u0_uk_K_r4_reg[9]/NET0131  ;
	input \u0_uk_K_r5_reg[0]/NET0131  ;
	input \u0_uk_K_r5_reg[10]/NET0131  ;
	input \u0_uk_K_r5_reg[11]/NET0131  ;
	input \u0_uk_K_r5_reg[12]/NET0131  ;
	input \u0_uk_K_r5_reg[13]/P0001  ;
	input \u0_uk_K_r5_reg[14]/NET0131  ;
	input \u0_uk_K_r5_reg[15]/NET0131  ;
	input \u0_uk_K_r5_reg[16]/NET0131  ;
	input \u0_uk_K_r5_reg[17]/NET0131  ;
	input \u0_uk_K_r5_reg[18]/NET0131  ;
	input \u0_uk_K_r5_reg[19]/NET0131  ;
	input \u0_uk_K_r5_reg[1]/NET0131  ;
	input \u0_uk_K_r5_reg[20]/NET0131  ;
	input \u0_uk_K_r5_reg[21]/NET0131  ;
	input \u0_uk_K_r5_reg[22]/NET0131  ;
	input \u0_uk_K_r5_reg[23]/NET0131  ;
	input \u0_uk_K_r5_reg[24]/NET0131  ;
	input \u0_uk_K_r5_reg[25]/NET0131  ;
	input \u0_uk_K_r5_reg[26]/NET0131  ;
	input \u0_uk_K_r5_reg[27]/NET0131  ;
	input \u0_uk_K_r5_reg[28]/NET0131  ;
	input \u0_uk_K_r5_reg[29]/NET0131  ;
	input \u0_uk_K_r5_reg[2]/NET0131  ;
	input \u0_uk_K_r5_reg[30]/NET0131  ;
	input \u0_uk_K_r5_reg[31]/NET0131  ;
	input \u0_uk_K_r5_reg[32]/NET0131  ;
	input \u0_uk_K_r5_reg[33]/NET0131  ;
	input \u0_uk_K_r5_reg[34]/NET0131  ;
	input \u0_uk_K_r5_reg[35]/NET0131  ;
	input \u0_uk_K_r5_reg[36]/NET0131  ;
	input \u0_uk_K_r5_reg[37]/P0001  ;
	input \u0_uk_K_r5_reg[38]/NET0131  ;
	input \u0_uk_K_r5_reg[39]/NET0131  ;
	input \u0_uk_K_r5_reg[3]/NET0131  ;
	input \u0_uk_K_r5_reg[40]/NET0131  ;
	input \u0_uk_K_r5_reg[41]/NET0131  ;
	input \u0_uk_K_r5_reg[42]/NET0131  ;
	input \u0_uk_K_r5_reg[43]/NET0131  ;
	input \u0_uk_K_r5_reg[44]/NET0131  ;
	input \u0_uk_K_r5_reg[46]/NET0131  ;
	input \u0_uk_K_r5_reg[47]/NET0131  ;
	input \u0_uk_K_r5_reg[48]/NET0131  ;
	input \u0_uk_K_r5_reg[49]/NET0131  ;
	input \u0_uk_K_r5_reg[4]/NET0131  ;
	input \u0_uk_K_r5_reg[50]/NET0131  ;
	input \u0_uk_K_r5_reg[51]/NET0131  ;
	input \u0_uk_K_r5_reg[52]/NET0131  ;
	input \u0_uk_K_r5_reg[53]/NET0131  ;
	input \u0_uk_K_r5_reg[54]/NET0131  ;
	input \u0_uk_K_r5_reg[55]/NET0131  ;
	input \u0_uk_K_r5_reg[5]/NET0131  ;
	input \u0_uk_K_r5_reg[6]/NET0131  ;
	input \u0_uk_K_r5_reg[7]/NET0131  ;
	input \u0_uk_K_r5_reg[8]/NET0131  ;
	input \u0_uk_K_r5_reg[9]/NET0131  ;
	input \u0_uk_K_r6_reg[0]/NET0131  ;
	input \u0_uk_K_r6_reg[10]/NET0131  ;
	input \u0_uk_K_r6_reg[11]/NET0131  ;
	input \u0_uk_K_r6_reg[12]/NET0131  ;
	input \u0_uk_K_r6_reg[13]/NET0131  ;
	input \u0_uk_K_r6_reg[14]/NET0131  ;
	input \u0_uk_K_r6_reg[15]/NET0131  ;
	input \u0_uk_K_r6_reg[16]/NET0131  ;
	input \u0_uk_K_r6_reg[17]/NET0131  ;
	input \u0_uk_K_r6_reg[18]/NET0131  ;
	input \u0_uk_K_r6_reg[19]/NET0131  ;
	input \u0_uk_K_r6_reg[1]/NET0131  ;
	input \u0_uk_K_r6_reg[20]/NET0131  ;
	input \u0_uk_K_r6_reg[21]/NET0131  ;
	input \u0_uk_K_r6_reg[22]/NET0131  ;
	input \u0_uk_K_r6_reg[23]/P0001  ;
	input \u0_uk_K_r6_reg[24]/NET0131  ;
	input \u0_uk_K_r6_reg[25]/NET0131  ;
	input \u0_uk_K_r6_reg[26]/P0001  ;
	input \u0_uk_K_r6_reg[27]/NET0131  ;
	input \u0_uk_K_r6_reg[28]/NET0131  ;
	input \u0_uk_K_r6_reg[29]/NET0131  ;
	input \u0_uk_K_r6_reg[2]/NET0131  ;
	input \u0_uk_K_r6_reg[30]/P0001  ;
	input \u0_uk_K_r6_reg[31]/NET0131  ;
	input \u0_uk_K_r6_reg[32]/NET0131  ;
	input \u0_uk_K_r6_reg[33]/NET0131  ;
	input \u0_uk_K_r6_reg[34]/NET0131  ;
	input \u0_uk_K_r6_reg[35]/NET0131  ;
	input \u0_uk_K_r6_reg[36]/NET0131  ;
	input \u0_uk_K_r6_reg[37]/NET0131  ;
	input \u0_uk_K_r6_reg[38]/NET0131  ;
	input \u0_uk_K_r6_reg[39]/NET0131  ;
	input \u0_uk_K_r6_reg[3]/NET0131  ;
	input \u0_uk_K_r6_reg[40]/NET0131  ;
	input \u0_uk_K_r6_reg[41]/NET0131  ;
	input \u0_uk_K_r6_reg[42]/NET0131  ;
	input \u0_uk_K_r6_reg[43]/NET0131  ;
	input \u0_uk_K_r6_reg[44]/NET0131  ;
	input \u0_uk_K_r6_reg[45]/NET0131  ;
	input \u0_uk_K_r6_reg[46]/NET0131  ;
	input \u0_uk_K_r6_reg[47]/NET0131  ;
	input \u0_uk_K_r6_reg[48]/NET0131  ;
	input \u0_uk_K_r6_reg[49]/NET0131  ;
	input \u0_uk_K_r6_reg[4]/NET0131  ;
	input \u0_uk_K_r6_reg[50]/NET0131  ;
	input \u0_uk_K_r6_reg[51]/NET0131  ;
	input \u0_uk_K_r6_reg[52]/NET0131  ;
	input \u0_uk_K_r6_reg[53]/NET0131  ;
	input \u0_uk_K_r6_reg[54]/NET0131  ;
	input \u0_uk_K_r6_reg[55]/P0001  ;
	input \u0_uk_K_r6_reg[5]/NET0131  ;
	input \u0_uk_K_r6_reg[6]/NET0131  ;
	input \u0_uk_K_r6_reg[7]/NET0131  ;
	input \u0_uk_K_r6_reg[8]/NET0131  ;
	input \u0_uk_K_r6_reg[9]/NET0131  ;
	input \u0_uk_K_r7_reg[0]/NET0131  ;
	input \u0_uk_K_r7_reg[10]/NET0131  ;
	input \u0_uk_K_r7_reg[11]/NET0131  ;
	input \u0_uk_K_r7_reg[12]/NET0131  ;
	input \u0_uk_K_r7_reg[13]/NET0131  ;
	input \u0_uk_K_r7_reg[14]/NET0131  ;
	input \u0_uk_K_r7_reg[15]/NET0131  ;
	input \u0_uk_K_r7_reg[16]/NET0131  ;
	input \u0_uk_K_r7_reg[17]/NET0131  ;
	input \u0_uk_K_r7_reg[18]/NET0131  ;
	input \u0_uk_K_r7_reg[19]/NET0131  ;
	input \u0_uk_K_r7_reg[1]/NET0131  ;
	input \u0_uk_K_r7_reg[20]/NET0131  ;
	input \u0_uk_K_r7_reg[21]/NET0131  ;
	input \u0_uk_K_r7_reg[22]/NET0131  ;
	input \u0_uk_K_r7_reg[23]/P0001  ;
	input \u0_uk_K_r7_reg[24]/NET0131  ;
	input \u0_uk_K_r7_reg[25]/NET0131  ;
	input \u0_uk_K_r7_reg[26]/P0001  ;
	input \u0_uk_K_r7_reg[27]/NET0131  ;
	input \u0_uk_K_r7_reg[28]/NET0131  ;
	input \u0_uk_K_r7_reg[29]/NET0131  ;
	input \u0_uk_K_r7_reg[2]/NET0131  ;
	input \u0_uk_K_r7_reg[30]/P0001  ;
	input \u0_uk_K_r7_reg[31]/NET0131  ;
	input \u0_uk_K_r7_reg[32]/NET0131  ;
	input \u0_uk_K_r7_reg[33]/NET0131  ;
	input \u0_uk_K_r7_reg[34]/NET0131  ;
	input \u0_uk_K_r7_reg[35]/NET0131  ;
	input \u0_uk_K_r7_reg[36]/NET0131  ;
	input \u0_uk_K_r7_reg[37]/NET0131  ;
	input \u0_uk_K_r7_reg[38]/NET0131  ;
	input \u0_uk_K_r7_reg[39]/NET0131  ;
	input \u0_uk_K_r7_reg[3]/NET0131  ;
	input \u0_uk_K_r7_reg[40]/NET0131  ;
	input \u0_uk_K_r7_reg[41]/NET0131  ;
	input \u0_uk_K_r7_reg[42]/NET0131  ;
	input \u0_uk_K_r7_reg[43]/NET0131  ;
	input \u0_uk_K_r7_reg[44]/NET0131  ;
	input \u0_uk_K_r7_reg[45]/NET0131  ;
	input \u0_uk_K_r7_reg[46]/NET0131  ;
	input \u0_uk_K_r7_reg[47]/NET0131  ;
	input \u0_uk_K_r7_reg[48]/NET0131  ;
	input \u0_uk_K_r7_reg[49]/NET0131  ;
	input \u0_uk_K_r7_reg[4]/NET0131  ;
	input \u0_uk_K_r7_reg[50]/NET0131  ;
	input \u0_uk_K_r7_reg[51]/NET0131  ;
	input \u0_uk_K_r7_reg[52]/NET0131  ;
	input \u0_uk_K_r7_reg[53]/NET0131  ;
	input \u0_uk_K_r7_reg[54]/NET0131  ;
	input \u0_uk_K_r7_reg[55]/P0001  ;
	input \u0_uk_K_r7_reg[5]/NET0131  ;
	input \u0_uk_K_r7_reg[6]/NET0131  ;
	input \u0_uk_K_r7_reg[7]/NET0131  ;
	input \u0_uk_K_r7_reg[8]/NET0131  ;
	input \u0_uk_K_r7_reg[9]/NET0131  ;
	input \u0_uk_K_r8_reg[0]/NET0131  ;
	input \u0_uk_K_r8_reg[10]/NET0131  ;
	input \u0_uk_K_r8_reg[11]/NET0131  ;
	input \u0_uk_K_r8_reg[12]/NET0131  ;
	input \u0_uk_K_r8_reg[13]/P0001  ;
	input \u0_uk_K_r8_reg[14]/NET0131  ;
	input \u0_uk_K_r8_reg[15]/NET0131  ;
	input \u0_uk_K_r8_reg[16]/NET0131  ;
	input \u0_uk_K_r8_reg[17]/NET0131  ;
	input \u0_uk_K_r8_reg[18]/NET0131  ;
	input \u0_uk_K_r8_reg[19]/NET0131  ;
	input \u0_uk_K_r8_reg[1]/NET0131  ;
	input \u0_uk_K_r8_reg[20]/NET0131  ;
	input \u0_uk_K_r8_reg[21]/NET0131  ;
	input \u0_uk_K_r8_reg[22]/NET0131  ;
	input \u0_uk_K_r8_reg[23]/NET0131  ;
	input \u0_uk_K_r8_reg[24]/NET0131  ;
	input \u0_uk_K_r8_reg[25]/NET0131  ;
	input \u0_uk_K_r8_reg[26]/NET0131  ;
	input \u0_uk_K_r8_reg[27]/NET0131  ;
	input \u0_uk_K_r8_reg[28]/NET0131  ;
	input \u0_uk_K_r8_reg[29]/NET0131  ;
	input \u0_uk_K_r8_reg[2]/NET0131  ;
	input \u0_uk_K_r8_reg[30]/NET0131  ;
	input \u0_uk_K_r8_reg[31]/NET0131  ;
	input \u0_uk_K_r8_reg[32]/NET0131  ;
	input \u0_uk_K_r8_reg[33]/NET0131  ;
	input \u0_uk_K_r8_reg[34]/NET0131  ;
	input \u0_uk_K_r8_reg[35]/NET0131  ;
	input \u0_uk_K_r8_reg[36]/NET0131  ;
	input \u0_uk_K_r8_reg[37]/P0001  ;
	input \u0_uk_K_r8_reg[38]/NET0131  ;
	input \u0_uk_K_r8_reg[39]/NET0131  ;
	input \u0_uk_K_r8_reg[3]/NET0131  ;
	input \u0_uk_K_r8_reg[40]/NET0131  ;
	input \u0_uk_K_r8_reg[41]/NET0131  ;
	input \u0_uk_K_r8_reg[42]/NET0131  ;
	input \u0_uk_K_r8_reg[43]/NET0131  ;
	input \u0_uk_K_r8_reg[44]/NET0131  ;
	input \u0_uk_K_r8_reg[46]/NET0131  ;
	input \u0_uk_K_r8_reg[47]/NET0131  ;
	input \u0_uk_K_r8_reg[48]/NET0131  ;
	input \u0_uk_K_r8_reg[49]/NET0131  ;
	input \u0_uk_K_r8_reg[4]/NET0131  ;
	input \u0_uk_K_r8_reg[50]/NET0131  ;
	input \u0_uk_K_r8_reg[51]/NET0131  ;
	input \u0_uk_K_r8_reg[52]/NET0131  ;
	input \u0_uk_K_r8_reg[53]/NET0131  ;
	input \u0_uk_K_r8_reg[54]/NET0131  ;
	input \u0_uk_K_r8_reg[55]/NET0131  ;
	input \u0_uk_K_r8_reg[5]/NET0131  ;
	input \u0_uk_K_r8_reg[6]/NET0131  ;
	input \u0_uk_K_r8_reg[7]/NET0131  ;
	input \u0_uk_K_r8_reg[8]/NET0131  ;
	input \u0_uk_K_r8_reg[9]/P0001  ;
	input \u0_uk_K_r9_reg[0]/P0001  ;
	input \u0_uk_K_r9_reg[10]/NET0131  ;
	input \u0_uk_K_r9_reg[11]/NET0131  ;
	input \u0_uk_K_r9_reg[12]/NET0131  ;
	input \u0_uk_K_r9_reg[13]/NET0131  ;
	input \u0_uk_K_r9_reg[14]/NET0131  ;
	input \u0_uk_K_r9_reg[15]/NET0131  ;
	input \u0_uk_K_r9_reg[16]/NET0131  ;
	input \u0_uk_K_r9_reg[17]/NET0131  ;
	input \u0_uk_K_r9_reg[18]/NET0131  ;
	input \u0_uk_K_r9_reg[19]/NET0131  ;
	input \u0_uk_K_r9_reg[1]/NET0131  ;
	input \u0_uk_K_r9_reg[20]/NET0131  ;
	input \u0_uk_K_r9_reg[21]/NET0131  ;
	input \u0_uk_K_r9_reg[22]/NET0131  ;
	input \u0_uk_K_r9_reg[23]/P0001  ;
	input \u0_uk_K_r9_reg[25]/NET0131  ;
	input \u0_uk_K_r9_reg[26]/NET0131  ;
	input \u0_uk_K_r9_reg[27]/P0001  ;
	input \u0_uk_K_r9_reg[28]/NET0131  ;
	input \u0_uk_K_r9_reg[29]/NET0131  ;
	input \u0_uk_K_r9_reg[30]/NET0131  ;
	input \u0_uk_K_r9_reg[31]/P0001  ;
	input \u0_uk_K_r9_reg[32]/NET0131  ;
	input \u0_uk_K_r9_reg[33]/NET0131  ;
	input \u0_uk_K_r9_reg[34]/NET0131  ;
	input \u0_uk_K_r9_reg[35]/NET0131  ;
	input \u0_uk_K_r9_reg[36]/NET0131  ;
	input \u0_uk_K_r9_reg[37]/NET0131  ;
	input \u0_uk_K_r9_reg[38]/NET0131  ;
	input \u0_uk_K_r9_reg[39]/NET0131  ;
	input \u0_uk_K_r9_reg[3]/NET0131  ;
	input \u0_uk_K_r9_reg[40]/NET0131  ;
	input \u0_uk_K_r9_reg[41]/NET0131  ;
	input \u0_uk_K_r9_reg[42]/NET0131  ;
	input \u0_uk_K_r9_reg[43]/NET0131  ;
	input \u0_uk_K_r9_reg[44]/NET0131  ;
	input \u0_uk_K_r9_reg[45]/NET0131  ;
	input \u0_uk_K_r9_reg[46]/NET0131  ;
	input \u0_uk_K_r9_reg[47]/NET0131  ;
	input \u0_uk_K_r9_reg[48]/NET0131  ;
	input \u0_uk_K_r9_reg[49]/NET0131  ;
	input \u0_uk_K_r9_reg[4]/NET0131  ;
	input \u0_uk_K_r9_reg[50]/NET0131  ;
	input \u0_uk_K_r9_reg[51]/NET0131  ;
	input \u0_uk_K_r9_reg[52]/NET0131  ;
	input \u0_uk_K_r9_reg[53]/NET0131  ;
	input \u0_uk_K_r9_reg[54]/NET0131  ;
	input \u0_uk_K_r9_reg[55]/NET0131  ;
	input \u0_uk_K_r9_reg[5]/NET0131  ;
	input \u0_uk_K_r9_reg[6]/NET0131  ;
	input \u0_uk_K_r9_reg[7]/NET0131  ;
	input \u0_uk_K_r9_reg[8]/NET0131  ;
	input \u0_uk_K_r9_reg[9]/NET0131  ;
	input \u1_L0_reg[10]/NET0131  ;
	input \u1_L0_reg[11]/NET0131  ;
	input \u1_L0_reg[12]/NET0131  ;
	input \u1_L0_reg[13]/NET0131  ;
	input \u1_L0_reg[14]/NET0131  ;
	input \u1_L0_reg[15]/P0001  ;
	input \u1_L0_reg[16]/NET0131  ;
	input \u1_L0_reg[17]/NET0131  ;
	input \u1_L0_reg[18]/NET0131  ;
	input \u1_L0_reg[19]/NET0131  ;
	input \u1_L0_reg[1]/NET0131  ;
	input \u1_L0_reg[20]/NET0131  ;
	input \u1_L0_reg[21]/NET0131  ;
	input \u1_L0_reg[22]/NET0131  ;
	input \u1_L0_reg[23]/NET0131  ;
	input \u1_L0_reg[24]/NET0131  ;
	input \u1_L0_reg[25]/NET0131  ;
	input \u1_L0_reg[26]/NET0131  ;
	input \u1_L0_reg[27]/NET0131  ;
	input \u1_L0_reg[28]/NET0131  ;
	input \u1_L0_reg[29]/NET0131  ;
	input \u1_L0_reg[2]/NET0131  ;
	input \u1_L0_reg[30]/NET0131  ;
	input \u1_L0_reg[31]/NET0131  ;
	input \u1_L0_reg[32]/NET0131  ;
	input \u1_L0_reg[3]/NET0131  ;
	input \u1_L0_reg[4]/NET0131  ;
	input \u1_L0_reg[5]/NET0131  ;
	input \u1_L0_reg[6]/NET0131  ;
	input \u1_L0_reg[7]/NET0131  ;
	input \u1_L0_reg[8]/NET0131  ;
	input \u1_L0_reg[9]/NET0131  ;
	input \u1_L10_reg[10]/NET0131  ;
	input \u1_L10_reg[11]/NET0131  ;
	input \u1_L10_reg[12]/NET0131  ;
	input \u1_L10_reg[13]/NET0131  ;
	input \u1_L10_reg[14]/NET0131  ;
	input \u1_L10_reg[15]/P0001  ;
	input \u1_L10_reg[16]/NET0131  ;
	input \u1_L10_reg[17]/NET0131  ;
	input \u1_L10_reg[18]/P0001  ;
	input \u1_L10_reg[19]/P0001  ;
	input \u1_L10_reg[1]/NET0131  ;
	input \u1_L10_reg[20]/NET0131  ;
	input \u1_L10_reg[21]/NET0131  ;
	input \u1_L10_reg[22]/NET0131  ;
	input \u1_L10_reg[23]/NET0131  ;
	input \u1_L10_reg[24]/NET0131  ;
	input \u1_L10_reg[25]/NET0131  ;
	input \u1_L10_reg[26]/NET0131  ;
	input \u1_L10_reg[27]/NET0131  ;
	input \u1_L10_reg[28]/NET0131  ;
	input \u1_L10_reg[29]/NET0131  ;
	input \u1_L10_reg[2]/NET0131  ;
	input \u1_L10_reg[30]/NET0131  ;
	input \u1_L10_reg[31]/NET0131  ;
	input \u1_L10_reg[32]/NET0131  ;
	input \u1_L10_reg[3]/NET0131  ;
	input \u1_L10_reg[4]/NET0131  ;
	input \u1_L10_reg[5]/NET0131  ;
	input \u1_L10_reg[6]/NET0131  ;
	input \u1_L10_reg[7]/NET0131  ;
	input \u1_L10_reg[8]/NET0131  ;
	input \u1_L10_reg[9]/NET0131  ;
	input \u1_L11_reg[10]/NET0131  ;
	input \u1_L11_reg[11]/NET0131  ;
	input \u1_L11_reg[12]/NET0131  ;
	input \u1_L11_reg[13]/NET0131  ;
	input \u1_L11_reg[14]/NET0131  ;
	input \u1_L11_reg[15]/P0001  ;
	input \u1_L11_reg[16]/NET0131  ;
	input \u1_L11_reg[17]/NET0131  ;
	input \u1_L11_reg[18]/P0001  ;
	input \u1_L11_reg[19]/P0001  ;
	input \u1_L11_reg[1]/NET0131  ;
	input \u1_L11_reg[20]/NET0131  ;
	input \u1_L11_reg[21]/NET0131  ;
	input \u1_L11_reg[22]/NET0131  ;
	input \u1_L11_reg[23]/NET0131  ;
	input \u1_L11_reg[24]/NET0131  ;
	input \u1_L11_reg[25]/NET0131  ;
	input \u1_L11_reg[26]/NET0131  ;
	input \u1_L11_reg[27]/NET0131  ;
	input \u1_L11_reg[28]/NET0131  ;
	input \u1_L11_reg[29]/NET0131  ;
	input \u1_L11_reg[2]/NET0131  ;
	input \u1_L11_reg[30]/NET0131  ;
	input \u1_L11_reg[31]/NET0131  ;
	input \u1_L11_reg[32]/NET0131  ;
	input \u1_L11_reg[3]/NET0131  ;
	input \u1_L11_reg[4]/NET0131  ;
	input \u1_L11_reg[5]/NET0131  ;
	input \u1_L11_reg[6]/NET0131  ;
	input \u1_L11_reg[7]/NET0131  ;
	input \u1_L11_reg[8]/NET0131  ;
	input \u1_L11_reg[9]/NET0131  ;
	input \u1_L12_reg[10]/NET0131  ;
	input \u1_L12_reg[11]/NET0131  ;
	input \u1_L12_reg[12]/NET0131  ;
	input \u1_L12_reg[13]/NET0131  ;
	input \u1_L12_reg[14]/NET0131  ;
	input \u1_L12_reg[15]/P0001  ;
	input \u1_L12_reg[16]/NET0131  ;
	input \u1_L12_reg[17]/NET0131  ;
	input \u1_L12_reg[18]/P0001  ;
	input \u1_L12_reg[19]/NET0131  ;
	input \u1_L12_reg[1]/NET0131  ;
	input \u1_L12_reg[20]/NET0131  ;
	input \u1_L12_reg[21]/NET0131  ;
	input \u1_L12_reg[22]/NET0131  ;
	input \u1_L12_reg[23]/P0001  ;
	input \u1_L12_reg[24]/NET0131  ;
	input \u1_L12_reg[25]/NET0131  ;
	input \u1_L12_reg[26]/NET0131  ;
	input \u1_L12_reg[27]/NET0131  ;
	input \u1_L12_reg[28]/NET0131  ;
	input \u1_L12_reg[29]/NET0131  ;
	input \u1_L12_reg[2]/NET0131  ;
	input \u1_L12_reg[30]/NET0131  ;
	input \u1_L12_reg[31]/NET0131  ;
	input \u1_L12_reg[32]/NET0131  ;
	input \u1_L12_reg[3]/NET0131  ;
	input \u1_L12_reg[4]/NET0131  ;
	input \u1_L12_reg[5]/NET0131  ;
	input \u1_L12_reg[6]/NET0131  ;
	input \u1_L12_reg[7]/NET0131  ;
	input \u1_L12_reg[8]/NET0131  ;
	input \u1_L12_reg[9]/NET0131  ;
	input \u1_L13_reg[10]/NET0131  ;
	input \u1_L13_reg[11]/NET0131  ;
	input \u1_L13_reg[12]/NET0131  ;
	input \u1_L13_reg[13]/NET0131  ;
	input \u1_L13_reg[14]/NET0131  ;
	input \u1_L13_reg[15]/P0001  ;
	input \u1_L13_reg[16]/NET0131  ;
	input \u1_L13_reg[17]/NET0131  ;
	input \u1_L13_reg[18]/P0001  ;
	input \u1_L13_reg[19]/P0001  ;
	input \u1_L13_reg[1]/NET0131  ;
	input \u1_L13_reg[20]/NET0131  ;
	input \u1_L13_reg[21]/NET0131  ;
	input \u1_L13_reg[22]/NET0131  ;
	input \u1_L13_reg[23]/P0001  ;
	input \u1_L13_reg[24]/NET0131  ;
	input \u1_L13_reg[25]/NET0131  ;
	input \u1_L13_reg[26]/NET0131  ;
	input \u1_L13_reg[27]/NET0131  ;
	input \u1_L13_reg[28]/NET0131  ;
	input \u1_L13_reg[29]/NET0131  ;
	input \u1_L13_reg[2]/NET0131  ;
	input \u1_L13_reg[30]/NET0131  ;
	input \u1_L13_reg[31]/NET0131  ;
	input \u1_L13_reg[32]/NET0131  ;
	input \u1_L13_reg[3]/NET0131  ;
	input \u1_L13_reg[4]/NET0131  ;
	input \u1_L13_reg[5]/NET0131  ;
	input \u1_L13_reg[6]/NET0131  ;
	input \u1_L13_reg[7]/NET0131  ;
	input \u1_L13_reg[8]/NET0131  ;
	input \u1_L13_reg[9]/NET0131  ;
	input \u1_L14_reg[10]/P0001  ;
	input \u1_L14_reg[11]/P0001  ;
	input \u1_L14_reg[12]/P0001  ;
	input \u1_L14_reg[13]/P0001  ;
	input \u1_L14_reg[14]/P0001  ;
	input \u1_L14_reg[15]/P0001  ;
	input \u1_L14_reg[16]/P0001  ;
	input \u1_L14_reg[17]/P0001  ;
	input \u1_L14_reg[18]/P0001  ;
	input \u1_L14_reg[19]/P0001  ;
	input \u1_L14_reg[1]/P0001  ;
	input \u1_L14_reg[20]/P0001  ;
	input \u1_L14_reg[21]/P0001  ;
	input \u1_L14_reg[22]/P0001  ;
	input \u1_L14_reg[23]/P0001  ;
	input \u1_L14_reg[24]/P0001  ;
	input \u1_L14_reg[25]/P0001  ;
	input \u1_L14_reg[26]/P0001  ;
	input \u1_L14_reg[27]/P0001  ;
	input \u1_L14_reg[28]/P0001  ;
	input \u1_L14_reg[29]/P0001  ;
	input \u1_L14_reg[2]/P0001  ;
	input \u1_L14_reg[30]/P0001  ;
	input \u1_L14_reg[31]/P0001  ;
	input \u1_L14_reg[32]/P0001  ;
	input \u1_L14_reg[3]/P0001  ;
	input \u1_L14_reg[4]/P0001  ;
	input \u1_L14_reg[5]/P0001  ;
	input \u1_L14_reg[6]/P0001  ;
	input \u1_L14_reg[7]/P0001  ;
	input \u1_L14_reg[8]/P0001  ;
	input \u1_L14_reg[9]/P0001  ;
	input \u1_L1_reg[10]/NET0131  ;
	input \u1_L1_reg[11]/NET0131  ;
	input \u1_L1_reg[12]/NET0131  ;
	input \u1_L1_reg[13]/NET0131  ;
	input \u1_L1_reg[14]/NET0131  ;
	input \u1_L1_reg[15]/P0001  ;
	input \u1_L1_reg[16]/NET0131  ;
	input \u1_L1_reg[17]/NET0131  ;
	input \u1_L1_reg[18]/NET0131  ;
	input \u1_L1_reg[19]/P0001  ;
	input \u1_L1_reg[1]/NET0131  ;
	input \u1_L1_reg[20]/NET0131  ;
	input \u1_L1_reg[21]/NET0131  ;
	input \u1_L1_reg[22]/NET0131  ;
	input \u1_L1_reg[23]/NET0131  ;
	input \u1_L1_reg[24]/NET0131  ;
	input \u1_L1_reg[25]/NET0131  ;
	input \u1_L1_reg[26]/NET0131  ;
	input \u1_L1_reg[27]/NET0131  ;
	input \u1_L1_reg[28]/NET0131  ;
	input \u1_L1_reg[29]/NET0131  ;
	input \u1_L1_reg[2]/NET0131  ;
	input \u1_L1_reg[30]/NET0131  ;
	input \u1_L1_reg[31]/NET0131  ;
	input \u1_L1_reg[32]/NET0131  ;
	input \u1_L1_reg[3]/NET0131  ;
	input \u1_L1_reg[4]/NET0131  ;
	input \u1_L1_reg[5]/NET0131  ;
	input \u1_L1_reg[6]/NET0131  ;
	input \u1_L1_reg[7]/NET0131  ;
	input \u1_L1_reg[8]/NET0131  ;
	input \u1_L1_reg[9]/NET0131  ;
	input \u1_L2_reg[10]/NET0131  ;
	input \u1_L2_reg[11]/NET0131  ;
	input \u1_L2_reg[12]/NET0131  ;
	input \u1_L2_reg[13]/NET0131  ;
	input \u1_L2_reg[14]/NET0131  ;
	input \u1_L2_reg[15]/P0001  ;
	input \u1_L2_reg[16]/NET0131  ;
	input \u1_L2_reg[17]/NET0131  ;
	input \u1_L2_reg[18]/NET0131  ;
	input \u1_L2_reg[19]/NET0131  ;
	input \u1_L2_reg[1]/NET0131  ;
	input \u1_L2_reg[20]/NET0131  ;
	input \u1_L2_reg[21]/NET0131  ;
	input \u1_L2_reg[22]/NET0131  ;
	input \u1_L2_reg[23]/NET0131  ;
	input \u1_L2_reg[24]/NET0131  ;
	input \u1_L2_reg[25]/NET0131  ;
	input \u1_L2_reg[26]/NET0131  ;
	input \u1_L2_reg[27]/NET0131  ;
	input \u1_L2_reg[28]/NET0131  ;
	input \u1_L2_reg[29]/NET0131  ;
	input \u1_L2_reg[2]/NET0131  ;
	input \u1_L2_reg[30]/NET0131  ;
	input \u1_L2_reg[31]/NET0131  ;
	input \u1_L2_reg[32]/NET0131  ;
	input \u1_L2_reg[3]/NET0131  ;
	input \u1_L2_reg[4]/NET0131  ;
	input \u1_L2_reg[5]/NET0131  ;
	input \u1_L2_reg[6]/NET0131  ;
	input \u1_L2_reg[7]/NET0131  ;
	input \u1_L2_reg[8]/NET0131  ;
	input \u1_L2_reg[9]/NET0131  ;
	input \u1_L3_reg[10]/NET0131  ;
	input \u1_L3_reg[11]/NET0131  ;
	input \u1_L3_reg[12]/NET0131  ;
	input \u1_L3_reg[13]/NET0131  ;
	input \u1_L3_reg[14]/NET0131  ;
	input \u1_L3_reg[15]/P0001  ;
	input \u1_L3_reg[16]/NET0131  ;
	input \u1_L3_reg[17]/NET0131  ;
	input \u1_L3_reg[18]/NET0131  ;
	input \u1_L3_reg[19]/NET0131  ;
	input \u1_L3_reg[1]/NET0131  ;
	input \u1_L3_reg[20]/NET0131  ;
	input \u1_L3_reg[21]/NET0131  ;
	input \u1_L3_reg[22]/NET0131  ;
	input \u1_L3_reg[23]/NET0131  ;
	input \u1_L3_reg[24]/NET0131  ;
	input \u1_L3_reg[25]/NET0131  ;
	input \u1_L3_reg[26]/NET0131  ;
	input \u1_L3_reg[27]/NET0131  ;
	input \u1_L3_reg[28]/NET0131  ;
	input \u1_L3_reg[29]/NET0131  ;
	input \u1_L3_reg[2]/NET0131  ;
	input \u1_L3_reg[30]/NET0131  ;
	input \u1_L3_reg[31]/NET0131  ;
	input \u1_L3_reg[32]/NET0131  ;
	input \u1_L3_reg[3]/NET0131  ;
	input \u1_L3_reg[4]/NET0131  ;
	input \u1_L3_reg[5]/NET0131  ;
	input \u1_L3_reg[6]/NET0131  ;
	input \u1_L3_reg[7]/NET0131  ;
	input \u1_L3_reg[8]/NET0131  ;
	input \u1_L3_reg[9]/NET0131  ;
	input \u1_L4_reg[10]/NET0131  ;
	input \u1_L4_reg[11]/P0001  ;
	input \u1_L4_reg[12]/NET0131  ;
	input \u1_L4_reg[13]/NET0131  ;
	input \u1_L4_reg[14]/NET0131  ;
	input \u1_L4_reg[15]/P0001  ;
	input \u1_L4_reg[16]/NET0131  ;
	input \u1_L4_reg[17]/NET0131  ;
	input \u1_L4_reg[18]/NET0131  ;
	input \u1_L4_reg[19]/P0001  ;
	input \u1_L4_reg[1]/NET0131  ;
	input \u1_L4_reg[20]/NET0131  ;
	input \u1_L4_reg[21]/NET0131  ;
	input \u1_L4_reg[22]/NET0131  ;
	input \u1_L4_reg[23]/NET0131  ;
	input \u1_L4_reg[24]/NET0131  ;
	input \u1_L4_reg[25]/NET0131  ;
	input \u1_L4_reg[26]/NET0131  ;
	input \u1_L4_reg[27]/NET0131  ;
	input \u1_L4_reg[28]/NET0131  ;
	input \u1_L4_reg[29]/NET0131  ;
	input \u1_L4_reg[2]/NET0131  ;
	input \u1_L4_reg[30]/NET0131  ;
	input \u1_L4_reg[31]/NET0131  ;
	input \u1_L4_reg[32]/NET0131  ;
	input \u1_L4_reg[3]/NET0131  ;
	input \u1_L4_reg[4]/NET0131  ;
	input \u1_L4_reg[5]/NET0131  ;
	input \u1_L4_reg[6]/NET0131  ;
	input \u1_L4_reg[7]/NET0131  ;
	input \u1_L4_reg[8]/NET0131  ;
	input \u1_L4_reg[9]/NET0131  ;
	input \u1_L5_reg[10]/NET0131  ;
	input \u1_L5_reg[11]/NET0131  ;
	input \u1_L5_reg[12]/NET0131  ;
	input \u1_L5_reg[13]/NET0131  ;
	input \u1_L5_reg[14]/NET0131  ;
	input \u1_L5_reg[15]/P0001  ;
	input \u1_L5_reg[16]/NET0131  ;
	input \u1_L5_reg[17]/NET0131  ;
	input \u1_L5_reg[18]/NET0131  ;
	input \u1_L5_reg[19]/NET0131  ;
	input \u1_L5_reg[1]/NET0131  ;
	input \u1_L5_reg[20]/NET0131  ;
	input \u1_L5_reg[21]/NET0131  ;
	input \u1_L5_reg[22]/NET0131  ;
	input \u1_L5_reg[23]/NET0131  ;
	input \u1_L5_reg[24]/NET0131  ;
	input \u1_L5_reg[25]/NET0131  ;
	input \u1_L5_reg[26]/NET0131  ;
	input \u1_L5_reg[27]/NET0131  ;
	input \u1_L5_reg[28]/NET0131  ;
	input \u1_L5_reg[29]/NET0131  ;
	input \u1_L5_reg[2]/NET0131  ;
	input \u1_L5_reg[30]/NET0131  ;
	input \u1_L5_reg[31]/NET0131  ;
	input \u1_L5_reg[32]/NET0131  ;
	input \u1_L5_reg[3]/NET0131  ;
	input \u1_L5_reg[4]/NET0131  ;
	input \u1_L5_reg[5]/NET0131  ;
	input \u1_L5_reg[6]/NET0131  ;
	input \u1_L5_reg[7]/NET0131  ;
	input \u1_L5_reg[8]/NET0131  ;
	input \u1_L5_reg[9]/NET0131  ;
	input \u1_L6_reg[10]/NET0131  ;
	input \u1_L6_reg[11]/NET0131  ;
	input \u1_L6_reg[12]/NET0131  ;
	input \u1_L6_reg[13]/NET0131  ;
	input \u1_L6_reg[14]/NET0131  ;
	input \u1_L6_reg[15]/P0001  ;
	input \u1_L6_reg[16]/NET0131  ;
	input \u1_L6_reg[17]/NET0131  ;
	input \u1_L6_reg[18]/NET0131  ;
	input \u1_L6_reg[19]/NET0131  ;
	input \u1_L6_reg[1]/NET0131  ;
	input \u1_L6_reg[20]/NET0131  ;
	input \u1_L6_reg[21]/NET0131  ;
	input \u1_L6_reg[22]/NET0131  ;
	input \u1_L6_reg[23]/NET0131  ;
	input \u1_L6_reg[24]/NET0131  ;
	input \u1_L6_reg[25]/NET0131  ;
	input \u1_L6_reg[26]/NET0131  ;
	input \u1_L6_reg[27]/NET0131  ;
	input \u1_L6_reg[28]/NET0131  ;
	input \u1_L6_reg[29]/NET0131  ;
	input \u1_L6_reg[2]/NET0131  ;
	input \u1_L6_reg[30]/NET0131  ;
	input \u1_L6_reg[31]/NET0131  ;
	input \u1_L6_reg[32]/NET0131  ;
	input \u1_L6_reg[3]/NET0131  ;
	input \u1_L6_reg[4]/NET0131  ;
	input \u1_L6_reg[5]/NET0131  ;
	input \u1_L6_reg[6]/NET0131  ;
	input \u1_L6_reg[7]/NET0131  ;
	input \u1_L6_reg[8]/NET0131  ;
	input \u1_L6_reg[9]/NET0131  ;
	input \u1_L7_reg[10]/NET0131  ;
	input \u1_L7_reg[11]/NET0131  ;
	input \u1_L7_reg[12]/NET0131  ;
	input \u1_L7_reg[13]/NET0131  ;
	input \u1_L7_reg[14]/NET0131  ;
	input \u1_L7_reg[15]/P0001  ;
	input \u1_L7_reg[16]/NET0131  ;
	input \u1_L7_reg[17]/NET0131  ;
	input \u1_L7_reg[18]/NET0131  ;
	input \u1_L7_reg[19]/P0001  ;
	input \u1_L7_reg[1]/NET0131  ;
	input \u1_L7_reg[20]/NET0131  ;
	input \u1_L7_reg[21]/NET0131  ;
	input \u1_L7_reg[22]/NET0131  ;
	input \u1_L7_reg[23]/NET0131  ;
	input \u1_L7_reg[24]/NET0131  ;
	input \u1_L7_reg[25]/NET0131  ;
	input \u1_L7_reg[26]/NET0131  ;
	input \u1_L7_reg[27]/NET0131  ;
	input \u1_L7_reg[28]/NET0131  ;
	input \u1_L7_reg[29]/NET0131  ;
	input \u1_L7_reg[2]/NET0131  ;
	input \u1_L7_reg[30]/NET0131  ;
	input \u1_L7_reg[31]/NET0131  ;
	input \u1_L7_reg[32]/NET0131  ;
	input \u1_L7_reg[3]/NET0131  ;
	input \u1_L7_reg[4]/NET0131  ;
	input \u1_L7_reg[5]/NET0131  ;
	input \u1_L7_reg[6]/NET0131  ;
	input \u1_L7_reg[7]/NET0131  ;
	input \u1_L7_reg[8]/NET0131  ;
	input \u1_L7_reg[9]/NET0131  ;
	input \u1_L8_reg[10]/NET0131  ;
	input \u1_L8_reg[11]/NET0131  ;
	input \u1_L8_reg[12]/NET0131  ;
	input \u1_L8_reg[13]/NET0131  ;
	input \u1_L8_reg[14]/NET0131  ;
	input \u1_L8_reg[15]/P0001  ;
	input \u1_L8_reg[16]/NET0131  ;
	input \u1_L8_reg[17]/NET0131  ;
	input \u1_L8_reg[18]/NET0131  ;
	input \u1_L8_reg[19]/P0001  ;
	input \u1_L8_reg[1]/NET0131  ;
	input \u1_L8_reg[20]/NET0131  ;
	input \u1_L8_reg[21]/NET0131  ;
	input \u1_L8_reg[22]/NET0131  ;
	input \u1_L8_reg[23]/NET0131  ;
	input \u1_L8_reg[24]/NET0131  ;
	input \u1_L8_reg[25]/NET0131  ;
	input \u1_L8_reg[26]/NET0131  ;
	input \u1_L8_reg[27]/NET0131  ;
	input \u1_L8_reg[28]/NET0131  ;
	input \u1_L8_reg[29]/NET0131  ;
	input \u1_L8_reg[2]/NET0131  ;
	input \u1_L8_reg[30]/NET0131  ;
	input \u1_L8_reg[31]/NET0131  ;
	input \u1_L8_reg[32]/NET0131  ;
	input \u1_L8_reg[3]/NET0131  ;
	input \u1_L8_reg[4]/NET0131  ;
	input \u1_L8_reg[5]/NET0131  ;
	input \u1_L8_reg[6]/NET0131  ;
	input \u1_L8_reg[7]/NET0131  ;
	input \u1_L8_reg[8]/NET0131  ;
	input \u1_L8_reg[9]/NET0131  ;
	input \u1_L9_reg[10]/NET0131  ;
	input \u1_L9_reg[11]/NET0131  ;
	input \u1_L9_reg[12]/NET0131  ;
	input \u1_L9_reg[13]/NET0131  ;
	input \u1_L9_reg[14]/NET0131  ;
	input \u1_L9_reg[15]/P0001  ;
	input \u1_L9_reg[16]/NET0131  ;
	input \u1_L9_reg[17]/NET0131  ;
	input \u1_L9_reg[18]/P0001  ;
	input \u1_L9_reg[19]/NET0131  ;
	input \u1_L9_reg[1]/NET0131  ;
	input \u1_L9_reg[20]/NET0131  ;
	input \u1_L9_reg[21]/NET0131  ;
	input \u1_L9_reg[22]/NET0131  ;
	input \u1_L9_reg[23]/NET0131  ;
	input \u1_L9_reg[24]/NET0131  ;
	input \u1_L9_reg[25]/NET0131  ;
	input \u1_L9_reg[26]/NET0131  ;
	input \u1_L9_reg[27]/NET0131  ;
	input \u1_L9_reg[28]/NET0131  ;
	input \u1_L9_reg[29]/NET0131  ;
	input \u1_L9_reg[2]/NET0131  ;
	input \u1_L9_reg[30]/NET0131  ;
	input \u1_L9_reg[31]/NET0131  ;
	input \u1_L9_reg[32]/NET0131  ;
	input \u1_L9_reg[3]/NET0131  ;
	input \u1_L9_reg[4]/NET0131  ;
	input \u1_L9_reg[5]/NET0131  ;
	input \u1_L9_reg[6]/NET0131  ;
	input \u1_L9_reg[7]/NET0131  ;
	input \u1_L9_reg[8]/NET0131  ;
	input \u1_L9_reg[9]/NET0131  ;
	input \u1_R0_reg[10]/NET0131  ;
	input \u1_R0_reg[11]/NET0131  ;
	input \u1_R0_reg[12]/NET0131  ;
	input \u1_R0_reg[13]/NET0131  ;
	input \u1_R0_reg[14]/NET0131  ;
	input \u1_R0_reg[15]/NET0131  ;
	input \u1_R0_reg[16]/NET0131  ;
	input \u1_R0_reg[17]/NET0131  ;
	input \u1_R0_reg[18]/NET0131  ;
	input \u1_R0_reg[19]/NET0131  ;
	input \u1_R0_reg[1]/NET0131  ;
	input \u1_R0_reg[20]/NET0131  ;
	input \u1_R0_reg[21]/NET0131  ;
	input \u1_R0_reg[22]/NET0131  ;
	input \u1_R0_reg[23]/NET0131  ;
	input \u1_R0_reg[24]/NET0131  ;
	input \u1_R0_reg[25]/NET0131  ;
	input \u1_R0_reg[26]/NET0131  ;
	input \u1_R0_reg[27]/NET0131  ;
	input \u1_R0_reg[28]/NET0131  ;
	input \u1_R0_reg[29]/NET0131  ;
	input \u1_R0_reg[2]/NET0131  ;
	input \u1_R0_reg[30]/NET0131  ;
	input \u1_R0_reg[31]/P0001  ;
	input \u1_R0_reg[32]/NET0131  ;
	input \u1_R0_reg[3]/NET0131  ;
	input \u1_R0_reg[4]/NET0131  ;
	input \u1_R0_reg[5]/NET0131  ;
	input \u1_R0_reg[6]/NET0131  ;
	input \u1_R0_reg[7]/NET0131  ;
	input \u1_R0_reg[8]/NET0131  ;
	input \u1_R0_reg[9]/NET0131  ;
	input \u1_R10_reg[10]/NET0131  ;
	input \u1_R10_reg[11]/NET0131  ;
	input \u1_R10_reg[12]/NET0131  ;
	input \u1_R10_reg[13]/NET0131  ;
	input \u1_R10_reg[14]/NET0131  ;
	input \u1_R10_reg[15]/NET0131  ;
	input \u1_R10_reg[16]/NET0131  ;
	input \u1_R10_reg[17]/NET0131  ;
	input \u1_R10_reg[18]/NET0131  ;
	input \u1_R10_reg[19]/NET0131  ;
	input \u1_R10_reg[1]/NET0131  ;
	input \u1_R10_reg[20]/NET0131  ;
	input \u1_R10_reg[21]/NET0131  ;
	input \u1_R10_reg[22]/NET0131  ;
	input \u1_R10_reg[23]/NET0131  ;
	input \u1_R10_reg[24]/NET0131  ;
	input \u1_R10_reg[25]/NET0131  ;
	input \u1_R10_reg[26]/NET0131  ;
	input \u1_R10_reg[27]/NET0131  ;
	input \u1_R10_reg[28]/NET0131  ;
	input \u1_R10_reg[29]/NET0131  ;
	input \u1_R10_reg[2]/NET0131  ;
	input \u1_R10_reg[30]/NET0131  ;
	input \u1_R10_reg[31]/P0001  ;
	input \u1_R10_reg[32]/NET0131  ;
	input \u1_R10_reg[3]/NET0131  ;
	input \u1_R10_reg[4]/NET0131  ;
	input \u1_R10_reg[5]/NET0131  ;
	input \u1_R10_reg[6]/NET0131  ;
	input \u1_R10_reg[7]/NET0131  ;
	input \u1_R10_reg[8]/NET0131  ;
	input \u1_R10_reg[9]/NET0131  ;
	input \u1_R11_reg[10]/NET0131  ;
	input \u1_R11_reg[11]/NET0131  ;
	input \u1_R11_reg[12]/NET0131  ;
	input \u1_R11_reg[13]/NET0131  ;
	input \u1_R11_reg[14]/NET0131  ;
	input \u1_R11_reg[15]/NET0131  ;
	input \u1_R11_reg[16]/NET0131  ;
	input \u1_R11_reg[17]/NET0131  ;
	input \u1_R11_reg[18]/NET0131  ;
	input \u1_R11_reg[19]/NET0131  ;
	input \u1_R11_reg[1]/NET0131  ;
	input \u1_R11_reg[20]/NET0131  ;
	input \u1_R11_reg[21]/NET0131  ;
	input \u1_R11_reg[22]/NET0131  ;
	input \u1_R11_reg[23]/NET0131  ;
	input \u1_R11_reg[24]/NET0131  ;
	input \u1_R11_reg[25]/NET0131  ;
	input \u1_R11_reg[26]/NET0131  ;
	input \u1_R11_reg[27]/NET0131  ;
	input \u1_R11_reg[28]/NET0131  ;
	input \u1_R11_reg[29]/NET0131  ;
	input \u1_R11_reg[2]/NET0131  ;
	input \u1_R11_reg[30]/NET0131  ;
	input \u1_R11_reg[31]/NET0131  ;
	input \u1_R11_reg[32]/NET0131  ;
	input \u1_R11_reg[3]/NET0131  ;
	input \u1_R11_reg[4]/NET0131  ;
	input \u1_R11_reg[5]/NET0131  ;
	input \u1_R11_reg[6]/NET0131  ;
	input \u1_R11_reg[7]/NET0131  ;
	input \u1_R11_reg[8]/NET0131  ;
	input \u1_R11_reg[9]/NET0131  ;
	input \u1_R12_reg[10]/NET0131  ;
	input \u1_R12_reg[11]/NET0131  ;
	input \u1_R12_reg[12]/NET0131  ;
	input \u1_R12_reg[13]/NET0131  ;
	input \u1_R12_reg[14]/NET0131  ;
	input \u1_R12_reg[15]/NET0131  ;
	input \u1_R12_reg[16]/NET0131  ;
	input \u1_R12_reg[17]/NET0131  ;
	input \u1_R12_reg[18]/NET0131  ;
	input \u1_R12_reg[19]/NET0131  ;
	input \u1_R12_reg[1]/NET0131  ;
	input \u1_R12_reg[20]/NET0131  ;
	input \u1_R12_reg[21]/NET0131  ;
	input \u1_R12_reg[22]/NET0131  ;
	input \u1_R12_reg[23]/NET0131  ;
	input \u1_R12_reg[24]/NET0131  ;
	input \u1_R12_reg[25]/NET0131  ;
	input \u1_R12_reg[26]/NET0131  ;
	input \u1_R12_reg[27]/NET0131  ;
	input \u1_R12_reg[28]/NET0131  ;
	input \u1_R12_reg[29]/NET0131  ;
	input \u1_R12_reg[2]/NET0131  ;
	input \u1_R12_reg[30]/NET0131  ;
	input \u1_R12_reg[31]/NET0131  ;
	input \u1_R12_reg[32]/NET0131  ;
	input \u1_R12_reg[3]/NET0131  ;
	input \u1_R12_reg[4]/NET0131  ;
	input \u1_R12_reg[5]/NET0131  ;
	input \u1_R12_reg[6]/NET0131  ;
	input \u1_R12_reg[7]/NET0131  ;
	input \u1_R12_reg[8]/NET0131  ;
	input \u1_R12_reg[9]/NET0131  ;
	input \u1_R13_reg[10]/NET0131  ;
	input \u1_R13_reg[11]/P0001  ;
	input \u1_R13_reg[12]/NET0131  ;
	input \u1_R13_reg[13]/NET0131  ;
	input \u1_R13_reg[14]/NET0131  ;
	input \u1_R13_reg[15]/NET0131  ;
	input \u1_R13_reg[16]/NET0131  ;
	input \u1_R13_reg[17]/NET0131  ;
	input \u1_R13_reg[18]/NET0131  ;
	input \u1_R13_reg[19]/NET0131  ;
	input \u1_R13_reg[1]/NET0131  ;
	input \u1_R13_reg[20]/NET0131  ;
	input \u1_R13_reg[21]/NET0131  ;
	input \u1_R13_reg[22]/NET0131  ;
	input \u1_R13_reg[23]/P0001  ;
	input \u1_R13_reg[24]/NET0131  ;
	input \u1_R13_reg[25]/NET0131  ;
	input \u1_R13_reg[26]/NET0131  ;
	input \u1_R13_reg[27]/P0001  ;
	input \u1_R13_reg[28]/NET0131  ;
	input \u1_R13_reg[29]/NET0131  ;
	input \u1_R13_reg[2]/NET0131  ;
	input \u1_R13_reg[30]/NET0131  ;
	input \u1_R13_reg[31]/P0001  ;
	input \u1_R13_reg[32]/NET0131  ;
	input \u1_R13_reg[3]/NET0131  ;
	input \u1_R13_reg[4]/NET0131  ;
	input \u1_R13_reg[5]/NET0131  ;
	input \u1_R13_reg[6]/NET0131  ;
	input \u1_R13_reg[7]/NET0131  ;
	input \u1_R13_reg[8]/NET0131  ;
	input \u1_R13_reg[9]/NET0131  ;
	input \u1_R14_reg[10]/P0001  ;
	input \u1_R14_reg[11]/P0001  ;
	input \u1_R14_reg[12]/NET0131  ;
	input \u1_R14_reg[13]/NET0131  ;
	input \u1_R14_reg[14]/NET0131  ;
	input \u1_R14_reg[15]/NET0131  ;
	input \u1_R14_reg[16]/NET0131  ;
	input \u1_R14_reg[17]/NET0131  ;
	input \u1_R14_reg[18]/NET0131  ;
	input \u1_R14_reg[19]/P0001  ;
	input \u1_R14_reg[1]/NET0131  ;
	input \u1_R14_reg[20]/NET0131  ;
	input \u1_R14_reg[21]/NET0131  ;
	input \u1_R14_reg[22]/P0001  ;
	input \u1_R14_reg[23]/P0001  ;
	input \u1_R14_reg[24]/NET0131  ;
	input \u1_R14_reg[25]/NET0131  ;
	input \u1_R14_reg[26]/NET0131  ;
	input \u1_R14_reg[27]/P0001  ;
	input \u1_R14_reg[28]/NET0131  ;
	input \u1_R14_reg[29]/NET0131  ;
	input \u1_R14_reg[2]/NET0131  ;
	input \u1_R14_reg[30]/NET0131  ;
	input \u1_R14_reg[31]/P0001  ;
	input \u1_R14_reg[32]/NET0131  ;
	input \u1_R14_reg[3]/NET0131  ;
	input \u1_R14_reg[4]/NET0131  ;
	input \u1_R14_reg[5]/NET0131  ;
	input \u1_R14_reg[6]/NET0131  ;
	input \u1_R14_reg[7]/P0001  ;
	input \u1_R14_reg[8]/NET0131  ;
	input \u1_R14_reg[9]/NET0131  ;
	input \u1_R1_reg[10]/NET0131  ;
	input \u1_R1_reg[11]/NET0131  ;
	input \u1_R1_reg[12]/NET0131  ;
	input \u1_R1_reg[13]/NET0131  ;
	input \u1_R1_reg[14]/NET0131  ;
	input \u1_R1_reg[15]/NET0131  ;
	input \u1_R1_reg[16]/NET0131  ;
	input \u1_R1_reg[17]/NET0131  ;
	input \u1_R1_reg[18]/NET0131  ;
	input \u1_R1_reg[19]/NET0131  ;
	input \u1_R1_reg[1]/NET0131  ;
	input \u1_R1_reg[20]/NET0131  ;
	input \u1_R1_reg[21]/NET0131  ;
	input \u1_R1_reg[22]/NET0131  ;
	input \u1_R1_reg[23]/NET0131  ;
	input \u1_R1_reg[24]/NET0131  ;
	input \u1_R1_reg[25]/NET0131  ;
	input \u1_R1_reg[26]/NET0131  ;
	input \u1_R1_reg[27]/NET0131  ;
	input \u1_R1_reg[28]/NET0131  ;
	input \u1_R1_reg[29]/NET0131  ;
	input \u1_R1_reg[2]/NET0131  ;
	input \u1_R1_reg[30]/NET0131  ;
	input \u1_R1_reg[31]/P0001  ;
	input \u1_R1_reg[32]/NET0131  ;
	input \u1_R1_reg[3]/NET0131  ;
	input \u1_R1_reg[4]/NET0131  ;
	input \u1_R1_reg[5]/NET0131  ;
	input \u1_R1_reg[6]/NET0131  ;
	input \u1_R1_reg[7]/NET0131  ;
	input \u1_R1_reg[8]/NET0131  ;
	input \u1_R1_reg[9]/NET0131  ;
	input \u1_R2_reg[10]/NET0131  ;
	input \u1_R2_reg[11]/NET0131  ;
	input \u1_R2_reg[12]/NET0131  ;
	input \u1_R2_reg[13]/NET0131  ;
	input \u1_R2_reg[14]/NET0131  ;
	input \u1_R2_reg[15]/NET0131  ;
	input \u1_R2_reg[16]/NET0131  ;
	input \u1_R2_reg[17]/NET0131  ;
	input \u1_R2_reg[18]/NET0131  ;
	input \u1_R2_reg[19]/NET0131  ;
	input \u1_R2_reg[1]/NET0131  ;
	input \u1_R2_reg[20]/NET0131  ;
	input \u1_R2_reg[21]/NET0131  ;
	input \u1_R2_reg[22]/NET0131  ;
	input \u1_R2_reg[23]/NET0131  ;
	input \u1_R2_reg[24]/NET0131  ;
	input \u1_R2_reg[25]/NET0131  ;
	input \u1_R2_reg[26]/NET0131  ;
	input \u1_R2_reg[27]/NET0131  ;
	input \u1_R2_reg[28]/NET0131  ;
	input \u1_R2_reg[29]/NET0131  ;
	input \u1_R2_reg[2]/NET0131  ;
	input \u1_R2_reg[30]/NET0131  ;
	input \u1_R2_reg[31]/P0001  ;
	input \u1_R2_reg[32]/NET0131  ;
	input \u1_R2_reg[3]/NET0131  ;
	input \u1_R2_reg[4]/NET0131  ;
	input \u1_R2_reg[5]/NET0131  ;
	input \u1_R2_reg[6]/NET0131  ;
	input \u1_R2_reg[7]/NET0131  ;
	input \u1_R2_reg[8]/NET0131  ;
	input \u1_R2_reg[9]/NET0131  ;
	input \u1_R3_reg[10]/NET0131  ;
	input \u1_R3_reg[11]/NET0131  ;
	input \u1_R3_reg[12]/NET0131  ;
	input \u1_R3_reg[13]/NET0131  ;
	input \u1_R3_reg[14]/NET0131  ;
	input \u1_R3_reg[15]/NET0131  ;
	input \u1_R3_reg[16]/NET0131  ;
	input \u1_R3_reg[17]/NET0131  ;
	input \u1_R3_reg[18]/NET0131  ;
	input \u1_R3_reg[19]/NET0131  ;
	input \u1_R3_reg[1]/NET0131  ;
	input \u1_R3_reg[20]/NET0131  ;
	input \u1_R3_reg[21]/NET0131  ;
	input \u1_R3_reg[22]/NET0131  ;
	input \u1_R3_reg[23]/NET0131  ;
	input \u1_R3_reg[24]/NET0131  ;
	input \u1_R3_reg[25]/NET0131  ;
	input \u1_R3_reg[26]/NET0131  ;
	input \u1_R3_reg[27]/NET0131  ;
	input \u1_R3_reg[28]/NET0131  ;
	input \u1_R3_reg[29]/NET0131  ;
	input \u1_R3_reg[2]/NET0131  ;
	input \u1_R3_reg[30]/NET0131  ;
	input \u1_R3_reg[31]/P0001  ;
	input \u1_R3_reg[32]/NET0131  ;
	input \u1_R3_reg[3]/NET0131  ;
	input \u1_R3_reg[4]/NET0131  ;
	input \u1_R3_reg[5]/NET0131  ;
	input \u1_R3_reg[6]/NET0131  ;
	input \u1_R3_reg[7]/NET0131  ;
	input \u1_R3_reg[8]/NET0131  ;
	input \u1_R3_reg[9]/NET0131  ;
	input \u1_R4_reg[10]/NET0131  ;
	input \u1_R4_reg[11]/P0001  ;
	input \u1_R4_reg[12]/NET0131  ;
	input \u1_R4_reg[13]/NET0131  ;
	input \u1_R4_reg[14]/NET0131  ;
	input \u1_R4_reg[15]/NET0131  ;
	input \u1_R4_reg[16]/NET0131  ;
	input \u1_R4_reg[17]/NET0131  ;
	input \u1_R4_reg[18]/NET0131  ;
	input \u1_R4_reg[19]/NET0131  ;
	input \u1_R4_reg[1]/NET0131  ;
	input \u1_R4_reg[20]/NET0131  ;
	input \u1_R4_reg[21]/NET0131  ;
	input \u1_R4_reg[22]/NET0131  ;
	input \u1_R4_reg[23]/NET0131  ;
	input \u1_R4_reg[24]/NET0131  ;
	input \u1_R4_reg[25]/NET0131  ;
	input \u1_R4_reg[26]/NET0131  ;
	input \u1_R4_reg[27]/NET0131  ;
	input \u1_R4_reg[28]/NET0131  ;
	input \u1_R4_reg[29]/NET0131  ;
	input \u1_R4_reg[2]/NET0131  ;
	input \u1_R4_reg[30]/NET0131  ;
	input \u1_R4_reg[31]/P0001  ;
	input \u1_R4_reg[32]/NET0131  ;
	input \u1_R4_reg[3]/NET0131  ;
	input \u1_R4_reg[4]/NET0131  ;
	input \u1_R4_reg[5]/NET0131  ;
	input \u1_R4_reg[6]/NET0131  ;
	input \u1_R4_reg[7]/NET0131  ;
	input \u1_R4_reg[8]/NET0131  ;
	input \u1_R4_reg[9]/NET0131  ;
	input \u1_R5_reg[10]/NET0131  ;
	input \u1_R5_reg[11]/NET0131  ;
	input \u1_R5_reg[12]/NET0131  ;
	input \u1_R5_reg[13]/NET0131  ;
	input \u1_R5_reg[14]/NET0131  ;
	input \u1_R5_reg[15]/NET0131  ;
	input \u1_R5_reg[16]/NET0131  ;
	input \u1_R5_reg[17]/NET0131  ;
	input \u1_R5_reg[18]/NET0131  ;
	input \u1_R5_reg[19]/NET0131  ;
	input \u1_R5_reg[1]/NET0131  ;
	input \u1_R5_reg[20]/NET0131  ;
	input \u1_R5_reg[21]/NET0131  ;
	input \u1_R5_reg[22]/NET0131  ;
	input \u1_R5_reg[23]/NET0131  ;
	input \u1_R5_reg[24]/NET0131  ;
	input \u1_R5_reg[25]/NET0131  ;
	input \u1_R5_reg[26]/NET0131  ;
	input \u1_R5_reg[27]/NET0131  ;
	input \u1_R5_reg[28]/NET0131  ;
	input \u1_R5_reg[29]/NET0131  ;
	input \u1_R5_reg[2]/NET0131  ;
	input \u1_R5_reg[30]/NET0131  ;
	input \u1_R5_reg[31]/P0001  ;
	input \u1_R5_reg[32]/NET0131  ;
	input \u1_R5_reg[3]/NET0131  ;
	input \u1_R5_reg[4]/NET0131  ;
	input \u1_R5_reg[5]/NET0131  ;
	input \u1_R5_reg[6]/NET0131  ;
	input \u1_R5_reg[7]/NET0131  ;
	input \u1_R5_reg[8]/NET0131  ;
	input \u1_R5_reg[9]/NET0131  ;
	input \u1_R6_reg[10]/NET0131  ;
	input \u1_R6_reg[11]/NET0131  ;
	input \u1_R6_reg[12]/NET0131  ;
	input \u1_R6_reg[13]/NET0131  ;
	input \u1_R6_reg[14]/NET0131  ;
	input \u1_R6_reg[15]/NET0131  ;
	input \u1_R6_reg[16]/NET0131  ;
	input \u1_R6_reg[17]/NET0131  ;
	input \u1_R6_reg[18]/NET0131  ;
	input \u1_R6_reg[19]/NET0131  ;
	input \u1_R6_reg[1]/NET0131  ;
	input \u1_R6_reg[20]/NET0131  ;
	input \u1_R6_reg[21]/NET0131  ;
	input \u1_R6_reg[22]/NET0131  ;
	input \u1_R6_reg[23]/NET0131  ;
	input \u1_R6_reg[24]/NET0131  ;
	input \u1_R6_reg[25]/NET0131  ;
	input \u1_R6_reg[26]/NET0131  ;
	input \u1_R6_reg[27]/NET0131  ;
	input \u1_R6_reg[28]/NET0131  ;
	input \u1_R6_reg[29]/NET0131  ;
	input \u1_R6_reg[2]/NET0131  ;
	input \u1_R6_reg[30]/NET0131  ;
	input \u1_R6_reg[31]/P0001  ;
	input \u1_R6_reg[32]/NET0131  ;
	input \u1_R6_reg[3]/NET0131  ;
	input \u1_R6_reg[4]/NET0131  ;
	input \u1_R6_reg[5]/NET0131  ;
	input \u1_R6_reg[6]/NET0131  ;
	input \u1_R6_reg[7]/NET0131  ;
	input \u1_R6_reg[8]/NET0131  ;
	input \u1_R6_reg[9]/NET0131  ;
	input \u1_R7_reg[10]/NET0131  ;
	input \u1_R7_reg[11]/NET0131  ;
	input \u1_R7_reg[12]/NET0131  ;
	input \u1_R7_reg[13]/NET0131  ;
	input \u1_R7_reg[14]/NET0131  ;
	input \u1_R7_reg[15]/NET0131  ;
	input \u1_R7_reg[16]/NET0131  ;
	input \u1_R7_reg[17]/NET0131  ;
	input \u1_R7_reg[18]/NET0131  ;
	input \u1_R7_reg[19]/NET0131  ;
	input \u1_R7_reg[1]/NET0131  ;
	input \u1_R7_reg[20]/NET0131  ;
	input \u1_R7_reg[21]/NET0131  ;
	input \u1_R7_reg[22]/NET0131  ;
	input \u1_R7_reg[23]/NET0131  ;
	input \u1_R7_reg[24]/NET0131  ;
	input \u1_R7_reg[25]/NET0131  ;
	input \u1_R7_reg[26]/NET0131  ;
	input \u1_R7_reg[27]/NET0131  ;
	input \u1_R7_reg[28]/NET0131  ;
	input \u1_R7_reg[29]/NET0131  ;
	input \u1_R7_reg[2]/NET0131  ;
	input \u1_R7_reg[30]/NET0131  ;
	input \u1_R7_reg[31]/P0001  ;
	input \u1_R7_reg[32]/NET0131  ;
	input \u1_R7_reg[3]/NET0131  ;
	input \u1_R7_reg[4]/NET0131  ;
	input \u1_R7_reg[5]/NET0131  ;
	input \u1_R7_reg[6]/NET0131  ;
	input \u1_R7_reg[7]/NET0131  ;
	input \u1_R7_reg[8]/NET0131  ;
	input \u1_R7_reg[9]/NET0131  ;
	input \u1_R8_reg[10]/NET0131  ;
	input \u1_R8_reg[11]/NET0131  ;
	input \u1_R8_reg[12]/NET0131  ;
	input \u1_R8_reg[13]/NET0131  ;
	input \u1_R8_reg[14]/NET0131  ;
	input \u1_R8_reg[15]/NET0131  ;
	input \u1_R8_reg[16]/NET0131  ;
	input \u1_R8_reg[17]/NET0131  ;
	input \u1_R8_reg[18]/NET0131  ;
	input \u1_R8_reg[19]/NET0131  ;
	input \u1_R8_reg[1]/NET0131  ;
	input \u1_R8_reg[20]/NET0131  ;
	input \u1_R8_reg[21]/NET0131  ;
	input \u1_R8_reg[22]/NET0131  ;
	input \u1_R8_reg[23]/NET0131  ;
	input \u1_R8_reg[24]/NET0131  ;
	input \u1_R8_reg[25]/NET0131  ;
	input \u1_R8_reg[26]/NET0131  ;
	input \u1_R8_reg[27]/NET0131  ;
	input \u1_R8_reg[28]/NET0131  ;
	input \u1_R8_reg[29]/NET0131  ;
	input \u1_R8_reg[2]/NET0131  ;
	input \u1_R8_reg[30]/NET0131  ;
	input \u1_R8_reg[31]/P0001  ;
	input \u1_R8_reg[32]/NET0131  ;
	input \u1_R8_reg[3]/NET0131  ;
	input \u1_R8_reg[4]/NET0131  ;
	input \u1_R8_reg[5]/NET0131  ;
	input \u1_R8_reg[6]/NET0131  ;
	input \u1_R8_reg[7]/NET0131  ;
	input \u1_R8_reg[8]/NET0131  ;
	input \u1_R8_reg[9]/NET0131  ;
	input \u1_R9_reg[10]/NET0131  ;
	input \u1_R9_reg[11]/NET0131  ;
	input \u1_R9_reg[12]/NET0131  ;
	input \u1_R9_reg[13]/NET0131  ;
	input \u1_R9_reg[14]/NET0131  ;
	input \u1_R9_reg[15]/NET0131  ;
	input \u1_R9_reg[16]/NET0131  ;
	input \u1_R9_reg[17]/NET0131  ;
	input \u1_R9_reg[18]/NET0131  ;
	input \u1_R9_reg[19]/NET0131  ;
	input \u1_R9_reg[1]/NET0131  ;
	input \u1_R9_reg[20]/NET0131  ;
	input \u1_R9_reg[21]/NET0131  ;
	input \u1_R9_reg[22]/NET0131  ;
	input \u1_R9_reg[23]/NET0131  ;
	input \u1_R9_reg[24]/NET0131  ;
	input \u1_R9_reg[25]/NET0131  ;
	input \u1_R9_reg[26]/NET0131  ;
	input \u1_R9_reg[27]/NET0131  ;
	input \u1_R9_reg[28]/NET0131  ;
	input \u1_R9_reg[29]/NET0131  ;
	input \u1_R9_reg[2]/NET0131  ;
	input \u1_R9_reg[30]/NET0131  ;
	input \u1_R9_reg[31]/NET0131  ;
	input \u1_R9_reg[32]/NET0131  ;
	input \u1_R9_reg[3]/NET0131  ;
	input \u1_R9_reg[4]/NET0131  ;
	input \u1_R9_reg[5]/NET0131  ;
	input \u1_R9_reg[6]/NET0131  ;
	input \u1_R9_reg[7]/NET0131  ;
	input \u1_R9_reg[8]/NET0131  ;
	input \u1_R9_reg[9]/NET0131  ;
	input \u1_desIn_r_reg[0]/NET0131  ;
	input \u1_desIn_r_reg[10]/NET0131  ;
	input \u1_desIn_r_reg[11]/NET0131  ;
	input \u1_desIn_r_reg[12]/NET0131  ;
	input \u1_desIn_r_reg[13]/NET0131  ;
	input \u1_desIn_r_reg[14]/NET0131  ;
	input \u1_desIn_r_reg[15]/NET0131  ;
	input \u1_desIn_r_reg[16]/NET0131  ;
	input \u1_desIn_r_reg[17]/NET0131  ;
	input \u1_desIn_r_reg[18]/P0001  ;
	input \u1_desIn_r_reg[19]/NET0131  ;
	input \u1_desIn_r_reg[1]/NET0131  ;
	input \u1_desIn_r_reg[20]/NET0131  ;
	input \u1_desIn_r_reg[21]/NET0131  ;
	input \u1_desIn_r_reg[22]/NET0131  ;
	input \u1_desIn_r_reg[23]/NET0131  ;
	input \u1_desIn_r_reg[24]/NET0131  ;
	input \u1_desIn_r_reg[25]/NET0131  ;
	input \u1_desIn_r_reg[26]/NET0131  ;
	input \u1_desIn_r_reg[27]/NET0131  ;
	input \u1_desIn_r_reg[28]/NET0131  ;
	input \u1_desIn_r_reg[29]/NET0131  ;
	input \u1_desIn_r_reg[2]/NET0131  ;
	input \u1_desIn_r_reg[30]/NET0131  ;
	input \u1_desIn_r_reg[31]/NET0131  ;
	input \u1_desIn_r_reg[32]/NET0131  ;
	input \u1_desIn_r_reg[33]/NET0131  ;
	input \u1_desIn_r_reg[34]/NET0131  ;
	input \u1_desIn_r_reg[35]/NET0131  ;
	input \u1_desIn_r_reg[36]/NET0131  ;
	input \u1_desIn_r_reg[37]/NET0131  ;
	input \u1_desIn_r_reg[38]/NET0131  ;
	input \u1_desIn_r_reg[39]/NET0131  ;
	input \u1_desIn_r_reg[3]/NET0131  ;
	input \u1_desIn_r_reg[40]/NET0131  ;
	input \u1_desIn_r_reg[41]/NET0131  ;
	input \u1_desIn_r_reg[42]/NET0131  ;
	input \u1_desIn_r_reg[43]/NET0131  ;
	input \u1_desIn_r_reg[44]/NET0131  ;
	input \u1_desIn_r_reg[45]/NET0131  ;
	input \u1_desIn_r_reg[46]/NET0131  ;
	input \u1_desIn_r_reg[47]/NET0131  ;
	input \u1_desIn_r_reg[48]/NET0131  ;
	input \u1_desIn_r_reg[49]/NET0131  ;
	input \u1_desIn_r_reg[4]/NET0131  ;
	input \u1_desIn_r_reg[50]/NET0131  ;
	input \u1_desIn_r_reg[51]/NET0131  ;
	input \u1_desIn_r_reg[52]/P0001  ;
	input \u1_desIn_r_reg[53]/NET0131  ;
	input \u1_desIn_r_reg[54]/NET0131  ;
	input \u1_desIn_r_reg[55]/NET0131  ;
	input \u1_desIn_r_reg[56]/NET0131  ;
	input \u1_desIn_r_reg[57]/NET0131  ;
	input \u1_desIn_r_reg[58]/NET0131  ;
	input \u1_desIn_r_reg[59]/NET0131  ;
	input \u1_desIn_r_reg[5]/NET0131  ;
	input \u1_desIn_r_reg[60]/NET0131  ;
	input \u1_desIn_r_reg[61]/NET0131  ;
	input \u1_desIn_r_reg[62]/NET0131  ;
	input \u1_desIn_r_reg[63]/NET0131  ;
	input \u1_desIn_r_reg[6]/NET0131  ;
	input \u1_desIn_r_reg[7]/NET0131  ;
	input \u1_desIn_r_reg[8]/NET0131  ;
	input \u1_desIn_r_reg[9]/NET0131  ;
	input \u1_key_r_reg[0]/NET0131  ;
	input \u1_key_r_reg[10]/NET0131  ;
	input \u1_key_r_reg[11]/NET0131  ;
	input \u1_key_r_reg[12]/NET0131  ;
	input \u1_key_r_reg[13]/NET0131  ;
	input \u1_key_r_reg[14]/NET0131  ;
	input \u1_key_r_reg[15]/NET0131  ;
	input \u1_key_r_reg[16]/NET0131  ;
	input \u1_key_r_reg[17]/NET0131  ;
	input \u1_key_r_reg[18]/NET0131  ;
	input \u1_key_r_reg[19]/NET0131  ;
	input \u1_key_r_reg[1]/NET0131  ;
	input \u1_key_r_reg[20]/NET0131  ;
	input \u1_key_r_reg[21]/NET0131  ;
	input \u1_key_r_reg[22]/NET0131  ;
	input \u1_key_r_reg[23]/NET0131  ;
	input \u1_key_r_reg[24]/NET0131  ;
	input \u1_key_r_reg[25]/NET0131  ;
	input \u1_key_r_reg[26]/NET0131  ;
	input \u1_key_r_reg[27]/NET0131  ;
	input \u1_key_r_reg[28]/NET0131  ;
	input \u1_key_r_reg[29]/NET0131  ;
	input \u1_key_r_reg[2]/NET0131  ;
	input \u1_key_r_reg[30]/NET0131  ;
	input \u1_key_r_reg[31]/NET0131  ;
	input \u1_key_r_reg[32]/NET0131  ;
	input \u1_key_r_reg[33]/NET0131  ;
	input \u1_key_r_reg[34]/NET0131  ;
	input \u1_key_r_reg[35]/P0001  ;
	input \u1_key_r_reg[36]/NET0131  ;
	input \u1_key_r_reg[37]/NET0131  ;
	input \u1_key_r_reg[38]/NET0131  ;
	input \u1_key_r_reg[39]/P0001  ;
	input \u1_key_r_reg[3]/NET0131  ;
	input \u1_key_r_reg[40]/NET0131  ;
	input \u1_key_r_reg[41]/NET0131  ;
	input \u1_key_r_reg[42]/P0001  ;
	input \u1_key_r_reg[43]/NET0131  ;
	input \u1_key_r_reg[44]/NET0131  ;
	input \u1_key_r_reg[45]/NET0131  ;
	input \u1_key_r_reg[46]/NET0131  ;
	input \u1_key_r_reg[47]/NET0131  ;
	input \u1_key_r_reg[48]/NET0131  ;
	input \u1_key_r_reg[49]/NET0131  ;
	input \u1_key_r_reg[4]/NET0131  ;
	input \u1_key_r_reg[50]/NET0131  ;
	input \u1_key_r_reg[51]/NET0131  ;
	input \u1_key_r_reg[52]/NET0131  ;
	input \u1_key_r_reg[53]/NET0131  ;
	input \u1_key_r_reg[54]/NET0131  ;
	input \u1_key_r_reg[55]/NET0131  ;
	input \u1_key_r_reg[5]/NET0131  ;
	input \u1_key_r_reg[6]/NET0131  ;
	input \u1_key_r_reg[7]/NET0131  ;
	input \u1_key_r_reg[8]/NET0131  ;
	input \u1_key_r_reg[9]/NET0131  ;
	input \u1_uk_K_r0_reg[0]/NET0131  ;
	input \u1_uk_K_r0_reg[10]/NET0131  ;
	input \u1_uk_K_r0_reg[11]/NET0131  ;
	input \u1_uk_K_r0_reg[12]/NET0131  ;
	input \u1_uk_K_r0_reg[13]/NET0131  ;
	input \u1_uk_K_r0_reg[14]/NET0131  ;
	input \u1_uk_K_r0_reg[15]/NET0131  ;
	input \u1_uk_K_r0_reg[16]/NET0131  ;
	input \u1_uk_K_r0_reg[17]/NET0131  ;
	input \u1_uk_K_r0_reg[18]/NET0131  ;
	input \u1_uk_K_r0_reg[19]/NET0131  ;
	input \u1_uk_K_r0_reg[20]/NET0131  ;
	input \u1_uk_K_r0_reg[21]/NET0131  ;
	input \u1_uk_K_r0_reg[22]/NET0131  ;
	input \u1_uk_K_r0_reg[23]/NET0131  ;
	input \u1_uk_K_r0_reg[24]/NET0131  ;
	input \u1_uk_K_r0_reg[25]/P0001  ;
	input \u1_uk_K_r0_reg[26]/NET0131  ;
	input \u1_uk_K_r0_reg[27]/NET0131  ;
	input \u1_uk_K_r0_reg[28]/NET0131  ;
	input \u1_uk_K_r0_reg[29]/NET0131  ;
	input \u1_uk_K_r0_reg[2]/NET0131  ;
	input \u1_uk_K_r0_reg[30]/NET0131  ;
	input \u1_uk_K_r0_reg[31]/NET0131  ;
	input \u1_uk_K_r0_reg[32]/NET0131  ;
	input \u1_uk_K_r0_reg[33]/NET0131  ;
	input \u1_uk_K_r0_reg[34]/NET0131  ;
	input \u1_uk_K_r0_reg[35]/NET0131  ;
	input \u1_uk_K_r0_reg[36]/NET0131  ;
	input \u1_uk_K_r0_reg[37]/NET0131  ;
	input \u1_uk_K_r0_reg[38]/NET0131  ;
	input \u1_uk_K_r0_reg[39]/NET0131  ;
	input \u1_uk_K_r0_reg[3]/NET0131  ;
	input \u1_uk_K_r0_reg[40]/NET0131  ;
	input \u1_uk_K_r0_reg[41]/NET0131  ;
	input \u1_uk_K_r0_reg[42]/NET0131  ;
	input \u1_uk_K_r0_reg[43]/NET0131  ;
	input \u1_uk_K_r0_reg[44]/NET0131  ;
	input \u1_uk_K_r0_reg[45]/NET0131  ;
	input \u1_uk_K_r0_reg[46]/NET0131  ;
	input \u1_uk_K_r0_reg[47]/NET0131  ;
	input \u1_uk_K_r0_reg[48]/NET0131  ;
	input \u1_uk_K_r0_reg[49]/NET0131  ;
	input \u1_uk_K_r0_reg[4]/NET0131  ;
	input \u1_uk_K_r0_reg[50]/NET0131  ;
	input \u1_uk_K_r0_reg[51]/NET0131  ;
	input \u1_uk_K_r0_reg[52]/P0001  ;
	input \u1_uk_K_r0_reg[54]/NET0131  ;
	input \u1_uk_K_r0_reg[55]/NET0131  ;
	input \u1_uk_K_r0_reg[5]/NET0131  ;
	input \u1_uk_K_r0_reg[6]/NET0131  ;
	input \u1_uk_K_r0_reg[7]/NET0131  ;
	input \u1_uk_K_r0_reg[8]/NET0131  ;
	input \u1_uk_K_r0_reg[9]/NET0131  ;
	input \u1_uk_K_r10_reg[0]/NET0131  ;
	input \u1_uk_K_r10_reg[10]/NET0131  ;
	input \u1_uk_K_r10_reg[11]/NET0131  ;
	input \u1_uk_K_r10_reg[12]/NET0131  ;
	input \u1_uk_K_r10_reg[14]/NET0131  ;
	input \u1_uk_K_r10_reg[15]/NET0131  ;
	input \u1_uk_K_r10_reg[16]/NET0131  ;
	input \u1_uk_K_r10_reg[17]/NET0131  ;
	input \u1_uk_K_r10_reg[18]/NET0131  ;
	input \u1_uk_K_r10_reg[19]/NET0131  ;
	input \u1_uk_K_r10_reg[1]/NET0131  ;
	input \u1_uk_K_r10_reg[20]/NET0131  ;
	input \u1_uk_K_r10_reg[21]/NET0131  ;
	input \u1_uk_K_r10_reg[22]/NET0131  ;
	input \u1_uk_K_r10_reg[23]/NET0131  ;
	input \u1_uk_K_r10_reg[24]/NET0131  ;
	input \u1_uk_K_r10_reg[25]/NET0131  ;
	input \u1_uk_K_r10_reg[26]/NET0131  ;
	input \u1_uk_K_r10_reg[27]/NET0131  ;
	input \u1_uk_K_r10_reg[28]/NET0131  ;
	input \u1_uk_K_r10_reg[29]/NET0131  ;
	input \u1_uk_K_r10_reg[2]/NET0131  ;
	input \u1_uk_K_r10_reg[30]/NET0131  ;
	input \u1_uk_K_r10_reg[31]/NET0131  ;
	input \u1_uk_K_r10_reg[32]/NET0131  ;
	input \u1_uk_K_r10_reg[33]/NET0131  ;
	input \u1_uk_K_r10_reg[34]/NET0131  ;
	input \u1_uk_K_r10_reg[35]/NET0131  ;
	input \u1_uk_K_r10_reg[36]/NET0131  ;
	input \u1_uk_K_r10_reg[37]/NET0131  ;
	input \u1_uk_K_r10_reg[38]/NET0131  ;
	input \u1_uk_K_r10_reg[39]/NET0131  ;
	input \u1_uk_K_r10_reg[3]/NET0131  ;
	input \u1_uk_K_r10_reg[40]/NET0131  ;
	input \u1_uk_K_r10_reg[41]/P0001  ;
	input \u1_uk_K_r10_reg[42]/NET0131  ;
	input \u1_uk_K_r10_reg[43]/NET0131  ;
	input \u1_uk_K_r10_reg[44]/NET0131  ;
	input \u1_uk_K_r10_reg[45]/P0001  ;
	input \u1_uk_K_r10_reg[46]/NET0131  ;
	input \u1_uk_K_r10_reg[47]/NET0131  ;
	input \u1_uk_K_r10_reg[48]/NET0131  ;
	input \u1_uk_K_r10_reg[49]/NET0131  ;
	input \u1_uk_K_r10_reg[4]/NET0131  ;
	input \u1_uk_K_r10_reg[50]/NET0131  ;
	input \u1_uk_K_r10_reg[51]/NET0131  ;
	input \u1_uk_K_r10_reg[52]/NET0131  ;
	input \u1_uk_K_r10_reg[53]/NET0131  ;
	input \u1_uk_K_r10_reg[54]/NET0131  ;
	input \u1_uk_K_r10_reg[55]/NET0131  ;
	input \u1_uk_K_r10_reg[5]/NET0131  ;
	input \u1_uk_K_r10_reg[6]/NET0131  ;
	input \u1_uk_K_r10_reg[7]/NET0131  ;
	input \u1_uk_K_r10_reg[8]/NET0131  ;
	input \u1_uk_K_r10_reg[9]/NET0131  ;
	input \u1_uk_K_r11_reg[0]/NET0131  ;
	input \u1_uk_K_r11_reg[10]/NET0131  ;
	input \u1_uk_K_r11_reg[11]/NET0131  ;
	input \u1_uk_K_r11_reg[12]/NET0131  ;
	input \u1_uk_K_r11_reg[13]/NET0131  ;
	input \u1_uk_K_r11_reg[14]/NET0131  ;
	input \u1_uk_K_r11_reg[15]/NET0131  ;
	input \u1_uk_K_r11_reg[16]/NET0131  ;
	input \u1_uk_K_r11_reg[17]/NET0131  ;
	input \u1_uk_K_r11_reg[18]/NET0131  ;
	input \u1_uk_K_r11_reg[19]/NET0131  ;
	input \u1_uk_K_r11_reg[1]/NET0131  ;
	input \u1_uk_K_r11_reg[20]/NET0131  ;
	input \u1_uk_K_r11_reg[21]/NET0131  ;
	input \u1_uk_K_r11_reg[22]/NET0131  ;
	input \u1_uk_K_r11_reg[23]/NET0131  ;
	input \u1_uk_K_r11_reg[24]/NET0131  ;
	input \u1_uk_K_r11_reg[25]/NET0131  ;
	input \u1_uk_K_r11_reg[26]/NET0131  ;
	input \u1_uk_K_r11_reg[27]/P0001  ;
	input \u1_uk_K_r11_reg[28]/NET0131  ;
	input \u1_uk_K_r11_reg[29]/NET0131  ;
	input \u1_uk_K_r11_reg[2]/NET0131  ;
	input \u1_uk_K_r11_reg[31]/NET0131  ;
	input \u1_uk_K_r11_reg[32]/NET0131  ;
	input \u1_uk_K_r11_reg[33]/NET0131  ;
	input \u1_uk_K_r11_reg[34]/NET0131  ;
	input \u1_uk_K_r11_reg[35]/NET0131  ;
	input \u1_uk_K_r11_reg[36]/NET0131  ;
	input \u1_uk_K_r11_reg[37]/NET0131  ;
	input \u1_uk_K_r11_reg[38]/NET0131  ;
	input \u1_uk_K_r11_reg[39]/NET0131  ;
	input \u1_uk_K_r11_reg[3]/NET0131  ;
	input \u1_uk_K_r11_reg[40]/NET0131  ;
	input \u1_uk_K_r11_reg[41]/NET0131  ;
	input \u1_uk_K_r11_reg[42]/NET0131  ;
	input \u1_uk_K_r11_reg[43]/NET0131  ;
	input \u1_uk_K_r11_reg[44]/NET0131  ;
	input \u1_uk_K_r11_reg[45]/NET0131  ;
	input \u1_uk_K_r11_reg[46]/NET0131  ;
	input \u1_uk_K_r11_reg[47]/NET0131  ;
	input \u1_uk_K_r11_reg[48]/NET0131  ;
	input \u1_uk_K_r11_reg[49]/NET0131  ;
	input \u1_uk_K_r11_reg[4]/NET0131  ;
	input \u1_uk_K_r11_reg[50]/NET0131  ;
	input \u1_uk_K_r11_reg[51]/NET0131  ;
	input \u1_uk_K_r11_reg[52]/NET0131  ;
	input \u1_uk_K_r11_reg[53]/P0001  ;
	input \u1_uk_K_r11_reg[54]/NET0131  ;
	input \u1_uk_K_r11_reg[55]/NET0131  ;
	input \u1_uk_K_r11_reg[5]/NET0131  ;
	input \u1_uk_K_r11_reg[6]/NET0131  ;
	input \u1_uk_K_r11_reg[7]/NET0131  ;
	input \u1_uk_K_r11_reg[8]/NET0131  ;
	input \u1_uk_K_r11_reg[9]/NET0131  ;
	input \u1_uk_K_r12_reg[0]/NET0131  ;
	input \u1_uk_K_r12_reg[10]/P0001  ;
	input \u1_uk_K_r12_reg[11]/NET0131  ;
	input \u1_uk_K_r12_reg[12]/NET0131  ;
	input \u1_uk_K_r12_reg[13]/NET0131  ;
	input \u1_uk_K_r12_reg[14]/NET0131  ;
	input \u1_uk_K_r12_reg[15]/NET0131  ;
	input \u1_uk_K_r12_reg[16]/NET0131  ;
	input \u1_uk_K_r12_reg[17]/NET0131  ;
	input \u1_uk_K_r12_reg[18]/NET0131  ;
	input \u1_uk_K_r12_reg[19]/NET0131  ;
	input \u1_uk_K_r12_reg[1]/NET0131  ;
	input \u1_uk_K_r12_reg[20]/NET0131  ;
	input \u1_uk_K_r12_reg[21]/NET0131  ;
	input \u1_uk_K_r12_reg[22]/NET0131  ;
	input \u1_uk_K_r12_reg[23]/NET0131  ;
	input \u1_uk_K_r12_reg[24]/NET0131  ;
	input \u1_uk_K_r12_reg[25]/NET0131  ;
	input \u1_uk_K_r12_reg[26]/NET0131  ;
	input \u1_uk_K_r12_reg[27]/NET0131  ;
	input \u1_uk_K_r12_reg[28]/NET0131  ;
	input \u1_uk_K_r12_reg[29]/NET0131  ;
	input \u1_uk_K_r12_reg[2]/NET0131  ;
	input \u1_uk_K_r12_reg[30]/NET0131  ;
	input \u1_uk_K_r12_reg[31]/NET0131  ;
	input \u1_uk_K_r12_reg[32]/NET0131  ;
	input \u1_uk_K_r12_reg[33]/NET0131  ;
	input \u1_uk_K_r12_reg[34]/NET0131  ;
	input \u1_uk_K_r12_reg[35]/NET0131  ;
	input \u1_uk_K_r12_reg[36]/NET0131  ;
	input \u1_uk_K_r12_reg[37]/NET0131  ;
	input \u1_uk_K_r12_reg[38]/NET0131  ;
	input \u1_uk_K_r12_reg[3]/NET0131  ;
	input \u1_uk_K_r12_reg[40]/NET0131  ;
	input \u1_uk_K_r12_reg[41]/NET0131  ;
	input \u1_uk_K_r12_reg[42]/NET0131  ;
	input \u1_uk_K_r12_reg[43]/NET0131  ;
	input \u1_uk_K_r12_reg[44]/P0001  ;
	input \u1_uk_K_r12_reg[45]/NET0131  ;
	input \u1_uk_K_r12_reg[46]/NET0131  ;
	input \u1_uk_K_r12_reg[47]/NET0131  ;
	input \u1_uk_K_r12_reg[48]/NET0131  ;
	input \u1_uk_K_r12_reg[49]/NET0131  ;
	input \u1_uk_K_r12_reg[4]/NET0131  ;
	input \u1_uk_K_r12_reg[50]/NET0131  ;
	input \u1_uk_K_r12_reg[51]/NET0131  ;
	input \u1_uk_K_r12_reg[52]/NET0131  ;
	input \u1_uk_K_r12_reg[53]/NET0131  ;
	input \u1_uk_K_r12_reg[54]/NET0131  ;
	input \u1_uk_K_r12_reg[55]/NET0131  ;
	input \u1_uk_K_r12_reg[5]/NET0131  ;
	input \u1_uk_K_r12_reg[6]/NET0131  ;
	input \u1_uk_K_r12_reg[7]/P0001  ;
	input \u1_uk_K_r12_reg[8]/NET0131  ;
	input \u1_uk_K_r12_reg[9]/NET0131  ;
	input \u1_uk_K_r13_reg[0]/NET0131  ;
	input \u1_uk_K_r13_reg[10]/NET0131  ;
	input \u1_uk_K_r13_reg[11]/NET0131  ;
	input \u1_uk_K_r13_reg[12]/NET0131  ;
	input \u1_uk_K_r13_reg[13]/NET0131  ;
	input \u1_uk_K_r13_reg[14]/NET0131  ;
	input \u1_uk_K_r13_reg[15]/NET0131  ;
	input \u1_uk_K_r13_reg[16]/NET0131  ;
	input \u1_uk_K_r13_reg[17]/NET0131  ;
	input \u1_uk_K_r13_reg[18]/NET0131  ;
	input \u1_uk_K_r13_reg[19]/NET0131  ;
	input \u1_uk_K_r13_reg[20]/NET0131  ;
	input \u1_uk_K_r13_reg[21]/NET0131  ;
	input \u1_uk_K_r13_reg[22]/NET0131  ;
	input \u1_uk_K_r13_reg[23]/NET0131  ;
	input \u1_uk_K_r13_reg[24]/NET0131  ;
	input \u1_uk_K_r13_reg[25]/P0001  ;
	input \u1_uk_K_r13_reg[26]/NET0131  ;
	input \u1_uk_K_r13_reg[27]/NET0131  ;
	input \u1_uk_K_r13_reg[28]/NET0131  ;
	input \u1_uk_K_r13_reg[29]/NET0131  ;
	input \u1_uk_K_r13_reg[2]/NET0131  ;
	input \u1_uk_K_r13_reg[30]/NET0131  ;
	input \u1_uk_K_r13_reg[31]/NET0131  ;
	input \u1_uk_K_r13_reg[32]/NET0131  ;
	input \u1_uk_K_r13_reg[33]/NET0131  ;
	input \u1_uk_K_r13_reg[34]/NET0131  ;
	input \u1_uk_K_r13_reg[35]/NET0131  ;
	input \u1_uk_K_r13_reg[36]/NET0131  ;
	input \u1_uk_K_r13_reg[37]/NET0131  ;
	input \u1_uk_K_r13_reg[38]/NET0131  ;
	input \u1_uk_K_r13_reg[39]/NET0131  ;
	input \u1_uk_K_r13_reg[3]/NET0131  ;
	input \u1_uk_K_r13_reg[40]/NET0131  ;
	input \u1_uk_K_r13_reg[41]/NET0131  ;
	input \u1_uk_K_r13_reg[42]/NET0131  ;
	input \u1_uk_K_r13_reg[43]/NET0131  ;
	input \u1_uk_K_r13_reg[44]/NET0131  ;
	input \u1_uk_K_r13_reg[45]/NET0131  ;
	input \u1_uk_K_r13_reg[46]/NET0131  ;
	input \u1_uk_K_r13_reg[47]/NET0131  ;
	input \u1_uk_K_r13_reg[48]/NET0131  ;
	input \u1_uk_K_r13_reg[49]/NET0131  ;
	input \u1_uk_K_r13_reg[4]/NET0131  ;
	input \u1_uk_K_r13_reg[50]/NET0131  ;
	input \u1_uk_K_r13_reg[51]/NET0131  ;
	input \u1_uk_K_r13_reg[52]/P0001  ;
	input \u1_uk_K_r13_reg[54]/NET0131  ;
	input \u1_uk_K_r13_reg[55]/NET0131  ;
	input \u1_uk_K_r13_reg[5]/NET0131  ;
	input \u1_uk_K_r13_reg[6]/NET0131  ;
	input \u1_uk_K_r13_reg[7]/NET0131  ;
	input \u1_uk_K_r13_reg[8]/NET0131  ;
	input \u1_uk_K_r13_reg[9]/NET0131  ;
	input \u1_uk_K_r14_reg[0]/P0001  ;
	input \u1_uk_K_r14_reg[10]/P0001  ;
	input \u1_uk_K_r14_reg[11]/NET0131  ;
	input \u1_uk_K_r14_reg[12]/NET0131  ;
	input \u1_uk_K_r14_reg[13]/NET0131  ;
	input \u1_uk_K_r14_reg[14]/NET0131  ;
	input \u1_uk_K_r14_reg[15]/NET0131  ;
	input \u1_uk_K_r14_reg[16]/NET0131  ;
	input \u1_uk_K_r14_reg[17]/NET0131  ;
	input \u1_uk_K_r14_reg[18]/NET0131  ;
	input \u1_uk_K_r14_reg[19]/NET0131  ;
	input \u1_uk_K_r14_reg[1]/NET0131  ;
	input \u1_uk_K_r14_reg[20]/NET0131  ;
	input \u1_uk_K_r14_reg[21]/NET0131  ;
	input \u1_uk_K_r14_reg[22]/NET0131  ;
	input \u1_uk_K_r14_reg[23]/NET0131  ;
	input \u1_uk_K_r14_reg[24]/NET0131  ;
	input \u1_uk_K_r14_reg[25]/NET0131  ;
	input \u1_uk_K_r14_reg[26]/NET0131  ;
	input \u1_uk_K_r14_reg[27]/NET0131  ;
	input \u1_uk_K_r14_reg[28]/NET0131  ;
	input \u1_uk_K_r14_reg[29]/NET0131  ;
	input \u1_uk_K_r14_reg[2]/NET0131  ;
	input \u1_uk_K_r14_reg[30]/NET0131  ;
	input \u1_uk_K_r14_reg[31]/NET0131  ;
	input \u1_uk_K_r14_reg[32]/NET0131  ;
	input \u1_uk_K_r14_reg[33]/NET0131  ;
	input \u1_uk_K_r14_reg[34]/NET0131  ;
	input \u1_uk_K_r14_reg[35]/P0001  ;
	input \u1_uk_K_r14_reg[36]/NET0131  ;
	input \u1_uk_K_r14_reg[37]/NET0131  ;
	input \u1_uk_K_r14_reg[38]/NET0131  ;
	input \u1_uk_K_r14_reg[39]/P0001  ;
	input \u1_uk_K_r14_reg[3]/NET0131  ;
	input \u1_uk_K_r14_reg[40]/NET0131  ;
	input \u1_uk_K_r14_reg[41]/NET0131  ;
	input \u1_uk_K_r14_reg[42]/P0001  ;
	input \u1_uk_K_r14_reg[43]/NET0131  ;
	input \u1_uk_K_r14_reg[44]/NET0131  ;
	input \u1_uk_K_r14_reg[45]/NET0131  ;
	input \u1_uk_K_r14_reg[46]/NET0131  ;
	input \u1_uk_K_r14_reg[47]/NET0131  ;
	input \u1_uk_K_r14_reg[48]/NET0131  ;
	input \u1_uk_K_r14_reg[49]/NET0131  ;
	input \u1_uk_K_r14_reg[4]/NET0131  ;
	input \u1_uk_K_r14_reg[50]/NET0131  ;
	input \u1_uk_K_r14_reg[51]/NET0131  ;
	input \u1_uk_K_r14_reg[52]/NET0131  ;
	input \u1_uk_K_r14_reg[53]/NET0131  ;
	input \u1_uk_K_r14_reg[54]/NET0131  ;
	input \u1_uk_K_r14_reg[55]/NET0131  ;
	input \u1_uk_K_r14_reg[5]/NET0131  ;
	input \u1_uk_K_r14_reg[6]/NET0131  ;
	input \u1_uk_K_r14_reg[7]/NET0131  ;
	input \u1_uk_K_r14_reg[8]/P0001  ;
	input \u1_uk_K_r14_reg[9]/NET0131  ;
	input \u1_uk_K_r1_reg[0]/NET0131  ;
	input \u1_uk_K_r1_reg[10]/P0001  ;
	input \u1_uk_K_r1_reg[11]/NET0131  ;
	input \u1_uk_K_r1_reg[12]/NET0131  ;
	input \u1_uk_K_r1_reg[13]/NET0131  ;
	input \u1_uk_K_r1_reg[14]/NET0131  ;
	input \u1_uk_K_r1_reg[15]/NET0131  ;
	input \u1_uk_K_r1_reg[16]/NET0131  ;
	input \u1_uk_K_r1_reg[17]/NET0131  ;
	input \u1_uk_K_r1_reg[18]/NET0131  ;
	input \u1_uk_K_r1_reg[19]/NET0131  ;
	input \u1_uk_K_r1_reg[1]/NET0131  ;
	input \u1_uk_K_r1_reg[20]/NET0131  ;
	input \u1_uk_K_r1_reg[21]/NET0131  ;
	input \u1_uk_K_r1_reg[22]/NET0131  ;
	input \u1_uk_K_r1_reg[23]/NET0131  ;
	input \u1_uk_K_r1_reg[24]/NET0131  ;
	input \u1_uk_K_r1_reg[25]/NET0131  ;
	input \u1_uk_K_r1_reg[26]/NET0131  ;
	input \u1_uk_K_r1_reg[27]/NET0131  ;
	input \u1_uk_K_r1_reg[28]/NET0131  ;
	input \u1_uk_K_r1_reg[29]/NET0131  ;
	input \u1_uk_K_r1_reg[2]/NET0131  ;
	input \u1_uk_K_r1_reg[30]/NET0131  ;
	input \u1_uk_K_r1_reg[31]/NET0131  ;
	input \u1_uk_K_r1_reg[32]/NET0131  ;
	input \u1_uk_K_r1_reg[33]/NET0131  ;
	input \u1_uk_K_r1_reg[34]/NET0131  ;
	input \u1_uk_K_r1_reg[35]/NET0131  ;
	input \u1_uk_K_r1_reg[36]/NET0131  ;
	input \u1_uk_K_r1_reg[37]/NET0131  ;
	input \u1_uk_K_r1_reg[38]/NET0131  ;
	input \u1_uk_K_r1_reg[3]/NET0131  ;
	input \u1_uk_K_r1_reg[40]/NET0131  ;
	input \u1_uk_K_r1_reg[41]/NET0131  ;
	input \u1_uk_K_r1_reg[42]/NET0131  ;
	input \u1_uk_K_r1_reg[43]/NET0131  ;
	input \u1_uk_K_r1_reg[44]/P0001  ;
	input \u1_uk_K_r1_reg[45]/NET0131  ;
	input \u1_uk_K_r1_reg[46]/NET0131  ;
	input \u1_uk_K_r1_reg[47]/NET0131  ;
	input \u1_uk_K_r1_reg[48]/NET0131  ;
	input \u1_uk_K_r1_reg[49]/NET0131  ;
	input \u1_uk_K_r1_reg[4]/NET0131  ;
	input \u1_uk_K_r1_reg[50]/NET0131  ;
	input \u1_uk_K_r1_reg[51]/NET0131  ;
	input \u1_uk_K_r1_reg[52]/NET0131  ;
	input \u1_uk_K_r1_reg[53]/NET0131  ;
	input \u1_uk_K_r1_reg[54]/NET0131  ;
	input \u1_uk_K_r1_reg[55]/NET0131  ;
	input \u1_uk_K_r1_reg[5]/NET0131  ;
	input \u1_uk_K_r1_reg[6]/NET0131  ;
	input \u1_uk_K_r1_reg[7]/P0001  ;
	input \u1_uk_K_r1_reg[8]/NET0131  ;
	input \u1_uk_K_r1_reg[9]/NET0131  ;
	input \u1_uk_K_r2_reg[0]/NET0131  ;
	input \u1_uk_K_r2_reg[10]/NET0131  ;
	input \u1_uk_K_r2_reg[11]/NET0131  ;
	input \u1_uk_K_r2_reg[12]/NET0131  ;
	input \u1_uk_K_r2_reg[13]/NET0131  ;
	input \u1_uk_K_r2_reg[14]/NET0131  ;
	input \u1_uk_K_r2_reg[15]/NET0131  ;
	input \u1_uk_K_r2_reg[16]/NET0131  ;
	input \u1_uk_K_r2_reg[17]/NET0131  ;
	input \u1_uk_K_r2_reg[18]/NET0131  ;
	input \u1_uk_K_r2_reg[19]/NET0131  ;
	input \u1_uk_K_r2_reg[1]/NET0131  ;
	input \u1_uk_K_r2_reg[20]/NET0131  ;
	input \u1_uk_K_r2_reg[21]/NET0131  ;
	input \u1_uk_K_r2_reg[22]/NET0131  ;
	input \u1_uk_K_r2_reg[23]/NET0131  ;
	input \u1_uk_K_r2_reg[24]/NET0131  ;
	input \u1_uk_K_r2_reg[25]/NET0131  ;
	input \u1_uk_K_r2_reg[26]/NET0131  ;
	input \u1_uk_K_r2_reg[27]/NET0131  ;
	input \u1_uk_K_r2_reg[28]/NET0131  ;
	input \u1_uk_K_r2_reg[29]/NET0131  ;
	input \u1_uk_K_r2_reg[2]/NET0131  ;
	input \u1_uk_K_r2_reg[31]/NET0131  ;
	input \u1_uk_K_r2_reg[32]/NET0131  ;
	input \u1_uk_K_r2_reg[33]/NET0131  ;
	input \u1_uk_K_r2_reg[34]/NET0131  ;
	input \u1_uk_K_r2_reg[35]/NET0131  ;
	input \u1_uk_K_r2_reg[36]/NET0131  ;
	input \u1_uk_K_r2_reg[37]/NET0131  ;
	input \u1_uk_K_r2_reg[38]/NET0131  ;
	input \u1_uk_K_r2_reg[39]/NET0131  ;
	input \u1_uk_K_r2_reg[3]/NET0131  ;
	input \u1_uk_K_r2_reg[40]/NET0131  ;
	input \u1_uk_K_r2_reg[41]/NET0131  ;
	input \u1_uk_K_r2_reg[42]/NET0131  ;
	input \u1_uk_K_r2_reg[43]/NET0131  ;
	input \u1_uk_K_r2_reg[44]/NET0131  ;
	input \u1_uk_K_r2_reg[45]/NET0131  ;
	input \u1_uk_K_r2_reg[46]/NET0131  ;
	input \u1_uk_K_r2_reg[47]/NET0131  ;
	input \u1_uk_K_r2_reg[48]/NET0131  ;
	input \u1_uk_K_r2_reg[49]/NET0131  ;
	input \u1_uk_K_r2_reg[4]/NET0131  ;
	input \u1_uk_K_r2_reg[50]/NET0131  ;
	input \u1_uk_K_r2_reg[51]/NET0131  ;
	input \u1_uk_K_r2_reg[52]/NET0131  ;
	input \u1_uk_K_r2_reg[53]/P0001  ;
	input \u1_uk_K_r2_reg[54]/NET0131  ;
	input \u1_uk_K_r2_reg[55]/NET0131  ;
	input \u1_uk_K_r2_reg[5]/NET0131  ;
	input \u1_uk_K_r2_reg[6]/NET0131  ;
	input \u1_uk_K_r2_reg[7]/NET0131  ;
	input \u1_uk_K_r2_reg[8]/NET0131  ;
	input \u1_uk_K_r2_reg[9]/NET0131  ;
	input \u1_uk_K_r3_reg[0]/NET0131  ;
	input \u1_uk_K_r3_reg[10]/NET0131  ;
	input \u1_uk_K_r3_reg[11]/NET0131  ;
	input \u1_uk_K_r3_reg[12]/NET0131  ;
	input \u1_uk_K_r3_reg[14]/NET0131  ;
	input \u1_uk_K_r3_reg[15]/NET0131  ;
	input \u1_uk_K_r3_reg[16]/NET0131  ;
	input \u1_uk_K_r3_reg[17]/NET0131  ;
	input \u1_uk_K_r3_reg[18]/NET0131  ;
	input \u1_uk_K_r3_reg[19]/NET0131  ;
	input \u1_uk_K_r3_reg[1]/NET0131  ;
	input \u1_uk_K_r3_reg[20]/NET0131  ;
	input \u1_uk_K_r3_reg[21]/NET0131  ;
	input \u1_uk_K_r3_reg[22]/NET0131  ;
	input \u1_uk_K_r3_reg[23]/NET0131  ;
	input \u1_uk_K_r3_reg[24]/NET0131  ;
	input \u1_uk_K_r3_reg[25]/NET0131  ;
	input \u1_uk_K_r3_reg[26]/NET0131  ;
	input \u1_uk_K_r3_reg[27]/NET0131  ;
	input \u1_uk_K_r3_reg[28]/NET0131  ;
	input \u1_uk_K_r3_reg[29]/NET0131  ;
	input \u1_uk_K_r3_reg[2]/NET0131  ;
	input \u1_uk_K_r3_reg[30]/NET0131  ;
	input \u1_uk_K_r3_reg[31]/NET0131  ;
	input \u1_uk_K_r3_reg[32]/NET0131  ;
	input \u1_uk_K_r3_reg[33]/NET0131  ;
	input \u1_uk_K_r3_reg[34]/NET0131  ;
	input \u1_uk_K_r3_reg[35]/NET0131  ;
	input \u1_uk_K_r3_reg[36]/NET0131  ;
	input \u1_uk_K_r3_reg[37]/NET0131  ;
	input \u1_uk_K_r3_reg[38]/NET0131  ;
	input \u1_uk_K_r3_reg[39]/NET0131  ;
	input \u1_uk_K_r3_reg[3]/NET0131  ;
	input \u1_uk_K_r3_reg[40]/NET0131  ;
	input \u1_uk_K_r3_reg[41]/NET0131  ;
	input \u1_uk_K_r3_reg[42]/NET0131  ;
	input \u1_uk_K_r3_reg[43]/NET0131  ;
	input \u1_uk_K_r3_reg[44]/NET0131  ;
	input \u1_uk_K_r3_reg[45]/NET0131  ;
	input \u1_uk_K_r3_reg[46]/NET0131  ;
	input \u1_uk_K_r3_reg[47]/NET0131  ;
	input \u1_uk_K_r3_reg[48]/NET0131  ;
	input \u1_uk_K_r3_reg[49]/NET0131  ;
	input \u1_uk_K_r3_reg[4]/NET0131  ;
	input \u1_uk_K_r3_reg[50]/NET0131  ;
	input \u1_uk_K_r3_reg[51]/NET0131  ;
	input \u1_uk_K_r3_reg[52]/NET0131  ;
	input \u1_uk_K_r3_reg[53]/NET0131  ;
	input \u1_uk_K_r3_reg[54]/NET0131  ;
	input \u1_uk_K_r3_reg[55]/NET0131  ;
	input \u1_uk_K_r3_reg[5]/NET0131  ;
	input \u1_uk_K_r3_reg[6]/NET0131  ;
	input \u1_uk_K_r3_reg[7]/NET0131  ;
	input \u1_uk_K_r3_reg[8]/NET0131  ;
	input \u1_uk_K_r3_reg[9]/NET0131  ;
	input \u1_uk_K_r4_reg[0]/P0001  ;
	input \u1_uk_K_r4_reg[10]/NET0131  ;
	input \u1_uk_K_r4_reg[11]/NET0131  ;
	input \u1_uk_K_r4_reg[12]/NET0131  ;
	input \u1_uk_K_r4_reg[13]/NET0131  ;
	input \u1_uk_K_r4_reg[14]/NET0131  ;
	input \u1_uk_K_r4_reg[15]/NET0131  ;
	input \u1_uk_K_r4_reg[16]/NET0131  ;
	input \u1_uk_K_r4_reg[17]/NET0131  ;
	input \u1_uk_K_r4_reg[18]/NET0131  ;
	input \u1_uk_K_r4_reg[19]/NET0131  ;
	input \u1_uk_K_r4_reg[1]/NET0131  ;
	input \u1_uk_K_r4_reg[20]/NET0131  ;
	input \u1_uk_K_r4_reg[21]/NET0131  ;
	input \u1_uk_K_r4_reg[22]/NET0131  ;
	input \u1_uk_K_r4_reg[23]/P0001  ;
	input \u1_uk_K_r4_reg[25]/NET0131  ;
	input \u1_uk_K_r4_reg[26]/NET0131  ;
	input \u1_uk_K_r4_reg[27]/P0001  ;
	input \u1_uk_K_r4_reg[28]/NET0131  ;
	input \u1_uk_K_r4_reg[29]/NET0131  ;
	input \u1_uk_K_r4_reg[30]/NET0131  ;
	input \u1_uk_K_r4_reg[31]/P0001  ;
	input \u1_uk_K_r4_reg[32]/NET0131  ;
	input \u1_uk_K_r4_reg[33]/NET0131  ;
	input \u1_uk_K_r4_reg[34]/NET0131  ;
	input \u1_uk_K_r4_reg[35]/NET0131  ;
	input \u1_uk_K_r4_reg[36]/NET0131  ;
	input \u1_uk_K_r4_reg[37]/NET0131  ;
	input \u1_uk_K_r4_reg[38]/NET0131  ;
	input \u1_uk_K_r4_reg[39]/NET0131  ;
	input \u1_uk_K_r4_reg[3]/NET0131  ;
	input \u1_uk_K_r4_reg[40]/NET0131  ;
	input \u1_uk_K_r4_reg[41]/NET0131  ;
	input \u1_uk_K_r4_reg[42]/NET0131  ;
	input \u1_uk_K_r4_reg[43]/NET0131  ;
	input \u1_uk_K_r4_reg[44]/NET0131  ;
	input \u1_uk_K_r4_reg[45]/NET0131  ;
	input \u1_uk_K_r4_reg[46]/NET0131  ;
	input \u1_uk_K_r4_reg[47]/NET0131  ;
	input \u1_uk_K_r4_reg[48]/NET0131  ;
	input \u1_uk_K_r4_reg[49]/NET0131  ;
	input \u1_uk_K_r4_reg[4]/NET0131  ;
	input \u1_uk_K_r4_reg[50]/NET0131  ;
	input \u1_uk_K_r4_reg[51]/NET0131  ;
	input \u1_uk_K_r4_reg[52]/NET0131  ;
	input \u1_uk_K_r4_reg[53]/NET0131  ;
	input \u1_uk_K_r4_reg[54]/NET0131  ;
	input \u1_uk_K_r4_reg[55]/NET0131  ;
	input \u1_uk_K_r4_reg[5]/NET0131  ;
	input \u1_uk_K_r4_reg[6]/NET0131  ;
	input \u1_uk_K_r4_reg[7]/NET0131  ;
	input \u1_uk_K_r4_reg[8]/NET0131  ;
	input \u1_uk_K_r4_reg[9]/NET0131  ;
	input \u1_uk_K_r5_reg[0]/NET0131  ;
	input \u1_uk_K_r5_reg[10]/NET0131  ;
	input \u1_uk_K_r5_reg[11]/NET0131  ;
	input \u1_uk_K_r5_reg[12]/P0001  ;
	input \u1_uk_K_r5_reg[13]/P0001  ;
	input \u1_uk_K_r5_reg[14]/NET0131  ;
	input \u1_uk_K_r5_reg[15]/NET0131  ;
	input \u1_uk_K_r5_reg[16]/NET0131  ;
	input \u1_uk_K_r5_reg[17]/NET0131  ;
	input \u1_uk_K_r5_reg[18]/NET0131  ;
	input \u1_uk_K_r5_reg[19]/NET0131  ;
	input \u1_uk_K_r5_reg[1]/NET0131  ;
	input \u1_uk_K_r5_reg[20]/NET0131  ;
	input \u1_uk_K_r5_reg[21]/NET0131  ;
	input \u1_uk_K_r5_reg[22]/NET0131  ;
	input \u1_uk_K_r5_reg[23]/NET0131  ;
	input \u1_uk_K_r5_reg[24]/NET0131  ;
	input \u1_uk_K_r5_reg[25]/NET0131  ;
	input \u1_uk_K_r5_reg[26]/NET0131  ;
	input \u1_uk_K_r5_reg[27]/NET0131  ;
	input \u1_uk_K_r5_reg[28]/NET0131  ;
	input \u1_uk_K_r5_reg[29]/NET0131  ;
	input \u1_uk_K_r5_reg[2]/NET0131  ;
	input \u1_uk_K_r5_reg[30]/NET0131  ;
	input \u1_uk_K_r5_reg[31]/NET0131  ;
	input \u1_uk_K_r5_reg[32]/NET0131  ;
	input \u1_uk_K_r5_reg[33]/NET0131  ;
	input \u1_uk_K_r5_reg[34]/NET0131  ;
	input \u1_uk_K_r5_reg[35]/NET0131  ;
	input \u1_uk_K_r5_reg[36]/NET0131  ;
	input \u1_uk_K_r5_reg[37]/P0001  ;
	input \u1_uk_K_r5_reg[38]/NET0131  ;
	input \u1_uk_K_r5_reg[39]/NET0131  ;
	input \u1_uk_K_r5_reg[3]/NET0131  ;
	input \u1_uk_K_r5_reg[40]/NET0131  ;
	input \u1_uk_K_r5_reg[41]/NET0131  ;
	input \u1_uk_K_r5_reg[42]/NET0131  ;
	input \u1_uk_K_r5_reg[43]/NET0131  ;
	input \u1_uk_K_r5_reg[44]/NET0131  ;
	input \u1_uk_K_r5_reg[46]/NET0131  ;
	input \u1_uk_K_r5_reg[47]/NET0131  ;
	input \u1_uk_K_r5_reg[48]/NET0131  ;
	input \u1_uk_K_r5_reg[49]/NET0131  ;
	input \u1_uk_K_r5_reg[4]/NET0131  ;
	input \u1_uk_K_r5_reg[50]/NET0131  ;
	input \u1_uk_K_r5_reg[51]/NET0131  ;
	input \u1_uk_K_r5_reg[52]/NET0131  ;
	input \u1_uk_K_r5_reg[53]/NET0131  ;
	input \u1_uk_K_r5_reg[54]/NET0131  ;
	input \u1_uk_K_r5_reg[55]/NET0131  ;
	input \u1_uk_K_r5_reg[5]/NET0131  ;
	input \u1_uk_K_r5_reg[6]/NET0131  ;
	input \u1_uk_K_r5_reg[7]/NET0131  ;
	input \u1_uk_K_r5_reg[8]/NET0131  ;
	input \u1_uk_K_r5_reg[9]/NET0131  ;
	input \u1_uk_K_r6_reg[0]/NET0131  ;
	input \u1_uk_K_r6_reg[10]/NET0131  ;
	input \u1_uk_K_r6_reg[11]/NET0131  ;
	input \u1_uk_K_r6_reg[12]/NET0131  ;
	input \u1_uk_K_r6_reg[13]/NET0131  ;
	input \u1_uk_K_r6_reg[14]/NET0131  ;
	input \u1_uk_K_r6_reg[15]/NET0131  ;
	input \u1_uk_K_r6_reg[16]/NET0131  ;
	input \u1_uk_K_r6_reg[17]/NET0131  ;
	input \u1_uk_K_r6_reg[18]/NET0131  ;
	input \u1_uk_K_r6_reg[19]/NET0131  ;
	input \u1_uk_K_r6_reg[1]/NET0131  ;
	input \u1_uk_K_r6_reg[20]/NET0131  ;
	input \u1_uk_K_r6_reg[21]/NET0131  ;
	input \u1_uk_K_r6_reg[22]/NET0131  ;
	input \u1_uk_K_r6_reg[23]/P0001  ;
	input \u1_uk_K_r6_reg[24]/NET0131  ;
	input \u1_uk_K_r6_reg[25]/NET0131  ;
	input \u1_uk_K_r6_reg[26]/NET0131  ;
	input \u1_uk_K_r6_reg[27]/NET0131  ;
	input \u1_uk_K_r6_reg[28]/NET0131  ;
	input \u1_uk_K_r6_reg[29]/NET0131  ;
	input \u1_uk_K_r6_reg[2]/NET0131  ;
	input \u1_uk_K_r6_reg[30]/P0001  ;
	input \u1_uk_K_r6_reg[31]/NET0131  ;
	input \u1_uk_K_r6_reg[32]/NET0131  ;
	input \u1_uk_K_r6_reg[33]/NET0131  ;
	input \u1_uk_K_r6_reg[34]/NET0131  ;
	input \u1_uk_K_r6_reg[35]/NET0131  ;
	input \u1_uk_K_r6_reg[36]/NET0131  ;
	input \u1_uk_K_r6_reg[37]/NET0131  ;
	input \u1_uk_K_r6_reg[38]/NET0131  ;
	input \u1_uk_K_r6_reg[39]/NET0131  ;
	input \u1_uk_K_r6_reg[3]/NET0131  ;
	input \u1_uk_K_r6_reg[40]/NET0131  ;
	input \u1_uk_K_r6_reg[41]/NET0131  ;
	input \u1_uk_K_r6_reg[42]/NET0131  ;
	input \u1_uk_K_r6_reg[43]/NET0131  ;
	input \u1_uk_K_r6_reg[44]/NET0131  ;
	input \u1_uk_K_r6_reg[45]/NET0131  ;
	input \u1_uk_K_r6_reg[46]/NET0131  ;
	input \u1_uk_K_r6_reg[47]/NET0131  ;
	input \u1_uk_K_r6_reg[48]/NET0131  ;
	input \u1_uk_K_r6_reg[49]/NET0131  ;
	input \u1_uk_K_r6_reg[4]/NET0131  ;
	input \u1_uk_K_r6_reg[50]/NET0131  ;
	input \u1_uk_K_r6_reg[51]/NET0131  ;
	input \u1_uk_K_r6_reg[52]/NET0131  ;
	input \u1_uk_K_r6_reg[53]/NET0131  ;
	input \u1_uk_K_r6_reg[54]/NET0131  ;
	input \u1_uk_K_r6_reg[55]/P0001  ;
	input \u1_uk_K_r6_reg[5]/NET0131  ;
	input \u1_uk_K_r6_reg[6]/NET0131  ;
	input \u1_uk_K_r6_reg[7]/NET0131  ;
	input \u1_uk_K_r6_reg[8]/NET0131  ;
	input \u1_uk_K_r6_reg[9]/NET0131  ;
	input \u1_uk_K_r7_reg[0]/NET0131  ;
	input \u1_uk_K_r7_reg[10]/NET0131  ;
	input \u1_uk_K_r7_reg[11]/NET0131  ;
	input \u1_uk_K_r7_reg[12]/NET0131  ;
	input \u1_uk_K_r7_reg[13]/NET0131  ;
	input \u1_uk_K_r7_reg[14]/NET0131  ;
	input \u1_uk_K_r7_reg[15]/NET0131  ;
	input \u1_uk_K_r7_reg[16]/NET0131  ;
	input \u1_uk_K_r7_reg[17]/NET0131  ;
	input \u1_uk_K_r7_reg[18]/NET0131  ;
	input \u1_uk_K_r7_reg[19]/NET0131  ;
	input \u1_uk_K_r7_reg[1]/NET0131  ;
	input \u1_uk_K_r7_reg[20]/NET0131  ;
	input \u1_uk_K_r7_reg[21]/NET0131  ;
	input \u1_uk_K_r7_reg[22]/NET0131  ;
	input \u1_uk_K_r7_reg[23]/P0001  ;
	input \u1_uk_K_r7_reg[24]/NET0131  ;
	input \u1_uk_K_r7_reg[25]/NET0131  ;
	input \u1_uk_K_r7_reg[26]/P0001  ;
	input \u1_uk_K_r7_reg[27]/NET0131  ;
	input \u1_uk_K_r7_reg[28]/NET0131  ;
	input \u1_uk_K_r7_reg[29]/NET0131  ;
	input \u1_uk_K_r7_reg[2]/NET0131  ;
	input \u1_uk_K_r7_reg[30]/P0001  ;
	input \u1_uk_K_r7_reg[31]/NET0131  ;
	input \u1_uk_K_r7_reg[32]/NET0131  ;
	input \u1_uk_K_r7_reg[33]/NET0131  ;
	input \u1_uk_K_r7_reg[34]/NET0131  ;
	input \u1_uk_K_r7_reg[35]/NET0131  ;
	input \u1_uk_K_r7_reg[36]/NET0131  ;
	input \u1_uk_K_r7_reg[37]/NET0131  ;
	input \u1_uk_K_r7_reg[38]/NET0131  ;
	input \u1_uk_K_r7_reg[39]/NET0131  ;
	input \u1_uk_K_r7_reg[3]/NET0131  ;
	input \u1_uk_K_r7_reg[40]/NET0131  ;
	input \u1_uk_K_r7_reg[41]/NET0131  ;
	input \u1_uk_K_r7_reg[42]/NET0131  ;
	input \u1_uk_K_r7_reg[43]/NET0131  ;
	input \u1_uk_K_r7_reg[44]/NET0131  ;
	input \u1_uk_K_r7_reg[45]/NET0131  ;
	input \u1_uk_K_r7_reg[46]/NET0131  ;
	input \u1_uk_K_r7_reg[47]/NET0131  ;
	input \u1_uk_K_r7_reg[48]/NET0131  ;
	input \u1_uk_K_r7_reg[49]/NET0131  ;
	input \u1_uk_K_r7_reg[4]/NET0131  ;
	input \u1_uk_K_r7_reg[50]/NET0131  ;
	input \u1_uk_K_r7_reg[51]/NET0131  ;
	input \u1_uk_K_r7_reg[52]/NET0131  ;
	input \u1_uk_K_r7_reg[53]/NET0131  ;
	input \u1_uk_K_r7_reg[54]/NET0131  ;
	input \u1_uk_K_r7_reg[55]/P0001  ;
	input \u1_uk_K_r7_reg[5]/NET0131  ;
	input \u1_uk_K_r7_reg[6]/NET0131  ;
	input \u1_uk_K_r7_reg[7]/NET0131  ;
	input \u1_uk_K_r7_reg[8]/NET0131  ;
	input \u1_uk_K_r7_reg[9]/NET0131  ;
	input \u1_uk_K_r8_reg[0]/NET0131  ;
	input \u1_uk_K_r8_reg[10]/NET0131  ;
	input \u1_uk_K_r8_reg[11]/NET0131  ;
	input \u1_uk_K_r8_reg[12]/NET0131  ;
	input \u1_uk_K_r8_reg[13]/P0001  ;
	input \u1_uk_K_r8_reg[14]/NET0131  ;
	input \u1_uk_K_r8_reg[15]/NET0131  ;
	input \u1_uk_K_r8_reg[16]/NET0131  ;
	input \u1_uk_K_r8_reg[17]/NET0131  ;
	input \u1_uk_K_r8_reg[18]/NET0131  ;
	input \u1_uk_K_r8_reg[19]/NET0131  ;
	input \u1_uk_K_r8_reg[1]/NET0131  ;
	input \u1_uk_K_r8_reg[20]/NET0131  ;
	input \u1_uk_K_r8_reg[21]/NET0131  ;
	input \u1_uk_K_r8_reg[22]/NET0131  ;
	input \u1_uk_K_r8_reg[23]/NET0131  ;
	input \u1_uk_K_r8_reg[24]/NET0131  ;
	input \u1_uk_K_r8_reg[25]/NET0131  ;
	input \u1_uk_K_r8_reg[26]/NET0131  ;
	input \u1_uk_K_r8_reg[27]/NET0131  ;
	input \u1_uk_K_r8_reg[28]/NET0131  ;
	input \u1_uk_K_r8_reg[29]/NET0131  ;
	input \u1_uk_K_r8_reg[2]/NET0131  ;
	input \u1_uk_K_r8_reg[30]/NET0131  ;
	input \u1_uk_K_r8_reg[31]/NET0131  ;
	input \u1_uk_K_r8_reg[32]/NET0131  ;
	input \u1_uk_K_r8_reg[33]/NET0131  ;
	input \u1_uk_K_r8_reg[34]/NET0131  ;
	input \u1_uk_K_r8_reg[35]/NET0131  ;
	input \u1_uk_K_r8_reg[36]/NET0131  ;
	input \u1_uk_K_r8_reg[37]/P0001  ;
	input \u1_uk_K_r8_reg[38]/NET0131  ;
	input \u1_uk_K_r8_reg[39]/NET0131  ;
	input \u1_uk_K_r8_reg[3]/NET0131  ;
	input \u1_uk_K_r8_reg[40]/NET0131  ;
	input \u1_uk_K_r8_reg[41]/NET0131  ;
	input \u1_uk_K_r8_reg[42]/NET0131  ;
	input \u1_uk_K_r8_reg[43]/NET0131  ;
	input \u1_uk_K_r8_reg[44]/NET0131  ;
	input \u1_uk_K_r8_reg[46]/NET0131  ;
	input \u1_uk_K_r8_reg[47]/NET0131  ;
	input \u1_uk_K_r8_reg[48]/NET0131  ;
	input \u1_uk_K_r8_reg[49]/NET0131  ;
	input \u1_uk_K_r8_reg[4]/NET0131  ;
	input \u1_uk_K_r8_reg[50]/NET0131  ;
	input \u1_uk_K_r8_reg[51]/NET0131  ;
	input \u1_uk_K_r8_reg[52]/NET0131  ;
	input \u1_uk_K_r8_reg[53]/NET0131  ;
	input \u1_uk_K_r8_reg[54]/NET0131  ;
	input \u1_uk_K_r8_reg[55]/NET0131  ;
	input \u1_uk_K_r8_reg[5]/NET0131  ;
	input \u1_uk_K_r8_reg[6]/NET0131  ;
	input \u1_uk_K_r8_reg[7]/NET0131  ;
	input \u1_uk_K_r8_reg[8]/NET0131  ;
	input \u1_uk_K_r8_reg[9]/NET0131  ;
	input \u1_uk_K_r9_reg[0]/P0001  ;
	input \u1_uk_K_r9_reg[10]/NET0131  ;
	input \u1_uk_K_r9_reg[11]/NET0131  ;
	input \u1_uk_K_r9_reg[12]/NET0131  ;
	input \u1_uk_K_r9_reg[13]/NET0131  ;
	input \u1_uk_K_r9_reg[14]/NET0131  ;
	input \u1_uk_K_r9_reg[15]/NET0131  ;
	input \u1_uk_K_r9_reg[16]/NET0131  ;
	input \u1_uk_K_r9_reg[17]/NET0131  ;
	input \u1_uk_K_r9_reg[18]/NET0131  ;
	input \u1_uk_K_r9_reg[19]/NET0131  ;
	input \u1_uk_K_r9_reg[1]/NET0131  ;
	input \u1_uk_K_r9_reg[20]/NET0131  ;
	input \u1_uk_K_r9_reg[21]/NET0131  ;
	input \u1_uk_K_r9_reg[22]/NET0131  ;
	input \u1_uk_K_r9_reg[23]/NET0131  ;
	input \u1_uk_K_r9_reg[25]/NET0131  ;
	input \u1_uk_K_r9_reg[26]/NET0131  ;
	input \u1_uk_K_r9_reg[27]/P0001  ;
	input \u1_uk_K_r9_reg[28]/NET0131  ;
	input \u1_uk_K_r9_reg[29]/NET0131  ;
	input \u1_uk_K_r9_reg[30]/NET0131  ;
	input \u1_uk_K_r9_reg[31]/P0001  ;
	input \u1_uk_K_r9_reg[32]/NET0131  ;
	input \u1_uk_K_r9_reg[33]/NET0131  ;
	input \u1_uk_K_r9_reg[34]/NET0131  ;
	input \u1_uk_K_r9_reg[35]/NET0131  ;
	input \u1_uk_K_r9_reg[36]/NET0131  ;
	input \u1_uk_K_r9_reg[37]/NET0131  ;
	input \u1_uk_K_r9_reg[38]/NET0131  ;
	input \u1_uk_K_r9_reg[39]/NET0131  ;
	input \u1_uk_K_r9_reg[3]/NET0131  ;
	input \u1_uk_K_r9_reg[40]/NET0131  ;
	input \u1_uk_K_r9_reg[41]/NET0131  ;
	input \u1_uk_K_r9_reg[42]/NET0131  ;
	input \u1_uk_K_r9_reg[43]/NET0131  ;
	input \u1_uk_K_r9_reg[44]/NET0131  ;
	input \u1_uk_K_r9_reg[45]/NET0131  ;
	input \u1_uk_K_r9_reg[46]/NET0131  ;
	input \u1_uk_K_r9_reg[47]/NET0131  ;
	input \u1_uk_K_r9_reg[48]/NET0131  ;
	input \u1_uk_K_r9_reg[49]/NET0131  ;
	input \u1_uk_K_r9_reg[4]/NET0131  ;
	input \u1_uk_K_r9_reg[50]/NET0131  ;
	input \u1_uk_K_r9_reg[51]/NET0131  ;
	input \u1_uk_K_r9_reg[52]/NET0131  ;
	input \u1_uk_K_r9_reg[53]/NET0131  ;
	input \u1_uk_K_r9_reg[54]/NET0131  ;
	input \u1_uk_K_r9_reg[55]/NET0131  ;
	input \u1_uk_K_r9_reg[5]/NET0131  ;
	input \u1_uk_K_r9_reg[6]/NET0131  ;
	input \u1_uk_K_r9_reg[7]/NET0131  ;
	input \u1_uk_K_r9_reg[8]/NET0131  ;
	input \u1_uk_K_r9_reg[9]/NET0131  ;
	input \u2_L0_reg[10]/NET0131  ;
	input \u2_L0_reg[11]/NET0131  ;
	input \u2_L0_reg[12]/NET0131  ;
	input \u2_L0_reg[13]/NET0131  ;
	input \u2_L0_reg[14]/NET0131  ;
	input \u2_L0_reg[15]/NET0131  ;
	input \u2_L0_reg[16]/NET0131  ;
	input \u2_L0_reg[17]/NET0131  ;
	input \u2_L0_reg[18]/P0001  ;
	input \u2_L0_reg[19]/NET0131  ;
	input \u2_L0_reg[1]/NET0131  ;
	input \u2_L0_reg[20]/NET0131  ;
	input \u2_L0_reg[21]/NET0131  ;
	input \u2_L0_reg[22]/NET0131  ;
	input \u2_L0_reg[23]/NET0131  ;
	input \u2_L0_reg[24]/NET0131  ;
	input \u2_L0_reg[25]/NET0131  ;
	input \u2_L0_reg[26]/NET0131  ;
	input \u2_L0_reg[27]/NET0131  ;
	input \u2_L0_reg[28]/NET0131  ;
	input \u2_L0_reg[29]/NET0131  ;
	input \u2_L0_reg[2]/NET0131  ;
	input \u2_L0_reg[30]/NET0131  ;
	input \u2_L0_reg[31]/NET0131  ;
	input \u2_L0_reg[32]/NET0131  ;
	input \u2_L0_reg[3]/NET0131  ;
	input \u2_L0_reg[4]/NET0131  ;
	input \u2_L0_reg[5]/NET0131  ;
	input \u2_L0_reg[6]/NET0131  ;
	input \u2_L0_reg[7]/NET0131  ;
	input \u2_L0_reg[8]/NET0131  ;
	input \u2_L0_reg[9]/NET0131  ;
	input \u2_L10_reg[10]/NET0131  ;
	input \u2_L10_reg[11]/NET0131  ;
	input \u2_L10_reg[12]/NET0131  ;
	input \u2_L10_reg[13]/NET0131  ;
	input \u2_L10_reg[14]/NET0131  ;
	input \u2_L10_reg[15]/NET0131  ;
	input \u2_L10_reg[16]/NET0131  ;
	input \u2_L10_reg[17]/NET0131  ;
	input \u2_L10_reg[18]/P0001  ;
	input \u2_L10_reg[19]/NET0131  ;
	input \u2_L10_reg[1]/NET0131  ;
	input \u2_L10_reg[20]/NET0131  ;
	input \u2_L10_reg[21]/NET0131  ;
	input \u2_L10_reg[22]/NET0131  ;
	input \u2_L10_reg[23]/NET0131  ;
	input \u2_L10_reg[24]/NET0131  ;
	input \u2_L10_reg[25]/NET0131  ;
	input \u2_L10_reg[26]/NET0131  ;
	input \u2_L10_reg[27]/NET0131  ;
	input \u2_L10_reg[28]/NET0131  ;
	input \u2_L10_reg[29]/NET0131  ;
	input \u2_L10_reg[2]/NET0131  ;
	input \u2_L10_reg[30]/NET0131  ;
	input \u2_L10_reg[31]/NET0131  ;
	input \u2_L10_reg[32]/NET0131  ;
	input \u2_L10_reg[3]/NET0131  ;
	input \u2_L10_reg[4]/NET0131  ;
	input \u2_L10_reg[5]/NET0131  ;
	input \u2_L10_reg[6]/NET0131  ;
	input \u2_L10_reg[7]/NET0131  ;
	input \u2_L10_reg[8]/NET0131  ;
	input \u2_L10_reg[9]/NET0131  ;
	input \u2_L11_reg[10]/NET0131  ;
	input \u2_L11_reg[11]/NET0131  ;
	input \u2_L11_reg[12]/NET0131  ;
	input \u2_L11_reg[13]/NET0131  ;
	input \u2_L11_reg[14]/NET0131  ;
	input \u2_L11_reg[15]/NET0131  ;
	input \u2_L11_reg[16]/NET0131  ;
	input \u2_L11_reg[17]/NET0131  ;
	input \u2_L11_reg[18]/P0001  ;
	input \u2_L11_reg[19]/NET0131  ;
	input \u2_L11_reg[1]/NET0131  ;
	input \u2_L11_reg[20]/NET0131  ;
	input \u2_L11_reg[21]/NET0131  ;
	input \u2_L11_reg[22]/NET0131  ;
	input \u2_L11_reg[23]/NET0131  ;
	input \u2_L11_reg[24]/NET0131  ;
	input \u2_L11_reg[25]/NET0131  ;
	input \u2_L11_reg[26]/NET0131  ;
	input \u2_L11_reg[27]/NET0131  ;
	input \u2_L11_reg[28]/NET0131  ;
	input \u2_L11_reg[29]/NET0131  ;
	input \u2_L11_reg[2]/NET0131  ;
	input \u2_L11_reg[30]/NET0131  ;
	input \u2_L11_reg[31]/NET0131  ;
	input \u2_L11_reg[32]/NET0131  ;
	input \u2_L11_reg[3]/NET0131  ;
	input \u2_L11_reg[4]/NET0131  ;
	input \u2_L11_reg[5]/NET0131  ;
	input \u2_L11_reg[6]/NET0131  ;
	input \u2_L11_reg[7]/NET0131  ;
	input \u2_L11_reg[8]/NET0131  ;
	input \u2_L11_reg[9]/NET0131  ;
	input \u2_L12_reg[10]/NET0131  ;
	input \u2_L12_reg[11]/NET0131  ;
	input \u2_L12_reg[12]/NET0131  ;
	input \u2_L12_reg[13]/NET0131  ;
	input \u2_L12_reg[14]/NET0131  ;
	input \u2_L12_reg[15]/NET0131  ;
	input \u2_L12_reg[16]/NET0131  ;
	input \u2_L12_reg[17]/NET0131  ;
	input \u2_L12_reg[18]/P0001  ;
	input \u2_L12_reg[19]/NET0131  ;
	input \u2_L12_reg[1]/NET0131  ;
	input \u2_L12_reg[20]/NET0131  ;
	input \u2_L12_reg[21]/NET0131  ;
	input \u2_L12_reg[22]/NET0131  ;
	input \u2_L12_reg[23]/NET0131  ;
	input \u2_L12_reg[24]/NET0131  ;
	input \u2_L12_reg[25]/NET0131  ;
	input \u2_L12_reg[26]/NET0131  ;
	input \u2_L12_reg[27]/NET0131  ;
	input \u2_L12_reg[28]/NET0131  ;
	input \u2_L12_reg[29]/NET0131  ;
	input \u2_L12_reg[2]/NET0131  ;
	input \u2_L12_reg[30]/NET0131  ;
	input \u2_L12_reg[31]/NET0131  ;
	input \u2_L12_reg[32]/NET0131  ;
	input \u2_L12_reg[3]/NET0131  ;
	input \u2_L12_reg[4]/NET0131  ;
	input \u2_L12_reg[5]/NET0131  ;
	input \u2_L12_reg[6]/NET0131  ;
	input \u2_L12_reg[7]/NET0131  ;
	input \u2_L12_reg[8]/NET0131  ;
	input \u2_L12_reg[9]/NET0131  ;
	input \u2_L13_reg[10]/NET0131  ;
	input \u2_L13_reg[11]/NET0131  ;
	input \u2_L13_reg[12]/NET0131  ;
	input \u2_L13_reg[13]/NET0131  ;
	input \u2_L13_reg[14]/NET0131  ;
	input \u2_L13_reg[15]/NET0131  ;
	input \u2_L13_reg[16]/NET0131  ;
	input \u2_L13_reg[17]/NET0131  ;
	input \u2_L13_reg[18]/P0001  ;
	input \u2_L13_reg[19]/P0001  ;
	input \u2_L13_reg[1]/NET0131  ;
	input \u2_L13_reg[20]/NET0131  ;
	input \u2_L13_reg[21]/NET0131  ;
	input \u2_L13_reg[22]/NET0131  ;
	input \u2_L13_reg[23]/P0001  ;
	input \u2_L13_reg[24]/NET0131  ;
	input \u2_L13_reg[25]/NET0131  ;
	input \u2_L13_reg[26]/NET0131  ;
	input \u2_L13_reg[27]/NET0131  ;
	input \u2_L13_reg[28]/NET0131  ;
	input \u2_L13_reg[29]/NET0131  ;
	input \u2_L13_reg[2]/NET0131  ;
	input \u2_L13_reg[30]/NET0131  ;
	input \u2_L13_reg[31]/NET0131  ;
	input \u2_L13_reg[32]/NET0131  ;
	input \u2_L13_reg[3]/NET0131  ;
	input \u2_L13_reg[4]/NET0131  ;
	input \u2_L13_reg[5]/NET0131  ;
	input \u2_L13_reg[6]/NET0131  ;
	input \u2_L13_reg[7]/NET0131  ;
	input \u2_L13_reg[8]/NET0131  ;
	input \u2_L13_reg[9]/NET0131  ;
	input \u2_L14_reg[10]/P0001  ;
	input \u2_L14_reg[11]/P0001  ;
	input \u2_L14_reg[12]/P0001  ;
	input \u2_L14_reg[13]/P0001  ;
	input \u2_L14_reg[14]/P0001  ;
	input \u2_L14_reg[15]/P0001  ;
	input \u2_L14_reg[16]/P0001  ;
	input \u2_L14_reg[17]/P0001  ;
	input \u2_L14_reg[18]/P0001  ;
	input \u2_L14_reg[19]/P0001  ;
	input \u2_L14_reg[1]/P0001  ;
	input \u2_L14_reg[20]/P0001  ;
	input \u2_L14_reg[21]/P0001  ;
	input \u2_L14_reg[22]/P0001  ;
	input \u2_L14_reg[23]/P0001  ;
	input \u2_L14_reg[24]/P0001  ;
	input \u2_L14_reg[25]/P0001  ;
	input \u2_L14_reg[26]/P0001  ;
	input \u2_L14_reg[27]/P0001  ;
	input \u2_L14_reg[28]/P0001  ;
	input \u2_L14_reg[29]/P0001  ;
	input \u2_L14_reg[2]/P0001  ;
	input \u2_L14_reg[30]/P0001  ;
	input \u2_L14_reg[31]/P0001  ;
	input \u2_L14_reg[32]/P0001  ;
	input \u2_L14_reg[3]/P0001  ;
	input \u2_L14_reg[4]/P0001  ;
	input \u2_L14_reg[5]/P0001  ;
	input \u2_L14_reg[6]/P0001  ;
	input \u2_L14_reg[7]/P0001  ;
	input \u2_L14_reg[8]/P0001  ;
	input \u2_L14_reg[9]/P0001  ;
	input \u2_L1_reg[10]/NET0131  ;
	input \u2_L1_reg[11]/NET0131  ;
	input \u2_L1_reg[12]/NET0131  ;
	input \u2_L1_reg[13]/NET0131  ;
	input \u2_L1_reg[14]/NET0131  ;
	input \u2_L1_reg[15]/NET0131  ;
	input \u2_L1_reg[16]/NET0131  ;
	input \u2_L1_reg[17]/NET0131  ;
	input \u2_L1_reg[18]/P0001  ;
	input \u2_L1_reg[19]/NET0131  ;
	input \u2_L1_reg[1]/NET0131  ;
	input \u2_L1_reg[20]/NET0131  ;
	input \u2_L1_reg[21]/NET0131  ;
	input \u2_L1_reg[22]/NET0131  ;
	input \u2_L1_reg[23]/NET0131  ;
	input \u2_L1_reg[24]/NET0131  ;
	input \u2_L1_reg[25]/NET0131  ;
	input \u2_L1_reg[26]/NET0131  ;
	input \u2_L1_reg[27]/NET0131  ;
	input \u2_L1_reg[28]/NET0131  ;
	input \u2_L1_reg[29]/NET0131  ;
	input \u2_L1_reg[2]/NET0131  ;
	input \u2_L1_reg[30]/NET0131  ;
	input \u2_L1_reg[31]/NET0131  ;
	input \u2_L1_reg[32]/NET0131  ;
	input \u2_L1_reg[3]/NET0131  ;
	input \u2_L1_reg[4]/NET0131  ;
	input \u2_L1_reg[5]/NET0131  ;
	input \u2_L1_reg[6]/NET0131  ;
	input \u2_L1_reg[7]/NET0131  ;
	input \u2_L1_reg[8]/NET0131  ;
	input \u2_L1_reg[9]/NET0131  ;
	input \u2_L2_reg[10]/NET0131  ;
	input \u2_L2_reg[11]/NET0131  ;
	input \u2_L2_reg[12]/NET0131  ;
	input \u2_L2_reg[13]/NET0131  ;
	input \u2_L2_reg[14]/NET0131  ;
	input \u2_L2_reg[15]/NET0131  ;
	input \u2_L2_reg[16]/NET0131  ;
	input \u2_L2_reg[17]/NET0131  ;
	input \u2_L2_reg[18]/P0001  ;
	input \u2_L2_reg[19]/NET0131  ;
	input \u2_L2_reg[1]/NET0131  ;
	input \u2_L2_reg[20]/NET0131  ;
	input \u2_L2_reg[21]/NET0131  ;
	input \u2_L2_reg[22]/NET0131  ;
	input \u2_L2_reg[23]/NET0131  ;
	input \u2_L2_reg[24]/NET0131  ;
	input \u2_L2_reg[25]/NET0131  ;
	input \u2_L2_reg[26]/NET0131  ;
	input \u2_L2_reg[27]/NET0131  ;
	input \u2_L2_reg[28]/NET0131  ;
	input \u2_L2_reg[29]/NET0131  ;
	input \u2_L2_reg[2]/NET0131  ;
	input \u2_L2_reg[30]/NET0131  ;
	input \u2_L2_reg[31]/NET0131  ;
	input \u2_L2_reg[32]/NET0131  ;
	input \u2_L2_reg[3]/NET0131  ;
	input \u2_L2_reg[4]/NET0131  ;
	input \u2_L2_reg[5]/NET0131  ;
	input \u2_L2_reg[6]/NET0131  ;
	input \u2_L2_reg[7]/NET0131  ;
	input \u2_L2_reg[8]/NET0131  ;
	input \u2_L2_reg[9]/NET0131  ;
	input \u2_L3_reg[10]/NET0131  ;
	input \u2_L3_reg[11]/NET0131  ;
	input \u2_L3_reg[12]/NET0131  ;
	input \u2_L3_reg[13]/NET0131  ;
	input \u2_L3_reg[14]/NET0131  ;
	input \u2_L3_reg[15]/NET0131  ;
	input \u2_L3_reg[16]/NET0131  ;
	input \u2_L3_reg[17]/NET0131  ;
	input \u2_L3_reg[18]/P0001  ;
	input \u2_L3_reg[19]/NET0131  ;
	input \u2_L3_reg[1]/NET0131  ;
	input \u2_L3_reg[20]/NET0131  ;
	input \u2_L3_reg[21]/NET0131  ;
	input \u2_L3_reg[22]/NET0131  ;
	input \u2_L3_reg[23]/NET0131  ;
	input \u2_L3_reg[24]/NET0131  ;
	input \u2_L3_reg[25]/NET0131  ;
	input \u2_L3_reg[26]/NET0131  ;
	input \u2_L3_reg[27]/NET0131  ;
	input \u2_L3_reg[28]/NET0131  ;
	input \u2_L3_reg[29]/NET0131  ;
	input \u2_L3_reg[2]/NET0131  ;
	input \u2_L3_reg[30]/NET0131  ;
	input \u2_L3_reg[31]/NET0131  ;
	input \u2_L3_reg[32]/NET0131  ;
	input \u2_L3_reg[3]/NET0131  ;
	input \u2_L3_reg[4]/NET0131  ;
	input \u2_L3_reg[5]/NET0131  ;
	input \u2_L3_reg[6]/NET0131  ;
	input \u2_L3_reg[7]/NET0131  ;
	input \u2_L3_reg[8]/NET0131  ;
	input \u2_L3_reg[9]/NET0131  ;
	input \u2_L4_reg[10]/NET0131  ;
	input \u2_L4_reg[11]/NET0131  ;
	input \u2_L4_reg[12]/NET0131  ;
	input \u2_L4_reg[13]/NET0131  ;
	input \u2_L4_reg[14]/NET0131  ;
	input \u2_L4_reg[15]/NET0131  ;
	input \u2_L4_reg[16]/NET0131  ;
	input \u2_L4_reg[17]/NET0131  ;
	input \u2_L4_reg[18]/P0001  ;
	input \u2_L4_reg[19]/NET0131  ;
	input \u2_L4_reg[1]/NET0131  ;
	input \u2_L4_reg[20]/NET0131  ;
	input \u2_L4_reg[21]/NET0131  ;
	input \u2_L4_reg[22]/NET0131  ;
	input \u2_L4_reg[23]/NET0131  ;
	input \u2_L4_reg[24]/NET0131  ;
	input \u2_L4_reg[25]/NET0131  ;
	input \u2_L4_reg[26]/NET0131  ;
	input \u2_L4_reg[27]/NET0131  ;
	input \u2_L4_reg[28]/NET0131  ;
	input \u2_L4_reg[29]/NET0131  ;
	input \u2_L4_reg[2]/NET0131  ;
	input \u2_L4_reg[30]/NET0131  ;
	input \u2_L4_reg[31]/NET0131  ;
	input \u2_L4_reg[32]/NET0131  ;
	input \u2_L4_reg[3]/NET0131  ;
	input \u2_L4_reg[4]/NET0131  ;
	input \u2_L4_reg[5]/NET0131  ;
	input \u2_L4_reg[6]/NET0131  ;
	input \u2_L4_reg[7]/NET0131  ;
	input \u2_L4_reg[8]/NET0131  ;
	input \u2_L4_reg[9]/NET0131  ;
	input \u2_L5_reg[10]/NET0131  ;
	input \u2_L5_reg[11]/NET0131  ;
	input \u2_L5_reg[12]/NET0131  ;
	input \u2_L5_reg[13]/NET0131  ;
	input \u2_L5_reg[14]/NET0131  ;
	input \u2_L5_reg[15]/NET0131  ;
	input \u2_L5_reg[16]/NET0131  ;
	input \u2_L5_reg[17]/NET0131  ;
	input \u2_L5_reg[18]/NET0131  ;
	input \u2_L5_reg[19]/NET0131  ;
	input \u2_L5_reg[1]/NET0131  ;
	input \u2_L5_reg[20]/NET0131  ;
	input \u2_L5_reg[21]/NET0131  ;
	input \u2_L5_reg[22]/NET0131  ;
	input \u2_L5_reg[23]/NET0131  ;
	input \u2_L5_reg[24]/NET0131  ;
	input \u2_L5_reg[25]/NET0131  ;
	input \u2_L5_reg[26]/NET0131  ;
	input \u2_L5_reg[27]/NET0131  ;
	input \u2_L5_reg[28]/NET0131  ;
	input \u2_L5_reg[29]/NET0131  ;
	input \u2_L5_reg[2]/NET0131  ;
	input \u2_L5_reg[30]/NET0131  ;
	input \u2_L5_reg[31]/NET0131  ;
	input \u2_L5_reg[32]/NET0131  ;
	input \u2_L5_reg[3]/NET0131  ;
	input \u2_L5_reg[4]/NET0131  ;
	input \u2_L5_reg[5]/NET0131  ;
	input \u2_L5_reg[6]/NET0131  ;
	input \u2_L5_reg[7]/NET0131  ;
	input \u2_L5_reg[8]/NET0131  ;
	input \u2_L5_reg[9]/NET0131  ;
	input \u2_L6_reg[10]/NET0131  ;
	input \u2_L6_reg[11]/NET0131  ;
	input \u2_L6_reg[12]/NET0131  ;
	input \u2_L6_reg[13]/NET0131  ;
	input \u2_L6_reg[14]/NET0131  ;
	input \u2_L6_reg[15]/NET0131  ;
	input \u2_L6_reg[16]/NET0131  ;
	input \u2_L6_reg[17]/NET0131  ;
	input \u2_L6_reg[18]/P0001  ;
	input \u2_L6_reg[19]/NET0131  ;
	input \u2_L6_reg[1]/NET0131  ;
	input \u2_L6_reg[20]/NET0131  ;
	input \u2_L6_reg[21]/NET0131  ;
	input \u2_L6_reg[22]/NET0131  ;
	input \u2_L6_reg[23]/NET0131  ;
	input \u2_L6_reg[24]/NET0131  ;
	input \u2_L6_reg[25]/NET0131  ;
	input \u2_L6_reg[26]/NET0131  ;
	input \u2_L6_reg[27]/NET0131  ;
	input \u2_L6_reg[28]/NET0131  ;
	input \u2_L6_reg[29]/NET0131  ;
	input \u2_L6_reg[2]/NET0131  ;
	input \u2_L6_reg[30]/NET0131  ;
	input \u2_L6_reg[31]/NET0131  ;
	input \u2_L6_reg[32]/NET0131  ;
	input \u2_L6_reg[3]/NET0131  ;
	input \u2_L6_reg[4]/NET0131  ;
	input \u2_L6_reg[5]/NET0131  ;
	input \u2_L6_reg[6]/NET0131  ;
	input \u2_L6_reg[7]/NET0131  ;
	input \u2_L6_reg[8]/NET0131  ;
	input \u2_L6_reg[9]/NET0131  ;
	input \u2_L7_reg[10]/NET0131  ;
	input \u2_L7_reg[11]/NET0131  ;
	input \u2_L7_reg[12]/NET0131  ;
	input \u2_L7_reg[13]/NET0131  ;
	input \u2_L7_reg[14]/NET0131  ;
	input \u2_L7_reg[15]/NET0131  ;
	input \u2_L7_reg[16]/NET0131  ;
	input \u2_L7_reg[17]/NET0131  ;
	input \u2_L7_reg[18]/P0001  ;
	input \u2_L7_reg[19]/NET0131  ;
	input \u2_L7_reg[1]/NET0131  ;
	input \u2_L7_reg[20]/NET0131  ;
	input \u2_L7_reg[21]/NET0131  ;
	input \u2_L7_reg[22]/NET0131  ;
	input \u2_L7_reg[23]/NET0131  ;
	input \u2_L7_reg[24]/NET0131  ;
	input \u2_L7_reg[25]/NET0131  ;
	input \u2_L7_reg[26]/NET0131  ;
	input \u2_L7_reg[27]/NET0131  ;
	input \u2_L7_reg[28]/NET0131  ;
	input \u2_L7_reg[29]/NET0131  ;
	input \u2_L7_reg[2]/NET0131  ;
	input \u2_L7_reg[30]/NET0131  ;
	input \u2_L7_reg[31]/NET0131  ;
	input \u2_L7_reg[32]/NET0131  ;
	input \u2_L7_reg[3]/NET0131  ;
	input \u2_L7_reg[4]/NET0131  ;
	input \u2_L7_reg[5]/NET0131  ;
	input \u2_L7_reg[6]/NET0131  ;
	input \u2_L7_reg[7]/NET0131  ;
	input \u2_L7_reg[8]/NET0131  ;
	input \u2_L7_reg[9]/NET0131  ;
	input \u2_L8_reg[10]/NET0131  ;
	input \u2_L8_reg[11]/NET0131  ;
	input \u2_L8_reg[12]/NET0131  ;
	input \u2_L8_reg[13]/NET0131  ;
	input \u2_L8_reg[14]/NET0131  ;
	input \u2_L8_reg[15]/NET0131  ;
	input \u2_L8_reg[16]/NET0131  ;
	input \u2_L8_reg[17]/NET0131  ;
	input \u2_L8_reg[18]/P0001  ;
	input \u2_L8_reg[19]/NET0131  ;
	input \u2_L8_reg[1]/NET0131  ;
	input \u2_L8_reg[20]/NET0131  ;
	input \u2_L8_reg[21]/NET0131  ;
	input \u2_L8_reg[22]/NET0131  ;
	input \u2_L8_reg[23]/NET0131  ;
	input \u2_L8_reg[24]/NET0131  ;
	input \u2_L8_reg[25]/NET0131  ;
	input \u2_L8_reg[26]/NET0131  ;
	input \u2_L8_reg[27]/NET0131  ;
	input \u2_L8_reg[28]/NET0131  ;
	input \u2_L8_reg[29]/NET0131  ;
	input \u2_L8_reg[2]/NET0131  ;
	input \u2_L8_reg[30]/NET0131  ;
	input \u2_L8_reg[31]/NET0131  ;
	input \u2_L8_reg[32]/NET0131  ;
	input \u2_L8_reg[3]/NET0131  ;
	input \u2_L8_reg[4]/NET0131  ;
	input \u2_L8_reg[5]/NET0131  ;
	input \u2_L8_reg[6]/NET0131  ;
	input \u2_L8_reg[7]/NET0131  ;
	input \u2_L8_reg[8]/NET0131  ;
	input \u2_L8_reg[9]/NET0131  ;
	input \u2_L9_reg[10]/NET0131  ;
	input \u2_L9_reg[11]/NET0131  ;
	input \u2_L9_reg[12]/NET0131  ;
	input \u2_L9_reg[13]/NET0131  ;
	input \u2_L9_reg[14]/NET0131  ;
	input \u2_L9_reg[15]/NET0131  ;
	input \u2_L9_reg[16]/NET0131  ;
	input \u2_L9_reg[17]/NET0131  ;
	input \u2_L9_reg[18]/P0001  ;
	input \u2_L9_reg[19]/NET0131  ;
	input \u2_L9_reg[1]/NET0131  ;
	input \u2_L9_reg[20]/NET0131  ;
	input \u2_L9_reg[21]/NET0131  ;
	input \u2_L9_reg[22]/NET0131  ;
	input \u2_L9_reg[23]/NET0131  ;
	input \u2_L9_reg[24]/NET0131  ;
	input \u2_L9_reg[25]/NET0131  ;
	input \u2_L9_reg[26]/NET0131  ;
	input \u2_L9_reg[27]/NET0131  ;
	input \u2_L9_reg[28]/NET0131  ;
	input \u2_L9_reg[29]/NET0131  ;
	input \u2_L9_reg[2]/NET0131  ;
	input \u2_L9_reg[30]/NET0131  ;
	input \u2_L9_reg[31]/NET0131  ;
	input \u2_L9_reg[32]/NET0131  ;
	input \u2_L9_reg[3]/NET0131  ;
	input \u2_L9_reg[4]/NET0131  ;
	input \u2_L9_reg[5]/NET0131  ;
	input \u2_L9_reg[6]/NET0131  ;
	input \u2_L9_reg[7]/NET0131  ;
	input \u2_L9_reg[8]/NET0131  ;
	input \u2_L9_reg[9]/NET0131  ;
	input \u2_R0_reg[10]/NET0131  ;
	input \u2_R0_reg[11]/P0001  ;
	input \u2_R0_reg[12]/NET0131  ;
	input \u2_R0_reg[13]/NET0131  ;
	input \u2_R0_reg[14]/NET0131  ;
	input \u2_R0_reg[15]/NET0131  ;
	input \u2_R0_reg[16]/NET0131  ;
	input \u2_R0_reg[17]/NET0131  ;
	input \u2_R0_reg[18]/NET0131  ;
	input \u2_R0_reg[19]/NET0131  ;
	input \u2_R0_reg[1]/NET0131  ;
	input \u2_R0_reg[20]/NET0131  ;
	input \u2_R0_reg[21]/NET0131  ;
	input \u2_R0_reg[22]/NET0131  ;
	input \u2_R0_reg[23]/NET0131  ;
	input \u2_R0_reg[24]/NET0131  ;
	input \u2_R0_reg[25]/NET0131  ;
	input \u2_R0_reg[26]/NET0131  ;
	input \u2_R0_reg[27]/NET0131  ;
	input \u2_R0_reg[28]/NET0131  ;
	input \u2_R0_reg[29]/NET0131  ;
	input \u2_R0_reg[2]/NET0131  ;
	input \u2_R0_reg[30]/NET0131  ;
	input \u2_R0_reg[31]/P0001  ;
	input \u2_R0_reg[32]/NET0131  ;
	input \u2_R0_reg[3]/NET0131  ;
	input \u2_R0_reg[4]/NET0131  ;
	input \u2_R0_reg[5]/NET0131  ;
	input \u2_R0_reg[6]/NET0131  ;
	input \u2_R0_reg[7]/NET0131  ;
	input \u2_R0_reg[8]/NET0131  ;
	input \u2_R0_reg[9]/NET0131  ;
	input \u2_R10_reg[10]/NET0131  ;
	input \u2_R10_reg[11]/NET0131  ;
	input \u2_R10_reg[12]/NET0131  ;
	input \u2_R10_reg[13]/NET0131  ;
	input \u2_R10_reg[14]/NET0131  ;
	input \u2_R10_reg[15]/NET0131  ;
	input \u2_R10_reg[16]/NET0131  ;
	input \u2_R10_reg[17]/NET0131  ;
	input \u2_R10_reg[18]/NET0131  ;
	input \u2_R10_reg[19]/NET0131  ;
	input \u2_R10_reg[1]/NET0131  ;
	input \u2_R10_reg[20]/NET0131  ;
	input \u2_R10_reg[21]/NET0131  ;
	input \u2_R10_reg[22]/NET0131  ;
	input \u2_R10_reg[23]/NET0131  ;
	input \u2_R10_reg[24]/NET0131  ;
	input \u2_R10_reg[25]/NET0131  ;
	input \u2_R10_reg[26]/NET0131  ;
	input \u2_R10_reg[27]/NET0131  ;
	input \u2_R10_reg[28]/NET0131  ;
	input \u2_R10_reg[29]/NET0131  ;
	input \u2_R10_reg[2]/NET0131  ;
	input \u2_R10_reg[30]/NET0131  ;
	input \u2_R10_reg[31]/P0001  ;
	input \u2_R10_reg[32]/NET0131  ;
	input \u2_R10_reg[3]/NET0131  ;
	input \u2_R10_reg[4]/NET0131  ;
	input \u2_R10_reg[5]/NET0131  ;
	input \u2_R10_reg[6]/NET0131  ;
	input \u2_R10_reg[7]/NET0131  ;
	input \u2_R10_reg[8]/NET0131  ;
	input \u2_R10_reg[9]/NET0131  ;
	input \u2_R11_reg[10]/NET0131  ;
	input \u2_R11_reg[11]/NET0131  ;
	input \u2_R11_reg[12]/NET0131  ;
	input \u2_R11_reg[13]/NET0131  ;
	input \u2_R11_reg[14]/NET0131  ;
	input \u2_R11_reg[15]/NET0131  ;
	input \u2_R11_reg[16]/NET0131  ;
	input \u2_R11_reg[17]/NET0131  ;
	input \u2_R11_reg[18]/NET0131  ;
	input \u2_R11_reg[19]/NET0131  ;
	input \u2_R11_reg[1]/NET0131  ;
	input \u2_R11_reg[20]/NET0131  ;
	input \u2_R11_reg[21]/NET0131  ;
	input \u2_R11_reg[22]/NET0131  ;
	input \u2_R11_reg[23]/NET0131  ;
	input \u2_R11_reg[24]/NET0131  ;
	input \u2_R11_reg[25]/NET0131  ;
	input \u2_R11_reg[26]/NET0131  ;
	input \u2_R11_reg[27]/NET0131  ;
	input \u2_R11_reg[28]/NET0131  ;
	input \u2_R11_reg[29]/NET0131  ;
	input \u2_R11_reg[2]/NET0131  ;
	input \u2_R11_reg[30]/NET0131  ;
	input \u2_R11_reg[31]/P0001  ;
	input \u2_R11_reg[32]/NET0131  ;
	input \u2_R11_reg[3]/NET0131  ;
	input \u2_R11_reg[4]/NET0131  ;
	input \u2_R11_reg[5]/NET0131  ;
	input \u2_R11_reg[6]/NET0131  ;
	input \u2_R11_reg[7]/NET0131  ;
	input \u2_R11_reg[8]/NET0131  ;
	input \u2_R11_reg[9]/NET0131  ;
	input \u2_R12_reg[10]/NET0131  ;
	input \u2_R12_reg[11]/NET0131  ;
	input \u2_R12_reg[12]/NET0131  ;
	input \u2_R12_reg[13]/NET0131  ;
	input \u2_R12_reg[14]/NET0131  ;
	input \u2_R12_reg[15]/NET0131  ;
	input \u2_R12_reg[16]/NET0131  ;
	input \u2_R12_reg[17]/NET0131  ;
	input \u2_R12_reg[18]/NET0131  ;
	input \u2_R12_reg[19]/NET0131  ;
	input \u2_R12_reg[1]/NET0131  ;
	input \u2_R12_reg[20]/NET0131  ;
	input \u2_R12_reg[21]/NET0131  ;
	input \u2_R12_reg[22]/NET0131  ;
	input \u2_R12_reg[23]/NET0131  ;
	input \u2_R12_reg[24]/NET0131  ;
	input \u2_R12_reg[25]/NET0131  ;
	input \u2_R12_reg[26]/NET0131  ;
	input \u2_R12_reg[27]/NET0131  ;
	input \u2_R12_reg[28]/NET0131  ;
	input \u2_R12_reg[29]/NET0131  ;
	input \u2_R12_reg[2]/NET0131  ;
	input \u2_R12_reg[30]/NET0131  ;
	input \u2_R12_reg[31]/P0001  ;
	input \u2_R12_reg[32]/NET0131  ;
	input \u2_R12_reg[3]/NET0131  ;
	input \u2_R12_reg[4]/NET0131  ;
	input \u2_R12_reg[5]/NET0131  ;
	input \u2_R12_reg[6]/NET0131  ;
	input \u2_R12_reg[7]/NET0131  ;
	input \u2_R12_reg[8]/NET0131  ;
	input \u2_R12_reg[9]/NET0131  ;
	input \u2_R13_reg[10]/NET0131  ;
	input \u2_R13_reg[11]/NET0131  ;
	input \u2_R13_reg[12]/NET0131  ;
	input \u2_R13_reg[13]/NET0131  ;
	input \u2_R13_reg[14]/NET0131  ;
	input \u2_R13_reg[15]/NET0131  ;
	input \u2_R13_reg[16]/NET0131  ;
	input \u2_R13_reg[17]/NET0131  ;
	input \u2_R13_reg[18]/NET0131  ;
	input \u2_R13_reg[19]/NET0131  ;
	input \u2_R13_reg[1]/NET0131  ;
	input \u2_R13_reg[20]/NET0131  ;
	input \u2_R13_reg[21]/NET0131  ;
	input \u2_R13_reg[22]/NET0131  ;
	input \u2_R13_reg[23]/NET0131  ;
	input \u2_R13_reg[24]/NET0131  ;
	input \u2_R13_reg[25]/NET0131  ;
	input \u2_R13_reg[26]/NET0131  ;
	input \u2_R13_reg[27]/P0001  ;
	input \u2_R13_reg[28]/NET0131  ;
	input \u2_R13_reg[29]/NET0131  ;
	input \u2_R13_reg[2]/NET0131  ;
	input \u2_R13_reg[30]/NET0131  ;
	input \u2_R13_reg[31]/P0001  ;
	input \u2_R13_reg[32]/NET0131  ;
	input \u2_R13_reg[3]/NET0131  ;
	input \u2_R13_reg[4]/NET0131  ;
	input \u2_R13_reg[5]/NET0131  ;
	input \u2_R13_reg[6]/NET0131  ;
	input \u2_R13_reg[7]/NET0131  ;
	input \u2_R13_reg[8]/NET0131  ;
	input \u2_R13_reg[9]/NET0131  ;
	input \u2_R14_reg[10]/P0001  ;
	input \u2_R14_reg[11]/P0001  ;
	input \u2_R14_reg[12]/NET0131  ;
	input \u2_R14_reg[13]/NET0131  ;
	input \u2_R14_reg[14]/NET0131  ;
	input \u2_R14_reg[15]/NET0131  ;
	input \u2_R14_reg[16]/NET0131  ;
	input \u2_R14_reg[17]/NET0131  ;
	input \u2_R14_reg[18]/NET0131  ;
	input \u2_R14_reg[19]/P0001  ;
	input \u2_R14_reg[1]/NET0131  ;
	input \u2_R14_reg[20]/NET0131  ;
	input \u2_R14_reg[21]/NET0131  ;
	input \u2_R14_reg[22]/P0001  ;
	input \u2_R14_reg[23]/P0001  ;
	input \u2_R14_reg[24]/NET0131  ;
	input \u2_R14_reg[25]/NET0131  ;
	input \u2_R14_reg[26]/P0001  ;
	input \u2_R14_reg[27]/P0001  ;
	input \u2_R14_reg[28]/NET0131  ;
	input \u2_R14_reg[29]/NET0131  ;
	input \u2_R14_reg[2]/NET0131  ;
	input \u2_R14_reg[30]/NET0131  ;
	input \u2_R14_reg[31]/P0001  ;
	input \u2_R14_reg[32]/NET0131  ;
	input \u2_R14_reg[3]/NET0131  ;
	input \u2_R14_reg[4]/NET0131  ;
	input \u2_R14_reg[5]/NET0131  ;
	input \u2_R14_reg[6]/NET0131  ;
	input \u2_R14_reg[7]/P0001  ;
	input \u2_R14_reg[8]/NET0131  ;
	input \u2_R14_reg[9]/NET0131  ;
	input \u2_R1_reg[10]/NET0131  ;
	input \u2_R1_reg[11]/P0001  ;
	input \u2_R1_reg[12]/NET0131  ;
	input \u2_R1_reg[13]/NET0131  ;
	input \u2_R1_reg[14]/NET0131  ;
	input \u2_R1_reg[15]/NET0131  ;
	input \u2_R1_reg[16]/NET0131  ;
	input \u2_R1_reg[17]/NET0131  ;
	input \u2_R1_reg[18]/NET0131  ;
	input \u2_R1_reg[19]/NET0131  ;
	input \u2_R1_reg[1]/NET0131  ;
	input \u2_R1_reg[20]/NET0131  ;
	input \u2_R1_reg[21]/NET0131  ;
	input \u2_R1_reg[22]/NET0131  ;
	input \u2_R1_reg[23]/NET0131  ;
	input \u2_R1_reg[24]/NET0131  ;
	input \u2_R1_reg[25]/NET0131  ;
	input \u2_R1_reg[26]/NET0131  ;
	input \u2_R1_reg[27]/NET0131  ;
	input \u2_R1_reg[28]/NET0131  ;
	input \u2_R1_reg[29]/NET0131  ;
	input \u2_R1_reg[2]/NET0131  ;
	input \u2_R1_reg[30]/NET0131  ;
	input \u2_R1_reg[31]/P0001  ;
	input \u2_R1_reg[32]/NET0131  ;
	input \u2_R1_reg[3]/NET0131  ;
	input \u2_R1_reg[4]/NET0131  ;
	input \u2_R1_reg[5]/NET0131  ;
	input \u2_R1_reg[6]/NET0131  ;
	input \u2_R1_reg[7]/NET0131  ;
	input \u2_R1_reg[8]/NET0131  ;
	input \u2_R1_reg[9]/NET0131  ;
	input \u2_R2_reg[10]/NET0131  ;
	input \u2_R2_reg[11]/NET0131  ;
	input \u2_R2_reg[12]/NET0131  ;
	input \u2_R2_reg[13]/NET0131  ;
	input \u2_R2_reg[14]/NET0131  ;
	input \u2_R2_reg[15]/NET0131  ;
	input \u2_R2_reg[16]/NET0131  ;
	input \u2_R2_reg[17]/NET0131  ;
	input \u2_R2_reg[18]/NET0131  ;
	input \u2_R2_reg[19]/NET0131  ;
	input \u2_R2_reg[1]/NET0131  ;
	input \u2_R2_reg[20]/NET0131  ;
	input \u2_R2_reg[21]/NET0131  ;
	input \u2_R2_reg[22]/NET0131  ;
	input \u2_R2_reg[23]/NET0131  ;
	input \u2_R2_reg[24]/NET0131  ;
	input \u2_R2_reg[25]/NET0131  ;
	input \u2_R2_reg[26]/NET0131  ;
	input \u2_R2_reg[27]/NET0131  ;
	input \u2_R2_reg[28]/NET0131  ;
	input \u2_R2_reg[29]/NET0131  ;
	input \u2_R2_reg[2]/NET0131  ;
	input \u2_R2_reg[30]/NET0131  ;
	input \u2_R2_reg[31]/P0001  ;
	input \u2_R2_reg[32]/NET0131  ;
	input \u2_R2_reg[3]/NET0131  ;
	input \u2_R2_reg[4]/NET0131  ;
	input \u2_R2_reg[5]/NET0131  ;
	input \u2_R2_reg[6]/NET0131  ;
	input \u2_R2_reg[7]/NET0131  ;
	input \u2_R2_reg[8]/NET0131  ;
	input \u2_R2_reg[9]/NET0131  ;
	input \u2_R3_reg[10]/NET0131  ;
	input \u2_R3_reg[11]/P0001  ;
	input \u2_R3_reg[12]/NET0131  ;
	input \u2_R3_reg[13]/NET0131  ;
	input \u2_R3_reg[14]/NET0131  ;
	input \u2_R3_reg[15]/NET0131  ;
	input \u2_R3_reg[16]/NET0131  ;
	input \u2_R3_reg[17]/NET0131  ;
	input \u2_R3_reg[18]/NET0131  ;
	input \u2_R3_reg[19]/NET0131  ;
	input \u2_R3_reg[1]/NET0131  ;
	input \u2_R3_reg[20]/NET0131  ;
	input \u2_R3_reg[21]/NET0131  ;
	input \u2_R3_reg[22]/NET0131  ;
	input \u2_R3_reg[23]/NET0131  ;
	input \u2_R3_reg[24]/NET0131  ;
	input \u2_R3_reg[25]/NET0131  ;
	input \u2_R3_reg[26]/NET0131  ;
	input \u2_R3_reg[27]/NET0131  ;
	input \u2_R3_reg[28]/NET0131  ;
	input \u2_R3_reg[29]/NET0131  ;
	input \u2_R3_reg[2]/NET0131  ;
	input \u2_R3_reg[30]/NET0131  ;
	input \u2_R3_reg[31]/P0001  ;
	input \u2_R3_reg[32]/NET0131  ;
	input \u2_R3_reg[3]/NET0131  ;
	input \u2_R3_reg[4]/NET0131  ;
	input \u2_R3_reg[5]/NET0131  ;
	input \u2_R3_reg[6]/NET0131  ;
	input \u2_R3_reg[7]/NET0131  ;
	input \u2_R3_reg[8]/NET0131  ;
	input \u2_R3_reg[9]/NET0131  ;
	input \u2_R4_reg[10]/NET0131  ;
	input \u2_R4_reg[11]/NET0131  ;
	input \u2_R4_reg[12]/NET0131  ;
	input \u2_R4_reg[13]/NET0131  ;
	input \u2_R4_reg[14]/NET0131  ;
	input \u2_R4_reg[15]/NET0131  ;
	input \u2_R4_reg[16]/NET0131  ;
	input \u2_R4_reg[17]/NET0131  ;
	input \u2_R4_reg[18]/NET0131  ;
	input \u2_R4_reg[19]/NET0131  ;
	input \u2_R4_reg[1]/NET0131  ;
	input \u2_R4_reg[20]/NET0131  ;
	input \u2_R4_reg[21]/NET0131  ;
	input \u2_R4_reg[22]/NET0131  ;
	input \u2_R4_reg[23]/NET0131  ;
	input \u2_R4_reg[24]/NET0131  ;
	input \u2_R4_reg[25]/NET0131  ;
	input \u2_R4_reg[26]/NET0131  ;
	input \u2_R4_reg[27]/NET0131  ;
	input \u2_R4_reg[28]/NET0131  ;
	input \u2_R4_reg[29]/NET0131  ;
	input \u2_R4_reg[2]/NET0131  ;
	input \u2_R4_reg[30]/NET0131  ;
	input \u2_R4_reg[31]/P0001  ;
	input \u2_R4_reg[32]/NET0131  ;
	input \u2_R4_reg[3]/NET0131  ;
	input \u2_R4_reg[4]/NET0131  ;
	input \u2_R4_reg[5]/NET0131  ;
	input \u2_R4_reg[6]/NET0131  ;
	input \u2_R4_reg[7]/NET0131  ;
	input \u2_R4_reg[8]/NET0131  ;
	input \u2_R4_reg[9]/NET0131  ;
	input \u2_R5_reg[10]/NET0131  ;
	input \u2_R5_reg[11]/NET0131  ;
	input \u2_R5_reg[12]/NET0131  ;
	input \u2_R5_reg[13]/NET0131  ;
	input \u2_R5_reg[14]/NET0131  ;
	input \u2_R5_reg[15]/NET0131  ;
	input \u2_R5_reg[16]/NET0131  ;
	input \u2_R5_reg[17]/NET0131  ;
	input \u2_R5_reg[18]/NET0131  ;
	input \u2_R5_reg[19]/NET0131  ;
	input \u2_R5_reg[1]/NET0131  ;
	input \u2_R5_reg[20]/NET0131  ;
	input \u2_R5_reg[21]/NET0131  ;
	input \u2_R5_reg[22]/NET0131  ;
	input \u2_R5_reg[23]/NET0131  ;
	input \u2_R5_reg[24]/NET0131  ;
	input \u2_R5_reg[25]/NET0131  ;
	input \u2_R5_reg[26]/NET0131  ;
	input \u2_R5_reg[27]/NET0131  ;
	input \u2_R5_reg[28]/NET0131  ;
	input \u2_R5_reg[29]/NET0131  ;
	input \u2_R5_reg[2]/NET0131  ;
	input \u2_R5_reg[30]/NET0131  ;
	input \u2_R5_reg[31]/P0001  ;
	input \u2_R5_reg[32]/NET0131  ;
	input \u2_R5_reg[3]/NET0131  ;
	input \u2_R5_reg[4]/NET0131  ;
	input \u2_R5_reg[5]/NET0131  ;
	input \u2_R5_reg[6]/NET0131  ;
	input \u2_R5_reg[7]/NET0131  ;
	input \u2_R5_reg[8]/NET0131  ;
	input \u2_R5_reg[9]/NET0131  ;
	input \u2_R6_reg[10]/NET0131  ;
	input \u2_R6_reg[11]/NET0131  ;
	input \u2_R6_reg[12]/NET0131  ;
	input \u2_R6_reg[13]/NET0131  ;
	input \u2_R6_reg[14]/NET0131  ;
	input \u2_R6_reg[15]/NET0131  ;
	input \u2_R6_reg[16]/NET0131  ;
	input \u2_R6_reg[17]/NET0131  ;
	input \u2_R6_reg[18]/NET0131  ;
	input \u2_R6_reg[19]/NET0131  ;
	input \u2_R6_reg[1]/NET0131  ;
	input \u2_R6_reg[20]/NET0131  ;
	input \u2_R6_reg[21]/NET0131  ;
	input \u2_R6_reg[22]/NET0131  ;
	input \u2_R6_reg[23]/NET0131  ;
	input \u2_R6_reg[24]/NET0131  ;
	input \u2_R6_reg[25]/NET0131  ;
	input \u2_R6_reg[26]/NET0131  ;
	input \u2_R6_reg[27]/NET0131  ;
	input \u2_R6_reg[28]/NET0131  ;
	input \u2_R6_reg[29]/NET0131  ;
	input \u2_R6_reg[2]/NET0131  ;
	input \u2_R6_reg[30]/NET0131  ;
	input \u2_R6_reg[31]/P0001  ;
	input \u2_R6_reg[32]/NET0131  ;
	input \u2_R6_reg[3]/NET0131  ;
	input \u2_R6_reg[4]/NET0131  ;
	input \u2_R6_reg[5]/NET0131  ;
	input \u2_R6_reg[6]/NET0131  ;
	input \u2_R6_reg[7]/NET0131  ;
	input \u2_R6_reg[8]/NET0131  ;
	input \u2_R6_reg[9]/NET0131  ;
	input \u2_R7_reg[10]/NET0131  ;
	input \u2_R7_reg[11]/NET0131  ;
	input \u2_R7_reg[12]/NET0131  ;
	input \u2_R7_reg[13]/NET0131  ;
	input \u2_R7_reg[14]/NET0131  ;
	input \u2_R7_reg[15]/NET0131  ;
	input \u2_R7_reg[16]/NET0131  ;
	input \u2_R7_reg[17]/NET0131  ;
	input \u2_R7_reg[18]/NET0131  ;
	input \u2_R7_reg[19]/NET0131  ;
	input \u2_R7_reg[1]/NET0131  ;
	input \u2_R7_reg[20]/NET0131  ;
	input \u2_R7_reg[21]/NET0131  ;
	input \u2_R7_reg[22]/NET0131  ;
	input \u2_R7_reg[23]/NET0131  ;
	input \u2_R7_reg[24]/NET0131  ;
	input \u2_R7_reg[25]/NET0131  ;
	input \u2_R7_reg[26]/NET0131  ;
	input \u2_R7_reg[27]/NET0131  ;
	input \u2_R7_reg[28]/NET0131  ;
	input \u2_R7_reg[29]/NET0131  ;
	input \u2_R7_reg[2]/NET0131  ;
	input \u2_R7_reg[30]/NET0131  ;
	input \u2_R7_reg[31]/P0001  ;
	input \u2_R7_reg[32]/NET0131  ;
	input \u2_R7_reg[3]/NET0131  ;
	input \u2_R7_reg[4]/NET0131  ;
	input \u2_R7_reg[5]/NET0131  ;
	input \u2_R7_reg[6]/NET0131  ;
	input \u2_R7_reg[7]/NET0131  ;
	input \u2_R7_reg[8]/NET0131  ;
	input \u2_R7_reg[9]/NET0131  ;
	input \u2_R8_reg[10]/NET0131  ;
	input \u2_R8_reg[11]/NET0131  ;
	input \u2_R8_reg[12]/NET0131  ;
	input \u2_R8_reg[13]/NET0131  ;
	input \u2_R8_reg[14]/NET0131  ;
	input \u2_R8_reg[15]/NET0131  ;
	input \u2_R8_reg[16]/NET0131  ;
	input \u2_R8_reg[17]/NET0131  ;
	input \u2_R8_reg[18]/NET0131  ;
	input \u2_R8_reg[19]/NET0131  ;
	input \u2_R8_reg[1]/NET0131  ;
	input \u2_R8_reg[20]/NET0131  ;
	input \u2_R8_reg[21]/NET0131  ;
	input \u2_R8_reg[22]/NET0131  ;
	input \u2_R8_reg[23]/NET0131  ;
	input \u2_R8_reg[24]/NET0131  ;
	input \u2_R8_reg[25]/NET0131  ;
	input \u2_R8_reg[26]/NET0131  ;
	input \u2_R8_reg[27]/NET0131  ;
	input \u2_R8_reg[28]/NET0131  ;
	input \u2_R8_reg[29]/NET0131  ;
	input \u2_R8_reg[2]/NET0131  ;
	input \u2_R8_reg[30]/NET0131  ;
	input \u2_R8_reg[31]/P0001  ;
	input \u2_R8_reg[32]/NET0131  ;
	input \u2_R8_reg[3]/NET0131  ;
	input \u2_R8_reg[4]/NET0131  ;
	input \u2_R8_reg[5]/NET0131  ;
	input \u2_R8_reg[6]/NET0131  ;
	input \u2_R8_reg[7]/NET0131  ;
	input \u2_R8_reg[8]/NET0131  ;
	input \u2_R8_reg[9]/NET0131  ;
	input \u2_R9_reg[10]/NET0131  ;
	input \u2_R9_reg[11]/NET0131  ;
	input \u2_R9_reg[12]/NET0131  ;
	input \u2_R9_reg[13]/NET0131  ;
	input \u2_R9_reg[14]/NET0131  ;
	input \u2_R9_reg[15]/NET0131  ;
	input \u2_R9_reg[16]/NET0131  ;
	input \u2_R9_reg[17]/NET0131  ;
	input \u2_R9_reg[18]/NET0131  ;
	input \u2_R9_reg[19]/NET0131  ;
	input \u2_R9_reg[1]/NET0131  ;
	input \u2_R9_reg[20]/NET0131  ;
	input \u2_R9_reg[21]/NET0131  ;
	input \u2_R9_reg[22]/NET0131  ;
	input \u2_R9_reg[23]/NET0131  ;
	input \u2_R9_reg[24]/NET0131  ;
	input \u2_R9_reg[25]/NET0131  ;
	input \u2_R9_reg[26]/NET0131  ;
	input \u2_R9_reg[27]/NET0131  ;
	input \u2_R9_reg[28]/NET0131  ;
	input \u2_R9_reg[29]/NET0131  ;
	input \u2_R9_reg[2]/NET0131  ;
	input \u2_R9_reg[30]/NET0131  ;
	input \u2_R9_reg[31]/P0001  ;
	input \u2_R9_reg[32]/NET0131  ;
	input \u2_R9_reg[3]/NET0131  ;
	input \u2_R9_reg[4]/NET0131  ;
	input \u2_R9_reg[5]/NET0131  ;
	input \u2_R9_reg[6]/NET0131  ;
	input \u2_R9_reg[7]/NET0131  ;
	input \u2_R9_reg[8]/NET0131  ;
	input \u2_R9_reg[9]/NET0131  ;
	input \u2_desIn_r_reg[0]/NET0131  ;
	input \u2_desIn_r_reg[10]/P0001  ;
	input \u2_desIn_r_reg[11]/NET0131  ;
	input \u2_desIn_r_reg[12]/NET0131  ;
	input \u2_desIn_r_reg[13]/NET0131  ;
	input \u2_desIn_r_reg[14]/NET0131  ;
	input \u2_desIn_r_reg[15]/NET0131  ;
	input \u2_desIn_r_reg[16]/NET0131  ;
	input \u2_desIn_r_reg[17]/NET0131  ;
	input \u2_desIn_r_reg[18]/NET0131  ;
	input \u2_desIn_r_reg[19]/NET0131  ;
	input \u2_desIn_r_reg[1]/NET0131  ;
	input \u2_desIn_r_reg[20]/NET0131  ;
	input \u2_desIn_r_reg[21]/NET0131  ;
	input \u2_desIn_r_reg[22]/NET0131  ;
	input \u2_desIn_r_reg[23]/NET0131  ;
	input \u2_desIn_r_reg[24]/NET0131  ;
	input \u2_desIn_r_reg[25]/NET0131  ;
	input \u2_desIn_r_reg[26]/NET0131  ;
	input \u2_desIn_r_reg[27]/NET0131  ;
	input \u2_desIn_r_reg[28]/NET0131  ;
	input \u2_desIn_r_reg[29]/NET0131  ;
	input \u2_desIn_r_reg[2]/NET0131  ;
	input \u2_desIn_r_reg[30]/NET0131  ;
	input \u2_desIn_r_reg[31]/NET0131  ;
	input \u2_desIn_r_reg[32]/NET0131  ;
	input \u2_desIn_r_reg[33]/NET0131  ;
	input \u2_desIn_r_reg[34]/NET0131  ;
	input \u2_desIn_r_reg[35]/NET0131  ;
	input \u2_desIn_r_reg[36]/NET0131  ;
	input \u2_desIn_r_reg[37]/NET0131  ;
	input \u2_desIn_r_reg[38]/NET0131  ;
	input \u2_desIn_r_reg[39]/NET0131  ;
	input \u2_desIn_r_reg[3]/NET0131  ;
	input \u2_desIn_r_reg[40]/NET0131  ;
	input \u2_desIn_r_reg[41]/NET0131  ;
	input \u2_desIn_r_reg[42]/NET0131  ;
	input \u2_desIn_r_reg[43]/NET0131  ;
	input \u2_desIn_r_reg[44]/NET0131  ;
	input \u2_desIn_r_reg[45]/NET0131  ;
	input \u2_desIn_r_reg[46]/NET0131  ;
	input \u2_desIn_r_reg[47]/NET0131  ;
	input \u2_desIn_r_reg[48]/NET0131  ;
	input \u2_desIn_r_reg[49]/NET0131  ;
	input \u2_desIn_r_reg[4]/NET0131  ;
	input \u2_desIn_r_reg[50]/NET0131  ;
	input \u2_desIn_r_reg[51]/NET0131  ;
	input \u2_desIn_r_reg[52]/NET0131  ;
	input \u2_desIn_r_reg[53]/NET0131  ;
	input \u2_desIn_r_reg[54]/NET0131  ;
	input \u2_desIn_r_reg[55]/NET0131  ;
	input \u2_desIn_r_reg[56]/NET0131  ;
	input \u2_desIn_r_reg[57]/NET0131  ;
	input \u2_desIn_r_reg[58]/NET0131  ;
	input \u2_desIn_r_reg[59]/NET0131  ;
	input \u2_desIn_r_reg[5]/NET0131  ;
	input \u2_desIn_r_reg[60]/NET0131  ;
	input \u2_desIn_r_reg[61]/NET0131  ;
	input \u2_desIn_r_reg[62]/NET0131  ;
	input \u2_desIn_r_reg[63]/NET0131  ;
	input \u2_desIn_r_reg[6]/NET0131  ;
	input \u2_desIn_r_reg[7]/NET0131  ;
	input \u2_desIn_r_reg[8]/NET0131  ;
	input \u2_desIn_r_reg[9]/NET0131  ;
	input \u2_key_r_reg[0]/NET0131  ;
	input \u2_key_r_reg[10]/NET0131  ;
	input \u2_key_r_reg[11]/NET0131  ;
	input \u2_key_r_reg[12]/NET0131  ;
	input \u2_key_r_reg[13]/NET0131  ;
	input \u2_key_r_reg[14]/NET0131  ;
	input \u2_key_r_reg[15]/NET0131  ;
	input \u2_key_r_reg[16]/NET0131  ;
	input \u2_key_r_reg[17]/NET0131  ;
	input \u2_key_r_reg[18]/NET0131  ;
	input \u2_key_r_reg[19]/NET0131  ;
	input \u2_key_r_reg[1]/NET0131  ;
	input \u2_key_r_reg[20]/NET0131  ;
	input \u2_key_r_reg[21]/NET0131  ;
	input \u2_key_r_reg[22]/NET0131  ;
	input \u2_key_r_reg[23]/NET0131  ;
	input \u2_key_r_reg[24]/NET0131  ;
	input \u2_key_r_reg[25]/NET0131  ;
	input \u2_key_r_reg[26]/NET0131  ;
	input \u2_key_r_reg[27]/NET0131  ;
	input \u2_key_r_reg[28]/NET0131  ;
	input \u2_key_r_reg[29]/NET0131  ;
	input \u2_key_r_reg[2]/NET0131  ;
	input \u2_key_r_reg[30]/NET0131  ;
	input \u2_key_r_reg[31]/NET0131  ;
	input \u2_key_r_reg[32]/NET0131  ;
	input \u2_key_r_reg[33]/NET0131  ;
	input \u2_key_r_reg[34]/NET0131  ;
	input \u2_key_r_reg[35]/P0001  ;
	input \u2_key_r_reg[36]/NET0131  ;
	input \u2_key_r_reg[37]/NET0131  ;
	input \u2_key_r_reg[38]/NET0131  ;
	input \u2_key_r_reg[39]/P0001  ;
	input \u2_key_r_reg[3]/NET0131  ;
	input \u2_key_r_reg[40]/NET0131  ;
	input \u2_key_r_reg[41]/NET0131  ;
	input \u2_key_r_reg[42]/P0001  ;
	input \u2_key_r_reg[43]/NET0131  ;
	input \u2_key_r_reg[44]/NET0131  ;
	input \u2_key_r_reg[45]/NET0131  ;
	input \u2_key_r_reg[46]/NET0131  ;
	input \u2_key_r_reg[47]/NET0131  ;
	input \u2_key_r_reg[48]/NET0131  ;
	input \u2_key_r_reg[49]/NET0131  ;
	input \u2_key_r_reg[4]/NET0131  ;
	input \u2_key_r_reg[50]/NET0131  ;
	input \u2_key_r_reg[51]/NET0131  ;
	input \u2_key_r_reg[52]/NET0131  ;
	input \u2_key_r_reg[53]/NET0131  ;
	input \u2_key_r_reg[54]/NET0131  ;
	input \u2_key_r_reg[55]/NET0131  ;
	input \u2_key_r_reg[5]/NET0131  ;
	input \u2_key_r_reg[6]/NET0131  ;
	input \u2_key_r_reg[7]/NET0131  ;
	input \u2_key_r_reg[8]/NET0131  ;
	input \u2_key_r_reg[9]/NET0131  ;
	input \u2_uk_K_r0_reg[0]/NET0131  ;
	input \u2_uk_K_r0_reg[10]/NET0131  ;
	input \u2_uk_K_r0_reg[11]/NET0131  ;
	input \u2_uk_K_r0_reg[12]/NET0131  ;
	input \u2_uk_K_r0_reg[13]/NET0131  ;
	input \u2_uk_K_r0_reg[14]/NET0131  ;
	input \u2_uk_K_r0_reg[15]/NET0131  ;
	input \u2_uk_K_r0_reg[16]/NET0131  ;
	input \u2_uk_K_r0_reg[17]/NET0131  ;
	input \u2_uk_K_r0_reg[18]/NET0131  ;
	input \u2_uk_K_r0_reg[19]/NET0131  ;
	input \u2_uk_K_r0_reg[20]/NET0131  ;
	input \u2_uk_K_r0_reg[21]/NET0131  ;
	input \u2_uk_K_r0_reg[22]/NET0131  ;
	input \u2_uk_K_r0_reg[23]/NET0131  ;
	input \u2_uk_K_r0_reg[24]/P0001  ;
	input \u2_uk_K_r0_reg[25]/P0001  ;
	input \u2_uk_K_r0_reg[26]/NET0131  ;
	input \u2_uk_K_r0_reg[27]/NET0131  ;
	input \u2_uk_K_r0_reg[28]/NET0131  ;
	input \u2_uk_K_r0_reg[29]/NET0131  ;
	input \u2_uk_K_r0_reg[2]/NET0131  ;
	input \u2_uk_K_r0_reg[30]/NET0131  ;
	input \u2_uk_K_r0_reg[31]/NET0131  ;
	input \u2_uk_K_r0_reg[32]/NET0131  ;
	input \u2_uk_K_r0_reg[33]/NET0131  ;
	input \u2_uk_K_r0_reg[34]/NET0131  ;
	input \u2_uk_K_r0_reg[35]/NET0131  ;
	input \u2_uk_K_r0_reg[36]/NET0131  ;
	input \u2_uk_K_r0_reg[37]/NET0131  ;
	input \u2_uk_K_r0_reg[38]/NET0131  ;
	input \u2_uk_K_r0_reg[39]/NET0131  ;
	input \u2_uk_K_r0_reg[3]/NET0131  ;
	input \u2_uk_K_r0_reg[40]/NET0131  ;
	input \u2_uk_K_r0_reg[41]/NET0131  ;
	input \u2_uk_K_r0_reg[42]/NET0131  ;
	input \u2_uk_K_r0_reg[43]/NET0131  ;
	input \u2_uk_K_r0_reg[44]/NET0131  ;
	input \u2_uk_K_r0_reg[45]/NET0131  ;
	input \u2_uk_K_r0_reg[46]/NET0131  ;
	input \u2_uk_K_r0_reg[47]/NET0131  ;
	input \u2_uk_K_r0_reg[48]/NET0131  ;
	input \u2_uk_K_r0_reg[49]/NET0131  ;
	input \u2_uk_K_r0_reg[4]/NET0131  ;
	input \u2_uk_K_r0_reg[50]/NET0131  ;
	input \u2_uk_K_r0_reg[51]/NET0131  ;
	input \u2_uk_K_r0_reg[52]/P0001  ;
	input \u2_uk_K_r0_reg[54]/NET0131  ;
	input \u2_uk_K_r0_reg[55]/NET0131  ;
	input \u2_uk_K_r0_reg[5]/NET0131  ;
	input \u2_uk_K_r0_reg[6]/NET0131  ;
	input \u2_uk_K_r0_reg[7]/NET0131  ;
	input \u2_uk_K_r0_reg[8]/NET0131  ;
	input \u2_uk_K_r0_reg[9]/NET0131  ;
	input \u2_uk_K_r10_reg[0]/NET0131  ;
	input \u2_uk_K_r10_reg[10]/NET0131  ;
	input \u2_uk_K_r10_reg[11]/NET0131  ;
	input \u2_uk_K_r10_reg[12]/NET0131  ;
	input \u2_uk_K_r10_reg[14]/NET0131  ;
	input \u2_uk_K_r10_reg[15]/NET0131  ;
	input \u2_uk_K_r10_reg[16]/NET0131  ;
	input \u2_uk_K_r10_reg[17]/NET0131  ;
	input \u2_uk_K_r10_reg[18]/NET0131  ;
	input \u2_uk_K_r10_reg[19]/NET0131  ;
	input \u2_uk_K_r10_reg[1]/NET0131  ;
	input \u2_uk_K_r10_reg[20]/NET0131  ;
	input \u2_uk_K_r10_reg[21]/NET0131  ;
	input \u2_uk_K_r10_reg[22]/NET0131  ;
	input \u2_uk_K_r10_reg[23]/NET0131  ;
	input \u2_uk_K_r10_reg[24]/NET0131  ;
	input \u2_uk_K_r10_reg[25]/NET0131  ;
	input \u2_uk_K_r10_reg[26]/NET0131  ;
	input \u2_uk_K_r10_reg[27]/NET0131  ;
	input \u2_uk_K_r10_reg[28]/NET0131  ;
	input \u2_uk_K_r10_reg[29]/NET0131  ;
	input \u2_uk_K_r10_reg[2]/NET0131  ;
	input \u2_uk_K_r10_reg[30]/NET0131  ;
	input \u2_uk_K_r10_reg[31]/NET0131  ;
	input \u2_uk_K_r10_reg[32]/NET0131  ;
	input \u2_uk_K_r10_reg[33]/NET0131  ;
	input \u2_uk_K_r10_reg[34]/NET0131  ;
	input \u2_uk_K_r10_reg[35]/NET0131  ;
	input \u2_uk_K_r10_reg[36]/NET0131  ;
	input \u2_uk_K_r10_reg[37]/NET0131  ;
	input \u2_uk_K_r10_reg[38]/NET0131  ;
	input \u2_uk_K_r10_reg[39]/NET0131  ;
	input \u2_uk_K_r10_reg[3]/NET0131  ;
	input \u2_uk_K_r10_reg[40]/NET0131  ;
	input \u2_uk_K_r10_reg[41]/NET0131  ;
	input \u2_uk_K_r10_reg[42]/NET0131  ;
	input \u2_uk_K_r10_reg[43]/NET0131  ;
	input \u2_uk_K_r10_reg[44]/NET0131  ;
	input \u2_uk_K_r10_reg[45]/P0001  ;
	input \u2_uk_K_r10_reg[46]/NET0131  ;
	input \u2_uk_K_r10_reg[47]/NET0131  ;
	input \u2_uk_K_r10_reg[48]/NET0131  ;
	input \u2_uk_K_r10_reg[49]/NET0131  ;
	input \u2_uk_K_r10_reg[4]/NET0131  ;
	input \u2_uk_K_r10_reg[50]/NET0131  ;
	input \u2_uk_K_r10_reg[51]/NET0131  ;
	input \u2_uk_K_r10_reg[52]/NET0131  ;
	input \u2_uk_K_r10_reg[53]/NET0131  ;
	input \u2_uk_K_r10_reg[54]/NET0131  ;
	input \u2_uk_K_r10_reg[55]/NET0131  ;
	input \u2_uk_K_r10_reg[5]/NET0131  ;
	input \u2_uk_K_r10_reg[6]/NET0131  ;
	input \u2_uk_K_r10_reg[7]/NET0131  ;
	input \u2_uk_K_r10_reg[8]/NET0131  ;
	input \u2_uk_K_r10_reg[9]/NET0131  ;
	input \u2_uk_K_r11_reg[0]/NET0131  ;
	input \u2_uk_K_r11_reg[10]/NET0131  ;
	input \u2_uk_K_r11_reg[11]/NET0131  ;
	input \u2_uk_K_r11_reg[12]/NET0131  ;
	input \u2_uk_K_r11_reg[13]/NET0131  ;
	input \u2_uk_K_r11_reg[14]/NET0131  ;
	input \u2_uk_K_r11_reg[15]/NET0131  ;
	input \u2_uk_K_r11_reg[16]/NET0131  ;
	input \u2_uk_K_r11_reg[17]/NET0131  ;
	input \u2_uk_K_r11_reg[18]/NET0131  ;
	input \u2_uk_K_r11_reg[19]/NET0131  ;
	input \u2_uk_K_r11_reg[1]/NET0131  ;
	input \u2_uk_K_r11_reg[20]/NET0131  ;
	input \u2_uk_K_r11_reg[21]/NET0131  ;
	input \u2_uk_K_r11_reg[22]/NET0131  ;
	input \u2_uk_K_r11_reg[23]/NET0131  ;
	input \u2_uk_K_r11_reg[24]/NET0131  ;
	input \u2_uk_K_r11_reg[25]/NET0131  ;
	input \u2_uk_K_r11_reg[26]/NET0131  ;
	input \u2_uk_K_r11_reg[27]/NET0131  ;
	input \u2_uk_K_r11_reg[28]/NET0131  ;
	input \u2_uk_K_r11_reg[29]/NET0131  ;
	input \u2_uk_K_r11_reg[2]/NET0131  ;
	input \u2_uk_K_r11_reg[31]/NET0131  ;
	input \u2_uk_K_r11_reg[32]/NET0131  ;
	input \u2_uk_K_r11_reg[33]/NET0131  ;
	input \u2_uk_K_r11_reg[34]/NET0131  ;
	input \u2_uk_K_r11_reg[35]/NET0131  ;
	input \u2_uk_K_r11_reg[36]/NET0131  ;
	input \u2_uk_K_r11_reg[37]/NET0131  ;
	input \u2_uk_K_r11_reg[38]/NET0131  ;
	input \u2_uk_K_r11_reg[39]/NET0131  ;
	input \u2_uk_K_r11_reg[3]/NET0131  ;
	input \u2_uk_K_r11_reg[40]/NET0131  ;
	input \u2_uk_K_r11_reg[41]/NET0131  ;
	input \u2_uk_K_r11_reg[42]/NET0131  ;
	input \u2_uk_K_r11_reg[43]/NET0131  ;
	input \u2_uk_K_r11_reg[44]/NET0131  ;
	input \u2_uk_K_r11_reg[45]/NET0131  ;
	input \u2_uk_K_r11_reg[46]/NET0131  ;
	input \u2_uk_K_r11_reg[47]/NET0131  ;
	input \u2_uk_K_r11_reg[48]/NET0131  ;
	input \u2_uk_K_r11_reg[49]/NET0131  ;
	input \u2_uk_K_r11_reg[4]/NET0131  ;
	input \u2_uk_K_r11_reg[50]/NET0131  ;
	input \u2_uk_K_r11_reg[51]/NET0131  ;
	input \u2_uk_K_r11_reg[52]/NET0131  ;
	input \u2_uk_K_r11_reg[53]/P0001  ;
	input \u2_uk_K_r11_reg[54]/NET0131  ;
	input \u2_uk_K_r11_reg[55]/NET0131  ;
	input \u2_uk_K_r11_reg[5]/NET0131  ;
	input \u2_uk_K_r11_reg[6]/NET0131  ;
	input \u2_uk_K_r11_reg[7]/NET0131  ;
	input \u2_uk_K_r11_reg[8]/NET0131  ;
	input \u2_uk_K_r11_reg[9]/NET0131  ;
	input \u2_uk_K_r12_reg[0]/NET0131  ;
	input \u2_uk_K_r12_reg[10]/P0001  ;
	input \u2_uk_K_r12_reg[11]/NET0131  ;
	input \u2_uk_K_r12_reg[12]/NET0131  ;
	input \u2_uk_K_r12_reg[13]/NET0131  ;
	input \u2_uk_K_r12_reg[14]/NET0131  ;
	input \u2_uk_K_r12_reg[15]/NET0131  ;
	input \u2_uk_K_r12_reg[16]/NET0131  ;
	input \u2_uk_K_r12_reg[17]/NET0131  ;
	input \u2_uk_K_r12_reg[18]/NET0131  ;
	input \u2_uk_K_r12_reg[19]/NET0131  ;
	input \u2_uk_K_r12_reg[1]/NET0131  ;
	input \u2_uk_K_r12_reg[20]/NET0131  ;
	input \u2_uk_K_r12_reg[21]/NET0131  ;
	input \u2_uk_K_r12_reg[22]/NET0131  ;
	input \u2_uk_K_r12_reg[23]/NET0131  ;
	input \u2_uk_K_r12_reg[24]/NET0131  ;
	input \u2_uk_K_r12_reg[25]/NET0131  ;
	input \u2_uk_K_r12_reg[26]/NET0131  ;
	input \u2_uk_K_r12_reg[27]/NET0131  ;
	input \u2_uk_K_r12_reg[28]/NET0131  ;
	input \u2_uk_K_r12_reg[29]/NET0131  ;
	input \u2_uk_K_r12_reg[2]/NET0131  ;
	input \u2_uk_K_r12_reg[30]/NET0131  ;
	input \u2_uk_K_r12_reg[31]/NET0131  ;
	input \u2_uk_K_r12_reg[32]/NET0131  ;
	input \u2_uk_K_r12_reg[33]/NET0131  ;
	input \u2_uk_K_r12_reg[34]/NET0131  ;
	input \u2_uk_K_r12_reg[35]/NET0131  ;
	input \u2_uk_K_r12_reg[36]/NET0131  ;
	input \u2_uk_K_r12_reg[37]/NET0131  ;
	input \u2_uk_K_r12_reg[38]/NET0131  ;
	input \u2_uk_K_r12_reg[3]/NET0131  ;
	input \u2_uk_K_r12_reg[40]/NET0131  ;
	input \u2_uk_K_r12_reg[41]/NET0131  ;
	input \u2_uk_K_r12_reg[42]/NET0131  ;
	input \u2_uk_K_r12_reg[43]/NET0131  ;
	input \u2_uk_K_r12_reg[44]/P0001  ;
	input \u2_uk_K_r12_reg[45]/NET0131  ;
	input \u2_uk_K_r12_reg[46]/NET0131  ;
	input \u2_uk_K_r12_reg[47]/NET0131  ;
	input \u2_uk_K_r12_reg[48]/NET0131  ;
	input \u2_uk_K_r12_reg[49]/NET0131  ;
	input \u2_uk_K_r12_reg[4]/NET0131  ;
	input \u2_uk_K_r12_reg[50]/NET0131  ;
	input \u2_uk_K_r12_reg[51]/NET0131  ;
	input \u2_uk_K_r12_reg[52]/NET0131  ;
	input \u2_uk_K_r12_reg[53]/NET0131  ;
	input \u2_uk_K_r12_reg[54]/NET0131  ;
	input \u2_uk_K_r12_reg[55]/NET0131  ;
	input \u2_uk_K_r12_reg[5]/NET0131  ;
	input \u2_uk_K_r12_reg[6]/NET0131  ;
	input \u2_uk_K_r12_reg[7]/P0001  ;
	input \u2_uk_K_r12_reg[8]/NET0131  ;
	input \u2_uk_K_r12_reg[9]/NET0131  ;
	input \u2_uk_K_r13_reg[0]/NET0131  ;
	input \u2_uk_K_r13_reg[10]/NET0131  ;
	input \u2_uk_K_r13_reg[11]/NET0131  ;
	input \u2_uk_K_r13_reg[12]/NET0131  ;
	input \u2_uk_K_r13_reg[13]/NET0131  ;
	input \u2_uk_K_r13_reg[14]/NET0131  ;
	input \u2_uk_K_r13_reg[15]/NET0131  ;
	input \u2_uk_K_r13_reg[16]/NET0131  ;
	input \u2_uk_K_r13_reg[17]/NET0131  ;
	input \u2_uk_K_r13_reg[18]/NET0131  ;
	input \u2_uk_K_r13_reg[19]/NET0131  ;
	input \u2_uk_K_r13_reg[20]/NET0131  ;
	input \u2_uk_K_r13_reg[21]/NET0131  ;
	input \u2_uk_K_r13_reg[22]/NET0131  ;
	input \u2_uk_K_r13_reg[23]/NET0131  ;
	input \u2_uk_K_r13_reg[24]/NET0131  ;
	input \u2_uk_K_r13_reg[25]/P0001  ;
	input \u2_uk_K_r13_reg[26]/NET0131  ;
	input \u2_uk_K_r13_reg[27]/NET0131  ;
	input \u2_uk_K_r13_reg[28]/NET0131  ;
	input \u2_uk_K_r13_reg[29]/NET0131  ;
	input \u2_uk_K_r13_reg[2]/NET0131  ;
	input \u2_uk_K_r13_reg[30]/NET0131  ;
	input \u2_uk_K_r13_reg[31]/NET0131  ;
	input \u2_uk_K_r13_reg[32]/NET0131  ;
	input \u2_uk_K_r13_reg[33]/NET0131  ;
	input \u2_uk_K_r13_reg[34]/NET0131  ;
	input \u2_uk_K_r13_reg[35]/NET0131  ;
	input \u2_uk_K_r13_reg[36]/NET0131  ;
	input \u2_uk_K_r13_reg[37]/NET0131  ;
	input \u2_uk_K_r13_reg[38]/NET0131  ;
	input \u2_uk_K_r13_reg[39]/NET0131  ;
	input \u2_uk_K_r13_reg[3]/NET0131  ;
	input \u2_uk_K_r13_reg[40]/NET0131  ;
	input \u2_uk_K_r13_reg[41]/NET0131  ;
	input \u2_uk_K_r13_reg[42]/NET0131  ;
	input \u2_uk_K_r13_reg[43]/NET0131  ;
	input \u2_uk_K_r13_reg[44]/NET0131  ;
	input \u2_uk_K_r13_reg[45]/NET0131  ;
	input \u2_uk_K_r13_reg[46]/NET0131  ;
	input \u2_uk_K_r13_reg[47]/NET0131  ;
	input \u2_uk_K_r13_reg[48]/NET0131  ;
	input \u2_uk_K_r13_reg[49]/NET0131  ;
	input \u2_uk_K_r13_reg[4]/NET0131  ;
	input \u2_uk_K_r13_reg[50]/NET0131  ;
	input \u2_uk_K_r13_reg[51]/NET0131  ;
	input \u2_uk_K_r13_reg[52]/NET0131  ;
	input \u2_uk_K_r13_reg[54]/NET0131  ;
	input \u2_uk_K_r13_reg[55]/NET0131  ;
	input \u2_uk_K_r13_reg[5]/NET0131  ;
	input \u2_uk_K_r13_reg[6]/NET0131  ;
	input \u2_uk_K_r13_reg[7]/NET0131  ;
	input \u2_uk_K_r13_reg[8]/NET0131  ;
	input \u2_uk_K_r13_reg[9]/NET0131  ;
	input \u2_uk_K_r14_reg[0]/NET0131  ;
	input \u2_uk_K_r14_reg[10]/P0001  ;
	input \u2_uk_K_r14_reg[11]/NET0131  ;
	input \u2_uk_K_r14_reg[12]/NET0131  ;
	input \u2_uk_K_r14_reg[13]/NET0131  ;
	input \u2_uk_K_r14_reg[14]/NET0131  ;
	input \u2_uk_K_r14_reg[15]/NET0131  ;
	input \u2_uk_K_r14_reg[16]/NET0131  ;
	input \u2_uk_K_r14_reg[17]/NET0131  ;
	input \u2_uk_K_r14_reg[18]/NET0131  ;
	input \u2_uk_K_r14_reg[19]/NET0131  ;
	input \u2_uk_K_r14_reg[1]/NET0131  ;
	input \u2_uk_K_r14_reg[20]/NET0131  ;
	input \u2_uk_K_r14_reg[21]/NET0131  ;
	input \u2_uk_K_r14_reg[22]/NET0131  ;
	input \u2_uk_K_r14_reg[23]/NET0131  ;
	input \u2_uk_K_r14_reg[24]/NET0131  ;
	input \u2_uk_K_r14_reg[25]/NET0131  ;
	input \u2_uk_K_r14_reg[26]/NET0131  ;
	input \u2_uk_K_r14_reg[27]/NET0131  ;
	input \u2_uk_K_r14_reg[28]/NET0131  ;
	input \u2_uk_K_r14_reg[29]/NET0131  ;
	input \u2_uk_K_r14_reg[2]/NET0131  ;
	input \u2_uk_K_r14_reg[30]/NET0131  ;
	input \u2_uk_K_r14_reg[31]/NET0131  ;
	input \u2_uk_K_r14_reg[32]/NET0131  ;
	input \u2_uk_K_r14_reg[33]/NET0131  ;
	input \u2_uk_K_r14_reg[34]/NET0131  ;
	input \u2_uk_K_r14_reg[35]/P0001  ;
	input \u2_uk_K_r14_reg[36]/NET0131  ;
	input \u2_uk_K_r14_reg[37]/NET0131  ;
	input \u2_uk_K_r14_reg[38]/NET0131  ;
	input \u2_uk_K_r14_reg[39]/P0001  ;
	input \u2_uk_K_r14_reg[3]/NET0131  ;
	input \u2_uk_K_r14_reg[40]/NET0131  ;
	input \u2_uk_K_r14_reg[41]/NET0131  ;
	input \u2_uk_K_r14_reg[42]/P0001  ;
	input \u2_uk_K_r14_reg[43]/NET0131  ;
	input \u2_uk_K_r14_reg[44]/NET0131  ;
	input \u2_uk_K_r14_reg[45]/NET0131  ;
	input \u2_uk_K_r14_reg[46]/NET0131  ;
	input \u2_uk_K_r14_reg[47]/NET0131  ;
	input \u2_uk_K_r14_reg[48]/NET0131  ;
	input \u2_uk_K_r14_reg[49]/P0001  ;
	input \u2_uk_K_r14_reg[4]/NET0131  ;
	input \u2_uk_K_r14_reg[50]/NET0131  ;
	input \u2_uk_K_r14_reg[51]/NET0131  ;
	input \u2_uk_K_r14_reg[52]/NET0131  ;
	input \u2_uk_K_r14_reg[53]/NET0131  ;
	input \u2_uk_K_r14_reg[54]/NET0131  ;
	input \u2_uk_K_r14_reg[55]/NET0131  ;
	input \u2_uk_K_r14_reg[5]/NET0131  ;
	input \u2_uk_K_r14_reg[6]/NET0131  ;
	input \u2_uk_K_r14_reg[7]/NET0131  ;
	input \u2_uk_K_r14_reg[8]/NET0131  ;
	input \u2_uk_K_r14_reg[9]/NET0131  ;
	input \u2_uk_K_r1_reg[0]/NET0131  ;
	input \u2_uk_K_r1_reg[10]/P0001  ;
	input \u2_uk_K_r1_reg[11]/NET0131  ;
	input \u2_uk_K_r1_reg[12]/NET0131  ;
	input \u2_uk_K_r1_reg[13]/NET0131  ;
	input \u2_uk_K_r1_reg[14]/NET0131  ;
	input \u2_uk_K_r1_reg[15]/NET0131  ;
	input \u2_uk_K_r1_reg[16]/NET0131  ;
	input \u2_uk_K_r1_reg[17]/NET0131  ;
	input \u2_uk_K_r1_reg[18]/NET0131  ;
	input \u2_uk_K_r1_reg[19]/NET0131  ;
	input \u2_uk_K_r1_reg[1]/NET0131  ;
	input \u2_uk_K_r1_reg[20]/NET0131  ;
	input \u2_uk_K_r1_reg[21]/NET0131  ;
	input \u2_uk_K_r1_reg[22]/NET0131  ;
	input \u2_uk_K_r1_reg[23]/NET0131  ;
	input \u2_uk_K_r1_reg[24]/NET0131  ;
	input \u2_uk_K_r1_reg[25]/NET0131  ;
	input \u2_uk_K_r1_reg[26]/NET0131  ;
	input \u2_uk_K_r1_reg[27]/NET0131  ;
	input \u2_uk_K_r1_reg[28]/NET0131  ;
	input \u2_uk_K_r1_reg[29]/NET0131  ;
	input \u2_uk_K_r1_reg[2]/NET0131  ;
	input \u2_uk_K_r1_reg[30]/NET0131  ;
	input \u2_uk_K_r1_reg[31]/NET0131  ;
	input \u2_uk_K_r1_reg[32]/NET0131  ;
	input \u2_uk_K_r1_reg[33]/NET0131  ;
	input \u2_uk_K_r1_reg[34]/NET0131  ;
	input \u2_uk_K_r1_reg[35]/NET0131  ;
	input \u2_uk_K_r1_reg[36]/NET0131  ;
	input \u2_uk_K_r1_reg[37]/NET0131  ;
	input \u2_uk_K_r1_reg[38]/NET0131  ;
	input \u2_uk_K_r1_reg[3]/NET0131  ;
	input \u2_uk_K_r1_reg[40]/NET0131  ;
	input \u2_uk_K_r1_reg[41]/NET0131  ;
	input \u2_uk_K_r1_reg[42]/NET0131  ;
	input \u2_uk_K_r1_reg[43]/NET0131  ;
	input \u2_uk_K_r1_reg[44]/P0001  ;
	input \u2_uk_K_r1_reg[45]/NET0131  ;
	input \u2_uk_K_r1_reg[46]/NET0131  ;
	input \u2_uk_K_r1_reg[47]/NET0131  ;
	input \u2_uk_K_r1_reg[48]/NET0131  ;
	input \u2_uk_K_r1_reg[49]/NET0131  ;
	input \u2_uk_K_r1_reg[4]/NET0131  ;
	input \u2_uk_K_r1_reg[50]/NET0131  ;
	input \u2_uk_K_r1_reg[51]/NET0131  ;
	input \u2_uk_K_r1_reg[52]/NET0131  ;
	input \u2_uk_K_r1_reg[53]/NET0131  ;
	input \u2_uk_K_r1_reg[54]/NET0131  ;
	input \u2_uk_K_r1_reg[55]/NET0131  ;
	input \u2_uk_K_r1_reg[5]/NET0131  ;
	input \u2_uk_K_r1_reg[6]/NET0131  ;
	input \u2_uk_K_r1_reg[7]/P0001  ;
	input \u2_uk_K_r1_reg[8]/NET0131  ;
	input \u2_uk_K_r1_reg[9]/NET0131  ;
	input \u2_uk_K_r2_reg[0]/NET0131  ;
	input \u2_uk_K_r2_reg[10]/NET0131  ;
	input \u2_uk_K_r2_reg[11]/NET0131  ;
	input \u2_uk_K_r2_reg[12]/NET0131  ;
	input \u2_uk_K_r2_reg[13]/NET0131  ;
	input \u2_uk_K_r2_reg[14]/NET0131  ;
	input \u2_uk_K_r2_reg[15]/NET0131  ;
	input \u2_uk_K_r2_reg[16]/NET0131  ;
	input \u2_uk_K_r2_reg[17]/NET0131  ;
	input \u2_uk_K_r2_reg[18]/NET0131  ;
	input \u2_uk_K_r2_reg[19]/NET0131  ;
	input \u2_uk_K_r2_reg[1]/NET0131  ;
	input \u2_uk_K_r2_reg[20]/NET0131  ;
	input \u2_uk_K_r2_reg[21]/NET0131  ;
	input \u2_uk_K_r2_reg[22]/NET0131  ;
	input \u2_uk_K_r2_reg[23]/NET0131  ;
	input \u2_uk_K_r2_reg[24]/NET0131  ;
	input \u2_uk_K_r2_reg[25]/NET0131  ;
	input \u2_uk_K_r2_reg[26]/NET0131  ;
	input \u2_uk_K_r2_reg[27]/NET0131  ;
	input \u2_uk_K_r2_reg[28]/NET0131  ;
	input \u2_uk_K_r2_reg[29]/NET0131  ;
	input \u2_uk_K_r2_reg[2]/NET0131  ;
	input \u2_uk_K_r2_reg[31]/NET0131  ;
	input \u2_uk_K_r2_reg[32]/NET0131  ;
	input \u2_uk_K_r2_reg[33]/NET0131  ;
	input \u2_uk_K_r2_reg[34]/NET0131  ;
	input \u2_uk_K_r2_reg[35]/NET0131  ;
	input \u2_uk_K_r2_reg[36]/NET0131  ;
	input \u2_uk_K_r2_reg[37]/NET0131  ;
	input \u2_uk_K_r2_reg[38]/NET0131  ;
	input \u2_uk_K_r2_reg[39]/NET0131  ;
	input \u2_uk_K_r2_reg[3]/NET0131  ;
	input \u2_uk_K_r2_reg[40]/NET0131  ;
	input \u2_uk_K_r2_reg[41]/NET0131  ;
	input \u2_uk_K_r2_reg[42]/NET0131  ;
	input \u2_uk_K_r2_reg[43]/NET0131  ;
	input \u2_uk_K_r2_reg[44]/NET0131  ;
	input \u2_uk_K_r2_reg[45]/NET0131  ;
	input \u2_uk_K_r2_reg[46]/NET0131  ;
	input \u2_uk_K_r2_reg[47]/NET0131  ;
	input \u2_uk_K_r2_reg[48]/NET0131  ;
	input \u2_uk_K_r2_reg[49]/NET0131  ;
	input \u2_uk_K_r2_reg[4]/NET0131  ;
	input \u2_uk_K_r2_reg[50]/NET0131  ;
	input \u2_uk_K_r2_reg[51]/NET0131  ;
	input \u2_uk_K_r2_reg[52]/NET0131  ;
	input \u2_uk_K_r2_reg[53]/P0001  ;
	input \u2_uk_K_r2_reg[54]/NET0131  ;
	input \u2_uk_K_r2_reg[55]/NET0131  ;
	input \u2_uk_K_r2_reg[5]/NET0131  ;
	input \u2_uk_K_r2_reg[6]/NET0131  ;
	input \u2_uk_K_r2_reg[7]/NET0131  ;
	input \u2_uk_K_r2_reg[8]/NET0131  ;
	input \u2_uk_K_r2_reg[9]/NET0131  ;
	input \u2_uk_K_r3_reg[0]/NET0131  ;
	input \u2_uk_K_r3_reg[10]/NET0131  ;
	input \u2_uk_K_r3_reg[11]/NET0131  ;
	input \u2_uk_K_r3_reg[12]/NET0131  ;
	input \u2_uk_K_r3_reg[14]/NET0131  ;
	input \u2_uk_K_r3_reg[15]/NET0131  ;
	input \u2_uk_K_r3_reg[16]/NET0131  ;
	input \u2_uk_K_r3_reg[17]/NET0131  ;
	input \u2_uk_K_r3_reg[18]/NET0131  ;
	input \u2_uk_K_r3_reg[19]/NET0131  ;
	input \u2_uk_K_r3_reg[1]/NET0131  ;
	input \u2_uk_K_r3_reg[20]/NET0131  ;
	input \u2_uk_K_r3_reg[21]/NET0131  ;
	input \u2_uk_K_r3_reg[22]/NET0131  ;
	input \u2_uk_K_r3_reg[23]/NET0131  ;
	input \u2_uk_K_r3_reg[24]/NET0131  ;
	input \u2_uk_K_r3_reg[25]/NET0131  ;
	input \u2_uk_K_r3_reg[26]/NET0131  ;
	input \u2_uk_K_r3_reg[27]/NET0131  ;
	input \u2_uk_K_r3_reg[28]/NET0131  ;
	input \u2_uk_K_r3_reg[29]/NET0131  ;
	input \u2_uk_K_r3_reg[2]/NET0131  ;
	input \u2_uk_K_r3_reg[30]/NET0131  ;
	input \u2_uk_K_r3_reg[31]/NET0131  ;
	input \u2_uk_K_r3_reg[32]/NET0131  ;
	input \u2_uk_K_r3_reg[33]/NET0131  ;
	input \u2_uk_K_r3_reg[34]/NET0131  ;
	input \u2_uk_K_r3_reg[35]/NET0131  ;
	input \u2_uk_K_r3_reg[36]/NET0131  ;
	input \u2_uk_K_r3_reg[37]/NET0131  ;
	input \u2_uk_K_r3_reg[38]/NET0131  ;
	input \u2_uk_K_r3_reg[39]/NET0131  ;
	input \u2_uk_K_r3_reg[3]/NET0131  ;
	input \u2_uk_K_r3_reg[40]/NET0131  ;
	input \u2_uk_K_r3_reg[41]/NET0131  ;
	input \u2_uk_K_r3_reg[42]/NET0131  ;
	input \u2_uk_K_r3_reg[43]/NET0131  ;
	input \u2_uk_K_r3_reg[44]/NET0131  ;
	input \u2_uk_K_r3_reg[45]/P0001  ;
	input \u2_uk_K_r3_reg[46]/NET0131  ;
	input \u2_uk_K_r3_reg[47]/NET0131  ;
	input \u2_uk_K_r3_reg[48]/NET0131  ;
	input \u2_uk_K_r3_reg[49]/NET0131  ;
	input \u2_uk_K_r3_reg[4]/NET0131  ;
	input \u2_uk_K_r3_reg[50]/NET0131  ;
	input \u2_uk_K_r3_reg[51]/NET0131  ;
	input \u2_uk_K_r3_reg[52]/NET0131  ;
	input \u2_uk_K_r3_reg[53]/NET0131  ;
	input \u2_uk_K_r3_reg[54]/NET0131  ;
	input \u2_uk_K_r3_reg[55]/NET0131  ;
	input \u2_uk_K_r3_reg[5]/NET0131  ;
	input \u2_uk_K_r3_reg[6]/NET0131  ;
	input \u2_uk_K_r3_reg[7]/NET0131  ;
	input \u2_uk_K_r3_reg[8]/NET0131  ;
	input \u2_uk_K_r3_reg[9]/NET0131  ;
	input \u2_uk_K_r4_reg[0]/P0001  ;
	input \u2_uk_K_r4_reg[10]/NET0131  ;
	input \u2_uk_K_r4_reg[11]/NET0131  ;
	input \u2_uk_K_r4_reg[12]/NET0131  ;
	input \u2_uk_K_r4_reg[13]/NET0131  ;
	input \u2_uk_K_r4_reg[14]/NET0131  ;
	input \u2_uk_K_r4_reg[15]/NET0131  ;
	input \u2_uk_K_r4_reg[16]/NET0131  ;
	input \u2_uk_K_r4_reg[17]/NET0131  ;
	input \u2_uk_K_r4_reg[18]/NET0131  ;
	input \u2_uk_K_r4_reg[19]/NET0131  ;
	input \u2_uk_K_r4_reg[1]/NET0131  ;
	input \u2_uk_K_r4_reg[20]/NET0131  ;
	input \u2_uk_K_r4_reg[21]/NET0131  ;
	input \u2_uk_K_r4_reg[22]/NET0131  ;
	input \u2_uk_K_r4_reg[23]/NET0131  ;
	input \u2_uk_K_r4_reg[25]/NET0131  ;
	input \u2_uk_K_r4_reg[26]/NET0131  ;
	input \u2_uk_K_r4_reg[27]/P0001  ;
	input \u2_uk_K_r4_reg[28]/NET0131  ;
	input \u2_uk_K_r4_reg[29]/NET0131  ;
	input \u2_uk_K_r4_reg[30]/NET0131  ;
	input \u2_uk_K_r4_reg[31]/P0001  ;
	input \u2_uk_K_r4_reg[32]/NET0131  ;
	input \u2_uk_K_r4_reg[33]/NET0131  ;
	input \u2_uk_K_r4_reg[34]/NET0131  ;
	input \u2_uk_K_r4_reg[35]/NET0131  ;
	input \u2_uk_K_r4_reg[36]/NET0131  ;
	input \u2_uk_K_r4_reg[37]/NET0131  ;
	input \u2_uk_K_r4_reg[38]/NET0131  ;
	input \u2_uk_K_r4_reg[39]/NET0131  ;
	input \u2_uk_K_r4_reg[3]/NET0131  ;
	input \u2_uk_K_r4_reg[40]/NET0131  ;
	input \u2_uk_K_r4_reg[41]/NET0131  ;
	input \u2_uk_K_r4_reg[42]/NET0131  ;
	input \u2_uk_K_r4_reg[43]/NET0131  ;
	input \u2_uk_K_r4_reg[44]/NET0131  ;
	input \u2_uk_K_r4_reg[45]/NET0131  ;
	input \u2_uk_K_r4_reg[46]/NET0131  ;
	input \u2_uk_K_r4_reg[47]/NET0131  ;
	input \u2_uk_K_r4_reg[48]/NET0131  ;
	input \u2_uk_K_r4_reg[49]/NET0131  ;
	input \u2_uk_K_r4_reg[4]/NET0131  ;
	input \u2_uk_K_r4_reg[50]/NET0131  ;
	input \u2_uk_K_r4_reg[51]/NET0131  ;
	input \u2_uk_K_r4_reg[52]/NET0131  ;
	input \u2_uk_K_r4_reg[53]/NET0131  ;
	input \u2_uk_K_r4_reg[54]/NET0131  ;
	input \u2_uk_K_r4_reg[55]/NET0131  ;
	input \u2_uk_K_r4_reg[5]/NET0131  ;
	input \u2_uk_K_r4_reg[6]/NET0131  ;
	input \u2_uk_K_r4_reg[7]/NET0131  ;
	input \u2_uk_K_r4_reg[8]/NET0131  ;
	input \u2_uk_K_r4_reg[9]/NET0131  ;
	input \u2_uk_K_r5_reg[0]/NET0131  ;
	input \u2_uk_K_r5_reg[10]/NET0131  ;
	input \u2_uk_K_r5_reg[11]/NET0131  ;
	input \u2_uk_K_r5_reg[12]/NET0131  ;
	input \u2_uk_K_r5_reg[13]/P0001  ;
	input \u2_uk_K_r5_reg[14]/NET0131  ;
	input \u2_uk_K_r5_reg[15]/NET0131  ;
	input \u2_uk_K_r5_reg[16]/NET0131  ;
	input \u2_uk_K_r5_reg[17]/NET0131  ;
	input \u2_uk_K_r5_reg[18]/NET0131  ;
	input \u2_uk_K_r5_reg[19]/NET0131  ;
	input \u2_uk_K_r5_reg[1]/NET0131  ;
	input \u2_uk_K_r5_reg[20]/NET0131  ;
	input \u2_uk_K_r5_reg[21]/NET0131  ;
	input \u2_uk_K_r5_reg[22]/NET0131  ;
	input \u2_uk_K_r5_reg[23]/NET0131  ;
	input \u2_uk_K_r5_reg[24]/NET0131  ;
	input \u2_uk_K_r5_reg[25]/NET0131  ;
	input \u2_uk_K_r5_reg[26]/NET0131  ;
	input \u2_uk_K_r5_reg[27]/NET0131  ;
	input \u2_uk_K_r5_reg[28]/NET0131  ;
	input \u2_uk_K_r5_reg[29]/NET0131  ;
	input \u2_uk_K_r5_reg[2]/NET0131  ;
	input \u2_uk_K_r5_reg[30]/NET0131  ;
	input \u2_uk_K_r5_reg[31]/NET0131  ;
	input \u2_uk_K_r5_reg[32]/NET0131  ;
	input \u2_uk_K_r5_reg[33]/NET0131  ;
	input \u2_uk_K_r5_reg[34]/NET0131  ;
	input \u2_uk_K_r5_reg[35]/NET0131  ;
	input \u2_uk_K_r5_reg[36]/NET0131  ;
	input \u2_uk_K_r5_reg[37]/P0001  ;
	input \u2_uk_K_r5_reg[38]/NET0131  ;
	input \u2_uk_K_r5_reg[39]/NET0131  ;
	input \u2_uk_K_r5_reg[3]/NET0131  ;
	input \u2_uk_K_r5_reg[40]/NET0131  ;
	input \u2_uk_K_r5_reg[41]/NET0131  ;
	input \u2_uk_K_r5_reg[42]/NET0131  ;
	input \u2_uk_K_r5_reg[43]/NET0131  ;
	input \u2_uk_K_r5_reg[44]/NET0131  ;
	input \u2_uk_K_r5_reg[46]/NET0131  ;
	input \u2_uk_K_r5_reg[47]/NET0131  ;
	input \u2_uk_K_r5_reg[48]/NET0131  ;
	input \u2_uk_K_r5_reg[49]/NET0131  ;
	input \u2_uk_K_r5_reg[4]/NET0131  ;
	input \u2_uk_K_r5_reg[50]/NET0131  ;
	input \u2_uk_K_r5_reg[51]/NET0131  ;
	input \u2_uk_K_r5_reg[52]/NET0131  ;
	input \u2_uk_K_r5_reg[53]/NET0131  ;
	input \u2_uk_K_r5_reg[54]/NET0131  ;
	input \u2_uk_K_r5_reg[55]/NET0131  ;
	input \u2_uk_K_r5_reg[5]/NET0131  ;
	input \u2_uk_K_r5_reg[6]/NET0131  ;
	input \u2_uk_K_r5_reg[7]/NET0131  ;
	input \u2_uk_K_r5_reg[8]/NET0131  ;
	input \u2_uk_K_r5_reg[9]/P0001  ;
	input \u2_uk_K_r6_reg[0]/NET0131  ;
	input \u2_uk_K_r6_reg[10]/NET0131  ;
	input \u2_uk_K_r6_reg[11]/NET0131  ;
	input \u2_uk_K_r6_reg[12]/NET0131  ;
	input \u2_uk_K_r6_reg[13]/NET0131  ;
	input \u2_uk_K_r6_reg[14]/NET0131  ;
	input \u2_uk_K_r6_reg[15]/NET0131  ;
	input \u2_uk_K_r6_reg[16]/NET0131  ;
	input \u2_uk_K_r6_reg[17]/NET0131  ;
	input \u2_uk_K_r6_reg[18]/NET0131  ;
	input \u2_uk_K_r6_reg[19]/NET0131  ;
	input \u2_uk_K_r6_reg[1]/NET0131  ;
	input \u2_uk_K_r6_reg[20]/NET0131  ;
	input \u2_uk_K_r6_reg[21]/NET0131  ;
	input \u2_uk_K_r6_reg[22]/NET0131  ;
	input \u2_uk_K_r6_reg[23]/P0001  ;
	input \u2_uk_K_r6_reg[24]/NET0131  ;
	input \u2_uk_K_r6_reg[25]/NET0131  ;
	input \u2_uk_K_r6_reg[26]/NET0131  ;
	input \u2_uk_K_r6_reg[27]/NET0131  ;
	input \u2_uk_K_r6_reg[28]/NET0131  ;
	input \u2_uk_K_r6_reg[29]/NET0131  ;
	input \u2_uk_K_r6_reg[2]/NET0131  ;
	input \u2_uk_K_r6_reg[30]/P0001  ;
	input \u2_uk_K_r6_reg[31]/NET0131  ;
	input \u2_uk_K_r6_reg[32]/NET0131  ;
	input \u2_uk_K_r6_reg[33]/NET0131  ;
	input \u2_uk_K_r6_reg[34]/NET0131  ;
	input \u2_uk_K_r6_reg[35]/NET0131  ;
	input \u2_uk_K_r6_reg[36]/NET0131  ;
	input \u2_uk_K_r6_reg[37]/NET0131  ;
	input \u2_uk_K_r6_reg[38]/NET0131  ;
	input \u2_uk_K_r6_reg[39]/NET0131  ;
	input \u2_uk_K_r6_reg[3]/NET0131  ;
	input \u2_uk_K_r6_reg[40]/NET0131  ;
	input \u2_uk_K_r6_reg[41]/NET0131  ;
	input \u2_uk_K_r6_reg[42]/NET0131  ;
	input \u2_uk_K_r6_reg[43]/NET0131  ;
	input \u2_uk_K_r6_reg[44]/NET0131  ;
	input \u2_uk_K_r6_reg[45]/NET0131  ;
	input \u2_uk_K_r6_reg[46]/NET0131  ;
	input \u2_uk_K_r6_reg[47]/NET0131  ;
	input \u2_uk_K_r6_reg[48]/NET0131  ;
	input \u2_uk_K_r6_reg[49]/NET0131  ;
	input \u2_uk_K_r6_reg[4]/NET0131  ;
	input \u2_uk_K_r6_reg[50]/NET0131  ;
	input \u2_uk_K_r6_reg[51]/NET0131  ;
	input \u2_uk_K_r6_reg[52]/NET0131  ;
	input \u2_uk_K_r6_reg[53]/NET0131  ;
	input \u2_uk_K_r6_reg[54]/NET0131  ;
	input \u2_uk_K_r6_reg[55]/P0001  ;
	input \u2_uk_K_r6_reg[5]/NET0131  ;
	input \u2_uk_K_r6_reg[6]/NET0131  ;
	input \u2_uk_K_r6_reg[7]/NET0131  ;
	input \u2_uk_K_r6_reg[8]/NET0131  ;
	input \u2_uk_K_r6_reg[9]/NET0131  ;
	input \u2_uk_K_r7_reg[0]/NET0131  ;
	input \u2_uk_K_r7_reg[10]/NET0131  ;
	input \u2_uk_K_r7_reg[11]/NET0131  ;
	input \u2_uk_K_r7_reg[12]/NET0131  ;
	input \u2_uk_K_r7_reg[13]/NET0131  ;
	input \u2_uk_K_r7_reg[14]/NET0131  ;
	input \u2_uk_K_r7_reg[15]/NET0131  ;
	input \u2_uk_K_r7_reg[16]/NET0131  ;
	input \u2_uk_K_r7_reg[17]/NET0131  ;
	input \u2_uk_K_r7_reg[18]/NET0131  ;
	input \u2_uk_K_r7_reg[19]/NET0131  ;
	input \u2_uk_K_r7_reg[1]/NET0131  ;
	input \u2_uk_K_r7_reg[20]/NET0131  ;
	input \u2_uk_K_r7_reg[21]/NET0131  ;
	input \u2_uk_K_r7_reg[22]/NET0131  ;
	input \u2_uk_K_r7_reg[23]/P0001  ;
	input \u2_uk_K_r7_reg[24]/NET0131  ;
	input \u2_uk_K_r7_reg[25]/NET0131  ;
	input \u2_uk_K_r7_reg[26]/NET0131  ;
	input \u2_uk_K_r7_reg[27]/NET0131  ;
	input \u2_uk_K_r7_reg[28]/NET0131  ;
	input \u2_uk_K_r7_reg[29]/NET0131  ;
	input \u2_uk_K_r7_reg[2]/NET0131  ;
	input \u2_uk_K_r7_reg[30]/P0001  ;
	input \u2_uk_K_r7_reg[31]/NET0131  ;
	input \u2_uk_K_r7_reg[32]/NET0131  ;
	input \u2_uk_K_r7_reg[33]/NET0131  ;
	input \u2_uk_K_r7_reg[34]/NET0131  ;
	input \u2_uk_K_r7_reg[35]/NET0131  ;
	input \u2_uk_K_r7_reg[36]/NET0131  ;
	input \u2_uk_K_r7_reg[37]/NET0131  ;
	input \u2_uk_K_r7_reg[38]/NET0131  ;
	input \u2_uk_K_r7_reg[39]/NET0131  ;
	input \u2_uk_K_r7_reg[3]/NET0131  ;
	input \u2_uk_K_r7_reg[40]/NET0131  ;
	input \u2_uk_K_r7_reg[41]/NET0131  ;
	input \u2_uk_K_r7_reg[42]/NET0131  ;
	input \u2_uk_K_r7_reg[43]/NET0131  ;
	input \u2_uk_K_r7_reg[44]/NET0131  ;
	input \u2_uk_K_r7_reg[45]/NET0131  ;
	input \u2_uk_K_r7_reg[46]/NET0131  ;
	input \u2_uk_K_r7_reg[47]/NET0131  ;
	input \u2_uk_K_r7_reg[48]/NET0131  ;
	input \u2_uk_K_r7_reg[49]/NET0131  ;
	input \u2_uk_K_r7_reg[4]/NET0131  ;
	input \u2_uk_K_r7_reg[50]/NET0131  ;
	input \u2_uk_K_r7_reg[51]/NET0131  ;
	input \u2_uk_K_r7_reg[52]/NET0131  ;
	input \u2_uk_K_r7_reg[53]/NET0131  ;
	input \u2_uk_K_r7_reg[54]/NET0131  ;
	input \u2_uk_K_r7_reg[55]/P0001  ;
	input \u2_uk_K_r7_reg[5]/NET0131  ;
	input \u2_uk_K_r7_reg[6]/NET0131  ;
	input \u2_uk_K_r7_reg[7]/NET0131  ;
	input \u2_uk_K_r7_reg[8]/NET0131  ;
	input \u2_uk_K_r7_reg[9]/NET0131  ;
	input \u2_uk_K_r8_reg[0]/NET0131  ;
	input \u2_uk_K_r8_reg[10]/NET0131  ;
	input \u2_uk_K_r8_reg[11]/NET0131  ;
	input \u2_uk_K_r8_reg[12]/NET0131  ;
	input \u2_uk_K_r8_reg[13]/P0001  ;
	input \u2_uk_K_r8_reg[14]/NET0131  ;
	input \u2_uk_K_r8_reg[15]/NET0131  ;
	input \u2_uk_K_r8_reg[16]/NET0131  ;
	input \u2_uk_K_r8_reg[17]/NET0131  ;
	input \u2_uk_K_r8_reg[18]/NET0131  ;
	input \u2_uk_K_r8_reg[19]/NET0131  ;
	input \u2_uk_K_r8_reg[1]/NET0131  ;
	input \u2_uk_K_r8_reg[20]/NET0131  ;
	input \u2_uk_K_r8_reg[21]/NET0131  ;
	input \u2_uk_K_r8_reg[22]/NET0131  ;
	input \u2_uk_K_r8_reg[23]/NET0131  ;
	input \u2_uk_K_r8_reg[24]/NET0131  ;
	input \u2_uk_K_r8_reg[25]/NET0131  ;
	input \u2_uk_K_r8_reg[26]/NET0131  ;
	input \u2_uk_K_r8_reg[27]/NET0131  ;
	input \u2_uk_K_r8_reg[28]/NET0131  ;
	input \u2_uk_K_r8_reg[29]/NET0131  ;
	input \u2_uk_K_r8_reg[2]/NET0131  ;
	input \u2_uk_K_r8_reg[30]/NET0131  ;
	input \u2_uk_K_r8_reg[31]/NET0131  ;
	input \u2_uk_K_r8_reg[32]/NET0131  ;
	input \u2_uk_K_r8_reg[33]/NET0131  ;
	input \u2_uk_K_r8_reg[34]/NET0131  ;
	input \u2_uk_K_r8_reg[35]/NET0131  ;
	input \u2_uk_K_r8_reg[36]/NET0131  ;
	input \u2_uk_K_r8_reg[37]/P0001  ;
	input \u2_uk_K_r8_reg[38]/NET0131  ;
	input \u2_uk_K_r8_reg[39]/NET0131  ;
	input \u2_uk_K_r8_reg[3]/NET0131  ;
	input \u2_uk_K_r8_reg[40]/NET0131  ;
	input \u2_uk_K_r8_reg[41]/NET0131  ;
	input \u2_uk_K_r8_reg[42]/NET0131  ;
	input \u2_uk_K_r8_reg[43]/NET0131  ;
	input \u2_uk_K_r8_reg[44]/NET0131  ;
	input \u2_uk_K_r8_reg[46]/NET0131  ;
	input \u2_uk_K_r8_reg[47]/NET0131  ;
	input \u2_uk_K_r8_reg[48]/NET0131  ;
	input \u2_uk_K_r8_reg[49]/NET0131  ;
	input \u2_uk_K_r8_reg[4]/NET0131  ;
	input \u2_uk_K_r8_reg[50]/NET0131  ;
	input \u2_uk_K_r8_reg[51]/NET0131  ;
	input \u2_uk_K_r8_reg[52]/NET0131  ;
	input \u2_uk_K_r8_reg[53]/NET0131  ;
	input \u2_uk_K_r8_reg[54]/NET0131  ;
	input \u2_uk_K_r8_reg[55]/NET0131  ;
	input \u2_uk_K_r8_reg[5]/NET0131  ;
	input \u2_uk_K_r8_reg[6]/NET0131  ;
	input \u2_uk_K_r8_reg[7]/NET0131  ;
	input \u2_uk_K_r8_reg[8]/NET0131  ;
	input \u2_uk_K_r8_reg[9]/NET0131  ;
	input \u2_uk_K_r9_reg[0]/P0001  ;
	input \u2_uk_K_r9_reg[10]/NET0131  ;
	input \u2_uk_K_r9_reg[11]/NET0131  ;
	input \u2_uk_K_r9_reg[12]/NET0131  ;
	input \u2_uk_K_r9_reg[13]/NET0131  ;
	input \u2_uk_K_r9_reg[14]/NET0131  ;
	input \u2_uk_K_r9_reg[15]/NET0131  ;
	input \u2_uk_K_r9_reg[16]/NET0131  ;
	input \u2_uk_K_r9_reg[17]/NET0131  ;
	input \u2_uk_K_r9_reg[18]/NET0131  ;
	input \u2_uk_K_r9_reg[19]/NET0131  ;
	input \u2_uk_K_r9_reg[1]/NET0131  ;
	input \u2_uk_K_r9_reg[20]/NET0131  ;
	input \u2_uk_K_r9_reg[21]/NET0131  ;
	input \u2_uk_K_r9_reg[22]/NET0131  ;
	input \u2_uk_K_r9_reg[23]/NET0131  ;
	input \u2_uk_K_r9_reg[25]/NET0131  ;
	input \u2_uk_K_r9_reg[26]/NET0131  ;
	input \u2_uk_K_r9_reg[27]/NET0131  ;
	input \u2_uk_K_r9_reg[28]/NET0131  ;
	input \u2_uk_K_r9_reg[29]/NET0131  ;
	input \u2_uk_K_r9_reg[30]/NET0131  ;
	input \u2_uk_K_r9_reg[31]/P0001  ;
	input \u2_uk_K_r9_reg[32]/NET0131  ;
	input \u2_uk_K_r9_reg[33]/NET0131  ;
	input \u2_uk_K_r9_reg[34]/NET0131  ;
	input \u2_uk_K_r9_reg[35]/NET0131  ;
	input \u2_uk_K_r9_reg[36]/NET0131  ;
	input \u2_uk_K_r9_reg[37]/NET0131  ;
	input \u2_uk_K_r9_reg[38]/NET0131  ;
	input \u2_uk_K_r9_reg[39]/NET0131  ;
	input \u2_uk_K_r9_reg[3]/NET0131  ;
	input \u2_uk_K_r9_reg[40]/NET0131  ;
	input \u2_uk_K_r9_reg[41]/NET0131  ;
	input \u2_uk_K_r9_reg[42]/NET0131  ;
	input \u2_uk_K_r9_reg[43]/NET0131  ;
	input \u2_uk_K_r9_reg[44]/NET0131  ;
	input \u2_uk_K_r9_reg[45]/NET0131  ;
	input \u2_uk_K_r9_reg[46]/NET0131  ;
	input \u2_uk_K_r9_reg[47]/NET0131  ;
	input \u2_uk_K_r9_reg[48]/NET0131  ;
	input \u2_uk_K_r9_reg[49]/NET0131  ;
	input \u2_uk_K_r9_reg[4]/NET0131  ;
	input \u2_uk_K_r9_reg[50]/NET0131  ;
	input \u2_uk_K_r9_reg[51]/NET0131  ;
	input \u2_uk_K_r9_reg[52]/NET0131  ;
	input \u2_uk_K_r9_reg[53]/NET0131  ;
	input \u2_uk_K_r9_reg[54]/NET0131  ;
	input \u2_uk_K_r9_reg[55]/NET0131  ;
	input \u2_uk_K_r9_reg[5]/NET0131  ;
	input \u2_uk_K_r9_reg[6]/NET0131  ;
	input \u2_uk_K_r9_reg[7]/NET0131  ;
	input \u2_uk_K_r9_reg[8]/NET0131  ;
	input \u2_uk_K_r9_reg[9]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g16/_0_  ;
	output \g191647/_3_  ;
	output \g191648/_3_  ;
	output \g191819/_3_  ;
	output \g191821/_0_  ;
	output \g191940/_3_  ;
	output \g191941/_0_  ;
	output \g191942/_0_  ;
	output \g191944/_0_  ;
	output \g191945/_0_  ;
	output \g191946/_0_  ;
	output \g191947/_3_  ;
	output \g191948/_0_  ;
	output \g191949/_0_  ;
	output \g191950/_0_  ;
	output \g191951/_3_  ;
	output \g191952/_0_  ;
	output \g192015/_3_  ;
	output \g192016/_3_  ;
	output \g192017/_3_  ;
	output \g192018/_3_  ;
	output \g192019/_3_  ;
	output \g192020/_0_  ;
	output \g192021/_3_  ;
	output \g192022/_0_  ;
	output \g192047/_0_  ;
	output \g192048/_0_  ;
	output \g192049/_0_  ;
	output \g192050/_0_  ;
	output \g192051/_0_  ;
	output \g192081/_0_  ;
	output \g193428/_3_  ;
	output \g193720/_0_  ;
	output \g193721/_0_  ;
	output \g193877/_0_  ;
	output \g193878/_0_  ;
	output \g193879/_0_  ;
	output \g193880/_3_  ;
	output \g193881/_0_  ;
	output \g193882/_0_  ;
	output \g193998/_0_  ;
	output \g193999/_0_  ;
	output \g194000/_3_  ;
	output \g194001/_0_  ;
	output \g194002/_0_  ;
	output \g194003/_0_  ;
	output \g194004/_0_  ;
	output \g194005/_0_  ;
	output \g194006/_0_  ;
	output \g194007/_0_  ;
	output \g194008/_0_  ;
	output \g194009/_0_  ;
	output \g194010/_0_  ;
	output \g194055/_3_  ;
	output \g194056/_3_  ;
	output \g194057/_0_  ;
	output \g194058/_0_  ;
	output \g194059/_0_  ;
	output \g194060/_0_  ;
	output \g194090/_0_  ;
	output \g194091/_0_  ;
	output \g194092/_0_  ;
	output \g194093/_0_  ;
	output \g195671/_0_  ;
	output \g195672/_3_  ;
	output \g195868/_0_  ;
	output \g195869/_0_  ;
	output \g195870/_0_  ;
	output \g196010/_0_  ;
	output \g196011/_0_  ;
	output \g196012/_0_  ;
	output \g196013/_0_  ;
	output \g196014/_0_  ;
	output \g196015/_0_  ;
	output \g196016/_0_  ;
	output \g196017/_0_  ;
	output \g196018/_0_  ;
	output \g196019/_3_  ;
	output \g196020/_0_  ;
	output \g196021/_0_  ;
	output \g196022/_0_  ;
	output \g196096/_3_  ;
	output \g196097/_0_  ;
	output \g196098/_0_  ;
	output \g196099/_0_  ;
	output \g196100/_3_  ;
	output \g196101/_0_  ;
	output \g196102/_0_  ;
	output \g196103/_0_  ;
	output \g196136/_0_  ;
	output \g196137/_0_  ;
	output \g196138/_0_  ;
	output \g196139/_0_  ;
	output \g196140/_0_  ;
	output \g196170/_0_  ;
	output \g197520/_3_  ;
	output \g197821/_0_  ;
	output \g197923/_0_  ;
	output \g197996/_0_  ;
	output \g197997/_3_  ;
	output \g197998/_0_  ;
	output \g197999/_0_  ;
	output \g198000/_0_  ;
	output \g198071/_0_  ;
	output \g198123/_0_  ;
	output \g198124/_0_  ;
	output \g198125/_0_  ;
	output \g198126/_0_  ;
	output \g198127/_0_  ;
	output \g198128/_0_  ;
	output \g198129/_0_  ;
	output \g198130/_0_  ;
	output \g198131/_0_  ;
	output \g198132/_0_  ;
	output \g198133/_0_  ;
	output \g198134/_3_  ;
	output \g198135/_0_  ;
	output \g198182/_0_  ;
	output \g198183/_3_  ;
	output \g198184/_0_  ;
	output \g198185/_0_  ;
	output \g198186/_0_  ;
	output \g198187/_0_  ;
	output \g198219/_0_  ;
	output \g198220/_0_  ;
	output \g198221/_0_  ;
	output \g198222/_0_  ;
	output \g199794/_0_  ;
	output \g199795/_3_  ;
	output \g200006/_0_  ;
	output \g200007/_0_  ;
	output \g200008/_0_  ;
	output \g200139/_0_  ;
	output \g200140/_0_  ;
	output \g200141/_0_  ;
	output \g200142/_0_  ;
	output \g200143/_0_  ;
	output \g200144/_0_  ;
	output \g200145/_0_  ;
	output \g200146/_0_  ;
	output \g200147/_0_  ;
	output \g200148/_0_  ;
	output \g200149/_0_  ;
	output \g200150/_3_  ;
	output \g200151/_0_  ;
	output \g200228/_3_  ;
	output \g200229/_0_  ;
	output \g200230/_0_  ;
	output \g200231/_0_  ;
	output \g200232/_3_  ;
	output \g200233/_0_  ;
	output \g200234/_0_  ;
	output \g200235/_0_  ;
	output \g200268/_0_  ;
	output \g200269/_0_  ;
	output \g200270/_0_  ;
	output \g200271/_0_  ;
	output \g200272/_0_  ;
	output \g200299/_0_  ;
	output \g201655/_3_  ;
	output \g201960/_0_  ;
	output \g201961/_0_  ;
	output \g202131/_0_  ;
	output \g202132/_0_  ;
	output \g202133/_3_  ;
	output \g202134/_0_  ;
	output \g202135/_0_  ;
	output \g202136/_0_  ;
	output \g202257/_0_  ;
	output \g202258/_0_  ;
	output \g202259/_3_  ;
	output \g202260/_0_  ;
	output \g202261/_0_  ;
	output \g202262/_0_  ;
	output \g202263/_0_  ;
	output \g202264/_0_  ;
	output \g202265/_0_  ;
	output \g202266/_0_  ;
	output \g202267/_0_  ;
	output \g202268/_0_  ;
	output \g202269/_0_  ;
	output \g202317/_0_  ;
	output \g202318/_3_  ;
	output \g202319/_0_  ;
	output \g202320/_0_  ;
	output \g202321/_0_  ;
	output \g202322/_0_  ;
	output \g202354/_0_  ;
	output \g202355/_0_  ;
	output \g202356/_0_  ;
	output \g202357/_0_  ;
	output \g203927/_0_  ;
	output \g203928/_3_  ;
	output \g204142/_0_  ;
	output \g204143/_0_  ;
	output \g204144/_0_  ;
	output \g204275/_0_  ;
	output \g204276/_0_  ;
	output \g204277/_0_  ;
	output \g204278/_0_  ;
	output \g204279/_0_  ;
	output \g204280/_0_  ;
	output \g204281/_0_  ;
	output \g204282/_0_  ;
	output \g204283/_0_  ;
	output \g204284/_0_  ;
	output \g204285/_0_  ;
	output \g204286/_3_  ;
	output \g204287/_0_  ;
	output \g204363/_3_  ;
	output \g204364/_0_  ;
	output \g204365/_0_  ;
	output \g204366/_0_  ;
	output \g204367/_3_  ;
	output \g204368/_0_  ;
	output \g204369/_0_  ;
	output \g204370/_0_  ;
	output \g204403/_0_  ;
	output \g204404/_0_  ;
	output \g204405/_0_  ;
	output \g204406/_0_  ;
	output \g204407/_0_  ;
	output \g204434/_0_  ;
	output \g205833/_3_  ;
	output \g206103/_0_  ;
	output \g206104/_0_  ;
	output \g206266/_0_  ;
	output \g206267/_0_  ;
	output \g206268/_0_  ;
	output \g206269/_3_  ;
	output \g206270/_0_  ;
	output \g206271/_0_  ;
	output \g206387/_0_  ;
	output \g206388/_0_  ;
	output \g206389/_3_  ;
	output \g206390/_0_  ;
	output \g206391/_0_  ;
	output \g206392/_0_  ;
	output \g206393/_0_  ;
	output \g206394/_0_  ;
	output \g206395/_0_  ;
	output \g206396/_0_  ;
	output \g206397/_0_  ;
	output \g206398/_0_  ;
	output \g206399/_0_  ;
	output \g206446/_0_  ;
	output \g206447/_3_  ;
	output \g206448/_0_  ;
	output \g206449/_0_  ;
	output \g206450/_0_  ;
	output \g206451/_0_  ;
	output \g206483/_0_  ;
	output \g206484/_0_  ;
	output \g206485/_0_  ;
	output \g206486/_0_  ;
	output \g208069/_0_  ;
	output \g208070/_3_  ;
	output \g208253/_0_  ;
	output \g208254/_0_  ;
	output \g208255/_0_  ;
	output \g208406/_0_  ;
	output \g208407/_0_  ;
	output \g208408/_0_  ;
	output \g208409/_0_  ;
	output \g208410/_0_  ;
	output \g208411/_0_  ;
	output \g208412/_0_  ;
	output \g208413/_0_  ;
	output \g208414/_0_  ;
	output \g208415/_3_  ;
	output \g208416/_0_  ;
	output \g208417/_0_  ;
	output \g208418/_0_  ;
	output \g208493/_3_  ;
	output \g208494/_0_  ;
	output \g208495/_0_  ;
	output \g208496/_0_  ;
	output \g208497/_3_  ;
	output \g208498/_0_  ;
	output \g208499/_0_  ;
	output \g208500/_0_  ;
	output \g208533/_0_  ;
	output \g208534/_0_  ;
	output \g208535/_0_  ;
	output \g208536/_0_  ;
	output \g208537/_0_  ;
	output \g208564/_0_  ;
	output \g209938/_3_  ;
	output \g210205/_0_  ;
	output \g210206/_0_  ;
	output \g210380/_0_  ;
	output \g210381/_0_  ;
	output \g210382/_0_  ;
	output \g210383/_3_  ;
	output \g210384/_0_  ;
	output \g210385/_0_  ;
	output \g210499/_0_  ;
	output \g210500/_0_  ;
	output \g210501/_3_  ;
	output \g210502/_0_  ;
	output \g210503/_0_  ;
	output \g210504/_0_  ;
	output \g210505/_0_  ;
	output \g210506/_0_  ;
	output \g210507/_0_  ;
	output \g210508/_0_  ;
	output \g210509/_0_  ;
	output \g210510/_0_  ;
	output \g210511/_0_  ;
	output \g210558/_0_  ;
	output \g210559/_3_  ;
	output \g210560/_0_  ;
	output \g210561/_0_  ;
	output \g210562/_0_  ;
	output \g210563/_0_  ;
	output \g210595/_0_  ;
	output \g210596/_0_  ;
	output \g210597/_0_  ;
	output \g210598/_0_  ;
	output \g212159/_0_  ;
	output \g212160/_3_  ;
	output \g212384/_0_  ;
	output \g212385/_0_  ;
	output \g212386/_0_  ;
	output \g212536/_0_  ;
	output \g212537/_0_  ;
	output \g212538/_0_  ;
	output \g212539/_0_  ;
	output \g212540/_0_  ;
	output \g212541/_0_  ;
	output \g212542/_0_  ;
	output \g212543/_0_  ;
	output \g212544/_0_  ;
	output \g212545/_0_  ;
	output \g212546/_3_  ;
	output \g212547/_0_  ;
	output \g212623/_3_  ;
	output \g212624/_0_  ;
	output \g212625/_0_  ;
	output \g212626/_0_  ;
	output \g212627/_0_  ;
	output \g212628/_3_  ;
	output \g212629/_0_  ;
	output \g212630/_0_  ;
	output \g212631/_0_  ;
	output \g212667/_0_  ;
	output \g212668/_0_  ;
	output \g212669/_0_  ;
	output \g212670/_0_  ;
	output \g212671/_0_  ;
	output \g212699/_0_  ;
	output \g214033/_3_  ;
	output \g214309/_3_  ;
	output \g214310/_0_  ;
	output \g214494/_0_  ;
	output \g214495/_0_  ;
	output \g214496/_0_  ;
	output \g214497/_3_  ;
	output \g214632/_0_  ;
	output \g214633/_0_  ;
	output \g214634/_3_  ;
	output \g214635/_0_  ;
	output \g214636/_0_  ;
	output \g214637/_0_  ;
	output \g214638/_0_  ;
	output \g214639/_0_  ;
	output \g214640/_0_  ;
	output \g214641/_0_  ;
	output \g214642/_0_  ;
	output \g214643/_0_  ;
	output \g214691/_0_  ;
	output \g214692/_0_  ;
	output \g214693/_3_  ;
	output \g214694/_0_  ;
	output \g214695/_0_  ;
	output \g214696/_0_  ;
	output \g214697/_0_  ;
	output \g214729/_0_  ;
	output \g214730/_0_  ;
	output \g214731/_0_  ;
	output \g214732/_0_  ;
	output \g214733/_0_  ;
	output \g216157/_0_  ;
	output \g216158/_3_  ;
	output \g216492/_0_  ;
	output \g216493/_0_  ;
	output \g216671/_0_  ;
	output \g216672/_0_  ;
	output \g216673/_0_  ;
	output \g216674/_0_  ;
	output \g216675/_0_  ;
	output \g216676/_3_  ;
	output \g216677/_0_  ;
	output \g216735/_0_  ;
	output \g216736/_3_  ;
	output \g216737/_0_  ;
	output \g216738/_0_  ;
	output \g216739/_0_  ;
	output \g216740/_0_  ;
	output \g216741/_0_  ;
	output \g216742/_0_  ;
	output \g216743/_0_  ;
	output \g216744/_0_  ;
	output \g216745/_0_  ;
	output \g216746/_3_  ;
	output \g216747/_0_  ;
	output \g216748/_0_  ;
	output \g216749/_0_  ;
	output \g216788/_0_  ;
	output \g216789/_0_  ;
	output \g216790/_0_  ;
	output \g216791/_0_  ;
	output \g216792/_0_  ;
	output \g216829/_0_  ;
	output \g218407/_3_  ;
	output \g218408/_0_  ;
	output \g218423/_3_  ;
	output \g218601/_0_  ;
	output \g218602/_0_  ;
	output \g218603/_0_  ;
	output \g218604/_0_  ;
	output \g218724/_0_  ;
	output \g218725/_0_  ;
	output \g218726/_0_  ;
	output \g218727/_0_  ;
	output \g218728/_0_  ;
	output \g218729/_0_  ;
	output \g218730/_0_  ;
	output \g218731/_0_  ;
	output \g218732/_0_  ;
	output \g218733/_0_  ;
	output \g218734/_0_  ;
	output \g218735/_3_  ;
	output \g218736/_0_  ;
	output \g218808/_3_  ;
	output \g218809/_0_  ;
	output \g218810/_0_  ;
	output \g218811/_3_  ;
	output \g218812/_0_  ;
	output \g218813/_0_  ;
	output \g218814/_0_  ;
	output \g218846/_0_  ;
	output \g218847/_0_  ;
	output \g218848/_0_  ;
	output \g218849/_0_  ;
	output \g218877/_0_  ;
	output \g22/_0_  ;
	output \g220545/_0_  ;
	output \g220546/_3_  ;
	output \g220725/_3_  ;
	output \g220726/_0_  ;
	output \g220793/_0_  ;
	output \g220794/_0_  ;
	output \g220795/_0_  ;
	output \g220796/_0_  ;
	output \g220797/_0_  ;
	output \g220798/_0_  ;
	output \g220799/_0_  ;
	output \g220800/_0_  ;
	output \g220801/_0_  ;
	output \g220802/_0_  ;
	output \g220803/_0_  ;
	output \g220804/_3_  ;
	output \g220805/_0_  ;
	output \g220806/_0_  ;
	output \g220807/_0_  ;
	output \g220872/_3_  ;
	output \g220873/_0_  ;
	output \g220874/_3_  ;
	output \g220875/_0_  ;
	output \g220876/_0_  ;
	output \g220877/_0_  ;
	output \g220921/_0_  ;
	output \g220922/_0_  ;
	output \g220923/_0_  ;
	output \g220924/_0_  ;
	output \g220925/_0_  ;
	output \g220926/_0_  ;
	output \g220969/_0_  ;
	output \g221011/_3_  ;
	output \g221039/_3_  ;
	output \g221086/_3_  ;
	output \g221131/_0_  ;
	output \g224010/_3_  ;
	output \g224368/_3_  ;
	output \g224369/_3_  ;
	output \g224532/_0_  ;
	output \g224533/_0_  ;
	output \g224534/_0_  ;
	output \g224535/_3_  ;
	output \g224536/_0_  ;
	output \g224537/_0_  ;
	output \g224640/_3_  ;
	output \g224641/_0_  ;
	output \g224642/_0_  ;
	output \g224643/_3_  ;
	output \g224644/_0_  ;
	output \g224645/_0_  ;
	output \g224646/_3_  ;
	output \g224647/_0_  ;
	output \g224648/_3_  ;
	output \g224649/_0_  ;
	output \g224650/_0_  ;
	output \g224651/_0_  ;
	output \g224652/_0_  ;
	output \g224690/_0_  ;
	output \g224691/_3_  ;
	output \g224692/_3_  ;
	output \g224693/_0_  ;
	output \g224694/_0_  ;
	output \g224695/_3_  ;
	output \g224723/_0_  ;
	output \g224724/_0_  ;
	output \g224725/_0_  ;
	output \g224726/_0_  ;
	output \g226372/_0_  ;
	output \g226373/_3_  ;
	output \g226549/_3_  ;
	output \g226550/_0_  ;
	output \g226616/_0_  ;
	output \g226635/_0_  ;
	output \g226636/_0_  ;
	output \g226637/_0_  ;
	output \g226638/_0_  ;
	output \g226639/_0_  ;
	output \g226640/_0_  ;
	output \g226641/_3_  ;
	output \g226642/_0_  ;
	output \g226643/_0_  ;
	output \g226644/_0_  ;
	output \g226645/_0_  ;
	output \g226646/_0_  ;
	output \g226692/_3_  ;
	output \g226693/_0_  ;
	output \g226694/_3_  ;
	output \g226695/_3_  ;
	output \g226696/_3_  ;
	output \g226697/_0_  ;
	output \g226698/_0_  ;
	output \g226699/_0_  ;
	output \g226728/_0_  ;
	output \g226729/_0_  ;
	output \g226730/_0_  ;
	output \g226731/_0_  ;
	output \g226732/_0_  ;
	output \g226759/_0_  ;
	output \g228250/_0_  ;
	output \g228396/_0_  ;
	output \g228397/_0_  ;
	output \g228566/_0_  ;
	output \g228567/_0_  ;
	output \g228568/_0_  ;
	output \g228609/_0_  ;
	output \g228610/_3_  ;
	output \g228688/_0_  ;
	output \g228689/_0_  ;
	output \g228690/_3_  ;
	output \g228691/_0_  ;
	output \g228692/_0_  ;
	output \g228693/_0_  ;
	output \g228694/_0_  ;
	output \g228695/_0_  ;
	output \g228696/_0_  ;
	output \g228697/_0_  ;
	output \g228698/_0_  ;
	output \g228699/_0_  ;
	output \g228700/_0_  ;
	output \g228748/_0_  ;
	output \g228749/_3_  ;
	output \g228750/_0_  ;
	output \g228751/_0_  ;
	output \g228752/_0_  ;
	output \g228753/_0_  ;
	output \g228784/_0_  ;
	output \g228785/_0_  ;
	output \g228786/_0_  ;
	output \g228787/_3_  ;
	output \g230339/_0_  ;
	output \g230340/_0_  ;
	output \g230546/_0_  ;
	output \g230580/_0_  ;
	output \g230679/_0_  ;
	output \g230680/_0_  ;
	output \g230681/_0_  ;
	output \g230682/_0_  ;
	output \g230683/_0_  ;
	output \g230684/_0_  ;
	output \g230685/_0_  ;
	output \g230686/_0_  ;
	output \g230687/_0_  ;
	output \g230688/_0_  ;
	output \g230689/_3_  ;
	output \g230690/_0_  ;
	output \g230710/_0_  ;
	output \g230766/_0_  ;
	output \g230767/_0_  ;
	output \g230768/_0_  ;
	output \g230769/_3_  ;
	output \g230770/_0_  ;
	output \g230771/_0_  ;
	output \g230772/_0_  ;
	output \g230773/_3_  ;
	output \g230810/_0_  ;
	output \g230811/_0_  ;
	output \g230812/_0_  ;
	output \g230813/_0_  ;
	output \g230814/_0_  ;
	output \g230840/_3_  ;
	output \g232196/_3_  ;
	output \g232469/_0_  ;
	output \g232470/_0_  ;
	output \g232633/_0_  ;
	output \g232635/_3_  ;
	output \g232636/_0_  ;
	output \g232637/_0_  ;
	output \g232691/_0_  ;
	output \g232747/_0_  ;
	output \g232748/_0_  ;
	output \g232749/_3_  ;
	output \g232750/_0_  ;
	output \g232751/_0_  ;
	output \g232752/_0_  ;
	output \g232753/_0_  ;
	output \g232754/_0_  ;
	output \g232755/_0_  ;
	output \g232756/_0_  ;
	output \g232757/_0_  ;
	output \g232758/_0_  ;
	output \g232759/_0_  ;
	output \g232804/_0_  ;
	output \g232805/_0_  ;
	output \g232806/_0_  ;
	output \g232807/_0_  ;
	output \g232808/_3_  ;
	output \g232809/_0_  ;
	output \g232841/_0_  ;
	output \g232842/_3_  ;
	output \g232843/_0_  ;
	output \g232844/_0_  ;
	output \g234520/_0_  ;
	output \g234687/_0_  ;
	output \g234688/_0_  ;
	output \g234689/_0_  ;
	output \g234764/_0_  ;
	output \g234765/_0_  ;
	output \g234766/_0_  ;
	output \g234767/_3_  ;
	output \g234768/_0_  ;
	output \g234769/_0_  ;
	output \g234770/_0_  ;
	output \g234771/_0_  ;
	output \g234772/_0_  ;
	output \g234773/_0_  ;
	output \g234774/_3_  ;
	output \g234775/_0_  ;
	output \g234776/_0_  ;
	output \g234824/_3_  ;
	output \g234825/_0_  ;
	output \g234826/_0_  ;
	output \g234827/_0_  ;
	output \g234828/_3_  ;
	output \g234829/_0_  ;
	output \g234830/_0_  ;
	output \g234831/_0_  ;
	output \g234867/_0_  ;
	output \g234868/_0_  ;
	output \g234869/_0_  ;
	output \g234870/_0_  ;
	output \g234896/_0_  ;
	output \g236294/_3_  ;
	output \g236541/_0_  ;
	output \g236542/_0_  ;
	output \g236724/_0_  ;
	output \g236725/_0_  ;
	output \g236726/_0_  ;
	output \g236727/_3_  ;
	output \g236728/_0_  ;
	output \g236729/_0_  ;
	output \g236821/_0_  ;
	output \g236822/_3_  ;
	output \g236823/_0_  ;
	output \g236824/_3_  ;
	output \g236825/_0_  ;
	output \g236826/_0_  ;
	output \g236827/_0_  ;
	output \g236828/_0_  ;
	output \g236829/_0_  ;
	output \g236830/_0_  ;
	output \g236831/_0_  ;
	output \g236832/_0_  ;
	output \g236877/_0_  ;
	output \g236878/_3_  ;
	output \g236879/_0_  ;
	output \g236880/_0_  ;
	output \g236881/_0_  ;
	output \g236882/_0_  ;
	output \g236914/_0_  ;
	output \g236915/_0_  ;
	output \g236916/_0_  ;
	output \g236917/_0_  ;
	output \g238530/_0_  ;
	output \g238531/_3_  ;
	output \g238723/_0_  ;
	output \g238724/_0_  ;
	output \g238725/_0_  ;
	output \g238840/_0_  ;
	output \g238841/_0_  ;
	output \g238842/_0_  ;
	output \g238843/_3_  ;
	output \g238844/_0_  ;
	output \g238845/_0_  ;
	output \g238846/_0_  ;
	output \g238847/_0_  ;
	output \g238848/_0_  ;
	output \g238849/_0_  ;
	output \g238850/_0_  ;
	output \g238851/_3_  ;
	output \g238852/_0_  ;
	output \g238924/_0_  ;
	output \g238925/_0_  ;
	output \g238926/_0_  ;
	output \g238927/_3_  ;
	output \g238928/_0_  ;
	output \g238929/_0_  ;
	output \g238930/_0_  ;
	output \g238965/_0_  ;
	output \g238966/_0_  ;
	output \g238967/_0_  ;
	output \g238968/_0_  ;
	output \g238969/_0_  ;
	output \g238996/_0_  ;
	output \g240353/_3_  ;
	output \g240640/_0_  ;
	output \g240641/_0_  ;
	output \g240813/_0_  ;
	output \g240814/_0_  ;
	output \g240815/_3_  ;
	output \g240816/_0_  ;
	output \g240817/_0_  ;
	output \g240818/_0_  ;
	output \g240925/_0_  ;
	output \g240926/_0_  ;
	output \g240927/_3_  ;
	output \g240928/_0_  ;
	output \g240929/_3_  ;
	output \g240930/_0_  ;
	output \g240931/_0_  ;
	output \g240932/_0_  ;
	output \g240933/_0_  ;
	output \g240934/_0_  ;
	output \g240935/_0_  ;
	output \g240936/_0_  ;
	output \g240937/_0_  ;
	output \g240984/_0_  ;
	output \g240985/_3_  ;
	output \g240986/_0_  ;
	output \g240987/_0_  ;
	output \g240988/_0_  ;
	output \g240989/_0_  ;
	output \g241021/_0_  ;
	output \g241022/_0_  ;
	output \g241023/_0_  ;
	output \g241024/_0_  ;
	output \g242616/_0_  ;
	output \g242617/_3_  ;
	output \g242815/_0_  ;
	output \g242816/_0_  ;
	output \g242817/_0_  ;
	output \g242955/_0_  ;
	output \g242956/_0_  ;
	output \g242957/_0_  ;
	output \g242958/_3_  ;
	output \g242959/_0_  ;
	output \g242960/_0_  ;
	output \g242961/_0_  ;
	output \g242962/_0_  ;
	output \g242963/_3_  ;
	output \g242964/_0_  ;
	output \g242965/_0_  ;
	output \g242966/_0_  ;
	output \g242967/_0_  ;
	output \g243037/_3_  ;
	output \g243038/_0_  ;
	output \g243039/_0_  ;
	output \g243040/_0_  ;
	output \g243041/_3_  ;
	output \g243042/_0_  ;
	output \g243043/_0_  ;
	output \g243044/_0_  ;
	output \g243078/_0_  ;
	output \g243079/_0_  ;
	output \g243080/_0_  ;
	output \g243081/_0_  ;
	output \g243082/_0_  ;
	output \g243109/_0_  ;
	output \g244465/_3_  ;
	output \g244753/_3_  ;
	output \g244754/_0_  ;
	output \g244924/_0_  ;
	output \g244925/_0_  ;
	output \g244926/_3_  ;
	output \g244927/_0_  ;
	output \g244928/_0_  ;
	output \g245035/_0_  ;
	output \g245036/_0_  ;
	output \g245037/_0_  ;
	output \g245038/_3_  ;
	output \g245039/_3_  ;
	output \g245040/_0_  ;
	output \g245041/_0_  ;
	output \g245043/_0_  ;
	output \g245045/_0_  ;
	output \g245046/_0_  ;
	output \g245047/_0_  ;
	output \g245092/_0_  ;
	output \g245093/_3_  ;
	output \g245094/_0_  ;
	output \g245095/_0_  ;
	output \g245096/_0_  ;
	output \g245097/_0_  ;
	output \g245129/_0_  ;
	output \g245130/_0_  ;
	output \g245131/_0_  ;
	output \g245132/_0_  ;
	output \g246715/_0_  ;
	output \g246716/_3_  ;
	output \g246911/_0_  ;
	output \g246912/_0_  ;
	output \g246913/_0_  ;
	output \g247057/_0_  ;
	output \g247058/_0_  ;
	output \g247059/_0_  ;
	output \g247060/_0_  ;
	output \g247061/_0_  ;
	output \g247062/_3_  ;
	output \g247063/_0_  ;
	output \g247064/_0_  ;
	output \g247065/_0_  ;
	output \g247066/_0_  ;
	output \g247067/_3_  ;
	output \g247068/_0_  ;
	output \g247069/_0_  ;
	output \g247137/_3_  ;
	output \g247138/_0_  ;
	output \g247139/_0_  ;
	output \g247140/_0_  ;
	output \g247141/_3_  ;
	output \g247142/_0_  ;
	output \g247143/_0_  ;
	output \g247144/_0_  ;
	output \g247179/_0_  ;
	output \g247180/_0_  ;
	output \g247181/_0_  ;
	output \g247182/_0_  ;
	output \g247183/_0_  ;
	output \g247210/_0_  ;
	output \g248581/_3_  ;
	output \g248828/_0_  ;
	output \g248829/_0_  ;
	output \g249033/_0_  ;
	output \g249035/_0_  ;
	output \g249036/_3_  ;
	output \g249037/_0_  ;
	output \g249038/_0_  ;
	output \g249147/_0_  ;
	output \g249148/_0_  ;
	output \g249149/_3_  ;
	output \g249150/_0_  ;
	output \g249152/_0_  ;
	output \g249153/_0_  ;
	output \g249155/_0_  ;
	output \g249156/_0_  ;
	output \g249157/_0_  ;
	output \g249200/_3_  ;
	output \g249201/_0_  ;
	output \g249202/_0_  ;
	output \g249203/_3_  ;
	output \g249204/_0_  ;
	output \g249205/_0_  ;
	output \g249206/_0_  ;
	output \g249207/_0_  ;
	output \g249239/_0_  ;
	output \g249240/_0_  ;
	output \g249241/_0_  ;
	output \g249242/_0_  ;
	output \g250815/_0_  ;
	output \g251006/_0_  ;
	output \g251007/_0_  ;
	output \g251008/_0_  ;
	output \g251009/_3_  ;
	output \g251160/_0_  ;
	output \g251161/_0_  ;
	output \g251162/_0_  ;
	output \g251163/_3_  ;
	output \g251164/_0_  ;
	output \g251165/_0_  ;
	output \g251166/_0_  ;
	output \g251167/_0_  ;
	output \g251168/_0_  ;
	output \g251169/_0_  ;
	output \g251170/_3_  ;
	output \g251171/_0_  ;
	output \g251245/_3_  ;
	output \g251246/_0_  ;
	output \g251247/_0_  ;
	output \g251248/_0_  ;
	output \g251249/_3_  ;
	output \g251250/_0_  ;
	output \g251251/_0_  ;
	output \g251252/_0_  ;
	output \g251286/_0_  ;
	output \g251287/_0_  ;
	output \g251288/_0_  ;
	output \g251289/_0_  ;
	output \g251290/_0_  ;
	output \g251291/_0_  ;
	output \g251318/_0_  ;
	output \g252698/_3_  ;
	output \g252942/_0_  ;
	output \g252943/_0_  ;
	output \g253118/_0_  ;
	output \g253119/_0_  ;
	output \g253120/_0_  ;
	output \g253121/_0_  ;
	output \g253122/_3_  ;
	output \g253123/_0_  ;
	output \g253236/_0_  ;
	output \g253237/_3_  ;
	output \g253238/_3_  ;
	output \g253239/_0_  ;
	output \g253240/_0_  ;
	output \g253241/_0_  ;
	output \g253242/_0_  ;
	output \g253243/_0_  ;
	output \g253244/_0_  ;
	output \g253245/_0_  ;
	output \g253246/_0_  ;
	output \g253247/_0_  ;
	output \g253248/_0_  ;
	output \g253306/_0_  ;
	output \g253307/_3_  ;
	output \g253308/_0_  ;
	output \g253309/_0_  ;
	output \g253310/_0_  ;
	output \g253311/_0_  ;
	output \g253356/_0_  ;
	output \g253357/_0_  ;
	output \g253358/_0_  ;
	output \g253359/_0_  ;
	output \g253436/_3_  ;
	output \g253437/_0_  ;
	output \g253438/_0_  ;
	output \g253469/_3_  ;
	output \g253470/_3_  ;
	output \g253471/_3_  ;
	output \g253521/_0_  ;
	output \g253522/_0_  ;
	output \g253523/_0_  ;
	output \g253524/_3_  ;
	output \g256730/_3_  ;
	output \g256731/_3_  ;
	output \g256927/_0_  ;
	output \g256928/_0_  ;
	output \g256929/_3_  ;
	output \g257049/_0_  ;
	output \g257050/_0_  ;
	output \g257051/_3_  ;
	output \g257052/_0_  ;
	output \g257053/_0_  ;
	output \g257054/_0_  ;
	output \g257055/_3_  ;
	output \g257056/_0_  ;
	output \g257057/_0_  ;
	output \g257058/_3_  ;
	output \g257059/_0_  ;
	output \g257060/_0_  ;
	output \g257082/_0_  ;
	output \g257125/_3_  ;
	output \g257126/_0_  ;
	output \g257127/_0_  ;
	output \g257128/_3_  ;
	output \g257129/_3_  ;
	output \g257130/_0_  ;
	output \g257131/_0_  ;
	output \g257132/_0_  ;
	output \g257163/_0_  ;
	output \g257164/_0_  ;
	output \g257165/_0_  ;
	output \g257166/_0_  ;
	output \g257167/_0_  ;
	output \g257194/_0_  ;
	output \g258552/_0_  ;
	output \g258850/_0_  ;
	output \g258851/_3_  ;
	output \g258993/_0_  ;
	output \g258994/_0_  ;
	output \g258995/_0_  ;
	output \g258996/_0_  ;
	output \g259026/_3_  ;
	output \g259027/_0_  ;
	output \g259105/_0_  ;
	output \g259106/_0_  ;
	output \g259107/_3_  ;
	output \g259108/_0_  ;
	output \g259109/_3_  ;
	output \g259110/_0_  ;
	output \g259111/_0_  ;
	output \g259112/_0_  ;
	output \g259113/_0_  ;
	output \g259114/_0_  ;
	output \g259115/_0_  ;
	output \g259116/_0_  ;
	output \g259117/_0_  ;
	output \g259163/_3_  ;
	output \g259164/_3_  ;
	output \g259165/_0_  ;
	output \g259166/_0_  ;
	output \g259167/_0_  ;
	output \g259168/_0_  ;
	output \g259197/_0_  ;
	output \g259198/_0_  ;
	output \g259199/_0_  ;
	output \g259200/_0_  ;
	output \g260774/_0_  ;
	output \g260792/_3_  ;
	output \g260991/_0_  ;
	output \g261013/_0_  ;
	output \g261070/_0_  ;
	output \g261125/_0_  ;
	output \g261126/_0_  ;
	output \g261128/_0_  ;
	output \g261129/_0_  ;
	output \g261130/_0_  ;
	output \g261131/_0_  ;
	output \g261132/_0_  ;
	output \g261133/_0_  ;
	output \g261134/_3_  ;
	output \g261135/_0_  ;
	output \g261136/_0_  ;
	output \g261158/_3_  ;
	output \g261206/_0_  ;
	output \g261207/_0_  ;
	output \g261208/_0_  ;
	output \g261209/_0_  ;
	output \g261210/_3_  ;
	output \g261211/_0_  ;
	output \g261212/_3_  ;
	output \g261213/_0_  ;
	output \g261248/_0_  ;
	output \g261249/_0_  ;
	output \g261250/_0_  ;
	output \g261251/_0_  ;
	output \g261252/_0_  ;
	output \g261279/_0_  ;
	output \g262658/_3_  ;
	output \g262949/_0_  ;
	output \g263008/_3_  ;
	output \g263092/_0_  ;
	output \g263093/_0_  ;
	output \g263099/_0_  ;
	output \g263100/_0_  ;
	output \g263101/_0_  ;
	output \g263159/_3_  ;
	output \g263204/_3_  ;
	output \g263205/_0_  ;
	output \g263206/_0_  ;
	output \g263208/_0_  ;
	output \g263209/_0_  ;
	output \g263210/_0_  ;
	output \g263211/_0_  ;
	output \g263212/_0_  ;
	output \g263213/_0_  ;
	output \g263214/_0_  ;
	output \g263215/_3_  ;
	output \g263216/_0_  ;
	output \g263260/_0_  ;
	output \g263261/_0_  ;
	output \g263262/_3_  ;
	output \g263263/_0_  ;
	output \g263264/_0_  ;
	output \g263265/_0_  ;
	output \g263297/_0_  ;
	output \g263298/_0_  ;
	output \g263299/_0_  ;
	output \g263300/_0_  ;
	output \g264930/_0_  ;
	output \g264946/_3_  ;
	output \g265143/_0_  ;
	output \g265144/_0_  ;
	output \g265152/_0_  ;
	output \g265222/_0_  ;
	output \g265223/_0_  ;
	output \g265224/_0_  ;
	output \g265225/_0_  ;
	output \g265226/_0_  ;
	output \g265227/_3_  ;
	output \g265228/_0_  ;
	output \g265229/_0_  ;
	output \g265230/_0_  ;
	output \g265231/_0_  ;
	output \g265232/_0_  ;
	output \g265233/_3_  ;
	output \g265234/_0_  ;
	output \g265306/_0_  ;
	output \g265307/_0_  ;
	output \g265308/_3_  ;
	output \g265309/_3_  ;
	output \g265310/_0_  ;
	output \g265311/_0_  ;
	output \g265312/_0_  ;
	output \g265313/_0_  ;
	output \g265348/_0_  ;
	output \g265349/_0_  ;
	output \g265350/_0_  ;
	output \g265351/_0_  ;
	output \g265379/_0_  ;
	output \g266965/_3_  ;
	output \g267049/_3_  ;
	output \g267050/_0_  ;
	output \g267215/_0_  ;
	output \g267216/_0_  ;
	output \g267263/_0_  ;
	output \g267264/_3_  ;
	output \g267265/_0_  ;
	output \g267266/_0_  ;
	output \g267314/_3_  ;
	output \g267315/_0_  ;
	output \g267316/_0_  ;
	output \g267317/_0_  ;
	output \g267318/_0_  ;
	output \g267319/_0_  ;
	output \g267320/_3_  ;
	output \g267321/_0_  ;
	output \g267322/_0_  ;
	output \g267324/_0_  ;
	output \g267325/_0_  ;
	output \g267326/_0_  ;
	output \g267372/_0_  ;
	output \g267373/_3_  ;
	output \g267374/_0_  ;
	output \g267375/_0_  ;
	output \g267376/_0_  ;
	output \g267377/_0_  ;
	output \g267409/_0_  ;
	output \g267410/_0_  ;
	output \g267411/_0_  ;
	output \g267412/_0_  ;
	output \g269004/_0_  ;
	output \g269099/_3_  ;
	output \g269202/_0_  ;
	output \g269226/_0_  ;
	output \g269333/_3_  ;
	output \g269334/_0_  ;
	output \g269335/_0_  ;
	output \g269355/_0_  ;
	output \g269356/_0_  ;
	output \g269357/_3_  ;
	output \g269358/_0_  ;
	output \g269359/_0_  ;
	output \g269360/_0_  ;
	output \g269361/_0_  ;
	output \g269362/_0_  ;
	output \g269363/_0_  ;
	output \g269364/_0_  ;
	output \g269414/_0_  ;
	output \g269415/_0_  ;
	output \g269416/_0_  ;
	output \g269417/_0_  ;
	output \g269418/_3_  ;
	output \g269419/_0_  ;
	output \g269420/_3_  ;
	output \g269421/_0_  ;
	output \g269456/_0_  ;
	output \g269457/_0_  ;
	output \g269458/_0_  ;
	output \g269459/_0_  ;
	output \g269460/_0_  ;
	output \g269487/_0_  ;
	output \g271006/_3_  ;
	output \g271186/_3_  ;
	output \g271187/_0_  ;
	output \g271299/_0_  ;
	output \g271300/_0_  ;
	output \g271301/_3_  ;
	output \g271302/_0_  ;
	output \g271303/_0_  ;
	output \g271352/_0_  ;
	output \g271410/_0_  ;
	output \g271411/_0_  ;
	output \g271412/_0_  ;
	output \g271413/_0_  ;
	output \g271414/_0_  ;
	output \g271415/_0_  ;
	output \g271416/_0_  ;
	output \g271417/_3_  ;
	output \g271418/_3_  ;
	output \g271419/_0_  ;
	output \g271420/_0_  ;
	output \g271421/_0_  ;
	output \g271422/_0_  ;
	output \g271468/_3_  ;
	output \g271469/_0_  ;
	output \g271470/_0_  ;
	output \g271471/_0_  ;
	output \g271472/_0_  ;
	output \g271473/_0_  ;
	output \g271505/_0_  ;
	output \g271506/_0_  ;
	output \g271507/_0_  ;
	output \g271508/_0_  ;
	output \g273135/_0_  ;
	output \g273136/_3_  ;
	output \g273362/_0_  ;
	output \g273373/_0_  ;
	output \g273374/_0_  ;
	output \g273431/_0_  ;
	output \g273432/_0_  ;
	output \g273433/_3_  ;
	output \g273434/_0_  ;
	output \g273435/_0_  ;
	output \g273436/_0_  ;
	output \g273437/_3_  ;
	output \g273438/_0_  ;
	output \g273439/_0_  ;
	output \g273441/_0_  ;
	output \g273442/_0_  ;
	output \g273443/_0_  ;
	output \g273515/_3_  ;
	output \g273516/_0_  ;
	output \g273517/_0_  ;
	output \g273518/_3_  ;
	output \g273519/_0_  ;
	output \g273520/_0_  ;
	output \g273521/_0_  ;
	output \g273522/_0_  ;
	output \g273557/_0_  ;
	output \g273558/_0_  ;
	output \g273559/_0_  ;
	output \g273560/_0_  ;
	output \g273561/_0_  ;
	output \g273588/_0_  ;
	output \g274960/_3_  ;
	output \g275266/_3_  ;
	output \g275327/_0_  ;
	output \g275396/_0_  ;
	output \g275397/_3_  ;
	output \g275398/_0_  ;
	output \g275455/_0_  ;
	output \g275456/_0_  ;
	output \g275463/_0_  ;
	output \g275510/_3_  ;
	output \g275511/_0_  ;
	output \g275512/_0_  ;
	output \g275513/_0_  ;
	output \g275514/_3_  ;
	output \g275515/_0_  ;
	output \g275516/_0_  ;
	output \g275517/_0_  ;
	output \g275518/_0_  ;
	output \g275519/_0_  ;
	output \g275520/_0_  ;
	output \g275521/_0_  ;
	output \g275522/_0_  ;
	output \g275568/_0_  ;
	output \g275569/_0_  ;
	output \g275570/_0_  ;
	output \g275571/_0_  ;
	output \g275572/_3_  ;
	output \g275573/_0_  ;
	output \g275605/_0_  ;
	output \g275606/_0_  ;
	output \g275607/_0_  ;
	output \g275608/_0_  ;
	output \g277189/_0_  ;
	output \g277294/_3_  ;
	output \g277367/_0_  ;
	output \g277456/_0_  ;
	output \g277457/_0_  ;
	output \g277512/_0_  ;
	output \g277513/_0_  ;
	output \g277514/_3_  ;
	output \g277515/_0_  ;
	output \g277516/_0_  ;
	output \g277517/_3_  ;
	output \g277518/_0_  ;
	output \g277519/_0_  ;
	output \g277520/_0_  ;
	output \g277521/_0_  ;
	output \g277594/_0_  ;
	output \g277595/_0_  ;
	output \g277596/_3_  ;
	output \g277597/_0_  ;
	output \g277598/_0_  ;
	output \g277599/_0_  ;
	output \g277600/_0_  ;
	output \g277601/_3_  ;
	output \g277635/_0_  ;
	output \g277636/_0_  ;
	output \g277637/_0_  ;
	output \g277638/_0_  ;
	output \g277639/_0_  ;
	output \g277666/_0_  ;
	output \g279090/_3_  ;
	output \g279330/_0_  ;
	output \g279331/_0_  ;
	output \g279493/_3_  ;
	output \g279494/_0_  ;
	output \g279495/_0_  ;
	output \g279502/_0_  ;
	output \g279503/_0_  ;
	output \g279504/_0_  ;
	output \g279590/_0_  ;
	output \g279591/_0_  ;
	output \g279592/_0_  ;
	output \g279593/_0_  ;
	output \g279594/_3_  ;
	output \g279595/_3_  ;
	output \g279596/_0_  ;
	output \g279597/_0_  ;
	output \g279598/_0_  ;
	output \g279599/_0_  ;
	output \g279600/_0_  ;
	output \g279601/_0_  ;
	output \g279602/_0_  ;
	output \g279649/_0_  ;
	output \g279650/_0_  ;
	output \g279651/_0_  ;
	output \g279652/_0_  ;
	output \g279653/_0_  ;
	output \g279654/_3_  ;
	output \g279686/_0_  ;
	output \g279687/_0_  ;
	output \g279688/_0_  ;
	output \g279689/_0_  ;
	output \g281329/_0_  ;
	output \g281394/_0_  ;
	output \g281483/_0_  ;
	output \g281498/_0_  ;
	output \g281532/_0_  ;
	output \g281616/_0_  ;
	output \g281617/_0_  ;
	output \g281618/_0_  ;
	output \g281619/_0_  ;
	output \g281620/_0_  ;
	output \g281621/_0_  ;
	output \g281622/_0_  ;
	output \g281623/_3_  ;
	output \g281624/_0_  ;
	output \g281642/_0_  ;
	output \g281643/_0_  ;
	output \g281644/_3_  ;
	output \g281645/_0_  ;
	output \g281696/_0_  ;
	output \g281697/_3_  ;
	output \g281698/_0_  ;
	output \g281699/_0_  ;
	output \g281700/_0_  ;
	output \g281701/_0_  ;
	output \g281702/_3_  ;
	output \g281703/_0_  ;
	output \g281799/_0_  ;
	output \g281800/_0_  ;
	output \g281801/_0_  ;
	output \g281802/_0_  ;
	output \g281803/_0_  ;
	output \g281965/_0_  ;
	output \g287377/_0_  ;
	output \g287867/_0_  ;
	output \g287899/_0_  ;
	output \g288304/_0_  ;
	output \g288334/_0_  ;
	output \g288350/_0_  ;
	output \g288351/_0_  ;
	output \g288352/_3_  ;
	output \g288353/_0_  ;
	output \g288668/_0_  ;
	output \g288669/_0_  ;
	output \g288670/_0_  ;
	output \g288671/_0_  ;
	output \g288673/_0_  ;
	output \g288674/_3_  ;
	output \g288675/_0_  ;
	output \g288676/_0_  ;
	output \g288677/_0_  ;
	output \g288678/_0_  ;
	output \g288679/_0_  ;
	output \g288680/_3_  ;
	output \g288889/_0_  ;
	output \g288890/_0_  ;
	output \g288891/_0_  ;
	output \g288892/_0_  ;
	output \g288893/_3_  ;
	output \g288894/_0_  ;
	output \g288895/_0_  ;
	output \g288984/_0_  ;
	output \g288985/_0_  ;
	output \g288986/_0_  ;
	output \g294974/_0_  ;
	output \g295054/_0_  ;
	output \g295601/_0_  ;
	output \g295607/_0_  ;
	output \g296036/_0_  ;
	output \g296037/_0_  ;
	output \g296038/_0_  ;
	output \g296039/_0_  ;
	output \g296040/_0_  ;
	output \g296041/_0_  ;
	output \g296042/_0_  ;
	output \g296043/_3_  ;
	output \g296044/_0_  ;
	output \g296045/_0_  ;
	output \g296046/_0_  ;
	output \g296047/_0_  ;
	output \g296048/_0_  ;
	output \g296049/_3_  ;
	output \g296522/_3_  ;
	output \g296523/_3_  ;
	output \g296524/_0_  ;
	output \g296525/_0_  ;
	output \g296526/_0_  ;
	output \g296527/_0_  ;
	output \g296528/_3_  ;
	output \g296529/_0_  ;
	output \g296530/_0_  ;
	output \g296531/_0_  ;
	output \g297026/_0_  ;
	output \g297027/_0_  ;
	output \g305620/_3_  ;
	output \g305621/_3_  ;
	output \g305622/_3_  ;
	output \g305623/_3_  ;
	output \g305624/_3_  ;
	output \g305625/_3_  ;
	output \g305626/_3_  ;
	output \g305627/_3_  ;
	output \g305628/_3_  ;
	output \g305629/_3_  ;
	output \g305630/_3_  ;
	output \g305631/_3_  ;
	output \g305632/_3_  ;
	output \g305633/_3_  ;
	output \g305634/_3_  ;
	output \g305635/_3_  ;
	output \g305636/_3_  ;
	output \g305637/_3_  ;
	output \g305638/_3_  ;
	output \g305639/_3_  ;
	output \g305640/_3_  ;
	output \g305641/_3_  ;
	output \g305642/_3_  ;
	output \g305643/_3_  ;
	output \g305644/_3_  ;
	output \g305645/_3_  ;
	output \g305646/_3_  ;
	output \g305647/_3_  ;
	output \g305648/_3_  ;
	output \g305649/_3_  ;
	output \g305650/_3_  ;
	output \g305651/_3_  ;
	output \g305652/_3_  ;
	output \g305653/_3_  ;
	output \g305654/_3_  ;
	output \g305655/_3_  ;
	output \g305656/_3_  ;
	output \g305657/_3_  ;
	output \g305658/_3_  ;
	output \g305659/_3_  ;
	output \g305660/_3_  ;
	output \g305661/_3_  ;
	output \g305662/_3_  ;
	output \g305663/_3_  ;
	output \g305664/_3_  ;
	output \g305665/_3_  ;
	output \g305666/_3_  ;
	output \g305667/_3_  ;
	output \g305668/_3_  ;
	output \g305669/_3_  ;
	output \g305670/_3_  ;
	output \g305671/_3_  ;
	output \g305672/_3_  ;
	output \g305673/_3_  ;
	output \g305674/_3_  ;
	output \g305675/_3_  ;
	output \g305676/_3_  ;
	output \g305677/_3_  ;
	output \g305678/_3_  ;
	output \g305679/_3_  ;
	output \g305680/_3_  ;
	output \g305681/_3_  ;
	output \g305682/_3_  ;
	output \g305683/_3_  ;
	output \g305684/_3_  ;
	output \g305685/_3_  ;
	output \g305686/_3_  ;
	output \g305687/_3_  ;
	output \g305688/_3_  ;
	output \g305689/_3_  ;
	output \g305690/_3_  ;
	output \g305691/_3_  ;
	output \g305692/_3_  ;
	output \g305693/_3_  ;
	output \g305694/_3_  ;
	output \g305695/_3_  ;
	output \g305696/_3_  ;
	output \g305697/_3_  ;
	output \g305698/_3_  ;
	output \g305699/_3_  ;
	output \g305700/_3_  ;
	output \g305701/_3_  ;
	output \g305702/_3_  ;
	output \g305703/_3_  ;
	output \g305704/_3_  ;
	output \g305705/_3_  ;
	output \g305706/_3_  ;
	output \g305707/_3_  ;
	output \g305708/_3_  ;
	output \g305709/_3_  ;
	output \g305710/_3_  ;
	output \g305711/_3_  ;
	output \g305712/_3_  ;
	output \g305713/_3_  ;
	output \g305714/_3_  ;
	output \g305715/_3_  ;
	output \g305716/_3_  ;
	output \g305717/_3_  ;
	output \g305718/_3_  ;
	output \g305719/_3_  ;
	output \g305720/_3_  ;
	output \g305721/_3_  ;
	output \g305722/_3_  ;
	output \g305723/_3_  ;
	output \g305724/_3_  ;
	output \g305725/_3_  ;
	output \g305726/_3_  ;
	output \g305727/_3_  ;
	output \g305728/_3_  ;
	output \g305729/_3_  ;
	output \g305730/_3_  ;
	output \g305731/_3_  ;
	output \g321371/_0_  ;
	output \g321424/_0_  ;
	output \g321474/_3_  ;
	output \g321637/_3_  ;
	output \g321688/_0_  ;
	output \g321712/_0_  ;
	output \g321772/_3_  ;
	output \g321832/_0_  ;
	output \g321999/_0_  ;
	output \g322013/_3_  ;
	output \g322109/_0_  ;
	output \g322184/_0_  ;
	output \g322250/_0_  ;
	output \g322274/_0_  ;
	output \g322293/_3_  ;
	output \g322437/_0_  ;
	output \g322537/_3_  ;
	output \g322584/_0_  ;
	output \g322830/_0_  ;
	output \g322871/_0_  ;
	output \g322882/_0_  ;
	output \g322933/_0_  ;
	output \g323004/_0_  ;
	output \g323104/_0_  ;
	output \g323125/_0_  ;
	output \g323138/_3_  ;
	output \g323273/_0_  ;
	output \u0_desOut_reg[0]/_05_  ;
	output \u0_desOut_reg[12]/_05_  ;
	output \u0_desOut_reg[14]/_05_  ;
	output \u0_desOut_reg[18]/_05_  ;
	output \u0_desOut_reg[20]/_05_  ;
	output \u0_desOut_reg[24]/_05_  ;
	output \u0_desOut_reg[26]/_05_  ;
	output \u0_desOut_reg[28]/_05_  ;
	output \u0_desOut_reg[2]/_05_  ;
	output \u0_desOut_reg[30]/_05_  ;
	output \u0_desOut_reg[32]/_05_  ;
	output \u0_desOut_reg[34]/_05_  ;
	output \u0_desOut_reg[36]/_05_  ;
	output \u0_desOut_reg[42]/_05_  ;
	output \u0_desOut_reg[44]/_05_  ;
	output \u0_desOut_reg[46]/_05_  ;
	output \u0_desOut_reg[48]/_05_  ;
	output \u0_desOut_reg[54]/_05_  ;
	output \u0_desOut_reg[56]/_05_  ;
	output \u0_desOut_reg[62]/_05_  ;
	output \u0_desOut_reg[6]/_05_  ;
	output \u0_desOut_reg[8]/_05_  ;
	output \u1_desOut_reg[0]/_05_  ;
	output \u1_desOut_reg[12]/_05_  ;
	output \u1_desOut_reg[14]/_05_  ;
	output \u1_desOut_reg[16]/_05_  ;
	output \u1_desOut_reg[18]/_05_  ;
	output \u1_desOut_reg[20]/_05_  ;
	output \u1_desOut_reg[22]/_05_  ;
	output \u1_desOut_reg[24]/_05_  ;
	output \u1_desOut_reg[26]/_05_  ;
	output \u1_desOut_reg[28]/_05_  ;
	output \u1_desOut_reg[2]/_05_  ;
	output \u1_desOut_reg[30]/_05_  ;
	output \u1_desOut_reg[32]/_05_  ;
	output \u1_desOut_reg[34]/_05_  ;
	output \u1_desOut_reg[36]/_05_  ;
	output \u1_desOut_reg[38]/_05_  ;
	output \u1_desOut_reg[42]/_05_  ;
	output \u1_desOut_reg[44]/_05_  ;
	output \u1_desOut_reg[46]/_05_  ;
	output \u1_desOut_reg[48]/_05_  ;
	output \u1_desOut_reg[4]/_05_  ;
	output \u1_desOut_reg[54]/_05_  ;
	output \u1_desOut_reg[56]/_05_  ;
	output \u1_desOut_reg[58]/_05_  ;
	output \u1_desOut_reg[60]/_05_  ;
	output \u1_desOut_reg[62]/_05_  ;
	output \u1_desOut_reg[6]/_05_  ;
	output \u1_desOut_reg[8]/_05_  ;
	output \u2_desOut_reg[0]/_05_  ;
	output \u2_desOut_reg[10]/_05_  ;
	output \u2_desOut_reg[12]/_05_  ;
	output \u2_desOut_reg[14]/_05_  ;
	output \u2_desOut_reg[16]/_05_  ;
	output \u2_desOut_reg[18]/_05_  ;
	output \u2_desOut_reg[20]/_05_  ;
	output \u2_desOut_reg[22]/_05_  ;
	output \u2_desOut_reg[24]/_05_  ;
	output \u2_desOut_reg[26]/_05_  ;
	output \u2_desOut_reg[28]/_05_  ;
	output \u2_desOut_reg[2]/_05_  ;
	output \u2_desOut_reg[30]/_05_  ;
	output \u2_desOut_reg[32]/_05_  ;
	output \u2_desOut_reg[34]/_05_  ;
	output \u2_desOut_reg[36]/_05_  ;
	output \u2_desOut_reg[38]/_05_  ;
	output \u2_desOut_reg[40]/_05_  ;
	output \u2_desOut_reg[42]/_05_  ;
	output \u2_desOut_reg[44]/_05_  ;
	output \u2_desOut_reg[46]/_05_  ;
	output \u2_desOut_reg[48]/_05_  ;
	output \u2_desOut_reg[4]/_05_  ;
	output \u2_desOut_reg[50]/_05_  ;
	output \u2_desOut_reg[52]/_05_  ;
	output \u2_desOut_reg[54]/_05_  ;
	output \u2_desOut_reg[56]/_05_  ;
	output \u2_desOut_reg[58]/_05_  ;
	output \u2_desOut_reg[60]/_05_  ;
	output \u2_desOut_reg[62]/_05_  ;
	output \u2_desOut_reg[6]/_05_  ;
	output \u2_desOut_reg[8]/_05_  ;
	wire _w36346_ ;
	wire _w36345_ ;
	wire _w36344_ ;
	wire _w36343_ ;
	wire _w36342_ ;
	wire _w36341_ ;
	wire _w36340_ ;
	wire _w36339_ ;
	wire _w36338_ ;
	wire _w36337_ ;
	wire _w36336_ ;
	wire _w36335_ ;
	wire _w36334_ ;
	wire _w36333_ ;
	wire _w36332_ ;
	wire _w36331_ ;
	wire _w36330_ ;
	wire _w36329_ ;
	wire _w36328_ ;
	wire _w36327_ ;
	wire _w36326_ ;
	wire _w36325_ ;
	wire _w36324_ ;
	wire _w36323_ ;
	wire _w36322_ ;
	wire _w36321_ ;
	wire _w36320_ ;
	wire _w36319_ ;
	wire _w36318_ ;
	wire _w36317_ ;
	wire _w36316_ ;
	wire _w36315_ ;
	wire _w36314_ ;
	wire _w36313_ ;
	wire _w36312_ ;
	wire _w36311_ ;
	wire _w36310_ ;
	wire _w36309_ ;
	wire _w36308_ ;
	wire _w36307_ ;
	wire _w36306_ ;
	wire _w36305_ ;
	wire _w36304_ ;
	wire _w36303_ ;
	wire _w36302_ ;
	wire _w36301_ ;
	wire _w36300_ ;
	wire _w36299_ ;
	wire _w36298_ ;
	wire _w36297_ ;
	wire _w36296_ ;
	wire _w36295_ ;
	wire _w36294_ ;
	wire _w36293_ ;
	wire _w36292_ ;
	wire _w36291_ ;
	wire _w36290_ ;
	wire _w36289_ ;
	wire _w36288_ ;
	wire _w36287_ ;
	wire _w36286_ ;
	wire _w36285_ ;
	wire _w36284_ ;
	wire _w36283_ ;
	wire _w36282_ ;
	wire _w36281_ ;
	wire _w36280_ ;
	wire _w36279_ ;
	wire _w36278_ ;
	wire _w36277_ ;
	wire _w36276_ ;
	wire _w36275_ ;
	wire _w36274_ ;
	wire _w36273_ ;
	wire _w36272_ ;
	wire _w36271_ ;
	wire _w36270_ ;
	wire _w36269_ ;
	wire _w36268_ ;
	wire _w36267_ ;
	wire _w36266_ ;
	wire _w36265_ ;
	wire _w36264_ ;
	wire _w36263_ ;
	wire _w36262_ ;
	wire _w36261_ ;
	wire _w36260_ ;
	wire _w36259_ ;
	wire _w36258_ ;
	wire _w36257_ ;
	wire _w36256_ ;
	wire _w36255_ ;
	wire _w36254_ ;
	wire _w36253_ ;
	wire _w36252_ ;
	wire _w36251_ ;
	wire _w36250_ ;
	wire _w36249_ ;
	wire _w36248_ ;
	wire _w36247_ ;
	wire _w36246_ ;
	wire _w36245_ ;
	wire _w36244_ ;
	wire _w36243_ ;
	wire _w36242_ ;
	wire _w36241_ ;
	wire _w36240_ ;
	wire _w36239_ ;
	wire _w36238_ ;
	wire _w36237_ ;
	wire _w36236_ ;
	wire _w36235_ ;
	wire _w36234_ ;
	wire _w36233_ ;
	wire _w36232_ ;
	wire _w36231_ ;
	wire _w36230_ ;
	wire _w36229_ ;
	wire _w36228_ ;
	wire _w36227_ ;
	wire _w36226_ ;
	wire _w36225_ ;
	wire _w36224_ ;
	wire _w36223_ ;
	wire _w36222_ ;
	wire _w36221_ ;
	wire _w36220_ ;
	wire _w36219_ ;
	wire _w36218_ ;
	wire _w36217_ ;
	wire _w36216_ ;
	wire _w36215_ ;
	wire _w36214_ ;
	wire _w36213_ ;
	wire _w36212_ ;
	wire _w36211_ ;
	wire _w36210_ ;
	wire _w36209_ ;
	wire _w36208_ ;
	wire _w36207_ ;
	wire _w36206_ ;
	wire _w36205_ ;
	wire _w36204_ ;
	wire _w36203_ ;
	wire _w36202_ ;
	wire _w36201_ ;
	wire _w36200_ ;
	wire _w36199_ ;
	wire _w36198_ ;
	wire _w36197_ ;
	wire _w36196_ ;
	wire _w36195_ ;
	wire _w36194_ ;
	wire _w36193_ ;
	wire _w36192_ ;
	wire _w36191_ ;
	wire _w36190_ ;
	wire _w36189_ ;
	wire _w36188_ ;
	wire _w36187_ ;
	wire _w36186_ ;
	wire _w36185_ ;
	wire _w36184_ ;
	wire _w36183_ ;
	wire _w36182_ ;
	wire _w36181_ ;
	wire _w36180_ ;
	wire _w36179_ ;
	wire _w36178_ ;
	wire _w36177_ ;
	wire _w36176_ ;
	wire _w36175_ ;
	wire _w36174_ ;
	wire _w36173_ ;
	wire _w36172_ ;
	wire _w36171_ ;
	wire _w36170_ ;
	wire _w36169_ ;
	wire _w36168_ ;
	wire _w36167_ ;
	wire _w36166_ ;
	wire _w36165_ ;
	wire _w36164_ ;
	wire _w36163_ ;
	wire _w36162_ ;
	wire _w36161_ ;
	wire _w36160_ ;
	wire _w36159_ ;
	wire _w36158_ ;
	wire _w36157_ ;
	wire _w36156_ ;
	wire _w36155_ ;
	wire _w36154_ ;
	wire _w36153_ ;
	wire _w36152_ ;
	wire _w36151_ ;
	wire _w36150_ ;
	wire _w36149_ ;
	wire _w36148_ ;
	wire _w36147_ ;
	wire _w36146_ ;
	wire _w36145_ ;
	wire _w36144_ ;
	wire _w36143_ ;
	wire _w36142_ ;
	wire _w36141_ ;
	wire _w36140_ ;
	wire _w36139_ ;
	wire _w36138_ ;
	wire _w36137_ ;
	wire _w36136_ ;
	wire _w36135_ ;
	wire _w36134_ ;
	wire _w36133_ ;
	wire _w36132_ ;
	wire _w36131_ ;
	wire _w36130_ ;
	wire _w36129_ ;
	wire _w36128_ ;
	wire _w36127_ ;
	wire _w36126_ ;
	wire _w36125_ ;
	wire _w36124_ ;
	wire _w36123_ ;
	wire _w36122_ ;
	wire _w36121_ ;
	wire _w36120_ ;
	wire _w36119_ ;
	wire _w36118_ ;
	wire _w36117_ ;
	wire _w36116_ ;
	wire _w36115_ ;
	wire _w36114_ ;
	wire _w36113_ ;
	wire _w36112_ ;
	wire _w36111_ ;
	wire _w36110_ ;
	wire _w36109_ ;
	wire _w36108_ ;
	wire _w36107_ ;
	wire _w36106_ ;
	wire _w36105_ ;
	wire _w36104_ ;
	wire _w36103_ ;
	wire _w36102_ ;
	wire _w36101_ ;
	wire _w36100_ ;
	wire _w36099_ ;
	wire _w36098_ ;
	wire _w36097_ ;
	wire _w36096_ ;
	wire _w36095_ ;
	wire _w36094_ ;
	wire _w36093_ ;
	wire _w36092_ ;
	wire _w36091_ ;
	wire _w36090_ ;
	wire _w36089_ ;
	wire _w36088_ ;
	wire _w36087_ ;
	wire _w36086_ ;
	wire _w36085_ ;
	wire _w36084_ ;
	wire _w36083_ ;
	wire _w36082_ ;
	wire _w36081_ ;
	wire _w36080_ ;
	wire _w36079_ ;
	wire _w36078_ ;
	wire _w36077_ ;
	wire _w36076_ ;
	wire _w36075_ ;
	wire _w36074_ ;
	wire _w36073_ ;
	wire _w36072_ ;
	wire _w36071_ ;
	wire _w36070_ ;
	wire _w36069_ ;
	wire _w36068_ ;
	wire _w36067_ ;
	wire _w36066_ ;
	wire _w36065_ ;
	wire _w36064_ ;
	wire _w36063_ ;
	wire _w36062_ ;
	wire _w36061_ ;
	wire _w36060_ ;
	wire _w36059_ ;
	wire _w36058_ ;
	wire _w36057_ ;
	wire _w36056_ ;
	wire _w36055_ ;
	wire _w36054_ ;
	wire _w36053_ ;
	wire _w36052_ ;
	wire _w36051_ ;
	wire _w36050_ ;
	wire _w36049_ ;
	wire _w36048_ ;
	wire _w36047_ ;
	wire _w36046_ ;
	wire _w36045_ ;
	wire _w36044_ ;
	wire _w36043_ ;
	wire _w36042_ ;
	wire _w36041_ ;
	wire _w36040_ ;
	wire _w36039_ ;
	wire _w36038_ ;
	wire _w36037_ ;
	wire _w36036_ ;
	wire _w36035_ ;
	wire _w36034_ ;
	wire _w36033_ ;
	wire _w36032_ ;
	wire _w36031_ ;
	wire _w36030_ ;
	wire _w36029_ ;
	wire _w36028_ ;
	wire _w36027_ ;
	wire _w36026_ ;
	wire _w36025_ ;
	wire _w36024_ ;
	wire _w36023_ ;
	wire _w36022_ ;
	wire _w36021_ ;
	wire _w36020_ ;
	wire _w36019_ ;
	wire _w36018_ ;
	wire _w36017_ ;
	wire _w36016_ ;
	wire _w36015_ ;
	wire _w36014_ ;
	wire _w36013_ ;
	wire _w36012_ ;
	wire _w36011_ ;
	wire _w36010_ ;
	wire _w36009_ ;
	wire _w36008_ ;
	wire _w36007_ ;
	wire _w36006_ ;
	wire _w36005_ ;
	wire _w36004_ ;
	wire _w36003_ ;
	wire _w36002_ ;
	wire _w36001_ ;
	wire _w36000_ ;
	wire _w35999_ ;
	wire _w35998_ ;
	wire _w35997_ ;
	wire _w35996_ ;
	wire _w35995_ ;
	wire _w35994_ ;
	wire _w35993_ ;
	wire _w35992_ ;
	wire _w35991_ ;
	wire _w35990_ ;
	wire _w35989_ ;
	wire _w35988_ ;
	wire _w35987_ ;
	wire _w35986_ ;
	wire _w35985_ ;
	wire _w35984_ ;
	wire _w35983_ ;
	wire _w35982_ ;
	wire _w35981_ ;
	wire _w35980_ ;
	wire _w35979_ ;
	wire _w35978_ ;
	wire _w35977_ ;
	wire _w35976_ ;
	wire _w35975_ ;
	wire _w35974_ ;
	wire _w35973_ ;
	wire _w35972_ ;
	wire _w35971_ ;
	wire _w35970_ ;
	wire _w35969_ ;
	wire _w35968_ ;
	wire _w35967_ ;
	wire _w35966_ ;
	wire _w35965_ ;
	wire _w35964_ ;
	wire _w35963_ ;
	wire _w35962_ ;
	wire _w35961_ ;
	wire _w35960_ ;
	wire _w35959_ ;
	wire _w35958_ ;
	wire _w35957_ ;
	wire _w35956_ ;
	wire _w35955_ ;
	wire _w35954_ ;
	wire _w35953_ ;
	wire _w35952_ ;
	wire _w35951_ ;
	wire _w35950_ ;
	wire _w35949_ ;
	wire _w35948_ ;
	wire _w35947_ ;
	wire _w35946_ ;
	wire _w35945_ ;
	wire _w35944_ ;
	wire _w35943_ ;
	wire _w35942_ ;
	wire _w35941_ ;
	wire _w35940_ ;
	wire _w35939_ ;
	wire _w35938_ ;
	wire _w35937_ ;
	wire _w35936_ ;
	wire _w35935_ ;
	wire _w35934_ ;
	wire _w35933_ ;
	wire _w35932_ ;
	wire _w35931_ ;
	wire _w35930_ ;
	wire _w35929_ ;
	wire _w35928_ ;
	wire _w35927_ ;
	wire _w35926_ ;
	wire _w35925_ ;
	wire _w35924_ ;
	wire _w35923_ ;
	wire _w35922_ ;
	wire _w35921_ ;
	wire _w35920_ ;
	wire _w35919_ ;
	wire _w35918_ ;
	wire _w35917_ ;
	wire _w35916_ ;
	wire _w35915_ ;
	wire _w35914_ ;
	wire _w35913_ ;
	wire _w35912_ ;
	wire _w35911_ ;
	wire _w35910_ ;
	wire _w35909_ ;
	wire _w35908_ ;
	wire _w35907_ ;
	wire _w35906_ ;
	wire _w35905_ ;
	wire _w35904_ ;
	wire _w35903_ ;
	wire _w35902_ ;
	wire _w35901_ ;
	wire _w35900_ ;
	wire _w35899_ ;
	wire _w35898_ ;
	wire _w35897_ ;
	wire _w35896_ ;
	wire _w35895_ ;
	wire _w35894_ ;
	wire _w35893_ ;
	wire _w35892_ ;
	wire _w35891_ ;
	wire _w35890_ ;
	wire _w35889_ ;
	wire _w35888_ ;
	wire _w35887_ ;
	wire _w35886_ ;
	wire _w35885_ ;
	wire _w35884_ ;
	wire _w35883_ ;
	wire _w35882_ ;
	wire _w35881_ ;
	wire _w35880_ ;
	wire _w35879_ ;
	wire _w35878_ ;
	wire _w35877_ ;
	wire _w35876_ ;
	wire _w35875_ ;
	wire _w35874_ ;
	wire _w35873_ ;
	wire _w35872_ ;
	wire _w35871_ ;
	wire _w35870_ ;
	wire _w35869_ ;
	wire _w35868_ ;
	wire _w35867_ ;
	wire _w35866_ ;
	wire _w35865_ ;
	wire _w35864_ ;
	wire _w35863_ ;
	wire _w35862_ ;
	wire _w35861_ ;
	wire _w35860_ ;
	wire _w35859_ ;
	wire _w35858_ ;
	wire _w35857_ ;
	wire _w35856_ ;
	wire _w35855_ ;
	wire _w35854_ ;
	wire _w35853_ ;
	wire _w35852_ ;
	wire _w35851_ ;
	wire _w35850_ ;
	wire _w35849_ ;
	wire _w35848_ ;
	wire _w35847_ ;
	wire _w35846_ ;
	wire _w35845_ ;
	wire _w35844_ ;
	wire _w35843_ ;
	wire _w35842_ ;
	wire _w35841_ ;
	wire _w35840_ ;
	wire _w35839_ ;
	wire _w35838_ ;
	wire _w35837_ ;
	wire _w35836_ ;
	wire _w35835_ ;
	wire _w35834_ ;
	wire _w35833_ ;
	wire _w35832_ ;
	wire _w35831_ ;
	wire _w35830_ ;
	wire _w35829_ ;
	wire _w35828_ ;
	wire _w35827_ ;
	wire _w35826_ ;
	wire _w35825_ ;
	wire _w35824_ ;
	wire _w35823_ ;
	wire _w35822_ ;
	wire _w35821_ ;
	wire _w35820_ ;
	wire _w35819_ ;
	wire _w35818_ ;
	wire _w35817_ ;
	wire _w35816_ ;
	wire _w35815_ ;
	wire _w35814_ ;
	wire _w35813_ ;
	wire _w35812_ ;
	wire _w35811_ ;
	wire _w35810_ ;
	wire _w35809_ ;
	wire _w35808_ ;
	wire _w35807_ ;
	wire _w35806_ ;
	wire _w35805_ ;
	wire _w35804_ ;
	wire _w35803_ ;
	wire _w35802_ ;
	wire _w35801_ ;
	wire _w35800_ ;
	wire _w35799_ ;
	wire _w35798_ ;
	wire _w35797_ ;
	wire _w35796_ ;
	wire _w35795_ ;
	wire _w35794_ ;
	wire _w35793_ ;
	wire _w35792_ ;
	wire _w35791_ ;
	wire _w35790_ ;
	wire _w35789_ ;
	wire _w35788_ ;
	wire _w35787_ ;
	wire _w35786_ ;
	wire _w35785_ ;
	wire _w35784_ ;
	wire _w35783_ ;
	wire _w35782_ ;
	wire _w35781_ ;
	wire _w35780_ ;
	wire _w35779_ ;
	wire _w35778_ ;
	wire _w35777_ ;
	wire _w35776_ ;
	wire _w35775_ ;
	wire _w35774_ ;
	wire _w35773_ ;
	wire _w35772_ ;
	wire _w35771_ ;
	wire _w35770_ ;
	wire _w35769_ ;
	wire _w35768_ ;
	wire _w35767_ ;
	wire _w35766_ ;
	wire _w35765_ ;
	wire _w35764_ ;
	wire _w35763_ ;
	wire _w35762_ ;
	wire _w35761_ ;
	wire _w35760_ ;
	wire _w35759_ ;
	wire _w35758_ ;
	wire _w35757_ ;
	wire _w35756_ ;
	wire _w35755_ ;
	wire _w35754_ ;
	wire _w35753_ ;
	wire _w35752_ ;
	wire _w35751_ ;
	wire _w35750_ ;
	wire _w35749_ ;
	wire _w35748_ ;
	wire _w35747_ ;
	wire _w35746_ ;
	wire _w35745_ ;
	wire _w35744_ ;
	wire _w35743_ ;
	wire _w35742_ ;
	wire _w35741_ ;
	wire _w35740_ ;
	wire _w35739_ ;
	wire _w35738_ ;
	wire _w35737_ ;
	wire _w35736_ ;
	wire _w35735_ ;
	wire _w35734_ ;
	wire _w35733_ ;
	wire _w35732_ ;
	wire _w35731_ ;
	wire _w35730_ ;
	wire _w35729_ ;
	wire _w35728_ ;
	wire _w35727_ ;
	wire _w35726_ ;
	wire _w35725_ ;
	wire _w35724_ ;
	wire _w35723_ ;
	wire _w35722_ ;
	wire _w35721_ ;
	wire _w35720_ ;
	wire _w35719_ ;
	wire _w35718_ ;
	wire _w35717_ ;
	wire _w35716_ ;
	wire _w35715_ ;
	wire _w35714_ ;
	wire _w35713_ ;
	wire _w35712_ ;
	wire _w35711_ ;
	wire _w35710_ ;
	wire _w35709_ ;
	wire _w35708_ ;
	wire _w35707_ ;
	wire _w35706_ ;
	wire _w35705_ ;
	wire _w35704_ ;
	wire _w35703_ ;
	wire _w35702_ ;
	wire _w35701_ ;
	wire _w35700_ ;
	wire _w35699_ ;
	wire _w35698_ ;
	wire _w35697_ ;
	wire _w35696_ ;
	wire _w35695_ ;
	wire _w35694_ ;
	wire _w35693_ ;
	wire _w35692_ ;
	wire _w35691_ ;
	wire _w35690_ ;
	wire _w35689_ ;
	wire _w35688_ ;
	wire _w35687_ ;
	wire _w35686_ ;
	wire _w35685_ ;
	wire _w35684_ ;
	wire _w35683_ ;
	wire _w35682_ ;
	wire _w35681_ ;
	wire _w35680_ ;
	wire _w35679_ ;
	wire _w35678_ ;
	wire _w35677_ ;
	wire _w35676_ ;
	wire _w35675_ ;
	wire _w35674_ ;
	wire _w35673_ ;
	wire _w35672_ ;
	wire _w35671_ ;
	wire _w35670_ ;
	wire _w35669_ ;
	wire _w35668_ ;
	wire _w35667_ ;
	wire _w35666_ ;
	wire _w35665_ ;
	wire _w35664_ ;
	wire _w35663_ ;
	wire _w35662_ ;
	wire _w35661_ ;
	wire _w35660_ ;
	wire _w35659_ ;
	wire _w35658_ ;
	wire _w35657_ ;
	wire _w35656_ ;
	wire _w35655_ ;
	wire _w35654_ ;
	wire _w35653_ ;
	wire _w35652_ ;
	wire _w35651_ ;
	wire _w35650_ ;
	wire _w35649_ ;
	wire _w35648_ ;
	wire _w35647_ ;
	wire _w35646_ ;
	wire _w35645_ ;
	wire _w35644_ ;
	wire _w35643_ ;
	wire _w35642_ ;
	wire _w35641_ ;
	wire _w35640_ ;
	wire _w35639_ ;
	wire _w35638_ ;
	wire _w35637_ ;
	wire _w35636_ ;
	wire _w35635_ ;
	wire _w35634_ ;
	wire _w35633_ ;
	wire _w35632_ ;
	wire _w35631_ ;
	wire _w35630_ ;
	wire _w35629_ ;
	wire _w35628_ ;
	wire _w35627_ ;
	wire _w35626_ ;
	wire _w35625_ ;
	wire _w35624_ ;
	wire _w35623_ ;
	wire _w35622_ ;
	wire _w35621_ ;
	wire _w35620_ ;
	wire _w35619_ ;
	wire _w35618_ ;
	wire _w35617_ ;
	wire _w35616_ ;
	wire _w35615_ ;
	wire _w35614_ ;
	wire _w35613_ ;
	wire _w35612_ ;
	wire _w35611_ ;
	wire _w35610_ ;
	wire _w35609_ ;
	wire _w35608_ ;
	wire _w35607_ ;
	wire _w35606_ ;
	wire _w35605_ ;
	wire _w35604_ ;
	wire _w35603_ ;
	wire _w35602_ ;
	wire _w35601_ ;
	wire _w35600_ ;
	wire _w35599_ ;
	wire _w35598_ ;
	wire _w35597_ ;
	wire _w35596_ ;
	wire _w35595_ ;
	wire _w35594_ ;
	wire _w35593_ ;
	wire _w35592_ ;
	wire _w35591_ ;
	wire _w35590_ ;
	wire _w35589_ ;
	wire _w35588_ ;
	wire _w35587_ ;
	wire _w35586_ ;
	wire _w35585_ ;
	wire _w35584_ ;
	wire _w35583_ ;
	wire _w35582_ ;
	wire _w35581_ ;
	wire _w35580_ ;
	wire _w35579_ ;
	wire _w35578_ ;
	wire _w35577_ ;
	wire _w35576_ ;
	wire _w35575_ ;
	wire _w35574_ ;
	wire _w35573_ ;
	wire _w35572_ ;
	wire _w35571_ ;
	wire _w35570_ ;
	wire _w35569_ ;
	wire _w35568_ ;
	wire _w35567_ ;
	wire _w35566_ ;
	wire _w35565_ ;
	wire _w35564_ ;
	wire _w35563_ ;
	wire _w35562_ ;
	wire _w35561_ ;
	wire _w35560_ ;
	wire _w35559_ ;
	wire _w35558_ ;
	wire _w35557_ ;
	wire _w35556_ ;
	wire _w35555_ ;
	wire _w35554_ ;
	wire _w35553_ ;
	wire _w35552_ ;
	wire _w35551_ ;
	wire _w35550_ ;
	wire _w35549_ ;
	wire _w35548_ ;
	wire _w35547_ ;
	wire _w35546_ ;
	wire _w35545_ ;
	wire _w35544_ ;
	wire _w35543_ ;
	wire _w35542_ ;
	wire _w35541_ ;
	wire _w35540_ ;
	wire _w35539_ ;
	wire _w35538_ ;
	wire _w35537_ ;
	wire _w35536_ ;
	wire _w35535_ ;
	wire _w35534_ ;
	wire _w35533_ ;
	wire _w35532_ ;
	wire _w35531_ ;
	wire _w35530_ ;
	wire _w35529_ ;
	wire _w35528_ ;
	wire _w35527_ ;
	wire _w35526_ ;
	wire _w35525_ ;
	wire _w35524_ ;
	wire _w35523_ ;
	wire _w35522_ ;
	wire _w35521_ ;
	wire _w35520_ ;
	wire _w35519_ ;
	wire _w35518_ ;
	wire _w35517_ ;
	wire _w35516_ ;
	wire _w35515_ ;
	wire _w35514_ ;
	wire _w35513_ ;
	wire _w35512_ ;
	wire _w35511_ ;
	wire _w35510_ ;
	wire _w35509_ ;
	wire _w35508_ ;
	wire _w35507_ ;
	wire _w35506_ ;
	wire _w35505_ ;
	wire _w35504_ ;
	wire _w35503_ ;
	wire _w35502_ ;
	wire _w35501_ ;
	wire _w35500_ ;
	wire _w35499_ ;
	wire _w35498_ ;
	wire _w35497_ ;
	wire _w35496_ ;
	wire _w35495_ ;
	wire _w35494_ ;
	wire _w35493_ ;
	wire _w35492_ ;
	wire _w35491_ ;
	wire _w35490_ ;
	wire _w35489_ ;
	wire _w35488_ ;
	wire _w35487_ ;
	wire _w35486_ ;
	wire _w35485_ ;
	wire _w35484_ ;
	wire _w35483_ ;
	wire _w35482_ ;
	wire _w35481_ ;
	wire _w35480_ ;
	wire _w35479_ ;
	wire _w35478_ ;
	wire _w35477_ ;
	wire _w35476_ ;
	wire _w35475_ ;
	wire _w35474_ ;
	wire _w35473_ ;
	wire _w35472_ ;
	wire _w35471_ ;
	wire _w35470_ ;
	wire _w35469_ ;
	wire _w35468_ ;
	wire _w35467_ ;
	wire _w35466_ ;
	wire _w35465_ ;
	wire _w35464_ ;
	wire _w35463_ ;
	wire _w35462_ ;
	wire _w35461_ ;
	wire _w35460_ ;
	wire _w35459_ ;
	wire _w35458_ ;
	wire _w35457_ ;
	wire _w35456_ ;
	wire _w35455_ ;
	wire _w35454_ ;
	wire _w35453_ ;
	wire _w35452_ ;
	wire _w35451_ ;
	wire _w35450_ ;
	wire _w35449_ ;
	wire _w35448_ ;
	wire _w35447_ ;
	wire _w35446_ ;
	wire _w35445_ ;
	wire _w35444_ ;
	wire _w35443_ ;
	wire _w35442_ ;
	wire _w35441_ ;
	wire _w35440_ ;
	wire _w35439_ ;
	wire _w35438_ ;
	wire _w35437_ ;
	wire _w35436_ ;
	wire _w35435_ ;
	wire _w35434_ ;
	wire _w35433_ ;
	wire _w35432_ ;
	wire _w35431_ ;
	wire _w35430_ ;
	wire _w35429_ ;
	wire _w35428_ ;
	wire _w35427_ ;
	wire _w35426_ ;
	wire _w35425_ ;
	wire _w35424_ ;
	wire _w35423_ ;
	wire _w35422_ ;
	wire _w35421_ ;
	wire _w35420_ ;
	wire _w35419_ ;
	wire _w35418_ ;
	wire _w35417_ ;
	wire _w35416_ ;
	wire _w35415_ ;
	wire _w35414_ ;
	wire _w35413_ ;
	wire _w35412_ ;
	wire _w35411_ ;
	wire _w35410_ ;
	wire _w35409_ ;
	wire _w35408_ ;
	wire _w35407_ ;
	wire _w35406_ ;
	wire _w35405_ ;
	wire _w35404_ ;
	wire _w35403_ ;
	wire _w35402_ ;
	wire _w35401_ ;
	wire _w35400_ ;
	wire _w35399_ ;
	wire _w35398_ ;
	wire _w35397_ ;
	wire _w35396_ ;
	wire _w35395_ ;
	wire _w35394_ ;
	wire _w35393_ ;
	wire _w35392_ ;
	wire _w35391_ ;
	wire _w35390_ ;
	wire _w35389_ ;
	wire _w35388_ ;
	wire _w35387_ ;
	wire _w35386_ ;
	wire _w35385_ ;
	wire _w35384_ ;
	wire _w35383_ ;
	wire _w35382_ ;
	wire _w35381_ ;
	wire _w35380_ ;
	wire _w35379_ ;
	wire _w35378_ ;
	wire _w35377_ ;
	wire _w35376_ ;
	wire _w35375_ ;
	wire _w35374_ ;
	wire _w35373_ ;
	wire _w35372_ ;
	wire _w35371_ ;
	wire _w35370_ ;
	wire _w35369_ ;
	wire _w35368_ ;
	wire _w35367_ ;
	wire _w35366_ ;
	wire _w35365_ ;
	wire _w35364_ ;
	wire _w35363_ ;
	wire _w35362_ ;
	wire _w35361_ ;
	wire _w35360_ ;
	wire _w35359_ ;
	wire _w35358_ ;
	wire _w35357_ ;
	wire _w35356_ ;
	wire _w35355_ ;
	wire _w35354_ ;
	wire _w35353_ ;
	wire _w35352_ ;
	wire _w35351_ ;
	wire _w35350_ ;
	wire _w35349_ ;
	wire _w35348_ ;
	wire _w35347_ ;
	wire _w35346_ ;
	wire _w35345_ ;
	wire _w35344_ ;
	wire _w35343_ ;
	wire _w35342_ ;
	wire _w35341_ ;
	wire _w35340_ ;
	wire _w35339_ ;
	wire _w35338_ ;
	wire _w35337_ ;
	wire _w35336_ ;
	wire _w35335_ ;
	wire _w35334_ ;
	wire _w35333_ ;
	wire _w35332_ ;
	wire _w35331_ ;
	wire _w35330_ ;
	wire _w35329_ ;
	wire _w35328_ ;
	wire _w35327_ ;
	wire _w35326_ ;
	wire _w35325_ ;
	wire _w35324_ ;
	wire _w35323_ ;
	wire _w35322_ ;
	wire _w35321_ ;
	wire _w35320_ ;
	wire _w35319_ ;
	wire _w35318_ ;
	wire _w35317_ ;
	wire _w35316_ ;
	wire _w35315_ ;
	wire _w35314_ ;
	wire _w35313_ ;
	wire _w35312_ ;
	wire _w35311_ ;
	wire _w35310_ ;
	wire _w35309_ ;
	wire _w35308_ ;
	wire _w35307_ ;
	wire _w35306_ ;
	wire _w35305_ ;
	wire _w35304_ ;
	wire _w35303_ ;
	wire _w35302_ ;
	wire _w35301_ ;
	wire _w35300_ ;
	wire _w35299_ ;
	wire _w35298_ ;
	wire _w35297_ ;
	wire _w35296_ ;
	wire _w35295_ ;
	wire _w35294_ ;
	wire _w35293_ ;
	wire _w35292_ ;
	wire _w35291_ ;
	wire _w35290_ ;
	wire _w35289_ ;
	wire _w35288_ ;
	wire _w35287_ ;
	wire _w35286_ ;
	wire _w35285_ ;
	wire _w35284_ ;
	wire _w35283_ ;
	wire _w35282_ ;
	wire _w35281_ ;
	wire _w35280_ ;
	wire _w35279_ ;
	wire _w35278_ ;
	wire _w35277_ ;
	wire _w35276_ ;
	wire _w35275_ ;
	wire _w35274_ ;
	wire _w35273_ ;
	wire _w35272_ ;
	wire _w35271_ ;
	wire _w35270_ ;
	wire _w35269_ ;
	wire _w35268_ ;
	wire _w35267_ ;
	wire _w35266_ ;
	wire _w35265_ ;
	wire _w35264_ ;
	wire _w35263_ ;
	wire _w35262_ ;
	wire _w35261_ ;
	wire _w35260_ ;
	wire _w35259_ ;
	wire _w35258_ ;
	wire _w35257_ ;
	wire _w35256_ ;
	wire _w35255_ ;
	wire _w35254_ ;
	wire _w35253_ ;
	wire _w35252_ ;
	wire _w35251_ ;
	wire _w35250_ ;
	wire _w35249_ ;
	wire _w35248_ ;
	wire _w35247_ ;
	wire _w35246_ ;
	wire _w35245_ ;
	wire _w35244_ ;
	wire _w35243_ ;
	wire _w35242_ ;
	wire _w35241_ ;
	wire _w35240_ ;
	wire _w35239_ ;
	wire _w35238_ ;
	wire _w35237_ ;
	wire _w35236_ ;
	wire _w35235_ ;
	wire _w35234_ ;
	wire _w35233_ ;
	wire _w35232_ ;
	wire _w35231_ ;
	wire _w35230_ ;
	wire _w35229_ ;
	wire _w35228_ ;
	wire _w35227_ ;
	wire _w35226_ ;
	wire _w35225_ ;
	wire _w35224_ ;
	wire _w35223_ ;
	wire _w35222_ ;
	wire _w35221_ ;
	wire _w35220_ ;
	wire _w35219_ ;
	wire _w35218_ ;
	wire _w35217_ ;
	wire _w35216_ ;
	wire _w35215_ ;
	wire _w35214_ ;
	wire _w35213_ ;
	wire _w35212_ ;
	wire _w35211_ ;
	wire _w35210_ ;
	wire _w35209_ ;
	wire _w35208_ ;
	wire _w35207_ ;
	wire _w35206_ ;
	wire _w35205_ ;
	wire _w35204_ ;
	wire _w35203_ ;
	wire _w35202_ ;
	wire _w35201_ ;
	wire _w35200_ ;
	wire _w35199_ ;
	wire _w35198_ ;
	wire _w35197_ ;
	wire _w35196_ ;
	wire _w35195_ ;
	wire _w35194_ ;
	wire _w35193_ ;
	wire _w35192_ ;
	wire _w35191_ ;
	wire _w35190_ ;
	wire _w35189_ ;
	wire _w35188_ ;
	wire _w35187_ ;
	wire _w35186_ ;
	wire _w35185_ ;
	wire _w35184_ ;
	wire _w35183_ ;
	wire _w35182_ ;
	wire _w35181_ ;
	wire _w35180_ ;
	wire _w35179_ ;
	wire _w35178_ ;
	wire _w35177_ ;
	wire _w35176_ ;
	wire _w35175_ ;
	wire _w35174_ ;
	wire _w35173_ ;
	wire _w35172_ ;
	wire _w35171_ ;
	wire _w35170_ ;
	wire _w35169_ ;
	wire _w35168_ ;
	wire _w35167_ ;
	wire _w35166_ ;
	wire _w35165_ ;
	wire _w35164_ ;
	wire _w35163_ ;
	wire _w35162_ ;
	wire _w35161_ ;
	wire _w35160_ ;
	wire _w35159_ ;
	wire _w35158_ ;
	wire _w35157_ ;
	wire _w35156_ ;
	wire _w35155_ ;
	wire _w35154_ ;
	wire _w35153_ ;
	wire _w35152_ ;
	wire _w35151_ ;
	wire _w35150_ ;
	wire _w35149_ ;
	wire _w35148_ ;
	wire _w35147_ ;
	wire _w35146_ ;
	wire _w35145_ ;
	wire _w35144_ ;
	wire _w35143_ ;
	wire _w35142_ ;
	wire _w35141_ ;
	wire _w35140_ ;
	wire _w35139_ ;
	wire _w35138_ ;
	wire _w35137_ ;
	wire _w35136_ ;
	wire _w35135_ ;
	wire _w35134_ ;
	wire _w35133_ ;
	wire _w35132_ ;
	wire _w35131_ ;
	wire _w35130_ ;
	wire _w35129_ ;
	wire _w35128_ ;
	wire _w35127_ ;
	wire _w35126_ ;
	wire _w35125_ ;
	wire _w35124_ ;
	wire _w35123_ ;
	wire _w35122_ ;
	wire _w35121_ ;
	wire _w35120_ ;
	wire _w35119_ ;
	wire _w35118_ ;
	wire _w35117_ ;
	wire _w35116_ ;
	wire _w35115_ ;
	wire _w35114_ ;
	wire _w35113_ ;
	wire _w35112_ ;
	wire _w35111_ ;
	wire _w35110_ ;
	wire _w35109_ ;
	wire _w35108_ ;
	wire _w35107_ ;
	wire _w35106_ ;
	wire _w35105_ ;
	wire _w35104_ ;
	wire _w35103_ ;
	wire _w35102_ ;
	wire _w35101_ ;
	wire _w35100_ ;
	wire _w35099_ ;
	wire _w35098_ ;
	wire _w35097_ ;
	wire _w35096_ ;
	wire _w35095_ ;
	wire _w35094_ ;
	wire _w35093_ ;
	wire _w35092_ ;
	wire _w35091_ ;
	wire _w35090_ ;
	wire _w35089_ ;
	wire _w35088_ ;
	wire _w35087_ ;
	wire _w35086_ ;
	wire _w35085_ ;
	wire _w35084_ ;
	wire _w35083_ ;
	wire _w35082_ ;
	wire _w35081_ ;
	wire _w35080_ ;
	wire _w35079_ ;
	wire _w35078_ ;
	wire _w35077_ ;
	wire _w35076_ ;
	wire _w35075_ ;
	wire _w35074_ ;
	wire _w35073_ ;
	wire _w35072_ ;
	wire _w35071_ ;
	wire _w35070_ ;
	wire _w35069_ ;
	wire _w35068_ ;
	wire _w35067_ ;
	wire _w35066_ ;
	wire _w35065_ ;
	wire _w35064_ ;
	wire _w35063_ ;
	wire _w35062_ ;
	wire _w35061_ ;
	wire _w35060_ ;
	wire _w35059_ ;
	wire _w35058_ ;
	wire _w35057_ ;
	wire _w35056_ ;
	wire _w35055_ ;
	wire _w35054_ ;
	wire _w35053_ ;
	wire _w35052_ ;
	wire _w35051_ ;
	wire _w35050_ ;
	wire _w35049_ ;
	wire _w35048_ ;
	wire _w35047_ ;
	wire _w35046_ ;
	wire _w35045_ ;
	wire _w35044_ ;
	wire _w35043_ ;
	wire _w35042_ ;
	wire _w35041_ ;
	wire _w35040_ ;
	wire _w35039_ ;
	wire _w35038_ ;
	wire _w35037_ ;
	wire _w35036_ ;
	wire _w35035_ ;
	wire _w35034_ ;
	wire _w35033_ ;
	wire _w35032_ ;
	wire _w35031_ ;
	wire _w35030_ ;
	wire _w35029_ ;
	wire _w35028_ ;
	wire _w35027_ ;
	wire _w35026_ ;
	wire _w35025_ ;
	wire _w35024_ ;
	wire _w35023_ ;
	wire _w35022_ ;
	wire _w35021_ ;
	wire _w35020_ ;
	wire _w35019_ ;
	wire _w35018_ ;
	wire _w35017_ ;
	wire _w35016_ ;
	wire _w35015_ ;
	wire _w35014_ ;
	wire _w35013_ ;
	wire _w35012_ ;
	wire _w35011_ ;
	wire _w35010_ ;
	wire _w35009_ ;
	wire _w35008_ ;
	wire _w35007_ ;
	wire _w35006_ ;
	wire _w35005_ ;
	wire _w35004_ ;
	wire _w35003_ ;
	wire _w35002_ ;
	wire _w35001_ ;
	wire _w35000_ ;
	wire _w34999_ ;
	wire _w34998_ ;
	wire _w34997_ ;
	wire _w34996_ ;
	wire _w34995_ ;
	wire _w34994_ ;
	wire _w34993_ ;
	wire _w34992_ ;
	wire _w34991_ ;
	wire _w34990_ ;
	wire _w34989_ ;
	wire _w34988_ ;
	wire _w34987_ ;
	wire _w34986_ ;
	wire _w34985_ ;
	wire _w34984_ ;
	wire _w34983_ ;
	wire _w34982_ ;
	wire _w34981_ ;
	wire _w34980_ ;
	wire _w34979_ ;
	wire _w34978_ ;
	wire _w34977_ ;
	wire _w34976_ ;
	wire _w34975_ ;
	wire _w34974_ ;
	wire _w34973_ ;
	wire _w34972_ ;
	wire _w34971_ ;
	wire _w34970_ ;
	wire _w34969_ ;
	wire _w34968_ ;
	wire _w34967_ ;
	wire _w34966_ ;
	wire _w34965_ ;
	wire _w34964_ ;
	wire _w34963_ ;
	wire _w34962_ ;
	wire _w34961_ ;
	wire _w34960_ ;
	wire _w34959_ ;
	wire _w34958_ ;
	wire _w34957_ ;
	wire _w34956_ ;
	wire _w34955_ ;
	wire _w34954_ ;
	wire _w34953_ ;
	wire _w34952_ ;
	wire _w34951_ ;
	wire _w34950_ ;
	wire _w34949_ ;
	wire _w34948_ ;
	wire _w34947_ ;
	wire _w34946_ ;
	wire _w34945_ ;
	wire _w34944_ ;
	wire _w34943_ ;
	wire _w34942_ ;
	wire _w34941_ ;
	wire _w34940_ ;
	wire _w34939_ ;
	wire _w34938_ ;
	wire _w34937_ ;
	wire _w34936_ ;
	wire _w34935_ ;
	wire _w34934_ ;
	wire _w34933_ ;
	wire _w34932_ ;
	wire _w34931_ ;
	wire _w34930_ ;
	wire _w34929_ ;
	wire _w34928_ ;
	wire _w34927_ ;
	wire _w34926_ ;
	wire _w34925_ ;
	wire _w34924_ ;
	wire _w34923_ ;
	wire _w34922_ ;
	wire _w34921_ ;
	wire _w34920_ ;
	wire _w34919_ ;
	wire _w34918_ ;
	wire _w34917_ ;
	wire _w34916_ ;
	wire _w34915_ ;
	wire _w34914_ ;
	wire _w34913_ ;
	wire _w34912_ ;
	wire _w34911_ ;
	wire _w34910_ ;
	wire _w34909_ ;
	wire _w34908_ ;
	wire _w34907_ ;
	wire _w34906_ ;
	wire _w34905_ ;
	wire _w34904_ ;
	wire _w34903_ ;
	wire _w34902_ ;
	wire _w34901_ ;
	wire _w34900_ ;
	wire _w34899_ ;
	wire _w34898_ ;
	wire _w34897_ ;
	wire _w34896_ ;
	wire _w34895_ ;
	wire _w34894_ ;
	wire _w34893_ ;
	wire _w34892_ ;
	wire _w34891_ ;
	wire _w34890_ ;
	wire _w34889_ ;
	wire _w34888_ ;
	wire _w34887_ ;
	wire _w34886_ ;
	wire _w34885_ ;
	wire _w34884_ ;
	wire _w34883_ ;
	wire _w34882_ ;
	wire _w34881_ ;
	wire _w34880_ ;
	wire _w34879_ ;
	wire _w34878_ ;
	wire _w34877_ ;
	wire _w34876_ ;
	wire _w34875_ ;
	wire _w34874_ ;
	wire _w34873_ ;
	wire _w34872_ ;
	wire _w34871_ ;
	wire _w34870_ ;
	wire _w34869_ ;
	wire _w34868_ ;
	wire _w34867_ ;
	wire _w34866_ ;
	wire _w34865_ ;
	wire _w34864_ ;
	wire _w34863_ ;
	wire _w34862_ ;
	wire _w34861_ ;
	wire _w34860_ ;
	wire _w34859_ ;
	wire _w34858_ ;
	wire _w34857_ ;
	wire _w34856_ ;
	wire _w34855_ ;
	wire _w34854_ ;
	wire _w34853_ ;
	wire _w34852_ ;
	wire _w34851_ ;
	wire _w34850_ ;
	wire _w34849_ ;
	wire _w34848_ ;
	wire _w34847_ ;
	wire _w34846_ ;
	wire _w34845_ ;
	wire _w34844_ ;
	wire _w34843_ ;
	wire _w34842_ ;
	wire _w34841_ ;
	wire _w34840_ ;
	wire _w34839_ ;
	wire _w34838_ ;
	wire _w34837_ ;
	wire _w34836_ ;
	wire _w34835_ ;
	wire _w34834_ ;
	wire _w34833_ ;
	wire _w34832_ ;
	wire _w34831_ ;
	wire _w34830_ ;
	wire _w34829_ ;
	wire _w34828_ ;
	wire _w34827_ ;
	wire _w34826_ ;
	wire _w34825_ ;
	wire _w34824_ ;
	wire _w34823_ ;
	wire _w34822_ ;
	wire _w34821_ ;
	wire _w34820_ ;
	wire _w34819_ ;
	wire _w34818_ ;
	wire _w34817_ ;
	wire _w34816_ ;
	wire _w34815_ ;
	wire _w34814_ ;
	wire _w34813_ ;
	wire _w34812_ ;
	wire _w34811_ ;
	wire _w34810_ ;
	wire _w34809_ ;
	wire _w34808_ ;
	wire _w34807_ ;
	wire _w34806_ ;
	wire _w34805_ ;
	wire _w34804_ ;
	wire _w34803_ ;
	wire _w34802_ ;
	wire _w34801_ ;
	wire _w34800_ ;
	wire _w34799_ ;
	wire _w34798_ ;
	wire _w34797_ ;
	wire _w34796_ ;
	wire _w34795_ ;
	wire _w34794_ ;
	wire _w34793_ ;
	wire _w34792_ ;
	wire _w34791_ ;
	wire _w34790_ ;
	wire _w34789_ ;
	wire _w34788_ ;
	wire _w34787_ ;
	wire _w34786_ ;
	wire _w34785_ ;
	wire _w34784_ ;
	wire _w34783_ ;
	wire _w34782_ ;
	wire _w34781_ ;
	wire _w34780_ ;
	wire _w34779_ ;
	wire _w34778_ ;
	wire _w34777_ ;
	wire _w34776_ ;
	wire _w34775_ ;
	wire _w34774_ ;
	wire _w34773_ ;
	wire _w34772_ ;
	wire _w34771_ ;
	wire _w34770_ ;
	wire _w34769_ ;
	wire _w34768_ ;
	wire _w34767_ ;
	wire _w34766_ ;
	wire _w34765_ ;
	wire _w34764_ ;
	wire _w34763_ ;
	wire _w34762_ ;
	wire _w34761_ ;
	wire _w34760_ ;
	wire _w34759_ ;
	wire _w34758_ ;
	wire _w34757_ ;
	wire _w34756_ ;
	wire _w34755_ ;
	wire _w34754_ ;
	wire _w34753_ ;
	wire _w34752_ ;
	wire _w34751_ ;
	wire _w34750_ ;
	wire _w34749_ ;
	wire _w34748_ ;
	wire _w34747_ ;
	wire _w34746_ ;
	wire _w34745_ ;
	wire _w34744_ ;
	wire _w34743_ ;
	wire _w34742_ ;
	wire _w34741_ ;
	wire _w34740_ ;
	wire _w34739_ ;
	wire _w34738_ ;
	wire _w34737_ ;
	wire _w34736_ ;
	wire _w34735_ ;
	wire _w34734_ ;
	wire _w34733_ ;
	wire _w34732_ ;
	wire _w34731_ ;
	wire _w34730_ ;
	wire _w34729_ ;
	wire _w34728_ ;
	wire _w34727_ ;
	wire _w34726_ ;
	wire _w34725_ ;
	wire _w34724_ ;
	wire _w34723_ ;
	wire _w34722_ ;
	wire _w34721_ ;
	wire _w34720_ ;
	wire _w34719_ ;
	wire _w34718_ ;
	wire _w34717_ ;
	wire _w34716_ ;
	wire _w34715_ ;
	wire _w34714_ ;
	wire _w34713_ ;
	wire _w34712_ ;
	wire _w34711_ ;
	wire _w34710_ ;
	wire _w34709_ ;
	wire _w34708_ ;
	wire _w34707_ ;
	wire _w34706_ ;
	wire _w34705_ ;
	wire _w34704_ ;
	wire _w34703_ ;
	wire _w34702_ ;
	wire _w34701_ ;
	wire _w34700_ ;
	wire _w34699_ ;
	wire _w34698_ ;
	wire _w34697_ ;
	wire _w34696_ ;
	wire _w34695_ ;
	wire _w34694_ ;
	wire _w34693_ ;
	wire _w34692_ ;
	wire _w34691_ ;
	wire _w34690_ ;
	wire _w34689_ ;
	wire _w34688_ ;
	wire _w34687_ ;
	wire _w34686_ ;
	wire _w34685_ ;
	wire _w34684_ ;
	wire _w34683_ ;
	wire _w34682_ ;
	wire _w34681_ ;
	wire _w34680_ ;
	wire _w34679_ ;
	wire _w34678_ ;
	wire _w34677_ ;
	wire _w34676_ ;
	wire _w34675_ ;
	wire _w34674_ ;
	wire _w34673_ ;
	wire _w34672_ ;
	wire _w34671_ ;
	wire _w34670_ ;
	wire _w34669_ ;
	wire _w34668_ ;
	wire _w34667_ ;
	wire _w34666_ ;
	wire _w34665_ ;
	wire _w34664_ ;
	wire _w34663_ ;
	wire _w34662_ ;
	wire _w34661_ ;
	wire _w34660_ ;
	wire _w34659_ ;
	wire _w34658_ ;
	wire _w34657_ ;
	wire _w34656_ ;
	wire _w34655_ ;
	wire _w34654_ ;
	wire _w34653_ ;
	wire _w34652_ ;
	wire _w34651_ ;
	wire _w34650_ ;
	wire _w34649_ ;
	wire _w34648_ ;
	wire _w34647_ ;
	wire _w34646_ ;
	wire _w34645_ ;
	wire _w34644_ ;
	wire _w34643_ ;
	wire _w34642_ ;
	wire _w34641_ ;
	wire _w34640_ ;
	wire _w34639_ ;
	wire _w34638_ ;
	wire _w34637_ ;
	wire _w34636_ ;
	wire _w34635_ ;
	wire _w34634_ ;
	wire _w34633_ ;
	wire _w34632_ ;
	wire _w34631_ ;
	wire _w34630_ ;
	wire _w34629_ ;
	wire _w34628_ ;
	wire _w34627_ ;
	wire _w34626_ ;
	wire _w34625_ ;
	wire _w34624_ ;
	wire _w34623_ ;
	wire _w34622_ ;
	wire _w34621_ ;
	wire _w34620_ ;
	wire _w34619_ ;
	wire _w34618_ ;
	wire _w34617_ ;
	wire _w34616_ ;
	wire _w34615_ ;
	wire _w34614_ ;
	wire _w34613_ ;
	wire _w34612_ ;
	wire _w34611_ ;
	wire _w34610_ ;
	wire _w34609_ ;
	wire _w34608_ ;
	wire _w34607_ ;
	wire _w34606_ ;
	wire _w34605_ ;
	wire _w34604_ ;
	wire _w34603_ ;
	wire _w34602_ ;
	wire _w34601_ ;
	wire _w34600_ ;
	wire _w34599_ ;
	wire _w34598_ ;
	wire _w34597_ ;
	wire _w34596_ ;
	wire _w34595_ ;
	wire _w34594_ ;
	wire _w34593_ ;
	wire _w34592_ ;
	wire _w34591_ ;
	wire _w34590_ ;
	wire _w34589_ ;
	wire _w34588_ ;
	wire _w34587_ ;
	wire _w34586_ ;
	wire _w34585_ ;
	wire _w34584_ ;
	wire _w34583_ ;
	wire _w34582_ ;
	wire _w34581_ ;
	wire _w34580_ ;
	wire _w34579_ ;
	wire _w34578_ ;
	wire _w34577_ ;
	wire _w34576_ ;
	wire _w34575_ ;
	wire _w34574_ ;
	wire _w34573_ ;
	wire _w34572_ ;
	wire _w34571_ ;
	wire _w34570_ ;
	wire _w34569_ ;
	wire _w34568_ ;
	wire _w34567_ ;
	wire _w34566_ ;
	wire _w34565_ ;
	wire _w34564_ ;
	wire _w34563_ ;
	wire _w34562_ ;
	wire _w34561_ ;
	wire _w34560_ ;
	wire _w34559_ ;
	wire _w34558_ ;
	wire _w34557_ ;
	wire _w34556_ ;
	wire _w34555_ ;
	wire _w34554_ ;
	wire _w34553_ ;
	wire _w34552_ ;
	wire _w34551_ ;
	wire _w34550_ ;
	wire _w34549_ ;
	wire _w34548_ ;
	wire _w34547_ ;
	wire _w34546_ ;
	wire _w34545_ ;
	wire _w34544_ ;
	wire _w34543_ ;
	wire _w34542_ ;
	wire _w34541_ ;
	wire _w34540_ ;
	wire _w34539_ ;
	wire _w34538_ ;
	wire _w34537_ ;
	wire _w34536_ ;
	wire _w34535_ ;
	wire _w34534_ ;
	wire _w34533_ ;
	wire _w34532_ ;
	wire _w34531_ ;
	wire _w34530_ ;
	wire _w34529_ ;
	wire _w34528_ ;
	wire _w34527_ ;
	wire _w34526_ ;
	wire _w34525_ ;
	wire _w34524_ ;
	wire _w34523_ ;
	wire _w34522_ ;
	wire _w34521_ ;
	wire _w34520_ ;
	wire _w34519_ ;
	wire _w34518_ ;
	wire _w34517_ ;
	wire _w34516_ ;
	wire _w34515_ ;
	wire _w34514_ ;
	wire _w34513_ ;
	wire _w34512_ ;
	wire _w34511_ ;
	wire _w34510_ ;
	wire _w34509_ ;
	wire _w34508_ ;
	wire _w34507_ ;
	wire _w34506_ ;
	wire _w34505_ ;
	wire _w34504_ ;
	wire _w34503_ ;
	wire _w34502_ ;
	wire _w34501_ ;
	wire _w34500_ ;
	wire _w34499_ ;
	wire _w34498_ ;
	wire _w34497_ ;
	wire _w34496_ ;
	wire _w34495_ ;
	wire _w34494_ ;
	wire _w34493_ ;
	wire _w34492_ ;
	wire _w34491_ ;
	wire _w34490_ ;
	wire _w34489_ ;
	wire _w34488_ ;
	wire _w34487_ ;
	wire _w34486_ ;
	wire _w34485_ ;
	wire _w34484_ ;
	wire _w34483_ ;
	wire _w34482_ ;
	wire _w34481_ ;
	wire _w34480_ ;
	wire _w34479_ ;
	wire _w34478_ ;
	wire _w34477_ ;
	wire _w34476_ ;
	wire _w34475_ ;
	wire _w34474_ ;
	wire _w34473_ ;
	wire _w34472_ ;
	wire _w34471_ ;
	wire _w34470_ ;
	wire _w34469_ ;
	wire _w34468_ ;
	wire _w34467_ ;
	wire _w34466_ ;
	wire _w34465_ ;
	wire _w34464_ ;
	wire _w34463_ ;
	wire _w34462_ ;
	wire _w34461_ ;
	wire _w34460_ ;
	wire _w34459_ ;
	wire _w34458_ ;
	wire _w34457_ ;
	wire _w34456_ ;
	wire _w34455_ ;
	wire _w34454_ ;
	wire _w34453_ ;
	wire _w34452_ ;
	wire _w34451_ ;
	wire _w34450_ ;
	wire _w34449_ ;
	wire _w34448_ ;
	wire _w34447_ ;
	wire _w34446_ ;
	wire _w34445_ ;
	wire _w34444_ ;
	wire _w34443_ ;
	wire _w34442_ ;
	wire _w34441_ ;
	wire _w34440_ ;
	wire _w34439_ ;
	wire _w34438_ ;
	wire _w34437_ ;
	wire _w34436_ ;
	wire _w34435_ ;
	wire _w34434_ ;
	wire _w34433_ ;
	wire _w34432_ ;
	wire _w34431_ ;
	wire _w34430_ ;
	wire _w34429_ ;
	wire _w34428_ ;
	wire _w34427_ ;
	wire _w34426_ ;
	wire _w34425_ ;
	wire _w34424_ ;
	wire _w34423_ ;
	wire _w34422_ ;
	wire _w34421_ ;
	wire _w34420_ ;
	wire _w34419_ ;
	wire _w34418_ ;
	wire _w34417_ ;
	wire _w34416_ ;
	wire _w34415_ ;
	wire _w34414_ ;
	wire _w34413_ ;
	wire _w34412_ ;
	wire _w34411_ ;
	wire _w34410_ ;
	wire _w34409_ ;
	wire _w34408_ ;
	wire _w34407_ ;
	wire _w34406_ ;
	wire _w34405_ ;
	wire _w34404_ ;
	wire _w34403_ ;
	wire _w34402_ ;
	wire _w34401_ ;
	wire _w34400_ ;
	wire _w34399_ ;
	wire _w34398_ ;
	wire _w34397_ ;
	wire _w34396_ ;
	wire _w34395_ ;
	wire _w34394_ ;
	wire _w34393_ ;
	wire _w34392_ ;
	wire _w34391_ ;
	wire _w34390_ ;
	wire _w34389_ ;
	wire _w34388_ ;
	wire _w34387_ ;
	wire _w34386_ ;
	wire _w34385_ ;
	wire _w34384_ ;
	wire _w34383_ ;
	wire _w34382_ ;
	wire _w34381_ ;
	wire _w34380_ ;
	wire _w34379_ ;
	wire _w34378_ ;
	wire _w34377_ ;
	wire _w34376_ ;
	wire _w34375_ ;
	wire _w34374_ ;
	wire _w34373_ ;
	wire _w34372_ ;
	wire _w34371_ ;
	wire _w34370_ ;
	wire _w34369_ ;
	wire _w34368_ ;
	wire _w34367_ ;
	wire _w34366_ ;
	wire _w34365_ ;
	wire _w34364_ ;
	wire _w34363_ ;
	wire _w34362_ ;
	wire _w34361_ ;
	wire _w34360_ ;
	wire _w34359_ ;
	wire _w34358_ ;
	wire _w34357_ ;
	wire _w34356_ ;
	wire _w34355_ ;
	wire _w34354_ ;
	wire _w34353_ ;
	wire _w34352_ ;
	wire _w34351_ ;
	wire _w34350_ ;
	wire _w34349_ ;
	wire _w34348_ ;
	wire _w34347_ ;
	wire _w34346_ ;
	wire _w34345_ ;
	wire _w34344_ ;
	wire _w34343_ ;
	wire _w34342_ ;
	wire _w34341_ ;
	wire _w34340_ ;
	wire _w34339_ ;
	wire _w34338_ ;
	wire _w34337_ ;
	wire _w34336_ ;
	wire _w34335_ ;
	wire _w34334_ ;
	wire _w34333_ ;
	wire _w34332_ ;
	wire _w34331_ ;
	wire _w34330_ ;
	wire _w34329_ ;
	wire _w34328_ ;
	wire _w34327_ ;
	wire _w34326_ ;
	wire _w34325_ ;
	wire _w34324_ ;
	wire _w34323_ ;
	wire _w34322_ ;
	wire _w34321_ ;
	wire _w34320_ ;
	wire _w34319_ ;
	wire _w34318_ ;
	wire _w34317_ ;
	wire _w34316_ ;
	wire _w34315_ ;
	wire _w34314_ ;
	wire _w34313_ ;
	wire _w34312_ ;
	wire _w34311_ ;
	wire _w34310_ ;
	wire _w34309_ ;
	wire _w34308_ ;
	wire _w34307_ ;
	wire _w34306_ ;
	wire _w34305_ ;
	wire _w34304_ ;
	wire _w34303_ ;
	wire _w34302_ ;
	wire _w34301_ ;
	wire _w34300_ ;
	wire _w34299_ ;
	wire _w34298_ ;
	wire _w34297_ ;
	wire _w34296_ ;
	wire _w34295_ ;
	wire _w34294_ ;
	wire _w34293_ ;
	wire _w34292_ ;
	wire _w34291_ ;
	wire _w34290_ ;
	wire _w34289_ ;
	wire _w34288_ ;
	wire _w34287_ ;
	wire _w34286_ ;
	wire _w34285_ ;
	wire _w34284_ ;
	wire _w34283_ ;
	wire _w34282_ ;
	wire _w34281_ ;
	wire _w34280_ ;
	wire _w34279_ ;
	wire _w34278_ ;
	wire _w34277_ ;
	wire _w34276_ ;
	wire _w34275_ ;
	wire _w34274_ ;
	wire _w34273_ ;
	wire _w34272_ ;
	wire _w34271_ ;
	wire _w34270_ ;
	wire _w34269_ ;
	wire _w34268_ ;
	wire _w34267_ ;
	wire _w34266_ ;
	wire _w34265_ ;
	wire _w34264_ ;
	wire _w34263_ ;
	wire _w34262_ ;
	wire _w34261_ ;
	wire _w34260_ ;
	wire _w34259_ ;
	wire _w34258_ ;
	wire _w34257_ ;
	wire _w34256_ ;
	wire _w34255_ ;
	wire _w34254_ ;
	wire _w34253_ ;
	wire _w34252_ ;
	wire _w34251_ ;
	wire _w34250_ ;
	wire _w34249_ ;
	wire _w34248_ ;
	wire _w34247_ ;
	wire _w34246_ ;
	wire _w34245_ ;
	wire _w34244_ ;
	wire _w34243_ ;
	wire _w34242_ ;
	wire _w34241_ ;
	wire _w34240_ ;
	wire _w34239_ ;
	wire _w34238_ ;
	wire _w34237_ ;
	wire _w34236_ ;
	wire _w34235_ ;
	wire _w34234_ ;
	wire _w34233_ ;
	wire _w34232_ ;
	wire _w34231_ ;
	wire _w34230_ ;
	wire _w34229_ ;
	wire _w34228_ ;
	wire _w34227_ ;
	wire _w34226_ ;
	wire _w34225_ ;
	wire _w34224_ ;
	wire _w34223_ ;
	wire _w34222_ ;
	wire _w34221_ ;
	wire _w34220_ ;
	wire _w34219_ ;
	wire _w34218_ ;
	wire _w34217_ ;
	wire _w34216_ ;
	wire _w34215_ ;
	wire _w34214_ ;
	wire _w34213_ ;
	wire _w34212_ ;
	wire _w34211_ ;
	wire _w34210_ ;
	wire _w34209_ ;
	wire _w34208_ ;
	wire _w34207_ ;
	wire _w34206_ ;
	wire _w34205_ ;
	wire _w34204_ ;
	wire _w34203_ ;
	wire _w34202_ ;
	wire _w34201_ ;
	wire _w34200_ ;
	wire _w34199_ ;
	wire _w34198_ ;
	wire _w34197_ ;
	wire _w34196_ ;
	wire _w34195_ ;
	wire _w34194_ ;
	wire _w34193_ ;
	wire _w34192_ ;
	wire _w34191_ ;
	wire _w34190_ ;
	wire _w34189_ ;
	wire _w34188_ ;
	wire _w34187_ ;
	wire _w34186_ ;
	wire _w34185_ ;
	wire _w34184_ ;
	wire _w34183_ ;
	wire _w34182_ ;
	wire _w34181_ ;
	wire _w34180_ ;
	wire _w34179_ ;
	wire _w34178_ ;
	wire _w34177_ ;
	wire _w34176_ ;
	wire _w34175_ ;
	wire _w34174_ ;
	wire _w34173_ ;
	wire _w34172_ ;
	wire _w34171_ ;
	wire _w34170_ ;
	wire _w34169_ ;
	wire _w34168_ ;
	wire _w34167_ ;
	wire _w34166_ ;
	wire _w34165_ ;
	wire _w34164_ ;
	wire _w34163_ ;
	wire _w34162_ ;
	wire _w34161_ ;
	wire _w34160_ ;
	wire _w34159_ ;
	wire _w34158_ ;
	wire _w34157_ ;
	wire _w34156_ ;
	wire _w34155_ ;
	wire _w34154_ ;
	wire _w34153_ ;
	wire _w34152_ ;
	wire _w34151_ ;
	wire _w34150_ ;
	wire _w34149_ ;
	wire _w34148_ ;
	wire _w34147_ ;
	wire _w34146_ ;
	wire _w34145_ ;
	wire _w34144_ ;
	wire _w34143_ ;
	wire _w34142_ ;
	wire _w34141_ ;
	wire _w34140_ ;
	wire _w34139_ ;
	wire _w34138_ ;
	wire _w34137_ ;
	wire _w34136_ ;
	wire _w34135_ ;
	wire _w34134_ ;
	wire _w34133_ ;
	wire _w34132_ ;
	wire _w34131_ ;
	wire _w34130_ ;
	wire _w34129_ ;
	wire _w34128_ ;
	wire _w34127_ ;
	wire _w34126_ ;
	wire _w34125_ ;
	wire _w34124_ ;
	wire _w34123_ ;
	wire _w34122_ ;
	wire _w34121_ ;
	wire _w34120_ ;
	wire _w34119_ ;
	wire _w34118_ ;
	wire _w34117_ ;
	wire _w34116_ ;
	wire _w34115_ ;
	wire _w34114_ ;
	wire _w34113_ ;
	wire _w34112_ ;
	wire _w34111_ ;
	wire _w34110_ ;
	wire _w34109_ ;
	wire _w34108_ ;
	wire _w34107_ ;
	wire _w34106_ ;
	wire _w34105_ ;
	wire _w34104_ ;
	wire _w34103_ ;
	wire _w34102_ ;
	wire _w34101_ ;
	wire _w34100_ ;
	wire _w34099_ ;
	wire _w34098_ ;
	wire _w34097_ ;
	wire _w34096_ ;
	wire _w34095_ ;
	wire _w34094_ ;
	wire _w34093_ ;
	wire _w34092_ ;
	wire _w34091_ ;
	wire _w34090_ ;
	wire _w34089_ ;
	wire _w34088_ ;
	wire _w34087_ ;
	wire _w34086_ ;
	wire _w34085_ ;
	wire _w34084_ ;
	wire _w34083_ ;
	wire _w34082_ ;
	wire _w34081_ ;
	wire _w34080_ ;
	wire _w34079_ ;
	wire _w34078_ ;
	wire _w34077_ ;
	wire _w34076_ ;
	wire _w34075_ ;
	wire _w34074_ ;
	wire _w34073_ ;
	wire _w34072_ ;
	wire _w34071_ ;
	wire _w34070_ ;
	wire _w34069_ ;
	wire _w34068_ ;
	wire _w34067_ ;
	wire _w34066_ ;
	wire _w34065_ ;
	wire _w34064_ ;
	wire _w34063_ ;
	wire _w34062_ ;
	wire _w34061_ ;
	wire _w34060_ ;
	wire _w34059_ ;
	wire _w34058_ ;
	wire _w34057_ ;
	wire _w34056_ ;
	wire _w34055_ ;
	wire _w34054_ ;
	wire _w34053_ ;
	wire _w34052_ ;
	wire _w34051_ ;
	wire _w34050_ ;
	wire _w34049_ ;
	wire _w34048_ ;
	wire _w34047_ ;
	wire _w34046_ ;
	wire _w34045_ ;
	wire _w34044_ ;
	wire _w34043_ ;
	wire _w34042_ ;
	wire _w34041_ ;
	wire _w34040_ ;
	wire _w34039_ ;
	wire _w34038_ ;
	wire _w34037_ ;
	wire _w34036_ ;
	wire _w34035_ ;
	wire _w34034_ ;
	wire _w34033_ ;
	wire _w34032_ ;
	wire _w34031_ ;
	wire _w34030_ ;
	wire _w34029_ ;
	wire _w34028_ ;
	wire _w34027_ ;
	wire _w34026_ ;
	wire _w34025_ ;
	wire _w34024_ ;
	wire _w34023_ ;
	wire _w34022_ ;
	wire _w34021_ ;
	wire _w34020_ ;
	wire _w34019_ ;
	wire _w34018_ ;
	wire _w34017_ ;
	wire _w34016_ ;
	wire _w34015_ ;
	wire _w34014_ ;
	wire _w34013_ ;
	wire _w34012_ ;
	wire _w34011_ ;
	wire _w34010_ ;
	wire _w34009_ ;
	wire _w34008_ ;
	wire _w34007_ ;
	wire _w34006_ ;
	wire _w34005_ ;
	wire _w34004_ ;
	wire _w34003_ ;
	wire _w34002_ ;
	wire _w34001_ ;
	wire _w34000_ ;
	wire _w33999_ ;
	wire _w33998_ ;
	wire _w33997_ ;
	wire _w33996_ ;
	wire _w33995_ ;
	wire _w33994_ ;
	wire _w33993_ ;
	wire _w33992_ ;
	wire _w33991_ ;
	wire _w33990_ ;
	wire _w33989_ ;
	wire _w33988_ ;
	wire _w33987_ ;
	wire _w33986_ ;
	wire _w33985_ ;
	wire _w33984_ ;
	wire _w33983_ ;
	wire _w33982_ ;
	wire _w33981_ ;
	wire _w33980_ ;
	wire _w33979_ ;
	wire _w33978_ ;
	wire _w33977_ ;
	wire _w33976_ ;
	wire _w33975_ ;
	wire _w33974_ ;
	wire _w33973_ ;
	wire _w33972_ ;
	wire _w33971_ ;
	wire _w33970_ ;
	wire _w33969_ ;
	wire _w33968_ ;
	wire _w33967_ ;
	wire _w33966_ ;
	wire _w33965_ ;
	wire _w33964_ ;
	wire _w33963_ ;
	wire _w33962_ ;
	wire _w33961_ ;
	wire _w33960_ ;
	wire _w33959_ ;
	wire _w33958_ ;
	wire _w33957_ ;
	wire _w33956_ ;
	wire _w33955_ ;
	wire _w33954_ ;
	wire _w33953_ ;
	wire _w33952_ ;
	wire _w33951_ ;
	wire _w33950_ ;
	wire _w33949_ ;
	wire _w33948_ ;
	wire _w33947_ ;
	wire _w33946_ ;
	wire _w33945_ ;
	wire _w33944_ ;
	wire _w33943_ ;
	wire _w33942_ ;
	wire _w33941_ ;
	wire _w33940_ ;
	wire _w33939_ ;
	wire _w33938_ ;
	wire _w33937_ ;
	wire _w33936_ ;
	wire _w33935_ ;
	wire _w33934_ ;
	wire _w33933_ ;
	wire _w33932_ ;
	wire _w33931_ ;
	wire _w33930_ ;
	wire _w33929_ ;
	wire _w33928_ ;
	wire _w33927_ ;
	wire _w33926_ ;
	wire _w33925_ ;
	wire _w33924_ ;
	wire _w33923_ ;
	wire _w33922_ ;
	wire _w33921_ ;
	wire _w33920_ ;
	wire _w33919_ ;
	wire _w33918_ ;
	wire _w33917_ ;
	wire _w33916_ ;
	wire _w33915_ ;
	wire _w33914_ ;
	wire _w33913_ ;
	wire _w33912_ ;
	wire _w33911_ ;
	wire _w33910_ ;
	wire _w33909_ ;
	wire _w33908_ ;
	wire _w33907_ ;
	wire _w33906_ ;
	wire _w33905_ ;
	wire _w33904_ ;
	wire _w33903_ ;
	wire _w33902_ ;
	wire _w33901_ ;
	wire _w33900_ ;
	wire _w33899_ ;
	wire _w33898_ ;
	wire _w33897_ ;
	wire _w33896_ ;
	wire _w33895_ ;
	wire _w33894_ ;
	wire _w33893_ ;
	wire _w33892_ ;
	wire _w33891_ ;
	wire _w33890_ ;
	wire _w33889_ ;
	wire _w33888_ ;
	wire _w33887_ ;
	wire _w33886_ ;
	wire _w33885_ ;
	wire _w33884_ ;
	wire _w33883_ ;
	wire _w33882_ ;
	wire _w33881_ ;
	wire _w33880_ ;
	wire _w33879_ ;
	wire _w33878_ ;
	wire _w33877_ ;
	wire _w33876_ ;
	wire _w33875_ ;
	wire _w33874_ ;
	wire _w33873_ ;
	wire _w33872_ ;
	wire _w33871_ ;
	wire _w33870_ ;
	wire _w33869_ ;
	wire _w33868_ ;
	wire _w33867_ ;
	wire _w33866_ ;
	wire _w33865_ ;
	wire _w33864_ ;
	wire _w33863_ ;
	wire _w33862_ ;
	wire _w33861_ ;
	wire _w33860_ ;
	wire _w33859_ ;
	wire _w33858_ ;
	wire _w33857_ ;
	wire _w33856_ ;
	wire _w33855_ ;
	wire _w33854_ ;
	wire _w33853_ ;
	wire _w33852_ ;
	wire _w33851_ ;
	wire _w33850_ ;
	wire _w33849_ ;
	wire _w33848_ ;
	wire _w33847_ ;
	wire _w33846_ ;
	wire _w33845_ ;
	wire _w33844_ ;
	wire _w33843_ ;
	wire _w33842_ ;
	wire _w33841_ ;
	wire _w33840_ ;
	wire _w33839_ ;
	wire _w33838_ ;
	wire _w33837_ ;
	wire _w33836_ ;
	wire _w33835_ ;
	wire _w33834_ ;
	wire _w33833_ ;
	wire _w33832_ ;
	wire _w33831_ ;
	wire _w33830_ ;
	wire _w33829_ ;
	wire _w33828_ ;
	wire _w33827_ ;
	wire _w33826_ ;
	wire _w33825_ ;
	wire _w33824_ ;
	wire _w33823_ ;
	wire _w33822_ ;
	wire _w33821_ ;
	wire _w33820_ ;
	wire _w33819_ ;
	wire _w33818_ ;
	wire _w33817_ ;
	wire _w33816_ ;
	wire _w33815_ ;
	wire _w33814_ ;
	wire _w33813_ ;
	wire _w33812_ ;
	wire _w33811_ ;
	wire _w33810_ ;
	wire _w33809_ ;
	wire _w33808_ ;
	wire _w33807_ ;
	wire _w33806_ ;
	wire _w33805_ ;
	wire _w33804_ ;
	wire _w33803_ ;
	wire _w33802_ ;
	wire _w33801_ ;
	wire _w33800_ ;
	wire _w33799_ ;
	wire _w33798_ ;
	wire _w33797_ ;
	wire _w33796_ ;
	wire _w33795_ ;
	wire _w33794_ ;
	wire _w33793_ ;
	wire _w33792_ ;
	wire _w33791_ ;
	wire _w33790_ ;
	wire _w33789_ ;
	wire _w33788_ ;
	wire _w33787_ ;
	wire _w33786_ ;
	wire _w33785_ ;
	wire _w33784_ ;
	wire _w33783_ ;
	wire _w33782_ ;
	wire _w33781_ ;
	wire _w33780_ ;
	wire _w33779_ ;
	wire _w33778_ ;
	wire _w33777_ ;
	wire _w33776_ ;
	wire _w33775_ ;
	wire _w33774_ ;
	wire _w33773_ ;
	wire _w33772_ ;
	wire _w33771_ ;
	wire _w33770_ ;
	wire _w33769_ ;
	wire _w33768_ ;
	wire _w33767_ ;
	wire _w33766_ ;
	wire _w33765_ ;
	wire _w33764_ ;
	wire _w33763_ ;
	wire _w33762_ ;
	wire _w33761_ ;
	wire _w33760_ ;
	wire _w33759_ ;
	wire _w33758_ ;
	wire _w33757_ ;
	wire _w33756_ ;
	wire _w33755_ ;
	wire _w33754_ ;
	wire _w33753_ ;
	wire _w33752_ ;
	wire _w33751_ ;
	wire _w33750_ ;
	wire _w33749_ ;
	wire _w33748_ ;
	wire _w33747_ ;
	wire _w33746_ ;
	wire _w33745_ ;
	wire _w33744_ ;
	wire _w33743_ ;
	wire _w33742_ ;
	wire _w33741_ ;
	wire _w33740_ ;
	wire _w33739_ ;
	wire _w33738_ ;
	wire _w33737_ ;
	wire _w33736_ ;
	wire _w33735_ ;
	wire _w33734_ ;
	wire _w33733_ ;
	wire _w33732_ ;
	wire _w33731_ ;
	wire _w33730_ ;
	wire _w33729_ ;
	wire _w33728_ ;
	wire _w33727_ ;
	wire _w33726_ ;
	wire _w33725_ ;
	wire _w33724_ ;
	wire _w33723_ ;
	wire _w33722_ ;
	wire _w33721_ ;
	wire _w33720_ ;
	wire _w33719_ ;
	wire _w33718_ ;
	wire _w33717_ ;
	wire _w33716_ ;
	wire _w33715_ ;
	wire _w33714_ ;
	wire _w33713_ ;
	wire _w33712_ ;
	wire _w33711_ ;
	wire _w33710_ ;
	wire _w33709_ ;
	wire _w33708_ ;
	wire _w33707_ ;
	wire _w33706_ ;
	wire _w33705_ ;
	wire _w33704_ ;
	wire _w33703_ ;
	wire _w33702_ ;
	wire _w33701_ ;
	wire _w33700_ ;
	wire _w33699_ ;
	wire _w33698_ ;
	wire _w33697_ ;
	wire _w33696_ ;
	wire _w33695_ ;
	wire _w33694_ ;
	wire _w33693_ ;
	wire _w33692_ ;
	wire _w33691_ ;
	wire _w33690_ ;
	wire _w33689_ ;
	wire _w33688_ ;
	wire _w33687_ ;
	wire _w33686_ ;
	wire _w33685_ ;
	wire _w33684_ ;
	wire _w33683_ ;
	wire _w33682_ ;
	wire _w33681_ ;
	wire _w33680_ ;
	wire _w33679_ ;
	wire _w33678_ ;
	wire _w33677_ ;
	wire _w33676_ ;
	wire _w33675_ ;
	wire _w33674_ ;
	wire _w33673_ ;
	wire _w33672_ ;
	wire _w33671_ ;
	wire _w33670_ ;
	wire _w33669_ ;
	wire _w33668_ ;
	wire _w33667_ ;
	wire _w33666_ ;
	wire _w33665_ ;
	wire _w33664_ ;
	wire _w33663_ ;
	wire _w33662_ ;
	wire _w33661_ ;
	wire _w33660_ ;
	wire _w33659_ ;
	wire _w33658_ ;
	wire _w33657_ ;
	wire _w33656_ ;
	wire _w33655_ ;
	wire _w33654_ ;
	wire _w33653_ ;
	wire _w33652_ ;
	wire _w33651_ ;
	wire _w33650_ ;
	wire _w33649_ ;
	wire _w33648_ ;
	wire _w33647_ ;
	wire _w33646_ ;
	wire _w33645_ ;
	wire _w33644_ ;
	wire _w33643_ ;
	wire _w33642_ ;
	wire _w33641_ ;
	wire _w33640_ ;
	wire _w33639_ ;
	wire _w33638_ ;
	wire _w33637_ ;
	wire _w33636_ ;
	wire _w33635_ ;
	wire _w33634_ ;
	wire _w33633_ ;
	wire _w33632_ ;
	wire _w33631_ ;
	wire _w33630_ ;
	wire _w33629_ ;
	wire _w33628_ ;
	wire _w33627_ ;
	wire _w33626_ ;
	wire _w33625_ ;
	wire _w33624_ ;
	wire _w33623_ ;
	wire _w33622_ ;
	wire _w33621_ ;
	wire _w33620_ ;
	wire _w33619_ ;
	wire _w33618_ ;
	wire _w33617_ ;
	wire _w33616_ ;
	wire _w33615_ ;
	wire _w33614_ ;
	wire _w33613_ ;
	wire _w33612_ ;
	wire _w33611_ ;
	wire _w33610_ ;
	wire _w33609_ ;
	wire _w33608_ ;
	wire _w33607_ ;
	wire _w33606_ ;
	wire _w33605_ ;
	wire _w33604_ ;
	wire _w33603_ ;
	wire _w33602_ ;
	wire _w33601_ ;
	wire _w33600_ ;
	wire _w33599_ ;
	wire _w33598_ ;
	wire _w33597_ ;
	wire _w33596_ ;
	wire _w33595_ ;
	wire _w33594_ ;
	wire _w33593_ ;
	wire _w33592_ ;
	wire _w33591_ ;
	wire _w33590_ ;
	wire _w33589_ ;
	wire _w33588_ ;
	wire _w33587_ ;
	wire _w33586_ ;
	wire _w33585_ ;
	wire _w33584_ ;
	wire _w33583_ ;
	wire _w33582_ ;
	wire _w33581_ ;
	wire _w33580_ ;
	wire _w33579_ ;
	wire _w33578_ ;
	wire _w33577_ ;
	wire _w33576_ ;
	wire _w33575_ ;
	wire _w33574_ ;
	wire _w33573_ ;
	wire _w33572_ ;
	wire _w33571_ ;
	wire _w33570_ ;
	wire _w33569_ ;
	wire _w33568_ ;
	wire _w33567_ ;
	wire _w33566_ ;
	wire _w33565_ ;
	wire _w33564_ ;
	wire _w33563_ ;
	wire _w33562_ ;
	wire _w33561_ ;
	wire _w33560_ ;
	wire _w33559_ ;
	wire _w33558_ ;
	wire _w33557_ ;
	wire _w33556_ ;
	wire _w33555_ ;
	wire _w33554_ ;
	wire _w33553_ ;
	wire _w33552_ ;
	wire _w33551_ ;
	wire _w33550_ ;
	wire _w33549_ ;
	wire _w33548_ ;
	wire _w33547_ ;
	wire _w33546_ ;
	wire _w33545_ ;
	wire _w33544_ ;
	wire _w33543_ ;
	wire _w33542_ ;
	wire _w33541_ ;
	wire _w33540_ ;
	wire _w33539_ ;
	wire _w33538_ ;
	wire _w33537_ ;
	wire _w33536_ ;
	wire _w33535_ ;
	wire _w33534_ ;
	wire _w33533_ ;
	wire _w33532_ ;
	wire _w33531_ ;
	wire _w33530_ ;
	wire _w33529_ ;
	wire _w33528_ ;
	wire _w33527_ ;
	wire _w33526_ ;
	wire _w33525_ ;
	wire _w33524_ ;
	wire _w33523_ ;
	wire _w33522_ ;
	wire _w33521_ ;
	wire _w33520_ ;
	wire _w33519_ ;
	wire _w33518_ ;
	wire _w33517_ ;
	wire _w33516_ ;
	wire _w33515_ ;
	wire _w33514_ ;
	wire _w33513_ ;
	wire _w33512_ ;
	wire _w33511_ ;
	wire _w33510_ ;
	wire _w33509_ ;
	wire _w33508_ ;
	wire _w33507_ ;
	wire _w33506_ ;
	wire _w33505_ ;
	wire _w33504_ ;
	wire _w33503_ ;
	wire _w33502_ ;
	wire _w33501_ ;
	wire _w33500_ ;
	wire _w33499_ ;
	wire _w33498_ ;
	wire _w33497_ ;
	wire _w33496_ ;
	wire _w33495_ ;
	wire _w33494_ ;
	wire _w33493_ ;
	wire _w33492_ ;
	wire _w33491_ ;
	wire _w33490_ ;
	wire _w33489_ ;
	wire _w33488_ ;
	wire _w33487_ ;
	wire _w33486_ ;
	wire _w33485_ ;
	wire _w33484_ ;
	wire _w33483_ ;
	wire _w33482_ ;
	wire _w33481_ ;
	wire _w33480_ ;
	wire _w33479_ ;
	wire _w33478_ ;
	wire _w33477_ ;
	wire _w33476_ ;
	wire _w33475_ ;
	wire _w33474_ ;
	wire _w33473_ ;
	wire _w33472_ ;
	wire _w33471_ ;
	wire _w33470_ ;
	wire _w33469_ ;
	wire _w33468_ ;
	wire _w33467_ ;
	wire _w33466_ ;
	wire _w33465_ ;
	wire _w33464_ ;
	wire _w33463_ ;
	wire _w33462_ ;
	wire _w33461_ ;
	wire _w33460_ ;
	wire _w33459_ ;
	wire _w33458_ ;
	wire _w33457_ ;
	wire _w33456_ ;
	wire _w33455_ ;
	wire _w33454_ ;
	wire _w33453_ ;
	wire _w33452_ ;
	wire _w33451_ ;
	wire _w33450_ ;
	wire _w33449_ ;
	wire _w33448_ ;
	wire _w33447_ ;
	wire _w33446_ ;
	wire _w33445_ ;
	wire _w33444_ ;
	wire _w33443_ ;
	wire _w33442_ ;
	wire _w33441_ ;
	wire _w33440_ ;
	wire _w33439_ ;
	wire _w33438_ ;
	wire _w33437_ ;
	wire _w33436_ ;
	wire _w33435_ ;
	wire _w33434_ ;
	wire _w33433_ ;
	wire _w33432_ ;
	wire _w33431_ ;
	wire _w33430_ ;
	wire _w33429_ ;
	wire _w33428_ ;
	wire _w33427_ ;
	wire _w33426_ ;
	wire _w33425_ ;
	wire _w33424_ ;
	wire _w33423_ ;
	wire _w33422_ ;
	wire _w33421_ ;
	wire _w33420_ ;
	wire _w33419_ ;
	wire _w33418_ ;
	wire _w33417_ ;
	wire _w33416_ ;
	wire _w33415_ ;
	wire _w33414_ ;
	wire _w33413_ ;
	wire _w33412_ ;
	wire _w33411_ ;
	wire _w33410_ ;
	wire _w33409_ ;
	wire _w33408_ ;
	wire _w33407_ ;
	wire _w33406_ ;
	wire _w33405_ ;
	wire _w33404_ ;
	wire _w33403_ ;
	wire _w33402_ ;
	wire _w33401_ ;
	wire _w33400_ ;
	wire _w33399_ ;
	wire _w33398_ ;
	wire _w33397_ ;
	wire _w33396_ ;
	wire _w33395_ ;
	wire _w33394_ ;
	wire _w33393_ ;
	wire _w33392_ ;
	wire _w33391_ ;
	wire _w33390_ ;
	wire _w33389_ ;
	wire _w33388_ ;
	wire _w33387_ ;
	wire _w33386_ ;
	wire _w33385_ ;
	wire _w33384_ ;
	wire _w33383_ ;
	wire _w33382_ ;
	wire _w33381_ ;
	wire _w33380_ ;
	wire _w33379_ ;
	wire _w33378_ ;
	wire _w33377_ ;
	wire _w33376_ ;
	wire _w33375_ ;
	wire _w33374_ ;
	wire _w33373_ ;
	wire _w33372_ ;
	wire _w33371_ ;
	wire _w33370_ ;
	wire _w33369_ ;
	wire _w33368_ ;
	wire _w33367_ ;
	wire _w33366_ ;
	wire _w33365_ ;
	wire _w33364_ ;
	wire _w33363_ ;
	wire _w33362_ ;
	wire _w33361_ ;
	wire _w33360_ ;
	wire _w33359_ ;
	wire _w33358_ ;
	wire _w33357_ ;
	wire _w33356_ ;
	wire _w33355_ ;
	wire _w33354_ ;
	wire _w33353_ ;
	wire _w33352_ ;
	wire _w33351_ ;
	wire _w33350_ ;
	wire _w33349_ ;
	wire _w33348_ ;
	wire _w33347_ ;
	wire _w33346_ ;
	wire _w33345_ ;
	wire _w33344_ ;
	wire _w33343_ ;
	wire _w33342_ ;
	wire _w33341_ ;
	wire _w33340_ ;
	wire _w33339_ ;
	wire _w33338_ ;
	wire _w33337_ ;
	wire _w33336_ ;
	wire _w33335_ ;
	wire _w33334_ ;
	wire _w33333_ ;
	wire _w33332_ ;
	wire _w33331_ ;
	wire _w33330_ ;
	wire _w33329_ ;
	wire _w33328_ ;
	wire _w33327_ ;
	wire _w33326_ ;
	wire _w33325_ ;
	wire _w33324_ ;
	wire _w33323_ ;
	wire _w33322_ ;
	wire _w33321_ ;
	wire _w33320_ ;
	wire _w33319_ ;
	wire _w33318_ ;
	wire _w33317_ ;
	wire _w33316_ ;
	wire _w33315_ ;
	wire _w33314_ ;
	wire _w33313_ ;
	wire _w33312_ ;
	wire _w33311_ ;
	wire _w33310_ ;
	wire _w33309_ ;
	wire _w33308_ ;
	wire _w33307_ ;
	wire _w33306_ ;
	wire _w33305_ ;
	wire _w33304_ ;
	wire _w33303_ ;
	wire _w33302_ ;
	wire _w33301_ ;
	wire _w33300_ ;
	wire _w33299_ ;
	wire _w33298_ ;
	wire _w33297_ ;
	wire _w33296_ ;
	wire _w33295_ ;
	wire _w33294_ ;
	wire _w33293_ ;
	wire _w33292_ ;
	wire _w33291_ ;
	wire _w33290_ ;
	wire _w33289_ ;
	wire _w33288_ ;
	wire _w33287_ ;
	wire _w33286_ ;
	wire _w33285_ ;
	wire _w33284_ ;
	wire _w33283_ ;
	wire _w33282_ ;
	wire _w33281_ ;
	wire _w33280_ ;
	wire _w33279_ ;
	wire _w33278_ ;
	wire _w33277_ ;
	wire _w33276_ ;
	wire _w33275_ ;
	wire _w33274_ ;
	wire _w33273_ ;
	wire _w33272_ ;
	wire _w33271_ ;
	wire _w33270_ ;
	wire _w33269_ ;
	wire _w33268_ ;
	wire _w33267_ ;
	wire _w33266_ ;
	wire _w33265_ ;
	wire _w33264_ ;
	wire _w33263_ ;
	wire _w33262_ ;
	wire _w33261_ ;
	wire _w33260_ ;
	wire _w33259_ ;
	wire _w33258_ ;
	wire _w33257_ ;
	wire _w33256_ ;
	wire _w33255_ ;
	wire _w33254_ ;
	wire _w33253_ ;
	wire _w33252_ ;
	wire _w33251_ ;
	wire _w33250_ ;
	wire _w33249_ ;
	wire _w33248_ ;
	wire _w33247_ ;
	wire _w33246_ ;
	wire _w33245_ ;
	wire _w33244_ ;
	wire _w33243_ ;
	wire _w33242_ ;
	wire _w33241_ ;
	wire _w33240_ ;
	wire _w33239_ ;
	wire _w33238_ ;
	wire _w33237_ ;
	wire _w33236_ ;
	wire _w33235_ ;
	wire _w33234_ ;
	wire _w33233_ ;
	wire _w33232_ ;
	wire _w33231_ ;
	wire _w33230_ ;
	wire _w33229_ ;
	wire _w33228_ ;
	wire _w33227_ ;
	wire _w33226_ ;
	wire _w33225_ ;
	wire _w33224_ ;
	wire _w33223_ ;
	wire _w33222_ ;
	wire _w33221_ ;
	wire _w33220_ ;
	wire _w33219_ ;
	wire _w33218_ ;
	wire _w33217_ ;
	wire _w33216_ ;
	wire _w33215_ ;
	wire _w33214_ ;
	wire _w33213_ ;
	wire _w33212_ ;
	wire _w33211_ ;
	wire _w33210_ ;
	wire _w33209_ ;
	wire _w33208_ ;
	wire _w33207_ ;
	wire _w33206_ ;
	wire _w33205_ ;
	wire _w33204_ ;
	wire _w33203_ ;
	wire _w33202_ ;
	wire _w33201_ ;
	wire _w33200_ ;
	wire _w33199_ ;
	wire _w33198_ ;
	wire _w33197_ ;
	wire _w33196_ ;
	wire _w33195_ ;
	wire _w33194_ ;
	wire _w33193_ ;
	wire _w33192_ ;
	wire _w33191_ ;
	wire _w33190_ ;
	wire _w33189_ ;
	wire _w33188_ ;
	wire _w33187_ ;
	wire _w33186_ ;
	wire _w33185_ ;
	wire _w33184_ ;
	wire _w33183_ ;
	wire _w33182_ ;
	wire _w33181_ ;
	wire _w33180_ ;
	wire _w33179_ ;
	wire _w33178_ ;
	wire _w33177_ ;
	wire _w33176_ ;
	wire _w33175_ ;
	wire _w33174_ ;
	wire _w33173_ ;
	wire _w33172_ ;
	wire _w33171_ ;
	wire _w33170_ ;
	wire _w33169_ ;
	wire _w33168_ ;
	wire _w33167_ ;
	wire _w33166_ ;
	wire _w33165_ ;
	wire _w33164_ ;
	wire _w33163_ ;
	wire _w33162_ ;
	wire _w33161_ ;
	wire _w33160_ ;
	wire _w33159_ ;
	wire _w33158_ ;
	wire _w33157_ ;
	wire _w33156_ ;
	wire _w33155_ ;
	wire _w33154_ ;
	wire _w33153_ ;
	wire _w33152_ ;
	wire _w33151_ ;
	wire _w33150_ ;
	wire _w33149_ ;
	wire _w33148_ ;
	wire _w33147_ ;
	wire _w33146_ ;
	wire _w33145_ ;
	wire _w33144_ ;
	wire _w33143_ ;
	wire _w33142_ ;
	wire _w33141_ ;
	wire _w33140_ ;
	wire _w33139_ ;
	wire _w33138_ ;
	wire _w33137_ ;
	wire _w33136_ ;
	wire _w33135_ ;
	wire _w33134_ ;
	wire _w33133_ ;
	wire _w33132_ ;
	wire _w33131_ ;
	wire _w33130_ ;
	wire _w33129_ ;
	wire _w33128_ ;
	wire _w33127_ ;
	wire _w33126_ ;
	wire _w33125_ ;
	wire _w33124_ ;
	wire _w33123_ ;
	wire _w33122_ ;
	wire _w33121_ ;
	wire _w33120_ ;
	wire _w33119_ ;
	wire _w33118_ ;
	wire _w33117_ ;
	wire _w33116_ ;
	wire _w33115_ ;
	wire _w33114_ ;
	wire _w33113_ ;
	wire _w33112_ ;
	wire _w33111_ ;
	wire _w33110_ ;
	wire _w33109_ ;
	wire _w33108_ ;
	wire _w33107_ ;
	wire _w33106_ ;
	wire _w33105_ ;
	wire _w33104_ ;
	wire _w33103_ ;
	wire _w33102_ ;
	wire _w33101_ ;
	wire _w33100_ ;
	wire _w33099_ ;
	wire _w33098_ ;
	wire _w33097_ ;
	wire _w33096_ ;
	wire _w33095_ ;
	wire _w33094_ ;
	wire _w33093_ ;
	wire _w33092_ ;
	wire _w33091_ ;
	wire _w33090_ ;
	wire _w33089_ ;
	wire _w33088_ ;
	wire _w33087_ ;
	wire _w33086_ ;
	wire _w33085_ ;
	wire _w33084_ ;
	wire _w33083_ ;
	wire _w33082_ ;
	wire _w33081_ ;
	wire _w33080_ ;
	wire _w33079_ ;
	wire _w33078_ ;
	wire _w33077_ ;
	wire _w33076_ ;
	wire _w33075_ ;
	wire _w33074_ ;
	wire _w33073_ ;
	wire _w33072_ ;
	wire _w33071_ ;
	wire _w33070_ ;
	wire _w33069_ ;
	wire _w33068_ ;
	wire _w33067_ ;
	wire _w33066_ ;
	wire _w33065_ ;
	wire _w33064_ ;
	wire _w33063_ ;
	wire _w33062_ ;
	wire _w33061_ ;
	wire _w33060_ ;
	wire _w33059_ ;
	wire _w33058_ ;
	wire _w33057_ ;
	wire _w33056_ ;
	wire _w33055_ ;
	wire _w33054_ ;
	wire _w33053_ ;
	wire _w33052_ ;
	wire _w33051_ ;
	wire _w33050_ ;
	wire _w33049_ ;
	wire _w33048_ ;
	wire _w33047_ ;
	wire _w33046_ ;
	wire _w33045_ ;
	wire _w33044_ ;
	wire _w33043_ ;
	wire _w33042_ ;
	wire _w33041_ ;
	wire _w33040_ ;
	wire _w33039_ ;
	wire _w33038_ ;
	wire _w33037_ ;
	wire _w33036_ ;
	wire _w33035_ ;
	wire _w33034_ ;
	wire _w33033_ ;
	wire _w33032_ ;
	wire _w33031_ ;
	wire _w33030_ ;
	wire _w33029_ ;
	wire _w33028_ ;
	wire _w33027_ ;
	wire _w33026_ ;
	wire _w33025_ ;
	wire _w33024_ ;
	wire _w33023_ ;
	wire _w33022_ ;
	wire _w33021_ ;
	wire _w33020_ ;
	wire _w33019_ ;
	wire _w33018_ ;
	wire _w33017_ ;
	wire _w33016_ ;
	wire _w33015_ ;
	wire _w33014_ ;
	wire _w33013_ ;
	wire _w33012_ ;
	wire _w33011_ ;
	wire _w33010_ ;
	wire _w33009_ ;
	wire _w33008_ ;
	wire _w33007_ ;
	wire _w33006_ ;
	wire _w33005_ ;
	wire _w33004_ ;
	wire _w33003_ ;
	wire _w33002_ ;
	wire _w33001_ ;
	wire _w33000_ ;
	wire _w32999_ ;
	wire _w32998_ ;
	wire _w32997_ ;
	wire _w32996_ ;
	wire _w32995_ ;
	wire _w32994_ ;
	wire _w32993_ ;
	wire _w32992_ ;
	wire _w32991_ ;
	wire _w32990_ ;
	wire _w32989_ ;
	wire _w32988_ ;
	wire _w32987_ ;
	wire _w32986_ ;
	wire _w32985_ ;
	wire _w32984_ ;
	wire _w32983_ ;
	wire _w32982_ ;
	wire _w32981_ ;
	wire _w32980_ ;
	wire _w32979_ ;
	wire _w32978_ ;
	wire _w32977_ ;
	wire _w32976_ ;
	wire _w32975_ ;
	wire _w32974_ ;
	wire _w32973_ ;
	wire _w32972_ ;
	wire _w32971_ ;
	wire _w32970_ ;
	wire _w32969_ ;
	wire _w32968_ ;
	wire _w32967_ ;
	wire _w32966_ ;
	wire _w32965_ ;
	wire _w32964_ ;
	wire _w32963_ ;
	wire _w32962_ ;
	wire _w32961_ ;
	wire _w32960_ ;
	wire _w32959_ ;
	wire _w32958_ ;
	wire _w32957_ ;
	wire _w32956_ ;
	wire _w32955_ ;
	wire _w32954_ ;
	wire _w32953_ ;
	wire _w32952_ ;
	wire _w32951_ ;
	wire _w32950_ ;
	wire _w32949_ ;
	wire _w32948_ ;
	wire _w32947_ ;
	wire _w32946_ ;
	wire _w32945_ ;
	wire _w32944_ ;
	wire _w32943_ ;
	wire _w32942_ ;
	wire _w32941_ ;
	wire _w32940_ ;
	wire _w32939_ ;
	wire _w32938_ ;
	wire _w32937_ ;
	wire _w32936_ ;
	wire _w32935_ ;
	wire _w32934_ ;
	wire _w32933_ ;
	wire _w32932_ ;
	wire _w32931_ ;
	wire _w32930_ ;
	wire _w32929_ ;
	wire _w32928_ ;
	wire _w32927_ ;
	wire _w32926_ ;
	wire _w32925_ ;
	wire _w32924_ ;
	wire _w32923_ ;
	wire _w32922_ ;
	wire _w32921_ ;
	wire _w32920_ ;
	wire _w32919_ ;
	wire _w32918_ ;
	wire _w32917_ ;
	wire _w32916_ ;
	wire _w32915_ ;
	wire _w32914_ ;
	wire _w32913_ ;
	wire _w32912_ ;
	wire _w32911_ ;
	wire _w32910_ ;
	wire _w32909_ ;
	wire _w32908_ ;
	wire _w32907_ ;
	wire _w32906_ ;
	wire _w32905_ ;
	wire _w32904_ ;
	wire _w32903_ ;
	wire _w32902_ ;
	wire _w32901_ ;
	wire _w32900_ ;
	wire _w32899_ ;
	wire _w32898_ ;
	wire _w32897_ ;
	wire _w32896_ ;
	wire _w32895_ ;
	wire _w32894_ ;
	wire _w32893_ ;
	wire _w32892_ ;
	wire _w32891_ ;
	wire _w32890_ ;
	wire _w32889_ ;
	wire _w32888_ ;
	wire _w32887_ ;
	wire _w32886_ ;
	wire _w32885_ ;
	wire _w32884_ ;
	wire _w32883_ ;
	wire _w32882_ ;
	wire _w32881_ ;
	wire _w32880_ ;
	wire _w32879_ ;
	wire _w32878_ ;
	wire _w32877_ ;
	wire _w32876_ ;
	wire _w32875_ ;
	wire _w32874_ ;
	wire _w32873_ ;
	wire _w32872_ ;
	wire _w32871_ ;
	wire _w32870_ ;
	wire _w32869_ ;
	wire _w32868_ ;
	wire _w32867_ ;
	wire _w32866_ ;
	wire _w32865_ ;
	wire _w32864_ ;
	wire _w32863_ ;
	wire _w32862_ ;
	wire _w32861_ ;
	wire _w32860_ ;
	wire _w32859_ ;
	wire _w32858_ ;
	wire _w32857_ ;
	wire _w32856_ ;
	wire _w32855_ ;
	wire _w32854_ ;
	wire _w32853_ ;
	wire _w32852_ ;
	wire _w32851_ ;
	wire _w32850_ ;
	wire _w32849_ ;
	wire _w32848_ ;
	wire _w32847_ ;
	wire _w32846_ ;
	wire _w32845_ ;
	wire _w32844_ ;
	wire _w32843_ ;
	wire _w32842_ ;
	wire _w32841_ ;
	wire _w32840_ ;
	wire _w32839_ ;
	wire _w32838_ ;
	wire _w32837_ ;
	wire _w32836_ ;
	wire _w32835_ ;
	wire _w32834_ ;
	wire _w32833_ ;
	wire _w32832_ ;
	wire _w32831_ ;
	wire _w32830_ ;
	wire _w32829_ ;
	wire _w32828_ ;
	wire _w32827_ ;
	wire _w32826_ ;
	wire _w32825_ ;
	wire _w32824_ ;
	wire _w32823_ ;
	wire _w32822_ ;
	wire _w32821_ ;
	wire _w32820_ ;
	wire _w32819_ ;
	wire _w32818_ ;
	wire _w32817_ ;
	wire _w32816_ ;
	wire _w32815_ ;
	wire _w32814_ ;
	wire _w32813_ ;
	wire _w32812_ ;
	wire _w32811_ ;
	wire _w32810_ ;
	wire _w32809_ ;
	wire _w32808_ ;
	wire _w32807_ ;
	wire _w32806_ ;
	wire _w32805_ ;
	wire _w32804_ ;
	wire _w32803_ ;
	wire _w32802_ ;
	wire _w32801_ ;
	wire _w32800_ ;
	wire _w32799_ ;
	wire _w32798_ ;
	wire _w32797_ ;
	wire _w32796_ ;
	wire _w32795_ ;
	wire _w32794_ ;
	wire _w32793_ ;
	wire _w32792_ ;
	wire _w32791_ ;
	wire _w32790_ ;
	wire _w32789_ ;
	wire _w32788_ ;
	wire _w32787_ ;
	wire _w32786_ ;
	wire _w32785_ ;
	wire _w32784_ ;
	wire _w32783_ ;
	wire _w32782_ ;
	wire _w32781_ ;
	wire _w32780_ ;
	wire _w32779_ ;
	wire _w32778_ ;
	wire _w32777_ ;
	wire _w32776_ ;
	wire _w32775_ ;
	wire _w32774_ ;
	wire _w32773_ ;
	wire _w32772_ ;
	wire _w32771_ ;
	wire _w32770_ ;
	wire _w32769_ ;
	wire _w32768_ ;
	wire _w32767_ ;
	wire _w32766_ ;
	wire _w32765_ ;
	wire _w32764_ ;
	wire _w32763_ ;
	wire _w32762_ ;
	wire _w32761_ ;
	wire _w32760_ ;
	wire _w32759_ ;
	wire _w32758_ ;
	wire _w32757_ ;
	wire _w32756_ ;
	wire _w32755_ ;
	wire _w32754_ ;
	wire _w32753_ ;
	wire _w32752_ ;
	wire _w32751_ ;
	wire _w32750_ ;
	wire _w32749_ ;
	wire _w32748_ ;
	wire _w32747_ ;
	wire _w32746_ ;
	wire _w32745_ ;
	wire _w32744_ ;
	wire _w32743_ ;
	wire _w32742_ ;
	wire _w32741_ ;
	wire _w32740_ ;
	wire _w32739_ ;
	wire _w32738_ ;
	wire _w32737_ ;
	wire _w32736_ ;
	wire _w32735_ ;
	wire _w32734_ ;
	wire _w32733_ ;
	wire _w32732_ ;
	wire _w32731_ ;
	wire _w32730_ ;
	wire _w32729_ ;
	wire _w32728_ ;
	wire _w32727_ ;
	wire _w32726_ ;
	wire _w32725_ ;
	wire _w32724_ ;
	wire _w32723_ ;
	wire _w32722_ ;
	wire _w32721_ ;
	wire _w32720_ ;
	wire _w32719_ ;
	wire _w32718_ ;
	wire _w32717_ ;
	wire _w32716_ ;
	wire _w32715_ ;
	wire _w32714_ ;
	wire _w32713_ ;
	wire _w32712_ ;
	wire _w32711_ ;
	wire _w32710_ ;
	wire _w32709_ ;
	wire _w32708_ ;
	wire _w32707_ ;
	wire _w32706_ ;
	wire _w32705_ ;
	wire _w32704_ ;
	wire _w32703_ ;
	wire _w32702_ ;
	wire _w32701_ ;
	wire _w32700_ ;
	wire _w32699_ ;
	wire _w32698_ ;
	wire _w32697_ ;
	wire _w32696_ ;
	wire _w32695_ ;
	wire _w32694_ ;
	wire _w32693_ ;
	wire _w32692_ ;
	wire _w32691_ ;
	wire _w32690_ ;
	wire _w32689_ ;
	wire _w32688_ ;
	wire _w32687_ ;
	wire _w32686_ ;
	wire _w32685_ ;
	wire _w32684_ ;
	wire _w32683_ ;
	wire _w32682_ ;
	wire _w32681_ ;
	wire _w32680_ ;
	wire _w32679_ ;
	wire _w32678_ ;
	wire _w32677_ ;
	wire _w32676_ ;
	wire _w32675_ ;
	wire _w32674_ ;
	wire _w32673_ ;
	wire _w32672_ ;
	wire _w32671_ ;
	wire _w32670_ ;
	wire _w32669_ ;
	wire _w32668_ ;
	wire _w32667_ ;
	wire _w32666_ ;
	wire _w32665_ ;
	wire _w32664_ ;
	wire _w32663_ ;
	wire _w32662_ ;
	wire _w32661_ ;
	wire _w32660_ ;
	wire _w32659_ ;
	wire _w32658_ ;
	wire _w32657_ ;
	wire _w32656_ ;
	wire _w32655_ ;
	wire _w32654_ ;
	wire _w32653_ ;
	wire _w32652_ ;
	wire _w32651_ ;
	wire _w32650_ ;
	wire _w32649_ ;
	wire _w32648_ ;
	wire _w32647_ ;
	wire _w32646_ ;
	wire _w32645_ ;
	wire _w32644_ ;
	wire _w32643_ ;
	wire _w32642_ ;
	wire _w32641_ ;
	wire _w32640_ ;
	wire _w32639_ ;
	wire _w32638_ ;
	wire _w32637_ ;
	wire _w32636_ ;
	wire _w32635_ ;
	wire _w32634_ ;
	wire _w32633_ ;
	wire _w32632_ ;
	wire _w32631_ ;
	wire _w32630_ ;
	wire _w32629_ ;
	wire _w32628_ ;
	wire _w32627_ ;
	wire _w32626_ ;
	wire _w32625_ ;
	wire _w32624_ ;
	wire _w32623_ ;
	wire _w32622_ ;
	wire _w32621_ ;
	wire _w32620_ ;
	wire _w32619_ ;
	wire _w32618_ ;
	wire _w32617_ ;
	wire _w32616_ ;
	wire _w32615_ ;
	wire _w32614_ ;
	wire _w32613_ ;
	wire _w32612_ ;
	wire _w32611_ ;
	wire _w32610_ ;
	wire _w32609_ ;
	wire _w32608_ ;
	wire _w32607_ ;
	wire _w32606_ ;
	wire _w32605_ ;
	wire _w32604_ ;
	wire _w32603_ ;
	wire _w32602_ ;
	wire _w32601_ ;
	wire _w32600_ ;
	wire _w32599_ ;
	wire _w32598_ ;
	wire _w32597_ ;
	wire _w32596_ ;
	wire _w32595_ ;
	wire _w32594_ ;
	wire _w32593_ ;
	wire _w32592_ ;
	wire _w32591_ ;
	wire _w32590_ ;
	wire _w32589_ ;
	wire _w32588_ ;
	wire _w32587_ ;
	wire _w32586_ ;
	wire _w32585_ ;
	wire _w32584_ ;
	wire _w32583_ ;
	wire _w32582_ ;
	wire _w32581_ ;
	wire _w32580_ ;
	wire _w32579_ ;
	wire _w32578_ ;
	wire _w32577_ ;
	wire _w32576_ ;
	wire _w32575_ ;
	wire _w32574_ ;
	wire _w32573_ ;
	wire _w32572_ ;
	wire _w32571_ ;
	wire _w32570_ ;
	wire _w32569_ ;
	wire _w32568_ ;
	wire _w32567_ ;
	wire _w32566_ ;
	wire _w32565_ ;
	wire _w32564_ ;
	wire _w32563_ ;
	wire _w32562_ ;
	wire _w32561_ ;
	wire _w32560_ ;
	wire _w32559_ ;
	wire _w32558_ ;
	wire _w32557_ ;
	wire _w32556_ ;
	wire _w32555_ ;
	wire _w32554_ ;
	wire _w32553_ ;
	wire _w32552_ ;
	wire _w32551_ ;
	wire _w32550_ ;
	wire _w32549_ ;
	wire _w32548_ ;
	wire _w32547_ ;
	wire _w32546_ ;
	wire _w32545_ ;
	wire _w32544_ ;
	wire _w32543_ ;
	wire _w32542_ ;
	wire _w32541_ ;
	wire _w32540_ ;
	wire _w32539_ ;
	wire _w32538_ ;
	wire _w32537_ ;
	wire _w32536_ ;
	wire _w32535_ ;
	wire _w32534_ ;
	wire _w32533_ ;
	wire _w32532_ ;
	wire _w32531_ ;
	wire _w32530_ ;
	wire _w32529_ ;
	wire _w32528_ ;
	wire _w32527_ ;
	wire _w32526_ ;
	wire _w32525_ ;
	wire _w32524_ ;
	wire _w32523_ ;
	wire _w32522_ ;
	wire _w32521_ ;
	wire _w32520_ ;
	wire _w32519_ ;
	wire _w32518_ ;
	wire _w32517_ ;
	wire _w32516_ ;
	wire _w32515_ ;
	wire _w32514_ ;
	wire _w32513_ ;
	wire _w32512_ ;
	wire _w32511_ ;
	wire _w32510_ ;
	wire _w32509_ ;
	wire _w32508_ ;
	wire _w32507_ ;
	wire _w32506_ ;
	wire _w32505_ ;
	wire _w32504_ ;
	wire _w32503_ ;
	wire _w32502_ ;
	wire _w32501_ ;
	wire _w32500_ ;
	wire _w32499_ ;
	wire _w32498_ ;
	wire _w32497_ ;
	wire _w32496_ ;
	wire _w32495_ ;
	wire _w32494_ ;
	wire _w32493_ ;
	wire _w32492_ ;
	wire _w32491_ ;
	wire _w32490_ ;
	wire _w32489_ ;
	wire _w32488_ ;
	wire _w32487_ ;
	wire _w32486_ ;
	wire _w32485_ ;
	wire _w32484_ ;
	wire _w32483_ ;
	wire _w32482_ ;
	wire _w32481_ ;
	wire _w32480_ ;
	wire _w32479_ ;
	wire _w32478_ ;
	wire _w32477_ ;
	wire _w32476_ ;
	wire _w32475_ ;
	wire _w32474_ ;
	wire _w32473_ ;
	wire _w32472_ ;
	wire _w32471_ ;
	wire _w32470_ ;
	wire _w32469_ ;
	wire _w32468_ ;
	wire _w32467_ ;
	wire _w32466_ ;
	wire _w32465_ ;
	wire _w32464_ ;
	wire _w32463_ ;
	wire _w32462_ ;
	wire _w32461_ ;
	wire _w32460_ ;
	wire _w32459_ ;
	wire _w32458_ ;
	wire _w32457_ ;
	wire _w32456_ ;
	wire _w32455_ ;
	wire _w32454_ ;
	wire _w32453_ ;
	wire _w32452_ ;
	wire _w32451_ ;
	wire _w32450_ ;
	wire _w32449_ ;
	wire _w32448_ ;
	wire _w32447_ ;
	wire _w32446_ ;
	wire _w32445_ ;
	wire _w32444_ ;
	wire _w32443_ ;
	wire _w32442_ ;
	wire _w32441_ ;
	wire _w32440_ ;
	wire _w32439_ ;
	wire _w32438_ ;
	wire _w32437_ ;
	wire _w32436_ ;
	wire _w32435_ ;
	wire _w32434_ ;
	wire _w32433_ ;
	wire _w32432_ ;
	wire _w32431_ ;
	wire _w32430_ ;
	wire _w32429_ ;
	wire _w32428_ ;
	wire _w32427_ ;
	wire _w32426_ ;
	wire _w32425_ ;
	wire _w32424_ ;
	wire _w32423_ ;
	wire _w32422_ ;
	wire _w32421_ ;
	wire _w32420_ ;
	wire _w32419_ ;
	wire _w32418_ ;
	wire _w32417_ ;
	wire _w32416_ ;
	wire _w32415_ ;
	wire _w32414_ ;
	wire _w32413_ ;
	wire _w32412_ ;
	wire _w32411_ ;
	wire _w32410_ ;
	wire _w32409_ ;
	wire _w32408_ ;
	wire _w32407_ ;
	wire _w32406_ ;
	wire _w32405_ ;
	wire _w32404_ ;
	wire _w32403_ ;
	wire _w32402_ ;
	wire _w32401_ ;
	wire _w32400_ ;
	wire _w32399_ ;
	wire _w32398_ ;
	wire _w32397_ ;
	wire _w32396_ ;
	wire _w32395_ ;
	wire _w32394_ ;
	wire _w32393_ ;
	wire _w32392_ ;
	wire _w32391_ ;
	wire _w32390_ ;
	wire _w32389_ ;
	wire _w32388_ ;
	wire _w32387_ ;
	wire _w32386_ ;
	wire _w32385_ ;
	wire _w32384_ ;
	wire _w32383_ ;
	wire _w32382_ ;
	wire _w32381_ ;
	wire _w32380_ ;
	wire _w32379_ ;
	wire _w32378_ ;
	wire _w32377_ ;
	wire _w32376_ ;
	wire _w32375_ ;
	wire _w32374_ ;
	wire _w32373_ ;
	wire _w32372_ ;
	wire _w32371_ ;
	wire _w32370_ ;
	wire _w32369_ ;
	wire _w32368_ ;
	wire _w32367_ ;
	wire _w32366_ ;
	wire _w32365_ ;
	wire _w32364_ ;
	wire _w32363_ ;
	wire _w32362_ ;
	wire _w32361_ ;
	wire _w32360_ ;
	wire _w32359_ ;
	wire _w32358_ ;
	wire _w32357_ ;
	wire _w32356_ ;
	wire _w32355_ ;
	wire _w32354_ ;
	wire _w32353_ ;
	wire _w32352_ ;
	wire _w32351_ ;
	wire _w32350_ ;
	wire _w32349_ ;
	wire _w32348_ ;
	wire _w32347_ ;
	wire _w32346_ ;
	wire _w32345_ ;
	wire _w32344_ ;
	wire _w32343_ ;
	wire _w32342_ ;
	wire _w32341_ ;
	wire _w32340_ ;
	wire _w32339_ ;
	wire _w32338_ ;
	wire _w32337_ ;
	wire _w32336_ ;
	wire _w32335_ ;
	wire _w32334_ ;
	wire _w32333_ ;
	wire _w32332_ ;
	wire _w32331_ ;
	wire _w32330_ ;
	wire _w32329_ ;
	wire _w32328_ ;
	wire _w32327_ ;
	wire _w32326_ ;
	wire _w32325_ ;
	wire _w32324_ ;
	wire _w32323_ ;
	wire _w32322_ ;
	wire _w32321_ ;
	wire _w32320_ ;
	wire _w32319_ ;
	wire _w32318_ ;
	wire _w32317_ ;
	wire _w32316_ ;
	wire _w32315_ ;
	wire _w32314_ ;
	wire _w32313_ ;
	wire _w32312_ ;
	wire _w32311_ ;
	wire _w32310_ ;
	wire _w32309_ ;
	wire _w32308_ ;
	wire _w32307_ ;
	wire _w32306_ ;
	wire _w32305_ ;
	wire _w32304_ ;
	wire _w32303_ ;
	wire _w32302_ ;
	wire _w32301_ ;
	wire _w32300_ ;
	wire _w32299_ ;
	wire _w32298_ ;
	wire _w32297_ ;
	wire _w32296_ ;
	wire _w32295_ ;
	wire _w32294_ ;
	wire _w32293_ ;
	wire _w32292_ ;
	wire _w32291_ ;
	wire _w32290_ ;
	wire _w32289_ ;
	wire _w32288_ ;
	wire _w32287_ ;
	wire _w32286_ ;
	wire _w32285_ ;
	wire _w32284_ ;
	wire _w32283_ ;
	wire _w32282_ ;
	wire _w32281_ ;
	wire _w32280_ ;
	wire _w32279_ ;
	wire _w32278_ ;
	wire _w32277_ ;
	wire _w32276_ ;
	wire _w32275_ ;
	wire _w32274_ ;
	wire _w32273_ ;
	wire _w32272_ ;
	wire _w32271_ ;
	wire _w32270_ ;
	wire _w32269_ ;
	wire _w32268_ ;
	wire _w32267_ ;
	wire _w32266_ ;
	wire _w32265_ ;
	wire _w32264_ ;
	wire _w32263_ ;
	wire _w32262_ ;
	wire _w32261_ ;
	wire _w32260_ ;
	wire _w32259_ ;
	wire _w32258_ ;
	wire _w32257_ ;
	wire _w32256_ ;
	wire _w32255_ ;
	wire _w32254_ ;
	wire _w32253_ ;
	wire _w32252_ ;
	wire _w32251_ ;
	wire _w32250_ ;
	wire _w32249_ ;
	wire _w32248_ ;
	wire _w32247_ ;
	wire _w32246_ ;
	wire _w32245_ ;
	wire _w32244_ ;
	wire _w32243_ ;
	wire _w32242_ ;
	wire _w32241_ ;
	wire _w32240_ ;
	wire _w32239_ ;
	wire _w32238_ ;
	wire _w32237_ ;
	wire _w32236_ ;
	wire _w32235_ ;
	wire _w32234_ ;
	wire _w32233_ ;
	wire _w32232_ ;
	wire _w32231_ ;
	wire _w32230_ ;
	wire _w32229_ ;
	wire _w32228_ ;
	wire _w32227_ ;
	wire _w32226_ ;
	wire _w32225_ ;
	wire _w32224_ ;
	wire _w32223_ ;
	wire _w32222_ ;
	wire _w32221_ ;
	wire _w32220_ ;
	wire _w32219_ ;
	wire _w32218_ ;
	wire _w32217_ ;
	wire _w32216_ ;
	wire _w32215_ ;
	wire _w32214_ ;
	wire _w32213_ ;
	wire _w32212_ ;
	wire _w32211_ ;
	wire _w32210_ ;
	wire _w32209_ ;
	wire _w32208_ ;
	wire _w32207_ ;
	wire _w32206_ ;
	wire _w32205_ ;
	wire _w32204_ ;
	wire _w32203_ ;
	wire _w32202_ ;
	wire _w32201_ ;
	wire _w32200_ ;
	wire _w32199_ ;
	wire _w32198_ ;
	wire _w32197_ ;
	wire _w32196_ ;
	wire _w32195_ ;
	wire _w32194_ ;
	wire _w32193_ ;
	wire _w32192_ ;
	wire _w32191_ ;
	wire _w32190_ ;
	wire _w32189_ ;
	wire _w32188_ ;
	wire _w32187_ ;
	wire _w32186_ ;
	wire _w32185_ ;
	wire _w32184_ ;
	wire _w32183_ ;
	wire _w32182_ ;
	wire _w32181_ ;
	wire _w32180_ ;
	wire _w32179_ ;
	wire _w32178_ ;
	wire _w32177_ ;
	wire _w32176_ ;
	wire _w32175_ ;
	wire _w32174_ ;
	wire _w32173_ ;
	wire _w32172_ ;
	wire _w32171_ ;
	wire _w32170_ ;
	wire _w32169_ ;
	wire _w32168_ ;
	wire _w32167_ ;
	wire _w32166_ ;
	wire _w32165_ ;
	wire _w32164_ ;
	wire _w32163_ ;
	wire _w32162_ ;
	wire _w32161_ ;
	wire _w32160_ ;
	wire _w32159_ ;
	wire _w32158_ ;
	wire _w32157_ ;
	wire _w32156_ ;
	wire _w32155_ ;
	wire _w32154_ ;
	wire _w32153_ ;
	wire _w32152_ ;
	wire _w32151_ ;
	wire _w32150_ ;
	wire _w32149_ ;
	wire _w32148_ ;
	wire _w32147_ ;
	wire _w32146_ ;
	wire _w32145_ ;
	wire _w32144_ ;
	wire _w32143_ ;
	wire _w32142_ ;
	wire _w32141_ ;
	wire _w32140_ ;
	wire _w32139_ ;
	wire _w32138_ ;
	wire _w32137_ ;
	wire _w32136_ ;
	wire _w32135_ ;
	wire _w32134_ ;
	wire _w32133_ ;
	wire _w32132_ ;
	wire _w32131_ ;
	wire _w32130_ ;
	wire _w32129_ ;
	wire _w32128_ ;
	wire _w32127_ ;
	wire _w32126_ ;
	wire _w32125_ ;
	wire _w32124_ ;
	wire _w32123_ ;
	wire _w32122_ ;
	wire _w32121_ ;
	wire _w32120_ ;
	wire _w32119_ ;
	wire _w32118_ ;
	wire _w32117_ ;
	wire _w32116_ ;
	wire _w32115_ ;
	wire _w32114_ ;
	wire _w32113_ ;
	wire _w32112_ ;
	wire _w32111_ ;
	wire _w32110_ ;
	wire _w32109_ ;
	wire _w32108_ ;
	wire _w32107_ ;
	wire _w32106_ ;
	wire _w32105_ ;
	wire _w32104_ ;
	wire _w32103_ ;
	wire _w32102_ ;
	wire _w32101_ ;
	wire _w32100_ ;
	wire _w32099_ ;
	wire _w32098_ ;
	wire _w32097_ ;
	wire _w32096_ ;
	wire _w32095_ ;
	wire _w32094_ ;
	wire _w32093_ ;
	wire _w32092_ ;
	wire _w32091_ ;
	wire _w32090_ ;
	wire _w32089_ ;
	wire _w32088_ ;
	wire _w32087_ ;
	wire _w32086_ ;
	wire _w32085_ ;
	wire _w32084_ ;
	wire _w32083_ ;
	wire _w32082_ ;
	wire _w32081_ ;
	wire _w32080_ ;
	wire _w32079_ ;
	wire _w32078_ ;
	wire _w32077_ ;
	wire _w32076_ ;
	wire _w32075_ ;
	wire _w32074_ ;
	wire _w32073_ ;
	wire _w32072_ ;
	wire _w32071_ ;
	wire _w32070_ ;
	wire _w32069_ ;
	wire _w32068_ ;
	wire _w32067_ ;
	wire _w32066_ ;
	wire _w32065_ ;
	wire _w32064_ ;
	wire _w32063_ ;
	wire _w32062_ ;
	wire _w32061_ ;
	wire _w32060_ ;
	wire _w32059_ ;
	wire _w32058_ ;
	wire _w32057_ ;
	wire _w32056_ ;
	wire _w32055_ ;
	wire _w32054_ ;
	wire _w32053_ ;
	wire _w32052_ ;
	wire _w32051_ ;
	wire _w32050_ ;
	wire _w32049_ ;
	wire _w32048_ ;
	wire _w32047_ ;
	wire _w32046_ ;
	wire _w32045_ ;
	wire _w32044_ ;
	wire _w32043_ ;
	wire _w32042_ ;
	wire _w32041_ ;
	wire _w32040_ ;
	wire _w32039_ ;
	wire _w32038_ ;
	wire _w32037_ ;
	wire _w32036_ ;
	wire _w32035_ ;
	wire _w32034_ ;
	wire _w32033_ ;
	wire _w32032_ ;
	wire _w32031_ ;
	wire _w32030_ ;
	wire _w32029_ ;
	wire _w32028_ ;
	wire _w32027_ ;
	wire _w32026_ ;
	wire _w32025_ ;
	wire _w32024_ ;
	wire _w32023_ ;
	wire _w32022_ ;
	wire _w32021_ ;
	wire _w32020_ ;
	wire _w32019_ ;
	wire _w32018_ ;
	wire _w32017_ ;
	wire _w32016_ ;
	wire _w32015_ ;
	wire _w32014_ ;
	wire _w32013_ ;
	wire _w32012_ ;
	wire _w32011_ ;
	wire _w32010_ ;
	wire _w32009_ ;
	wire _w32008_ ;
	wire _w32007_ ;
	wire _w32006_ ;
	wire _w32005_ ;
	wire _w32004_ ;
	wire _w32003_ ;
	wire _w32002_ ;
	wire _w32001_ ;
	wire _w32000_ ;
	wire _w31999_ ;
	wire _w31998_ ;
	wire _w31997_ ;
	wire _w31996_ ;
	wire _w31995_ ;
	wire _w31994_ ;
	wire _w31993_ ;
	wire _w31992_ ;
	wire _w31991_ ;
	wire _w31990_ ;
	wire _w31989_ ;
	wire _w31988_ ;
	wire _w31987_ ;
	wire _w31986_ ;
	wire _w31985_ ;
	wire _w31984_ ;
	wire _w31983_ ;
	wire _w31982_ ;
	wire _w31981_ ;
	wire _w31980_ ;
	wire _w31979_ ;
	wire _w31978_ ;
	wire _w31977_ ;
	wire _w31976_ ;
	wire _w31975_ ;
	wire _w31974_ ;
	wire _w31973_ ;
	wire _w31972_ ;
	wire _w31971_ ;
	wire _w31970_ ;
	wire _w31969_ ;
	wire _w31968_ ;
	wire _w31967_ ;
	wire _w31966_ ;
	wire _w31965_ ;
	wire _w31964_ ;
	wire _w31963_ ;
	wire _w31962_ ;
	wire _w31961_ ;
	wire _w31960_ ;
	wire _w31959_ ;
	wire _w31958_ ;
	wire _w31957_ ;
	wire _w31956_ ;
	wire _w31955_ ;
	wire _w31954_ ;
	wire _w31953_ ;
	wire _w31952_ ;
	wire _w31951_ ;
	wire _w31950_ ;
	wire _w31949_ ;
	wire _w31948_ ;
	wire _w31947_ ;
	wire _w31946_ ;
	wire _w31945_ ;
	wire _w31944_ ;
	wire _w31943_ ;
	wire _w31942_ ;
	wire _w31941_ ;
	wire _w31940_ ;
	wire _w31939_ ;
	wire _w31938_ ;
	wire _w31937_ ;
	wire _w31936_ ;
	wire _w31935_ ;
	wire _w31934_ ;
	wire _w31933_ ;
	wire _w31932_ ;
	wire _w31931_ ;
	wire _w31930_ ;
	wire _w31929_ ;
	wire _w31928_ ;
	wire _w31927_ ;
	wire _w31926_ ;
	wire _w31925_ ;
	wire _w31924_ ;
	wire _w31923_ ;
	wire _w31922_ ;
	wire _w31921_ ;
	wire _w31920_ ;
	wire _w31919_ ;
	wire _w31918_ ;
	wire _w31917_ ;
	wire _w31916_ ;
	wire _w31915_ ;
	wire _w31914_ ;
	wire _w31913_ ;
	wire _w31912_ ;
	wire _w31911_ ;
	wire _w31910_ ;
	wire _w31909_ ;
	wire _w31908_ ;
	wire _w31907_ ;
	wire _w31906_ ;
	wire _w31905_ ;
	wire _w31904_ ;
	wire _w31903_ ;
	wire _w31902_ ;
	wire _w31901_ ;
	wire _w31900_ ;
	wire _w31899_ ;
	wire _w31898_ ;
	wire _w31897_ ;
	wire _w31896_ ;
	wire _w31895_ ;
	wire _w31894_ ;
	wire _w31893_ ;
	wire _w31892_ ;
	wire _w31891_ ;
	wire _w31890_ ;
	wire _w31889_ ;
	wire _w31888_ ;
	wire _w31887_ ;
	wire _w31886_ ;
	wire _w31885_ ;
	wire _w31884_ ;
	wire _w31883_ ;
	wire _w31882_ ;
	wire _w31881_ ;
	wire _w31880_ ;
	wire _w31879_ ;
	wire _w31878_ ;
	wire _w31877_ ;
	wire _w31876_ ;
	wire _w31875_ ;
	wire _w31874_ ;
	wire _w31873_ ;
	wire _w31872_ ;
	wire _w31871_ ;
	wire _w31870_ ;
	wire _w31869_ ;
	wire _w31868_ ;
	wire _w31867_ ;
	wire _w31866_ ;
	wire _w31865_ ;
	wire _w31864_ ;
	wire _w31863_ ;
	wire _w31862_ ;
	wire _w31861_ ;
	wire _w31860_ ;
	wire _w31859_ ;
	wire _w31858_ ;
	wire _w31857_ ;
	wire _w31856_ ;
	wire _w31855_ ;
	wire _w31854_ ;
	wire _w31853_ ;
	wire _w31852_ ;
	wire _w31851_ ;
	wire _w31850_ ;
	wire _w31849_ ;
	wire _w31848_ ;
	wire _w31847_ ;
	wire _w31846_ ;
	wire _w31845_ ;
	wire _w31844_ ;
	wire _w31843_ ;
	wire _w31842_ ;
	wire _w31841_ ;
	wire _w31840_ ;
	wire _w31839_ ;
	wire _w31838_ ;
	wire _w31837_ ;
	wire _w31836_ ;
	wire _w31835_ ;
	wire _w31834_ ;
	wire _w31833_ ;
	wire _w31832_ ;
	wire _w31831_ ;
	wire _w31830_ ;
	wire _w31829_ ;
	wire _w31828_ ;
	wire _w31827_ ;
	wire _w31826_ ;
	wire _w31825_ ;
	wire _w31824_ ;
	wire _w31823_ ;
	wire _w31822_ ;
	wire _w31821_ ;
	wire _w31820_ ;
	wire _w31819_ ;
	wire _w31818_ ;
	wire _w31817_ ;
	wire _w31816_ ;
	wire _w31815_ ;
	wire _w31814_ ;
	wire _w31813_ ;
	wire _w31812_ ;
	wire _w31811_ ;
	wire _w31810_ ;
	wire _w31809_ ;
	wire _w31808_ ;
	wire _w31807_ ;
	wire _w31806_ ;
	wire _w31805_ ;
	wire _w31804_ ;
	wire _w31803_ ;
	wire _w31802_ ;
	wire _w31801_ ;
	wire _w31800_ ;
	wire _w31799_ ;
	wire _w31798_ ;
	wire _w31797_ ;
	wire _w31796_ ;
	wire _w31795_ ;
	wire _w31794_ ;
	wire _w31793_ ;
	wire _w31792_ ;
	wire _w31791_ ;
	wire _w31790_ ;
	wire _w31789_ ;
	wire _w31788_ ;
	wire _w31787_ ;
	wire _w31786_ ;
	wire _w31785_ ;
	wire _w31784_ ;
	wire _w31783_ ;
	wire _w31782_ ;
	wire _w31781_ ;
	wire _w31780_ ;
	wire _w31779_ ;
	wire _w31778_ ;
	wire _w31777_ ;
	wire _w31776_ ;
	wire _w31775_ ;
	wire _w31774_ ;
	wire _w31773_ ;
	wire _w31772_ ;
	wire _w31771_ ;
	wire _w31770_ ;
	wire _w31769_ ;
	wire _w31768_ ;
	wire _w31767_ ;
	wire _w31766_ ;
	wire _w31765_ ;
	wire _w31764_ ;
	wire _w31763_ ;
	wire _w31762_ ;
	wire _w31761_ ;
	wire _w31760_ ;
	wire _w31759_ ;
	wire _w31758_ ;
	wire _w31757_ ;
	wire _w31756_ ;
	wire _w31755_ ;
	wire _w31754_ ;
	wire _w31753_ ;
	wire _w31752_ ;
	wire _w31751_ ;
	wire _w31750_ ;
	wire _w31749_ ;
	wire _w31748_ ;
	wire _w31747_ ;
	wire _w31746_ ;
	wire _w31745_ ;
	wire _w31744_ ;
	wire _w31743_ ;
	wire _w31742_ ;
	wire _w31741_ ;
	wire _w31740_ ;
	wire _w31739_ ;
	wire _w31738_ ;
	wire _w31737_ ;
	wire _w31736_ ;
	wire _w31735_ ;
	wire _w31734_ ;
	wire _w31733_ ;
	wire _w31732_ ;
	wire _w31731_ ;
	wire _w31730_ ;
	wire _w31729_ ;
	wire _w31728_ ;
	wire _w31727_ ;
	wire _w31726_ ;
	wire _w31725_ ;
	wire _w31724_ ;
	wire _w31723_ ;
	wire _w31722_ ;
	wire _w31721_ ;
	wire _w31720_ ;
	wire _w31719_ ;
	wire _w31718_ ;
	wire _w31717_ ;
	wire _w31716_ ;
	wire _w31715_ ;
	wire _w31714_ ;
	wire _w31713_ ;
	wire _w31712_ ;
	wire _w31711_ ;
	wire _w31710_ ;
	wire _w31709_ ;
	wire _w31708_ ;
	wire _w31707_ ;
	wire _w31706_ ;
	wire _w31705_ ;
	wire _w31704_ ;
	wire _w31703_ ;
	wire _w31702_ ;
	wire _w31701_ ;
	wire _w31700_ ;
	wire _w31699_ ;
	wire _w31698_ ;
	wire _w31697_ ;
	wire _w31696_ ;
	wire _w31695_ ;
	wire _w31694_ ;
	wire _w31693_ ;
	wire _w31692_ ;
	wire _w31691_ ;
	wire _w31690_ ;
	wire _w31689_ ;
	wire _w31688_ ;
	wire _w31687_ ;
	wire _w31686_ ;
	wire _w31685_ ;
	wire _w31684_ ;
	wire _w31683_ ;
	wire _w31682_ ;
	wire _w31681_ ;
	wire _w31680_ ;
	wire _w31679_ ;
	wire _w31678_ ;
	wire _w31677_ ;
	wire _w31676_ ;
	wire _w31675_ ;
	wire _w31674_ ;
	wire _w31673_ ;
	wire _w31672_ ;
	wire _w31671_ ;
	wire _w31670_ ;
	wire _w31669_ ;
	wire _w31668_ ;
	wire _w31667_ ;
	wire _w31666_ ;
	wire _w31665_ ;
	wire _w31664_ ;
	wire _w31663_ ;
	wire _w31662_ ;
	wire _w31661_ ;
	wire _w31660_ ;
	wire _w31659_ ;
	wire _w31658_ ;
	wire _w31657_ ;
	wire _w31656_ ;
	wire _w31655_ ;
	wire _w31654_ ;
	wire _w31653_ ;
	wire _w31652_ ;
	wire _w31651_ ;
	wire _w31650_ ;
	wire _w31649_ ;
	wire _w31648_ ;
	wire _w31647_ ;
	wire _w31646_ ;
	wire _w31645_ ;
	wire _w31644_ ;
	wire _w31643_ ;
	wire _w31642_ ;
	wire _w31641_ ;
	wire _w31640_ ;
	wire _w31639_ ;
	wire _w31638_ ;
	wire _w31637_ ;
	wire _w31636_ ;
	wire _w31635_ ;
	wire _w31634_ ;
	wire _w31633_ ;
	wire _w31632_ ;
	wire _w31631_ ;
	wire _w31630_ ;
	wire _w31629_ ;
	wire _w31628_ ;
	wire _w31627_ ;
	wire _w31626_ ;
	wire _w31625_ ;
	wire _w31624_ ;
	wire _w31623_ ;
	wire _w31622_ ;
	wire _w31621_ ;
	wire _w31620_ ;
	wire _w31619_ ;
	wire _w31618_ ;
	wire _w31617_ ;
	wire _w31616_ ;
	wire _w31615_ ;
	wire _w31614_ ;
	wire _w31613_ ;
	wire _w31612_ ;
	wire _w31611_ ;
	wire _w31610_ ;
	wire _w31609_ ;
	wire _w31608_ ;
	wire _w31607_ ;
	wire _w31606_ ;
	wire _w31605_ ;
	wire _w31604_ ;
	wire _w31603_ ;
	wire _w31602_ ;
	wire _w31601_ ;
	wire _w31600_ ;
	wire _w31599_ ;
	wire _w31598_ ;
	wire _w31597_ ;
	wire _w31596_ ;
	wire _w31595_ ;
	wire _w31594_ ;
	wire _w31593_ ;
	wire _w31592_ ;
	wire _w31591_ ;
	wire _w31590_ ;
	wire _w31589_ ;
	wire _w31588_ ;
	wire _w31587_ ;
	wire _w31586_ ;
	wire _w31585_ ;
	wire _w31584_ ;
	wire _w31583_ ;
	wire _w31582_ ;
	wire _w31581_ ;
	wire _w31580_ ;
	wire _w31579_ ;
	wire _w31578_ ;
	wire _w31577_ ;
	wire _w31576_ ;
	wire _w31575_ ;
	wire _w31574_ ;
	wire _w31573_ ;
	wire _w31572_ ;
	wire _w31571_ ;
	wire _w31570_ ;
	wire _w31569_ ;
	wire _w31568_ ;
	wire _w31567_ ;
	wire _w31566_ ;
	wire _w31565_ ;
	wire _w31564_ ;
	wire _w31563_ ;
	wire _w31562_ ;
	wire _w31561_ ;
	wire _w31560_ ;
	wire _w31559_ ;
	wire _w31558_ ;
	wire _w31557_ ;
	wire _w31556_ ;
	wire _w31555_ ;
	wire _w31554_ ;
	wire _w31553_ ;
	wire _w31552_ ;
	wire _w31551_ ;
	wire _w31550_ ;
	wire _w31549_ ;
	wire _w31548_ ;
	wire _w31547_ ;
	wire _w31546_ ;
	wire _w31545_ ;
	wire _w31544_ ;
	wire _w31543_ ;
	wire _w31542_ ;
	wire _w31541_ ;
	wire _w31540_ ;
	wire _w31539_ ;
	wire _w31538_ ;
	wire _w31537_ ;
	wire _w31536_ ;
	wire _w31535_ ;
	wire _w31534_ ;
	wire _w31533_ ;
	wire _w31532_ ;
	wire _w31531_ ;
	wire _w31530_ ;
	wire _w31529_ ;
	wire _w31528_ ;
	wire _w31527_ ;
	wire _w31526_ ;
	wire _w31525_ ;
	wire _w31524_ ;
	wire _w31523_ ;
	wire _w31522_ ;
	wire _w31521_ ;
	wire _w31520_ ;
	wire _w31519_ ;
	wire _w31518_ ;
	wire _w31517_ ;
	wire _w31516_ ;
	wire _w31515_ ;
	wire _w31514_ ;
	wire _w31513_ ;
	wire _w31512_ ;
	wire _w31511_ ;
	wire _w31510_ ;
	wire _w31509_ ;
	wire _w31508_ ;
	wire _w31507_ ;
	wire _w31506_ ;
	wire _w31505_ ;
	wire _w31504_ ;
	wire _w31503_ ;
	wire _w31502_ ;
	wire _w31501_ ;
	wire _w31500_ ;
	wire _w31499_ ;
	wire _w31498_ ;
	wire _w31497_ ;
	wire _w31496_ ;
	wire _w31495_ ;
	wire _w31494_ ;
	wire _w31493_ ;
	wire _w31492_ ;
	wire _w31491_ ;
	wire _w31490_ ;
	wire _w31489_ ;
	wire _w31488_ ;
	wire _w31487_ ;
	wire _w31486_ ;
	wire _w31485_ ;
	wire _w31484_ ;
	wire _w31483_ ;
	wire _w31482_ ;
	wire _w31481_ ;
	wire _w31480_ ;
	wire _w31479_ ;
	wire _w31478_ ;
	wire _w31477_ ;
	wire _w31476_ ;
	wire _w31475_ ;
	wire _w31474_ ;
	wire _w31473_ ;
	wire _w31472_ ;
	wire _w31471_ ;
	wire _w31470_ ;
	wire _w31469_ ;
	wire _w31468_ ;
	wire _w31467_ ;
	wire _w31466_ ;
	wire _w31465_ ;
	wire _w31464_ ;
	wire _w31463_ ;
	wire _w31462_ ;
	wire _w31461_ ;
	wire _w31460_ ;
	wire _w31459_ ;
	wire _w31458_ ;
	wire _w31457_ ;
	wire _w31456_ ;
	wire _w31455_ ;
	wire _w31454_ ;
	wire _w31453_ ;
	wire _w31452_ ;
	wire _w31451_ ;
	wire _w31450_ ;
	wire _w31449_ ;
	wire _w31448_ ;
	wire _w31447_ ;
	wire _w31446_ ;
	wire _w31445_ ;
	wire _w31444_ ;
	wire _w31443_ ;
	wire _w31442_ ;
	wire _w31441_ ;
	wire _w31440_ ;
	wire _w31439_ ;
	wire _w31438_ ;
	wire _w31437_ ;
	wire _w31436_ ;
	wire _w31435_ ;
	wire _w31434_ ;
	wire _w31433_ ;
	wire _w31432_ ;
	wire _w31431_ ;
	wire _w31430_ ;
	wire _w31429_ ;
	wire _w31428_ ;
	wire _w31427_ ;
	wire _w31426_ ;
	wire _w31425_ ;
	wire _w31424_ ;
	wire _w31423_ ;
	wire _w31422_ ;
	wire _w31421_ ;
	wire _w31420_ ;
	wire _w31419_ ;
	wire _w31418_ ;
	wire _w31417_ ;
	wire _w31416_ ;
	wire _w31415_ ;
	wire _w31414_ ;
	wire _w31413_ ;
	wire _w31412_ ;
	wire _w31411_ ;
	wire _w31410_ ;
	wire _w31409_ ;
	wire _w31408_ ;
	wire _w31407_ ;
	wire _w31406_ ;
	wire _w31405_ ;
	wire _w31404_ ;
	wire _w31403_ ;
	wire _w31402_ ;
	wire _w31401_ ;
	wire _w31400_ ;
	wire _w31399_ ;
	wire _w31398_ ;
	wire _w31397_ ;
	wire _w31396_ ;
	wire _w31395_ ;
	wire _w31394_ ;
	wire _w31393_ ;
	wire _w31392_ ;
	wire _w31391_ ;
	wire _w31390_ ;
	wire _w31389_ ;
	wire _w31388_ ;
	wire _w31387_ ;
	wire _w31386_ ;
	wire _w31385_ ;
	wire _w31384_ ;
	wire _w31383_ ;
	wire _w31382_ ;
	wire _w31381_ ;
	wire _w31380_ ;
	wire _w31379_ ;
	wire _w31378_ ;
	wire _w31377_ ;
	wire _w31376_ ;
	wire _w31375_ ;
	wire _w31374_ ;
	wire _w31373_ ;
	wire _w31372_ ;
	wire _w31371_ ;
	wire _w31370_ ;
	wire _w31369_ ;
	wire _w31368_ ;
	wire _w31367_ ;
	wire _w31366_ ;
	wire _w31365_ ;
	wire _w31364_ ;
	wire _w31363_ ;
	wire _w31362_ ;
	wire _w31361_ ;
	wire _w31360_ ;
	wire _w31359_ ;
	wire _w31358_ ;
	wire _w31357_ ;
	wire _w31356_ ;
	wire _w31355_ ;
	wire _w31354_ ;
	wire _w31353_ ;
	wire _w31352_ ;
	wire _w31351_ ;
	wire _w31350_ ;
	wire _w31349_ ;
	wire _w31348_ ;
	wire _w31347_ ;
	wire _w31346_ ;
	wire _w31345_ ;
	wire _w31344_ ;
	wire _w31343_ ;
	wire _w31342_ ;
	wire _w31341_ ;
	wire _w31340_ ;
	wire _w31339_ ;
	wire _w31338_ ;
	wire _w31337_ ;
	wire _w31336_ ;
	wire _w31335_ ;
	wire _w31334_ ;
	wire _w31333_ ;
	wire _w31332_ ;
	wire _w31331_ ;
	wire _w31330_ ;
	wire _w31329_ ;
	wire _w31328_ ;
	wire _w31327_ ;
	wire _w31326_ ;
	wire _w31325_ ;
	wire _w31324_ ;
	wire _w31323_ ;
	wire _w31322_ ;
	wire _w31321_ ;
	wire _w31320_ ;
	wire _w31319_ ;
	wire _w31318_ ;
	wire _w31317_ ;
	wire _w31316_ ;
	wire _w31315_ ;
	wire _w31314_ ;
	wire _w31313_ ;
	wire _w31312_ ;
	wire _w31311_ ;
	wire _w31310_ ;
	wire _w31309_ ;
	wire _w31308_ ;
	wire _w31307_ ;
	wire _w31306_ ;
	wire _w31305_ ;
	wire _w31304_ ;
	wire _w31303_ ;
	wire _w31302_ ;
	wire _w31301_ ;
	wire _w31300_ ;
	wire _w31299_ ;
	wire _w31298_ ;
	wire _w31297_ ;
	wire _w31296_ ;
	wire _w31295_ ;
	wire _w31294_ ;
	wire _w31293_ ;
	wire _w31292_ ;
	wire _w31291_ ;
	wire _w31290_ ;
	wire _w31289_ ;
	wire _w31288_ ;
	wire _w31287_ ;
	wire _w31286_ ;
	wire _w31285_ ;
	wire _w31284_ ;
	wire _w31283_ ;
	wire _w31282_ ;
	wire _w31281_ ;
	wire _w31280_ ;
	wire _w31279_ ;
	wire _w31278_ ;
	wire _w31277_ ;
	wire _w31276_ ;
	wire _w31275_ ;
	wire _w31274_ ;
	wire _w31273_ ;
	wire _w31272_ ;
	wire _w31271_ ;
	wire _w31270_ ;
	wire _w31269_ ;
	wire _w31268_ ;
	wire _w31267_ ;
	wire _w31266_ ;
	wire _w31265_ ;
	wire _w31264_ ;
	wire _w31263_ ;
	wire _w31262_ ;
	wire _w31261_ ;
	wire _w31260_ ;
	wire _w31259_ ;
	wire _w31258_ ;
	wire _w31257_ ;
	wire _w31256_ ;
	wire _w31255_ ;
	wire _w31254_ ;
	wire _w31253_ ;
	wire _w31252_ ;
	wire _w31251_ ;
	wire _w31250_ ;
	wire _w31249_ ;
	wire _w31248_ ;
	wire _w31247_ ;
	wire _w31246_ ;
	wire _w31245_ ;
	wire _w31244_ ;
	wire _w31243_ ;
	wire _w31242_ ;
	wire _w31241_ ;
	wire _w31240_ ;
	wire _w31239_ ;
	wire _w31238_ ;
	wire _w31237_ ;
	wire _w31236_ ;
	wire _w31235_ ;
	wire _w31234_ ;
	wire _w31233_ ;
	wire _w31232_ ;
	wire _w31231_ ;
	wire _w31230_ ;
	wire _w31229_ ;
	wire _w31228_ ;
	wire _w31227_ ;
	wire _w31226_ ;
	wire _w31225_ ;
	wire _w31224_ ;
	wire _w31223_ ;
	wire _w31222_ ;
	wire _w31221_ ;
	wire _w31220_ ;
	wire _w31219_ ;
	wire _w31218_ ;
	wire _w31217_ ;
	wire _w31216_ ;
	wire _w31215_ ;
	wire _w31214_ ;
	wire _w31213_ ;
	wire _w31212_ ;
	wire _w31211_ ;
	wire _w31210_ ;
	wire _w31209_ ;
	wire _w31208_ ;
	wire _w31207_ ;
	wire _w31206_ ;
	wire _w31205_ ;
	wire _w31204_ ;
	wire _w31203_ ;
	wire _w31202_ ;
	wire _w31201_ ;
	wire _w31200_ ;
	wire _w31199_ ;
	wire _w31198_ ;
	wire _w31197_ ;
	wire _w31196_ ;
	wire _w31195_ ;
	wire _w31194_ ;
	wire _w31193_ ;
	wire _w31192_ ;
	wire _w31191_ ;
	wire _w31190_ ;
	wire _w31189_ ;
	wire _w31188_ ;
	wire _w31187_ ;
	wire _w31186_ ;
	wire _w31185_ ;
	wire _w31184_ ;
	wire _w31183_ ;
	wire _w31182_ ;
	wire _w31181_ ;
	wire _w31180_ ;
	wire _w31179_ ;
	wire _w31178_ ;
	wire _w31177_ ;
	wire _w31176_ ;
	wire _w31175_ ;
	wire _w31174_ ;
	wire _w31173_ ;
	wire _w31172_ ;
	wire _w31171_ ;
	wire _w31170_ ;
	wire _w31169_ ;
	wire _w31168_ ;
	wire _w31167_ ;
	wire _w31166_ ;
	wire _w31165_ ;
	wire _w31164_ ;
	wire _w31163_ ;
	wire _w31162_ ;
	wire _w31161_ ;
	wire _w31160_ ;
	wire _w31159_ ;
	wire _w31158_ ;
	wire _w31157_ ;
	wire _w31156_ ;
	wire _w31155_ ;
	wire _w31154_ ;
	wire _w31153_ ;
	wire _w31152_ ;
	wire _w31151_ ;
	wire _w31150_ ;
	wire _w31149_ ;
	wire _w31148_ ;
	wire _w31147_ ;
	wire _w31146_ ;
	wire _w31145_ ;
	wire _w31144_ ;
	wire _w31143_ ;
	wire _w31142_ ;
	wire _w31141_ ;
	wire _w31140_ ;
	wire _w31139_ ;
	wire _w31138_ ;
	wire _w31137_ ;
	wire _w31136_ ;
	wire _w31135_ ;
	wire _w31134_ ;
	wire _w31133_ ;
	wire _w31132_ ;
	wire _w31131_ ;
	wire _w31130_ ;
	wire _w31129_ ;
	wire _w31128_ ;
	wire _w31127_ ;
	wire _w31126_ ;
	wire _w31125_ ;
	wire _w31124_ ;
	wire _w31123_ ;
	wire _w31122_ ;
	wire _w31121_ ;
	wire _w31120_ ;
	wire _w31119_ ;
	wire _w31118_ ;
	wire _w31117_ ;
	wire _w31116_ ;
	wire _w31115_ ;
	wire _w31114_ ;
	wire _w31113_ ;
	wire _w31112_ ;
	wire _w31111_ ;
	wire _w31110_ ;
	wire _w31109_ ;
	wire _w31108_ ;
	wire _w31107_ ;
	wire _w31106_ ;
	wire _w31105_ ;
	wire _w31104_ ;
	wire _w31103_ ;
	wire _w31102_ ;
	wire _w31101_ ;
	wire _w31100_ ;
	wire _w31099_ ;
	wire _w31098_ ;
	wire _w31097_ ;
	wire _w31096_ ;
	wire _w31095_ ;
	wire _w31094_ ;
	wire _w31093_ ;
	wire _w31092_ ;
	wire _w31091_ ;
	wire _w31090_ ;
	wire _w31089_ ;
	wire _w31088_ ;
	wire _w31087_ ;
	wire _w31086_ ;
	wire _w31085_ ;
	wire _w31084_ ;
	wire _w31083_ ;
	wire _w31082_ ;
	wire _w31081_ ;
	wire _w31080_ ;
	wire _w31079_ ;
	wire _w31078_ ;
	wire _w31077_ ;
	wire _w31076_ ;
	wire _w31075_ ;
	wire _w31074_ ;
	wire _w31073_ ;
	wire _w31072_ ;
	wire _w31071_ ;
	wire _w31070_ ;
	wire _w31069_ ;
	wire _w31068_ ;
	wire _w31067_ ;
	wire _w31066_ ;
	wire _w31065_ ;
	wire _w31064_ ;
	wire _w31063_ ;
	wire _w31062_ ;
	wire _w31061_ ;
	wire _w31060_ ;
	wire _w31059_ ;
	wire _w31058_ ;
	wire _w31057_ ;
	wire _w31056_ ;
	wire _w31055_ ;
	wire _w31054_ ;
	wire _w31053_ ;
	wire _w31052_ ;
	wire _w31051_ ;
	wire _w31050_ ;
	wire _w31049_ ;
	wire _w31048_ ;
	wire _w31047_ ;
	wire _w31046_ ;
	wire _w31045_ ;
	wire _w31044_ ;
	wire _w31043_ ;
	wire _w31042_ ;
	wire _w31041_ ;
	wire _w31040_ ;
	wire _w31039_ ;
	wire _w31038_ ;
	wire _w31037_ ;
	wire _w31036_ ;
	wire _w31035_ ;
	wire _w31034_ ;
	wire _w31033_ ;
	wire _w31032_ ;
	wire _w31031_ ;
	wire _w31030_ ;
	wire _w31029_ ;
	wire _w31028_ ;
	wire _w31027_ ;
	wire _w31026_ ;
	wire _w31025_ ;
	wire _w31024_ ;
	wire _w31023_ ;
	wire _w31022_ ;
	wire _w31021_ ;
	wire _w31020_ ;
	wire _w31019_ ;
	wire _w31018_ ;
	wire _w31017_ ;
	wire _w31016_ ;
	wire _w31015_ ;
	wire _w31014_ ;
	wire _w31013_ ;
	wire _w31012_ ;
	wire _w31011_ ;
	wire _w31010_ ;
	wire _w31009_ ;
	wire _w31008_ ;
	wire _w31007_ ;
	wire _w31006_ ;
	wire _w31005_ ;
	wire _w31004_ ;
	wire _w31003_ ;
	wire _w31002_ ;
	wire _w31001_ ;
	wire _w31000_ ;
	wire _w30999_ ;
	wire _w30998_ ;
	wire _w30997_ ;
	wire _w30996_ ;
	wire _w30995_ ;
	wire _w30994_ ;
	wire _w30993_ ;
	wire _w30992_ ;
	wire _w30991_ ;
	wire _w30990_ ;
	wire _w30989_ ;
	wire _w30988_ ;
	wire _w30987_ ;
	wire _w30986_ ;
	wire _w30985_ ;
	wire _w30984_ ;
	wire _w30983_ ;
	wire _w30982_ ;
	wire _w30981_ ;
	wire _w30980_ ;
	wire _w30979_ ;
	wire _w30978_ ;
	wire _w30977_ ;
	wire _w30976_ ;
	wire _w30975_ ;
	wire _w30974_ ;
	wire _w30973_ ;
	wire _w30972_ ;
	wire _w30971_ ;
	wire _w30970_ ;
	wire _w30969_ ;
	wire _w30968_ ;
	wire _w30967_ ;
	wire _w30966_ ;
	wire _w30965_ ;
	wire _w30964_ ;
	wire _w30963_ ;
	wire _w30962_ ;
	wire _w30961_ ;
	wire _w30960_ ;
	wire _w30959_ ;
	wire _w30958_ ;
	wire _w30957_ ;
	wire _w30956_ ;
	wire _w30955_ ;
	wire _w30954_ ;
	wire _w30953_ ;
	wire _w30952_ ;
	wire _w30951_ ;
	wire _w30950_ ;
	wire _w30949_ ;
	wire _w30948_ ;
	wire _w30947_ ;
	wire _w30946_ ;
	wire _w30945_ ;
	wire _w30944_ ;
	wire _w30943_ ;
	wire _w30942_ ;
	wire _w30941_ ;
	wire _w30940_ ;
	wire _w30939_ ;
	wire _w30938_ ;
	wire _w30937_ ;
	wire _w30936_ ;
	wire _w30935_ ;
	wire _w30934_ ;
	wire _w30933_ ;
	wire _w30932_ ;
	wire _w30931_ ;
	wire _w30930_ ;
	wire _w30929_ ;
	wire _w30928_ ;
	wire _w30927_ ;
	wire _w30926_ ;
	wire _w30925_ ;
	wire _w30924_ ;
	wire _w30923_ ;
	wire _w30922_ ;
	wire _w30921_ ;
	wire _w30920_ ;
	wire _w30919_ ;
	wire _w30918_ ;
	wire _w30917_ ;
	wire _w30916_ ;
	wire _w30915_ ;
	wire _w30914_ ;
	wire _w30913_ ;
	wire _w30912_ ;
	wire _w30911_ ;
	wire _w30910_ ;
	wire _w30909_ ;
	wire _w30908_ ;
	wire _w30907_ ;
	wire _w30906_ ;
	wire _w30905_ ;
	wire _w30904_ ;
	wire _w30903_ ;
	wire _w30902_ ;
	wire _w30901_ ;
	wire _w30900_ ;
	wire _w30899_ ;
	wire _w30898_ ;
	wire _w30897_ ;
	wire _w30896_ ;
	wire _w30895_ ;
	wire _w30894_ ;
	wire _w30893_ ;
	wire _w30892_ ;
	wire _w30891_ ;
	wire _w30890_ ;
	wire _w30889_ ;
	wire _w30888_ ;
	wire _w30887_ ;
	wire _w30886_ ;
	wire _w30885_ ;
	wire _w30884_ ;
	wire _w30883_ ;
	wire _w30882_ ;
	wire _w30881_ ;
	wire _w30880_ ;
	wire _w30879_ ;
	wire _w30878_ ;
	wire _w30877_ ;
	wire _w30876_ ;
	wire _w30875_ ;
	wire _w30874_ ;
	wire _w30873_ ;
	wire _w30872_ ;
	wire _w30871_ ;
	wire _w30870_ ;
	wire _w30869_ ;
	wire _w30868_ ;
	wire _w30867_ ;
	wire _w30866_ ;
	wire _w30865_ ;
	wire _w30864_ ;
	wire _w30863_ ;
	wire _w30862_ ;
	wire _w30861_ ;
	wire _w30860_ ;
	wire _w30859_ ;
	wire _w30858_ ;
	wire _w30857_ ;
	wire _w30856_ ;
	wire _w30855_ ;
	wire _w30854_ ;
	wire _w30853_ ;
	wire _w30852_ ;
	wire _w30851_ ;
	wire _w30850_ ;
	wire _w30849_ ;
	wire _w30848_ ;
	wire _w30847_ ;
	wire _w30846_ ;
	wire _w30845_ ;
	wire _w30844_ ;
	wire _w30843_ ;
	wire _w30842_ ;
	wire _w30841_ ;
	wire _w30840_ ;
	wire _w30839_ ;
	wire _w30838_ ;
	wire _w30837_ ;
	wire _w30836_ ;
	wire _w30835_ ;
	wire _w30834_ ;
	wire _w30833_ ;
	wire _w30832_ ;
	wire _w30831_ ;
	wire _w30830_ ;
	wire _w30829_ ;
	wire _w30828_ ;
	wire _w30827_ ;
	wire _w30826_ ;
	wire _w30825_ ;
	wire _w30824_ ;
	wire _w30823_ ;
	wire _w30822_ ;
	wire _w30821_ ;
	wire _w30820_ ;
	wire _w30819_ ;
	wire _w30818_ ;
	wire _w30817_ ;
	wire _w30816_ ;
	wire _w30815_ ;
	wire _w30814_ ;
	wire _w30813_ ;
	wire _w30812_ ;
	wire _w30811_ ;
	wire _w30810_ ;
	wire _w30809_ ;
	wire _w30808_ ;
	wire _w30807_ ;
	wire _w30806_ ;
	wire _w30805_ ;
	wire _w30804_ ;
	wire _w30803_ ;
	wire _w30802_ ;
	wire _w30801_ ;
	wire _w30800_ ;
	wire _w30799_ ;
	wire _w30798_ ;
	wire _w30797_ ;
	wire _w30796_ ;
	wire _w30795_ ;
	wire _w30794_ ;
	wire _w30793_ ;
	wire _w30792_ ;
	wire _w30791_ ;
	wire _w30790_ ;
	wire _w30789_ ;
	wire _w30788_ ;
	wire _w30787_ ;
	wire _w30786_ ;
	wire _w30785_ ;
	wire _w30784_ ;
	wire _w30783_ ;
	wire _w30782_ ;
	wire _w30781_ ;
	wire _w30780_ ;
	wire _w30779_ ;
	wire _w30778_ ;
	wire _w30777_ ;
	wire _w30776_ ;
	wire _w30775_ ;
	wire _w30774_ ;
	wire _w30773_ ;
	wire _w30772_ ;
	wire _w30771_ ;
	wire _w30770_ ;
	wire _w30769_ ;
	wire _w30768_ ;
	wire _w30767_ ;
	wire _w30766_ ;
	wire _w30765_ ;
	wire _w30764_ ;
	wire _w30763_ ;
	wire _w30762_ ;
	wire _w30761_ ;
	wire _w30760_ ;
	wire _w30759_ ;
	wire _w30758_ ;
	wire _w30757_ ;
	wire _w30756_ ;
	wire _w30755_ ;
	wire _w30754_ ;
	wire _w30753_ ;
	wire _w30752_ ;
	wire _w30751_ ;
	wire _w30750_ ;
	wire _w30749_ ;
	wire _w30748_ ;
	wire _w30747_ ;
	wire _w30746_ ;
	wire _w30745_ ;
	wire _w30744_ ;
	wire _w30743_ ;
	wire _w30742_ ;
	wire _w30741_ ;
	wire _w30740_ ;
	wire _w30739_ ;
	wire _w30738_ ;
	wire _w30737_ ;
	wire _w30736_ ;
	wire _w30735_ ;
	wire _w30734_ ;
	wire _w30733_ ;
	wire _w30732_ ;
	wire _w30731_ ;
	wire _w30730_ ;
	wire _w30729_ ;
	wire _w30728_ ;
	wire _w30727_ ;
	wire _w30726_ ;
	wire _w30725_ ;
	wire _w30724_ ;
	wire _w30723_ ;
	wire _w30722_ ;
	wire _w30721_ ;
	wire _w30720_ ;
	wire _w30719_ ;
	wire _w30718_ ;
	wire _w30717_ ;
	wire _w30716_ ;
	wire _w30715_ ;
	wire _w30714_ ;
	wire _w30713_ ;
	wire _w30712_ ;
	wire _w30711_ ;
	wire _w30710_ ;
	wire _w30709_ ;
	wire _w30708_ ;
	wire _w30707_ ;
	wire _w30706_ ;
	wire _w30705_ ;
	wire _w30704_ ;
	wire _w30703_ ;
	wire _w30702_ ;
	wire _w30701_ ;
	wire _w30700_ ;
	wire _w30699_ ;
	wire _w30698_ ;
	wire _w30697_ ;
	wire _w30696_ ;
	wire _w30695_ ;
	wire _w30694_ ;
	wire _w30693_ ;
	wire _w30692_ ;
	wire _w30691_ ;
	wire _w30690_ ;
	wire _w30689_ ;
	wire _w30688_ ;
	wire _w30687_ ;
	wire _w30686_ ;
	wire _w30685_ ;
	wire _w30684_ ;
	wire _w30683_ ;
	wire _w30682_ ;
	wire _w30681_ ;
	wire _w30680_ ;
	wire _w30679_ ;
	wire _w30678_ ;
	wire _w30677_ ;
	wire _w30676_ ;
	wire _w30675_ ;
	wire _w30674_ ;
	wire _w30673_ ;
	wire _w30672_ ;
	wire _w30671_ ;
	wire _w30670_ ;
	wire _w30669_ ;
	wire _w30668_ ;
	wire _w30667_ ;
	wire _w30666_ ;
	wire _w30665_ ;
	wire _w30664_ ;
	wire _w30663_ ;
	wire _w30662_ ;
	wire _w30661_ ;
	wire _w30660_ ;
	wire _w30659_ ;
	wire _w30658_ ;
	wire _w30657_ ;
	wire _w30656_ ;
	wire _w30655_ ;
	wire _w30654_ ;
	wire _w30653_ ;
	wire _w30652_ ;
	wire _w30651_ ;
	wire _w30650_ ;
	wire _w30649_ ;
	wire _w30648_ ;
	wire _w30647_ ;
	wire _w30646_ ;
	wire _w30645_ ;
	wire _w30644_ ;
	wire _w30643_ ;
	wire _w30642_ ;
	wire _w30641_ ;
	wire _w30640_ ;
	wire _w30639_ ;
	wire _w30638_ ;
	wire _w30637_ ;
	wire _w30636_ ;
	wire _w30635_ ;
	wire _w30634_ ;
	wire _w30633_ ;
	wire _w30632_ ;
	wire _w30631_ ;
	wire _w30630_ ;
	wire _w30629_ ;
	wire _w30628_ ;
	wire _w30627_ ;
	wire _w30626_ ;
	wire _w30625_ ;
	wire _w30624_ ;
	wire _w30623_ ;
	wire _w30622_ ;
	wire _w30621_ ;
	wire _w30620_ ;
	wire _w30619_ ;
	wire _w30618_ ;
	wire _w30617_ ;
	wire _w30616_ ;
	wire _w30615_ ;
	wire _w30614_ ;
	wire _w30613_ ;
	wire _w30612_ ;
	wire _w30611_ ;
	wire _w30610_ ;
	wire _w30609_ ;
	wire _w30608_ ;
	wire _w30607_ ;
	wire _w30606_ ;
	wire _w30605_ ;
	wire _w30604_ ;
	wire _w30603_ ;
	wire _w30602_ ;
	wire _w30601_ ;
	wire _w30600_ ;
	wire _w30599_ ;
	wire _w30598_ ;
	wire _w30597_ ;
	wire _w30596_ ;
	wire _w30595_ ;
	wire _w30594_ ;
	wire _w30593_ ;
	wire _w30592_ ;
	wire _w30591_ ;
	wire _w30590_ ;
	wire _w30589_ ;
	wire _w30588_ ;
	wire _w30587_ ;
	wire _w30586_ ;
	wire _w30585_ ;
	wire _w30584_ ;
	wire _w30583_ ;
	wire _w30582_ ;
	wire _w30581_ ;
	wire _w30580_ ;
	wire _w30579_ ;
	wire _w30578_ ;
	wire _w30577_ ;
	wire _w30576_ ;
	wire _w30575_ ;
	wire _w30574_ ;
	wire _w30573_ ;
	wire _w30572_ ;
	wire _w30571_ ;
	wire _w30570_ ;
	wire _w30569_ ;
	wire _w30568_ ;
	wire _w30567_ ;
	wire _w30566_ ;
	wire _w30565_ ;
	wire _w30564_ ;
	wire _w30563_ ;
	wire _w30562_ ;
	wire _w30561_ ;
	wire _w30560_ ;
	wire _w30559_ ;
	wire _w30558_ ;
	wire _w30557_ ;
	wire _w30556_ ;
	wire _w30555_ ;
	wire _w30554_ ;
	wire _w30553_ ;
	wire _w30552_ ;
	wire _w30551_ ;
	wire _w30550_ ;
	wire _w30549_ ;
	wire _w30548_ ;
	wire _w30547_ ;
	wire _w30546_ ;
	wire _w30545_ ;
	wire _w30544_ ;
	wire _w30543_ ;
	wire _w30542_ ;
	wire _w30541_ ;
	wire _w30540_ ;
	wire _w30539_ ;
	wire _w30538_ ;
	wire _w30537_ ;
	wire _w30536_ ;
	wire _w30535_ ;
	wire _w30534_ ;
	wire _w30533_ ;
	wire _w30532_ ;
	wire _w30531_ ;
	wire _w30530_ ;
	wire _w30529_ ;
	wire _w30528_ ;
	wire _w30527_ ;
	wire _w30526_ ;
	wire _w30525_ ;
	wire _w30524_ ;
	wire _w30523_ ;
	wire _w30522_ ;
	wire _w30521_ ;
	wire _w30520_ ;
	wire _w30519_ ;
	wire _w30518_ ;
	wire _w30517_ ;
	wire _w30516_ ;
	wire _w30515_ ;
	wire _w30514_ ;
	wire _w30513_ ;
	wire _w30512_ ;
	wire _w30511_ ;
	wire _w30510_ ;
	wire _w30509_ ;
	wire _w30508_ ;
	wire _w30507_ ;
	wire _w30506_ ;
	wire _w30505_ ;
	wire _w30504_ ;
	wire _w30503_ ;
	wire _w30502_ ;
	wire _w30501_ ;
	wire _w30500_ ;
	wire _w30499_ ;
	wire _w30498_ ;
	wire _w30497_ ;
	wire _w30496_ ;
	wire _w30495_ ;
	wire _w30494_ ;
	wire _w30493_ ;
	wire _w30492_ ;
	wire _w30491_ ;
	wire _w30490_ ;
	wire _w30489_ ;
	wire _w30488_ ;
	wire _w30487_ ;
	wire _w30486_ ;
	wire _w30485_ ;
	wire _w30484_ ;
	wire _w30483_ ;
	wire _w30482_ ;
	wire _w30481_ ;
	wire _w30480_ ;
	wire _w30479_ ;
	wire _w30478_ ;
	wire _w30477_ ;
	wire _w30476_ ;
	wire _w30475_ ;
	wire _w30474_ ;
	wire _w30473_ ;
	wire _w30472_ ;
	wire _w30471_ ;
	wire _w30470_ ;
	wire _w30469_ ;
	wire _w30468_ ;
	wire _w30467_ ;
	wire _w30466_ ;
	wire _w30465_ ;
	wire _w30464_ ;
	wire _w30463_ ;
	wire _w30462_ ;
	wire _w30461_ ;
	wire _w30460_ ;
	wire _w30459_ ;
	wire _w30458_ ;
	wire _w30457_ ;
	wire _w30456_ ;
	wire _w30455_ ;
	wire _w30454_ ;
	wire _w30453_ ;
	wire _w30452_ ;
	wire _w30451_ ;
	wire _w30450_ ;
	wire _w30449_ ;
	wire _w30448_ ;
	wire _w30447_ ;
	wire _w30446_ ;
	wire _w30445_ ;
	wire _w30444_ ;
	wire _w30443_ ;
	wire _w30442_ ;
	wire _w30441_ ;
	wire _w30440_ ;
	wire _w30439_ ;
	wire _w30438_ ;
	wire _w30437_ ;
	wire _w30436_ ;
	wire _w30435_ ;
	wire _w30434_ ;
	wire _w30433_ ;
	wire _w30432_ ;
	wire _w30431_ ;
	wire _w30430_ ;
	wire _w30429_ ;
	wire _w30428_ ;
	wire _w30427_ ;
	wire _w30426_ ;
	wire _w30425_ ;
	wire _w30424_ ;
	wire _w30423_ ;
	wire _w30422_ ;
	wire _w30421_ ;
	wire _w30420_ ;
	wire _w30419_ ;
	wire _w30418_ ;
	wire _w30417_ ;
	wire _w30416_ ;
	wire _w30415_ ;
	wire _w30414_ ;
	wire _w30413_ ;
	wire _w30412_ ;
	wire _w30411_ ;
	wire _w30410_ ;
	wire _w30409_ ;
	wire _w30408_ ;
	wire _w30407_ ;
	wire _w30406_ ;
	wire _w30405_ ;
	wire _w30404_ ;
	wire _w30403_ ;
	wire _w30402_ ;
	wire _w30401_ ;
	wire _w30400_ ;
	wire _w30399_ ;
	wire _w30398_ ;
	wire _w30397_ ;
	wire _w30396_ ;
	wire _w30395_ ;
	wire _w30394_ ;
	wire _w30393_ ;
	wire _w30392_ ;
	wire _w30391_ ;
	wire _w30390_ ;
	wire _w30389_ ;
	wire _w30388_ ;
	wire _w30387_ ;
	wire _w30386_ ;
	wire _w30385_ ;
	wire _w30384_ ;
	wire _w30383_ ;
	wire _w30382_ ;
	wire _w30381_ ;
	wire _w30380_ ;
	wire _w30379_ ;
	wire _w30378_ ;
	wire _w30377_ ;
	wire _w30376_ ;
	wire _w30375_ ;
	wire _w30374_ ;
	wire _w30373_ ;
	wire _w30372_ ;
	wire _w30371_ ;
	wire _w30370_ ;
	wire _w30369_ ;
	wire _w30368_ ;
	wire _w30367_ ;
	wire _w30366_ ;
	wire _w30365_ ;
	wire _w30364_ ;
	wire _w30363_ ;
	wire _w30362_ ;
	wire _w30361_ ;
	wire _w30360_ ;
	wire _w30359_ ;
	wire _w30358_ ;
	wire _w30357_ ;
	wire _w30356_ ;
	wire _w30355_ ;
	wire _w30354_ ;
	wire _w30353_ ;
	wire _w30352_ ;
	wire _w30351_ ;
	wire _w30350_ ;
	wire _w30349_ ;
	wire _w30348_ ;
	wire _w30347_ ;
	wire _w30346_ ;
	wire _w30345_ ;
	wire _w30344_ ;
	wire _w30343_ ;
	wire _w30342_ ;
	wire _w30341_ ;
	wire _w30340_ ;
	wire _w30339_ ;
	wire _w30338_ ;
	wire _w30337_ ;
	wire _w30336_ ;
	wire _w30335_ ;
	wire _w30334_ ;
	wire _w30333_ ;
	wire _w30332_ ;
	wire _w30331_ ;
	wire _w30330_ ;
	wire _w30329_ ;
	wire _w30328_ ;
	wire _w30327_ ;
	wire _w30326_ ;
	wire _w30325_ ;
	wire _w30324_ ;
	wire _w30323_ ;
	wire _w30322_ ;
	wire _w30321_ ;
	wire _w30320_ ;
	wire _w30319_ ;
	wire _w30318_ ;
	wire _w30317_ ;
	wire _w30316_ ;
	wire _w30315_ ;
	wire _w30314_ ;
	wire _w30313_ ;
	wire _w30312_ ;
	wire _w30311_ ;
	wire _w30310_ ;
	wire _w30309_ ;
	wire _w30308_ ;
	wire _w30307_ ;
	wire _w30306_ ;
	wire _w30305_ ;
	wire _w30304_ ;
	wire _w30303_ ;
	wire _w30302_ ;
	wire _w30301_ ;
	wire _w30300_ ;
	wire _w30299_ ;
	wire _w30298_ ;
	wire _w30297_ ;
	wire _w30296_ ;
	wire _w30295_ ;
	wire _w30294_ ;
	wire _w30293_ ;
	wire _w30292_ ;
	wire _w30291_ ;
	wire _w30290_ ;
	wire _w30289_ ;
	wire _w30288_ ;
	wire _w30287_ ;
	wire _w30286_ ;
	wire _w30285_ ;
	wire _w30284_ ;
	wire _w30283_ ;
	wire _w30282_ ;
	wire _w30281_ ;
	wire _w30280_ ;
	wire _w30279_ ;
	wire _w30278_ ;
	wire _w30277_ ;
	wire _w30276_ ;
	wire _w30275_ ;
	wire _w30274_ ;
	wire _w30273_ ;
	wire _w30272_ ;
	wire _w30271_ ;
	wire _w30270_ ;
	wire _w30269_ ;
	wire _w30268_ ;
	wire _w30267_ ;
	wire _w30266_ ;
	wire _w30265_ ;
	wire _w30264_ ;
	wire _w30263_ ;
	wire _w30262_ ;
	wire _w30261_ ;
	wire _w30260_ ;
	wire _w30259_ ;
	wire _w30258_ ;
	wire _w30257_ ;
	wire _w30256_ ;
	wire _w30255_ ;
	wire _w30254_ ;
	wire _w30253_ ;
	wire _w30252_ ;
	wire _w30251_ ;
	wire _w30250_ ;
	wire _w30249_ ;
	wire _w30248_ ;
	wire _w30247_ ;
	wire _w30246_ ;
	wire _w30245_ ;
	wire _w30244_ ;
	wire _w30243_ ;
	wire _w30242_ ;
	wire _w30241_ ;
	wire _w30240_ ;
	wire _w30239_ ;
	wire _w30238_ ;
	wire _w30237_ ;
	wire _w30236_ ;
	wire _w30235_ ;
	wire _w30234_ ;
	wire _w30233_ ;
	wire _w30232_ ;
	wire _w30231_ ;
	wire _w30230_ ;
	wire _w30229_ ;
	wire _w30228_ ;
	wire _w30227_ ;
	wire _w30226_ ;
	wire _w30225_ ;
	wire _w30224_ ;
	wire _w30223_ ;
	wire _w30222_ ;
	wire _w30221_ ;
	wire _w30220_ ;
	wire _w30219_ ;
	wire _w30218_ ;
	wire _w30217_ ;
	wire _w30216_ ;
	wire _w30215_ ;
	wire _w30214_ ;
	wire _w30213_ ;
	wire _w30212_ ;
	wire _w30211_ ;
	wire _w30210_ ;
	wire _w30209_ ;
	wire _w30208_ ;
	wire _w30207_ ;
	wire _w30206_ ;
	wire _w30205_ ;
	wire _w30204_ ;
	wire _w30203_ ;
	wire _w30202_ ;
	wire _w30201_ ;
	wire _w30200_ ;
	wire _w30199_ ;
	wire _w30198_ ;
	wire _w30197_ ;
	wire _w30196_ ;
	wire _w30195_ ;
	wire _w30194_ ;
	wire _w30193_ ;
	wire _w30192_ ;
	wire _w30191_ ;
	wire _w30190_ ;
	wire _w30189_ ;
	wire _w30188_ ;
	wire _w30187_ ;
	wire _w30186_ ;
	wire _w30185_ ;
	wire _w30184_ ;
	wire _w30183_ ;
	wire _w30182_ ;
	wire _w30181_ ;
	wire _w30180_ ;
	wire _w30179_ ;
	wire _w30178_ ;
	wire _w30177_ ;
	wire _w30176_ ;
	wire _w30175_ ;
	wire _w30174_ ;
	wire _w30173_ ;
	wire _w30172_ ;
	wire _w30171_ ;
	wire _w30170_ ;
	wire _w30169_ ;
	wire _w30168_ ;
	wire _w30167_ ;
	wire _w30166_ ;
	wire _w30165_ ;
	wire _w30164_ ;
	wire _w30163_ ;
	wire _w30162_ ;
	wire _w30161_ ;
	wire _w30160_ ;
	wire _w30159_ ;
	wire _w30158_ ;
	wire _w30157_ ;
	wire _w30156_ ;
	wire _w30155_ ;
	wire _w30154_ ;
	wire _w30153_ ;
	wire _w30152_ ;
	wire _w30151_ ;
	wire _w30150_ ;
	wire _w30149_ ;
	wire _w30148_ ;
	wire _w30147_ ;
	wire _w30146_ ;
	wire _w30145_ ;
	wire _w30144_ ;
	wire _w30143_ ;
	wire _w30142_ ;
	wire _w30141_ ;
	wire _w30140_ ;
	wire _w30139_ ;
	wire _w30138_ ;
	wire _w30137_ ;
	wire _w30136_ ;
	wire _w30135_ ;
	wire _w30134_ ;
	wire _w30133_ ;
	wire _w30132_ ;
	wire _w30131_ ;
	wire _w30130_ ;
	wire _w30129_ ;
	wire _w30128_ ;
	wire _w30127_ ;
	wire _w30126_ ;
	wire _w30125_ ;
	wire _w30124_ ;
	wire _w30123_ ;
	wire _w30122_ ;
	wire _w30121_ ;
	wire _w30120_ ;
	wire _w30119_ ;
	wire _w30118_ ;
	wire _w30117_ ;
	wire _w30116_ ;
	wire _w30115_ ;
	wire _w30114_ ;
	wire _w30113_ ;
	wire _w30112_ ;
	wire _w30111_ ;
	wire _w30110_ ;
	wire _w30109_ ;
	wire _w30108_ ;
	wire _w30107_ ;
	wire _w30106_ ;
	wire _w30105_ ;
	wire _w30104_ ;
	wire _w30103_ ;
	wire _w30102_ ;
	wire _w30101_ ;
	wire _w30100_ ;
	wire _w30099_ ;
	wire _w30098_ ;
	wire _w30097_ ;
	wire _w30096_ ;
	wire _w30095_ ;
	wire _w30094_ ;
	wire _w30093_ ;
	wire _w30092_ ;
	wire _w30091_ ;
	wire _w30090_ ;
	wire _w30089_ ;
	wire _w30088_ ;
	wire _w30087_ ;
	wire _w30086_ ;
	wire _w30085_ ;
	wire _w30084_ ;
	wire _w30083_ ;
	wire _w30082_ ;
	wire _w30081_ ;
	wire _w30080_ ;
	wire _w30079_ ;
	wire _w30078_ ;
	wire _w30077_ ;
	wire _w30076_ ;
	wire _w30075_ ;
	wire _w30074_ ;
	wire _w30073_ ;
	wire _w30072_ ;
	wire _w30071_ ;
	wire _w30070_ ;
	wire _w30069_ ;
	wire _w30068_ ;
	wire _w30067_ ;
	wire _w30066_ ;
	wire _w30065_ ;
	wire _w30064_ ;
	wire _w30063_ ;
	wire _w30062_ ;
	wire _w30061_ ;
	wire _w30060_ ;
	wire _w30059_ ;
	wire _w30058_ ;
	wire _w30057_ ;
	wire _w30056_ ;
	wire _w30055_ ;
	wire _w30054_ ;
	wire _w30053_ ;
	wire _w30052_ ;
	wire _w30051_ ;
	wire _w30050_ ;
	wire _w30049_ ;
	wire _w30048_ ;
	wire _w30047_ ;
	wire _w30046_ ;
	wire _w30045_ ;
	wire _w30044_ ;
	wire _w30043_ ;
	wire _w30042_ ;
	wire _w30041_ ;
	wire _w30040_ ;
	wire _w30039_ ;
	wire _w30038_ ;
	wire _w30037_ ;
	wire _w30036_ ;
	wire _w30035_ ;
	wire _w30034_ ;
	wire _w30033_ ;
	wire _w30032_ ;
	wire _w30031_ ;
	wire _w30030_ ;
	wire _w30029_ ;
	wire _w30028_ ;
	wire _w30027_ ;
	wire _w30026_ ;
	wire _w30025_ ;
	wire _w30024_ ;
	wire _w30023_ ;
	wire _w30022_ ;
	wire _w30021_ ;
	wire _w30020_ ;
	wire _w30019_ ;
	wire _w30018_ ;
	wire _w30017_ ;
	wire _w30016_ ;
	wire _w30015_ ;
	wire _w30014_ ;
	wire _w30013_ ;
	wire _w30012_ ;
	wire _w30011_ ;
	wire _w30010_ ;
	wire _w30009_ ;
	wire _w30008_ ;
	wire _w30007_ ;
	wire _w30006_ ;
	wire _w30005_ ;
	wire _w30004_ ;
	wire _w30003_ ;
	wire _w30002_ ;
	wire _w30001_ ;
	wire _w30000_ ;
	wire _w29999_ ;
	wire _w29998_ ;
	wire _w29997_ ;
	wire _w29996_ ;
	wire _w29995_ ;
	wire _w29994_ ;
	wire _w29993_ ;
	wire _w29992_ ;
	wire _w29991_ ;
	wire _w29990_ ;
	wire _w29989_ ;
	wire _w29988_ ;
	wire _w29987_ ;
	wire _w29986_ ;
	wire _w29985_ ;
	wire _w29984_ ;
	wire _w29983_ ;
	wire _w29982_ ;
	wire _w29981_ ;
	wire _w29980_ ;
	wire _w29979_ ;
	wire _w29978_ ;
	wire _w29977_ ;
	wire _w29976_ ;
	wire _w29975_ ;
	wire _w29974_ ;
	wire _w29973_ ;
	wire _w29972_ ;
	wire _w29971_ ;
	wire _w29970_ ;
	wire _w29969_ ;
	wire _w29968_ ;
	wire _w29967_ ;
	wire _w29966_ ;
	wire _w29965_ ;
	wire _w29964_ ;
	wire _w29963_ ;
	wire _w29962_ ;
	wire _w29961_ ;
	wire _w29960_ ;
	wire _w29959_ ;
	wire _w29958_ ;
	wire _w29957_ ;
	wire _w29956_ ;
	wire _w29955_ ;
	wire _w29954_ ;
	wire _w29953_ ;
	wire _w29952_ ;
	wire _w29951_ ;
	wire _w29950_ ;
	wire _w29949_ ;
	wire _w29948_ ;
	wire _w29947_ ;
	wire _w29946_ ;
	wire _w29945_ ;
	wire _w29944_ ;
	wire _w29943_ ;
	wire _w29942_ ;
	wire _w29941_ ;
	wire _w29940_ ;
	wire _w29939_ ;
	wire _w29938_ ;
	wire _w29937_ ;
	wire _w29936_ ;
	wire _w29935_ ;
	wire _w29934_ ;
	wire _w29933_ ;
	wire _w29932_ ;
	wire _w29931_ ;
	wire _w29930_ ;
	wire _w29929_ ;
	wire _w29928_ ;
	wire _w29927_ ;
	wire _w29926_ ;
	wire _w29925_ ;
	wire _w29924_ ;
	wire _w29923_ ;
	wire _w29922_ ;
	wire _w29921_ ;
	wire _w29920_ ;
	wire _w29919_ ;
	wire _w29918_ ;
	wire _w29917_ ;
	wire _w29916_ ;
	wire _w29915_ ;
	wire _w29914_ ;
	wire _w29913_ ;
	wire _w29912_ ;
	wire _w29911_ ;
	wire _w29910_ ;
	wire _w29909_ ;
	wire _w29908_ ;
	wire _w29907_ ;
	wire _w29906_ ;
	wire _w29905_ ;
	wire _w29904_ ;
	wire _w29903_ ;
	wire _w29902_ ;
	wire _w29901_ ;
	wire _w29900_ ;
	wire _w29899_ ;
	wire _w29898_ ;
	wire _w29897_ ;
	wire _w29896_ ;
	wire _w29895_ ;
	wire _w29894_ ;
	wire _w29893_ ;
	wire _w29892_ ;
	wire _w29891_ ;
	wire _w29890_ ;
	wire _w29889_ ;
	wire _w29888_ ;
	wire _w29887_ ;
	wire _w29886_ ;
	wire _w29885_ ;
	wire _w29884_ ;
	wire _w29883_ ;
	wire _w29882_ ;
	wire _w29881_ ;
	wire _w29880_ ;
	wire _w29879_ ;
	wire _w29878_ ;
	wire _w29877_ ;
	wire _w29876_ ;
	wire _w29875_ ;
	wire _w29874_ ;
	wire _w29873_ ;
	wire _w29872_ ;
	wire _w29871_ ;
	wire _w29870_ ;
	wire _w29869_ ;
	wire _w29868_ ;
	wire _w29867_ ;
	wire _w29866_ ;
	wire _w29865_ ;
	wire _w29864_ ;
	wire _w29863_ ;
	wire _w29862_ ;
	wire _w29861_ ;
	wire _w29860_ ;
	wire _w29859_ ;
	wire _w29858_ ;
	wire _w29857_ ;
	wire _w29856_ ;
	wire _w29855_ ;
	wire _w29854_ ;
	wire _w29853_ ;
	wire _w29852_ ;
	wire _w29851_ ;
	wire _w29850_ ;
	wire _w29849_ ;
	wire _w29848_ ;
	wire _w29847_ ;
	wire _w29846_ ;
	wire _w29845_ ;
	wire _w29844_ ;
	wire _w29843_ ;
	wire _w29842_ ;
	wire _w29841_ ;
	wire _w29840_ ;
	wire _w29839_ ;
	wire _w29838_ ;
	wire _w29837_ ;
	wire _w29836_ ;
	wire _w29835_ ;
	wire _w29834_ ;
	wire _w29833_ ;
	wire _w29832_ ;
	wire _w29831_ ;
	wire _w29830_ ;
	wire _w29829_ ;
	wire _w29828_ ;
	wire _w29827_ ;
	wire _w29826_ ;
	wire _w29825_ ;
	wire _w29824_ ;
	wire _w29823_ ;
	wire _w29822_ ;
	wire _w29821_ ;
	wire _w29820_ ;
	wire _w29819_ ;
	wire _w29818_ ;
	wire _w29817_ ;
	wire _w29816_ ;
	wire _w29815_ ;
	wire _w29814_ ;
	wire _w29813_ ;
	wire _w29812_ ;
	wire _w29811_ ;
	wire _w29810_ ;
	wire _w29809_ ;
	wire _w29808_ ;
	wire _w29807_ ;
	wire _w29806_ ;
	wire _w29805_ ;
	wire _w29804_ ;
	wire _w29803_ ;
	wire _w29802_ ;
	wire _w29801_ ;
	wire _w29800_ ;
	wire _w29799_ ;
	wire _w29798_ ;
	wire _w29797_ ;
	wire _w29796_ ;
	wire _w29795_ ;
	wire _w29794_ ;
	wire _w29793_ ;
	wire _w29792_ ;
	wire _w29791_ ;
	wire _w29790_ ;
	wire _w29789_ ;
	wire _w29788_ ;
	wire _w29787_ ;
	wire _w29786_ ;
	wire _w29785_ ;
	wire _w29784_ ;
	wire _w29783_ ;
	wire _w29782_ ;
	wire _w29781_ ;
	wire _w29780_ ;
	wire _w29779_ ;
	wire _w29778_ ;
	wire _w29777_ ;
	wire _w29776_ ;
	wire _w29775_ ;
	wire _w29774_ ;
	wire _w29773_ ;
	wire _w29772_ ;
	wire _w29771_ ;
	wire _w29770_ ;
	wire _w29769_ ;
	wire _w29768_ ;
	wire _w29767_ ;
	wire _w29766_ ;
	wire _w29765_ ;
	wire _w29764_ ;
	wire _w29763_ ;
	wire _w29762_ ;
	wire _w29761_ ;
	wire _w29760_ ;
	wire _w29759_ ;
	wire _w29758_ ;
	wire _w29757_ ;
	wire _w29756_ ;
	wire _w29755_ ;
	wire _w29754_ ;
	wire _w29753_ ;
	wire _w29752_ ;
	wire _w29751_ ;
	wire _w29750_ ;
	wire _w29749_ ;
	wire _w29748_ ;
	wire _w29747_ ;
	wire _w29746_ ;
	wire _w29745_ ;
	wire _w29744_ ;
	wire _w29743_ ;
	wire _w29742_ ;
	wire _w29741_ ;
	wire _w29740_ ;
	wire _w29739_ ;
	wire _w29738_ ;
	wire _w29737_ ;
	wire _w29736_ ;
	wire _w29735_ ;
	wire _w29734_ ;
	wire _w29733_ ;
	wire _w29732_ ;
	wire _w29731_ ;
	wire _w29730_ ;
	wire _w29729_ ;
	wire _w29728_ ;
	wire _w29727_ ;
	wire _w29726_ ;
	wire _w29725_ ;
	wire _w29724_ ;
	wire _w29723_ ;
	wire _w29722_ ;
	wire _w29721_ ;
	wire _w29720_ ;
	wire _w29719_ ;
	wire _w29718_ ;
	wire _w29717_ ;
	wire _w29716_ ;
	wire _w29715_ ;
	wire _w29714_ ;
	wire _w29713_ ;
	wire _w29712_ ;
	wire _w29711_ ;
	wire _w29710_ ;
	wire _w29709_ ;
	wire _w29708_ ;
	wire _w29707_ ;
	wire _w29706_ ;
	wire _w29705_ ;
	wire _w29704_ ;
	wire _w29703_ ;
	wire _w29702_ ;
	wire _w29701_ ;
	wire _w29700_ ;
	wire _w29699_ ;
	wire _w29698_ ;
	wire _w29697_ ;
	wire _w29696_ ;
	wire _w29695_ ;
	wire _w29694_ ;
	wire _w29693_ ;
	wire _w29692_ ;
	wire _w29691_ ;
	wire _w29690_ ;
	wire _w29689_ ;
	wire _w29688_ ;
	wire _w29687_ ;
	wire _w29686_ ;
	wire _w29685_ ;
	wire _w29684_ ;
	wire _w29683_ ;
	wire _w29682_ ;
	wire _w29681_ ;
	wire _w29680_ ;
	wire _w29679_ ;
	wire _w29678_ ;
	wire _w29677_ ;
	wire _w29676_ ;
	wire _w29675_ ;
	wire _w29674_ ;
	wire _w29673_ ;
	wire _w29672_ ;
	wire _w29671_ ;
	wire _w29670_ ;
	wire _w29669_ ;
	wire _w29668_ ;
	wire _w29667_ ;
	wire _w29666_ ;
	wire _w29665_ ;
	wire _w29664_ ;
	wire _w29663_ ;
	wire _w29662_ ;
	wire _w29661_ ;
	wire _w29660_ ;
	wire _w29659_ ;
	wire _w29658_ ;
	wire _w29657_ ;
	wire _w29656_ ;
	wire _w29655_ ;
	wire _w29654_ ;
	wire _w29653_ ;
	wire _w29652_ ;
	wire _w29651_ ;
	wire _w29650_ ;
	wire _w29649_ ;
	wire _w29648_ ;
	wire _w29647_ ;
	wire _w29646_ ;
	wire _w29645_ ;
	wire _w29644_ ;
	wire _w29643_ ;
	wire _w29642_ ;
	wire _w29641_ ;
	wire _w29640_ ;
	wire _w29639_ ;
	wire _w29638_ ;
	wire _w29637_ ;
	wire _w29636_ ;
	wire _w29635_ ;
	wire _w29634_ ;
	wire _w29633_ ;
	wire _w29632_ ;
	wire _w29631_ ;
	wire _w29630_ ;
	wire _w29629_ ;
	wire _w29628_ ;
	wire _w29627_ ;
	wire _w29626_ ;
	wire _w29625_ ;
	wire _w29624_ ;
	wire _w29623_ ;
	wire _w29622_ ;
	wire _w29621_ ;
	wire _w29620_ ;
	wire _w29619_ ;
	wire _w29618_ ;
	wire _w29617_ ;
	wire _w29616_ ;
	wire _w29615_ ;
	wire _w29614_ ;
	wire _w29613_ ;
	wire _w29612_ ;
	wire _w29611_ ;
	wire _w29610_ ;
	wire _w29609_ ;
	wire _w29608_ ;
	wire _w29607_ ;
	wire _w29606_ ;
	wire _w29605_ ;
	wire _w29604_ ;
	wire _w29603_ ;
	wire _w29602_ ;
	wire _w29601_ ;
	wire _w29600_ ;
	wire _w29599_ ;
	wire _w29598_ ;
	wire _w29597_ ;
	wire _w29596_ ;
	wire _w29595_ ;
	wire _w29594_ ;
	wire _w29593_ ;
	wire _w29592_ ;
	wire _w29591_ ;
	wire _w29590_ ;
	wire _w29589_ ;
	wire _w29588_ ;
	wire _w29587_ ;
	wire _w29586_ ;
	wire _w29585_ ;
	wire _w29584_ ;
	wire _w29583_ ;
	wire _w29582_ ;
	wire _w29581_ ;
	wire _w29580_ ;
	wire _w29579_ ;
	wire _w29578_ ;
	wire _w29577_ ;
	wire _w29576_ ;
	wire _w29575_ ;
	wire _w29574_ ;
	wire _w29573_ ;
	wire _w29572_ ;
	wire _w29571_ ;
	wire _w29570_ ;
	wire _w29569_ ;
	wire _w29568_ ;
	wire _w29567_ ;
	wire _w29566_ ;
	wire _w29565_ ;
	wire _w29564_ ;
	wire _w29563_ ;
	wire _w29562_ ;
	wire _w29561_ ;
	wire _w29560_ ;
	wire _w29559_ ;
	wire _w29558_ ;
	wire _w29557_ ;
	wire _w29556_ ;
	wire _w29555_ ;
	wire _w29554_ ;
	wire _w29553_ ;
	wire _w29552_ ;
	wire _w29551_ ;
	wire _w29550_ ;
	wire _w29549_ ;
	wire _w29548_ ;
	wire _w29547_ ;
	wire _w29546_ ;
	wire _w29545_ ;
	wire _w29544_ ;
	wire _w29543_ ;
	wire _w29542_ ;
	wire _w29541_ ;
	wire _w29540_ ;
	wire _w29539_ ;
	wire _w29538_ ;
	wire _w29537_ ;
	wire _w29536_ ;
	wire _w29535_ ;
	wire _w29534_ ;
	wire _w29533_ ;
	wire _w29532_ ;
	wire _w29531_ ;
	wire _w29530_ ;
	wire _w29529_ ;
	wire _w29528_ ;
	wire _w29527_ ;
	wire _w29526_ ;
	wire _w29525_ ;
	wire _w29524_ ;
	wire _w29523_ ;
	wire _w29522_ ;
	wire _w29521_ ;
	wire _w29520_ ;
	wire _w29519_ ;
	wire _w29518_ ;
	wire _w29517_ ;
	wire _w29516_ ;
	wire _w29515_ ;
	wire _w29514_ ;
	wire _w29513_ ;
	wire _w29512_ ;
	wire _w29511_ ;
	wire _w29510_ ;
	wire _w29509_ ;
	wire _w29508_ ;
	wire _w29507_ ;
	wire _w29506_ ;
	wire _w29505_ ;
	wire _w29504_ ;
	wire _w29503_ ;
	wire _w29502_ ;
	wire _w29501_ ;
	wire _w29500_ ;
	wire _w29499_ ;
	wire _w29498_ ;
	wire _w29497_ ;
	wire _w29496_ ;
	wire _w29495_ ;
	wire _w29494_ ;
	wire _w29493_ ;
	wire _w29492_ ;
	wire _w29491_ ;
	wire _w29490_ ;
	wire _w29489_ ;
	wire _w29488_ ;
	wire _w29487_ ;
	wire _w29486_ ;
	wire _w29485_ ;
	wire _w29484_ ;
	wire _w29483_ ;
	wire _w29482_ ;
	wire _w29481_ ;
	wire _w29480_ ;
	wire _w29479_ ;
	wire _w29478_ ;
	wire _w29477_ ;
	wire _w29476_ ;
	wire _w29475_ ;
	wire _w29474_ ;
	wire _w29473_ ;
	wire _w29472_ ;
	wire _w29471_ ;
	wire _w29470_ ;
	wire _w29469_ ;
	wire _w29468_ ;
	wire _w29467_ ;
	wire _w29466_ ;
	wire _w29465_ ;
	wire _w29464_ ;
	wire _w29463_ ;
	wire _w29462_ ;
	wire _w29461_ ;
	wire _w29460_ ;
	wire _w29459_ ;
	wire _w29458_ ;
	wire _w29457_ ;
	wire _w29456_ ;
	wire _w29455_ ;
	wire _w29454_ ;
	wire _w29453_ ;
	wire _w29452_ ;
	wire _w29451_ ;
	wire _w29450_ ;
	wire _w29449_ ;
	wire _w29448_ ;
	wire _w29447_ ;
	wire _w29446_ ;
	wire _w29445_ ;
	wire _w29444_ ;
	wire _w29443_ ;
	wire _w29442_ ;
	wire _w29441_ ;
	wire _w29440_ ;
	wire _w29439_ ;
	wire _w29438_ ;
	wire _w29437_ ;
	wire _w29436_ ;
	wire _w29435_ ;
	wire _w29434_ ;
	wire _w29433_ ;
	wire _w29432_ ;
	wire _w29431_ ;
	wire _w29430_ ;
	wire _w29429_ ;
	wire _w29428_ ;
	wire _w29427_ ;
	wire _w29426_ ;
	wire _w29425_ ;
	wire _w29424_ ;
	wire _w29423_ ;
	wire _w29422_ ;
	wire _w29421_ ;
	wire _w29420_ ;
	wire _w29419_ ;
	wire _w29418_ ;
	wire _w29417_ ;
	wire _w29416_ ;
	wire _w29415_ ;
	wire _w29414_ ;
	wire _w29413_ ;
	wire _w29412_ ;
	wire _w29411_ ;
	wire _w29410_ ;
	wire _w29409_ ;
	wire _w29408_ ;
	wire _w29407_ ;
	wire _w29406_ ;
	wire _w29405_ ;
	wire _w29404_ ;
	wire _w29403_ ;
	wire _w29402_ ;
	wire _w29401_ ;
	wire _w29400_ ;
	wire _w29399_ ;
	wire _w29398_ ;
	wire _w29397_ ;
	wire _w29396_ ;
	wire _w29395_ ;
	wire _w29394_ ;
	wire _w29393_ ;
	wire _w29392_ ;
	wire _w29391_ ;
	wire _w29390_ ;
	wire _w29389_ ;
	wire _w29388_ ;
	wire _w29387_ ;
	wire _w29386_ ;
	wire _w29385_ ;
	wire _w29384_ ;
	wire _w29383_ ;
	wire _w29382_ ;
	wire _w29381_ ;
	wire _w29380_ ;
	wire _w29379_ ;
	wire _w29378_ ;
	wire _w29377_ ;
	wire _w29376_ ;
	wire _w29375_ ;
	wire _w29374_ ;
	wire _w29373_ ;
	wire _w29372_ ;
	wire _w29371_ ;
	wire _w29370_ ;
	wire _w29369_ ;
	wire _w29368_ ;
	wire _w29367_ ;
	wire _w29366_ ;
	wire _w29365_ ;
	wire _w29364_ ;
	wire _w29363_ ;
	wire _w29362_ ;
	wire _w29361_ ;
	wire _w29360_ ;
	wire _w29359_ ;
	wire _w29358_ ;
	wire _w29357_ ;
	wire _w29356_ ;
	wire _w29355_ ;
	wire _w29354_ ;
	wire _w29353_ ;
	wire _w29352_ ;
	wire _w29351_ ;
	wire _w29350_ ;
	wire _w29349_ ;
	wire _w29348_ ;
	wire _w29347_ ;
	wire _w29346_ ;
	wire _w29345_ ;
	wire _w29344_ ;
	wire _w29343_ ;
	wire _w29342_ ;
	wire _w29341_ ;
	wire _w29340_ ;
	wire _w29339_ ;
	wire _w29338_ ;
	wire _w29337_ ;
	wire _w29336_ ;
	wire _w29335_ ;
	wire _w29334_ ;
	wire _w29333_ ;
	wire _w29332_ ;
	wire _w29331_ ;
	wire _w29330_ ;
	wire _w29329_ ;
	wire _w29328_ ;
	wire _w29327_ ;
	wire _w29326_ ;
	wire _w29325_ ;
	wire _w29324_ ;
	wire _w29323_ ;
	wire _w29322_ ;
	wire _w29321_ ;
	wire _w29320_ ;
	wire _w29319_ ;
	wire _w29318_ ;
	wire _w29317_ ;
	wire _w29316_ ;
	wire _w29315_ ;
	wire _w29314_ ;
	wire _w29313_ ;
	wire _w29312_ ;
	wire _w29311_ ;
	wire _w29310_ ;
	wire _w29309_ ;
	wire _w29308_ ;
	wire _w29307_ ;
	wire _w29306_ ;
	wire _w29305_ ;
	wire _w29304_ ;
	wire _w29303_ ;
	wire _w29302_ ;
	wire _w29301_ ;
	wire _w29300_ ;
	wire _w29299_ ;
	wire _w29298_ ;
	wire _w29297_ ;
	wire _w29296_ ;
	wire _w29295_ ;
	wire _w29294_ ;
	wire _w29293_ ;
	wire _w29292_ ;
	wire _w29291_ ;
	wire _w29290_ ;
	wire _w29289_ ;
	wire _w29288_ ;
	wire _w29287_ ;
	wire _w29286_ ;
	wire _w29285_ ;
	wire _w29284_ ;
	wire _w29283_ ;
	wire _w29282_ ;
	wire _w29281_ ;
	wire _w29280_ ;
	wire _w29279_ ;
	wire _w29278_ ;
	wire _w29277_ ;
	wire _w29276_ ;
	wire _w29275_ ;
	wire _w29274_ ;
	wire _w29273_ ;
	wire _w29272_ ;
	wire _w29271_ ;
	wire _w29270_ ;
	wire _w29269_ ;
	wire _w29268_ ;
	wire _w29267_ ;
	wire _w29266_ ;
	wire _w29265_ ;
	wire _w29264_ ;
	wire _w29263_ ;
	wire _w29262_ ;
	wire _w29261_ ;
	wire _w29260_ ;
	wire _w29259_ ;
	wire _w29258_ ;
	wire _w29257_ ;
	wire _w29256_ ;
	wire _w29255_ ;
	wire _w29254_ ;
	wire _w29253_ ;
	wire _w29252_ ;
	wire _w29251_ ;
	wire _w29250_ ;
	wire _w29249_ ;
	wire _w29248_ ;
	wire _w29247_ ;
	wire _w29246_ ;
	wire _w29245_ ;
	wire _w29244_ ;
	wire _w29243_ ;
	wire _w29242_ ;
	wire _w29241_ ;
	wire _w29240_ ;
	wire _w29239_ ;
	wire _w29238_ ;
	wire _w29237_ ;
	wire _w29236_ ;
	wire _w29235_ ;
	wire _w29234_ ;
	wire _w29233_ ;
	wire _w29232_ ;
	wire _w29231_ ;
	wire _w29230_ ;
	wire _w29229_ ;
	wire _w29228_ ;
	wire _w29227_ ;
	wire _w29226_ ;
	wire _w29225_ ;
	wire _w29224_ ;
	wire _w29223_ ;
	wire _w29222_ ;
	wire _w29221_ ;
	wire _w29220_ ;
	wire _w29219_ ;
	wire _w29218_ ;
	wire _w29217_ ;
	wire _w29216_ ;
	wire _w29215_ ;
	wire _w29214_ ;
	wire _w29213_ ;
	wire _w29212_ ;
	wire _w29211_ ;
	wire _w29210_ ;
	wire _w29209_ ;
	wire _w29208_ ;
	wire _w29207_ ;
	wire _w29206_ ;
	wire _w29205_ ;
	wire _w29204_ ;
	wire _w29203_ ;
	wire _w29202_ ;
	wire _w29201_ ;
	wire _w29200_ ;
	wire _w29199_ ;
	wire _w29198_ ;
	wire _w29197_ ;
	wire _w29196_ ;
	wire _w29195_ ;
	wire _w29194_ ;
	wire _w29193_ ;
	wire _w29192_ ;
	wire _w29191_ ;
	wire _w29190_ ;
	wire _w29189_ ;
	wire _w29188_ ;
	wire _w29187_ ;
	wire _w29186_ ;
	wire _w29185_ ;
	wire _w29184_ ;
	wire _w29183_ ;
	wire _w29182_ ;
	wire _w29181_ ;
	wire _w29180_ ;
	wire _w29179_ ;
	wire _w29178_ ;
	wire _w29177_ ;
	wire _w29176_ ;
	wire _w29175_ ;
	wire _w29174_ ;
	wire _w29173_ ;
	wire _w29172_ ;
	wire _w29171_ ;
	wire _w29170_ ;
	wire _w29169_ ;
	wire _w29168_ ;
	wire _w29167_ ;
	wire _w29166_ ;
	wire _w29165_ ;
	wire _w29164_ ;
	wire _w29163_ ;
	wire _w29162_ ;
	wire _w29161_ ;
	wire _w29160_ ;
	wire _w29159_ ;
	wire _w29158_ ;
	wire _w29157_ ;
	wire _w29156_ ;
	wire _w29155_ ;
	wire _w29154_ ;
	wire _w29153_ ;
	wire _w29152_ ;
	wire _w29151_ ;
	wire _w29150_ ;
	wire _w29149_ ;
	wire _w29148_ ;
	wire _w29147_ ;
	wire _w29146_ ;
	wire _w29145_ ;
	wire _w29144_ ;
	wire _w29143_ ;
	wire _w29142_ ;
	wire _w29141_ ;
	wire _w29140_ ;
	wire _w29139_ ;
	wire _w29138_ ;
	wire _w29137_ ;
	wire _w29136_ ;
	wire _w29135_ ;
	wire _w29134_ ;
	wire _w29133_ ;
	wire _w29132_ ;
	wire _w29131_ ;
	wire _w29130_ ;
	wire _w29129_ ;
	wire _w29128_ ;
	wire _w29127_ ;
	wire _w29126_ ;
	wire _w29125_ ;
	wire _w29124_ ;
	wire _w29123_ ;
	wire _w29122_ ;
	wire _w29121_ ;
	wire _w29120_ ;
	wire _w29119_ ;
	wire _w29118_ ;
	wire _w29117_ ;
	wire _w29116_ ;
	wire _w29115_ ;
	wire _w29114_ ;
	wire _w29113_ ;
	wire _w29112_ ;
	wire _w29111_ ;
	wire _w29110_ ;
	wire _w29109_ ;
	wire _w29108_ ;
	wire _w29107_ ;
	wire _w29106_ ;
	wire _w29105_ ;
	wire _w29104_ ;
	wire _w29103_ ;
	wire _w29102_ ;
	wire _w29101_ ;
	wire _w29100_ ;
	wire _w29099_ ;
	wire _w29098_ ;
	wire _w29097_ ;
	wire _w29096_ ;
	wire _w29095_ ;
	wire _w29094_ ;
	wire _w29093_ ;
	wire _w29092_ ;
	wire _w29091_ ;
	wire _w29090_ ;
	wire _w29089_ ;
	wire _w29088_ ;
	wire _w29087_ ;
	wire _w29086_ ;
	wire _w29085_ ;
	wire _w29084_ ;
	wire _w29083_ ;
	wire _w29082_ ;
	wire _w29081_ ;
	wire _w29080_ ;
	wire _w29079_ ;
	wire _w29078_ ;
	wire _w29077_ ;
	wire _w29076_ ;
	wire _w29075_ ;
	wire _w29074_ ;
	wire _w29073_ ;
	wire _w29072_ ;
	wire _w29071_ ;
	wire _w29070_ ;
	wire _w29069_ ;
	wire _w29068_ ;
	wire _w29067_ ;
	wire _w29066_ ;
	wire _w29065_ ;
	wire _w29064_ ;
	wire _w29063_ ;
	wire _w29062_ ;
	wire _w29061_ ;
	wire _w29060_ ;
	wire _w29059_ ;
	wire _w29058_ ;
	wire _w29057_ ;
	wire _w29056_ ;
	wire _w29055_ ;
	wire _w29054_ ;
	wire _w29053_ ;
	wire _w29052_ ;
	wire _w29051_ ;
	wire _w29050_ ;
	wire _w29049_ ;
	wire _w29048_ ;
	wire _w29047_ ;
	wire _w29046_ ;
	wire _w29045_ ;
	wire _w29044_ ;
	wire _w29043_ ;
	wire _w29042_ ;
	wire _w29041_ ;
	wire _w29040_ ;
	wire _w29039_ ;
	wire _w29038_ ;
	wire _w29037_ ;
	wire _w29036_ ;
	wire _w29035_ ;
	wire _w29034_ ;
	wire _w29033_ ;
	wire _w29032_ ;
	wire _w29031_ ;
	wire _w29030_ ;
	wire _w29029_ ;
	wire _w29028_ ;
	wire _w29027_ ;
	wire _w29026_ ;
	wire _w29025_ ;
	wire _w29024_ ;
	wire _w29023_ ;
	wire _w29022_ ;
	wire _w29021_ ;
	wire _w29020_ ;
	wire _w29019_ ;
	wire _w29018_ ;
	wire _w29017_ ;
	wire _w29016_ ;
	wire _w29015_ ;
	wire _w29014_ ;
	wire _w29013_ ;
	wire _w29012_ ;
	wire _w29011_ ;
	wire _w29010_ ;
	wire _w29009_ ;
	wire _w29008_ ;
	wire _w29007_ ;
	wire _w29006_ ;
	wire _w29005_ ;
	wire _w29004_ ;
	wire _w29003_ ;
	wire _w29002_ ;
	wire _w29001_ ;
	wire _w29000_ ;
	wire _w28999_ ;
	wire _w28998_ ;
	wire _w28997_ ;
	wire _w28996_ ;
	wire _w28995_ ;
	wire _w28994_ ;
	wire _w28993_ ;
	wire _w28992_ ;
	wire _w28991_ ;
	wire _w28990_ ;
	wire _w28989_ ;
	wire _w28988_ ;
	wire _w28987_ ;
	wire _w28986_ ;
	wire _w28985_ ;
	wire _w28984_ ;
	wire _w28983_ ;
	wire _w28982_ ;
	wire _w28981_ ;
	wire _w28980_ ;
	wire _w28979_ ;
	wire _w28978_ ;
	wire _w28977_ ;
	wire _w28976_ ;
	wire _w28975_ ;
	wire _w28974_ ;
	wire _w28973_ ;
	wire _w28972_ ;
	wire _w28971_ ;
	wire _w28970_ ;
	wire _w28969_ ;
	wire _w28968_ ;
	wire _w28967_ ;
	wire _w28966_ ;
	wire _w28965_ ;
	wire _w28964_ ;
	wire _w28963_ ;
	wire _w28962_ ;
	wire _w28961_ ;
	wire _w28960_ ;
	wire _w28959_ ;
	wire _w28958_ ;
	wire _w28957_ ;
	wire _w28956_ ;
	wire _w28955_ ;
	wire _w28954_ ;
	wire _w28953_ ;
	wire _w28952_ ;
	wire _w28951_ ;
	wire _w28950_ ;
	wire _w28949_ ;
	wire _w28948_ ;
	wire _w28947_ ;
	wire _w28946_ ;
	wire _w28945_ ;
	wire _w28944_ ;
	wire _w28943_ ;
	wire _w28942_ ;
	wire _w28941_ ;
	wire _w28940_ ;
	wire _w28939_ ;
	wire _w28938_ ;
	wire _w28937_ ;
	wire _w28936_ ;
	wire _w28935_ ;
	wire _w28934_ ;
	wire _w28933_ ;
	wire _w28932_ ;
	wire _w28931_ ;
	wire _w28930_ ;
	wire _w28929_ ;
	wire _w28928_ ;
	wire _w28927_ ;
	wire _w28926_ ;
	wire _w28925_ ;
	wire _w28924_ ;
	wire _w28923_ ;
	wire _w28922_ ;
	wire _w28921_ ;
	wire _w28920_ ;
	wire _w28919_ ;
	wire _w28918_ ;
	wire _w28917_ ;
	wire _w28916_ ;
	wire _w28915_ ;
	wire _w28914_ ;
	wire _w28913_ ;
	wire _w28912_ ;
	wire _w28911_ ;
	wire _w28910_ ;
	wire _w28909_ ;
	wire _w28908_ ;
	wire _w28907_ ;
	wire _w28906_ ;
	wire _w28905_ ;
	wire _w28904_ ;
	wire _w28903_ ;
	wire _w28902_ ;
	wire _w28901_ ;
	wire _w28900_ ;
	wire _w28899_ ;
	wire _w28898_ ;
	wire _w28897_ ;
	wire _w28896_ ;
	wire _w28895_ ;
	wire _w28894_ ;
	wire _w28893_ ;
	wire _w28892_ ;
	wire _w28891_ ;
	wire _w28890_ ;
	wire _w28889_ ;
	wire _w28888_ ;
	wire _w28887_ ;
	wire _w28886_ ;
	wire _w28885_ ;
	wire _w28884_ ;
	wire _w28883_ ;
	wire _w28882_ ;
	wire _w28881_ ;
	wire _w28880_ ;
	wire _w28879_ ;
	wire _w28878_ ;
	wire _w28877_ ;
	wire _w28876_ ;
	wire _w28875_ ;
	wire _w28874_ ;
	wire _w28873_ ;
	wire _w28872_ ;
	wire _w28871_ ;
	wire _w28870_ ;
	wire _w28869_ ;
	wire _w28868_ ;
	wire _w28867_ ;
	wire _w28866_ ;
	wire _w28865_ ;
	wire _w28864_ ;
	wire _w28863_ ;
	wire _w28862_ ;
	wire _w28861_ ;
	wire _w28860_ ;
	wire _w28859_ ;
	wire _w28858_ ;
	wire _w28857_ ;
	wire _w28856_ ;
	wire _w28855_ ;
	wire _w28854_ ;
	wire _w28853_ ;
	wire _w28852_ ;
	wire _w28851_ ;
	wire _w28850_ ;
	wire _w28849_ ;
	wire _w28848_ ;
	wire _w28847_ ;
	wire _w28846_ ;
	wire _w28845_ ;
	wire _w28844_ ;
	wire _w28843_ ;
	wire _w28842_ ;
	wire _w28841_ ;
	wire _w28840_ ;
	wire _w28839_ ;
	wire _w28838_ ;
	wire _w28837_ ;
	wire _w28836_ ;
	wire _w28835_ ;
	wire _w28834_ ;
	wire _w28833_ ;
	wire _w28832_ ;
	wire _w28831_ ;
	wire _w28830_ ;
	wire _w28829_ ;
	wire _w28828_ ;
	wire _w28827_ ;
	wire _w28826_ ;
	wire _w28825_ ;
	wire _w28824_ ;
	wire _w28823_ ;
	wire _w28822_ ;
	wire _w28821_ ;
	wire _w28820_ ;
	wire _w28819_ ;
	wire _w28818_ ;
	wire _w28817_ ;
	wire _w28816_ ;
	wire _w28815_ ;
	wire _w28814_ ;
	wire _w28813_ ;
	wire _w28812_ ;
	wire _w28811_ ;
	wire _w28810_ ;
	wire _w28809_ ;
	wire _w28808_ ;
	wire _w28807_ ;
	wire _w28806_ ;
	wire _w28805_ ;
	wire _w28804_ ;
	wire _w28803_ ;
	wire _w28802_ ;
	wire _w28801_ ;
	wire _w28800_ ;
	wire _w28799_ ;
	wire _w28798_ ;
	wire _w28797_ ;
	wire _w28796_ ;
	wire _w28795_ ;
	wire _w28794_ ;
	wire _w28793_ ;
	wire _w28792_ ;
	wire _w28791_ ;
	wire _w28790_ ;
	wire _w28789_ ;
	wire _w28788_ ;
	wire _w28787_ ;
	wire _w28786_ ;
	wire _w28785_ ;
	wire _w28784_ ;
	wire _w28783_ ;
	wire _w28782_ ;
	wire _w28781_ ;
	wire _w28780_ ;
	wire _w28779_ ;
	wire _w28778_ ;
	wire _w28777_ ;
	wire _w28776_ ;
	wire _w28775_ ;
	wire _w28774_ ;
	wire _w28773_ ;
	wire _w28772_ ;
	wire _w28771_ ;
	wire _w28770_ ;
	wire _w28769_ ;
	wire _w28768_ ;
	wire _w28767_ ;
	wire _w28766_ ;
	wire _w28765_ ;
	wire _w28764_ ;
	wire _w28763_ ;
	wire _w28762_ ;
	wire _w28761_ ;
	wire _w28760_ ;
	wire _w28759_ ;
	wire _w28758_ ;
	wire _w28757_ ;
	wire _w28756_ ;
	wire _w28755_ ;
	wire _w28754_ ;
	wire _w28753_ ;
	wire _w28752_ ;
	wire _w28751_ ;
	wire _w28750_ ;
	wire _w28749_ ;
	wire _w28748_ ;
	wire _w28747_ ;
	wire _w28746_ ;
	wire _w28745_ ;
	wire _w28744_ ;
	wire _w28743_ ;
	wire _w28742_ ;
	wire _w28741_ ;
	wire _w28740_ ;
	wire _w28739_ ;
	wire _w28738_ ;
	wire _w28737_ ;
	wire _w28736_ ;
	wire _w28735_ ;
	wire _w28734_ ;
	wire _w28733_ ;
	wire _w28732_ ;
	wire _w28731_ ;
	wire _w28730_ ;
	wire _w28729_ ;
	wire _w28728_ ;
	wire _w28727_ ;
	wire _w28726_ ;
	wire _w28725_ ;
	wire _w28724_ ;
	wire _w28723_ ;
	wire _w28722_ ;
	wire _w28721_ ;
	wire _w28720_ ;
	wire _w28719_ ;
	wire _w28718_ ;
	wire _w28717_ ;
	wire _w28716_ ;
	wire _w28715_ ;
	wire _w28714_ ;
	wire _w28713_ ;
	wire _w28712_ ;
	wire _w28711_ ;
	wire _w28710_ ;
	wire _w28709_ ;
	wire _w28708_ ;
	wire _w28707_ ;
	wire _w28706_ ;
	wire _w28705_ ;
	wire _w28704_ ;
	wire _w28703_ ;
	wire _w28702_ ;
	wire _w28701_ ;
	wire _w28700_ ;
	wire _w28699_ ;
	wire _w28698_ ;
	wire _w28697_ ;
	wire _w28696_ ;
	wire _w28695_ ;
	wire _w28694_ ;
	wire _w28693_ ;
	wire _w28692_ ;
	wire _w28691_ ;
	wire _w28690_ ;
	wire _w28689_ ;
	wire _w28688_ ;
	wire _w28687_ ;
	wire _w28686_ ;
	wire _w28685_ ;
	wire _w28684_ ;
	wire _w28683_ ;
	wire _w28682_ ;
	wire _w28681_ ;
	wire _w28680_ ;
	wire _w28679_ ;
	wire _w28678_ ;
	wire _w28677_ ;
	wire _w28676_ ;
	wire _w28675_ ;
	wire _w28674_ ;
	wire _w28673_ ;
	wire _w28672_ ;
	wire _w28671_ ;
	wire _w28670_ ;
	wire _w28669_ ;
	wire _w28668_ ;
	wire _w28667_ ;
	wire _w28666_ ;
	wire _w28665_ ;
	wire _w28664_ ;
	wire _w28663_ ;
	wire _w28662_ ;
	wire _w28661_ ;
	wire _w28660_ ;
	wire _w28659_ ;
	wire _w28658_ ;
	wire _w28657_ ;
	wire _w28656_ ;
	wire _w28655_ ;
	wire _w28654_ ;
	wire _w28653_ ;
	wire _w28652_ ;
	wire _w28651_ ;
	wire _w28650_ ;
	wire _w28649_ ;
	wire _w28648_ ;
	wire _w28647_ ;
	wire _w28646_ ;
	wire _w28645_ ;
	wire _w28644_ ;
	wire _w28643_ ;
	wire _w28642_ ;
	wire _w28641_ ;
	wire _w28640_ ;
	wire _w28639_ ;
	wire _w28638_ ;
	wire _w28637_ ;
	wire _w28636_ ;
	wire _w28635_ ;
	wire _w28634_ ;
	wire _w28633_ ;
	wire _w28632_ ;
	wire _w28631_ ;
	wire _w28630_ ;
	wire _w28629_ ;
	wire _w28628_ ;
	wire _w28627_ ;
	wire _w28626_ ;
	wire _w28625_ ;
	wire _w28624_ ;
	wire _w28623_ ;
	wire _w28622_ ;
	wire _w28621_ ;
	wire _w28620_ ;
	wire _w28619_ ;
	wire _w28618_ ;
	wire _w28617_ ;
	wire _w28616_ ;
	wire _w28615_ ;
	wire _w28614_ ;
	wire _w28613_ ;
	wire _w28612_ ;
	wire _w28611_ ;
	wire _w28610_ ;
	wire _w28609_ ;
	wire _w28608_ ;
	wire _w28607_ ;
	wire _w28606_ ;
	wire _w28605_ ;
	wire _w28604_ ;
	wire _w28603_ ;
	wire _w28602_ ;
	wire _w28601_ ;
	wire _w28600_ ;
	wire _w28599_ ;
	wire _w28598_ ;
	wire _w28597_ ;
	wire _w28596_ ;
	wire _w28595_ ;
	wire _w28594_ ;
	wire _w28593_ ;
	wire _w28592_ ;
	wire _w28591_ ;
	wire _w28590_ ;
	wire _w28589_ ;
	wire _w28588_ ;
	wire _w28587_ ;
	wire _w28586_ ;
	wire _w28585_ ;
	wire _w28584_ ;
	wire _w28583_ ;
	wire _w28582_ ;
	wire _w28581_ ;
	wire _w28580_ ;
	wire _w28579_ ;
	wire _w28578_ ;
	wire _w28577_ ;
	wire _w28576_ ;
	wire _w28575_ ;
	wire _w28574_ ;
	wire _w28573_ ;
	wire _w28572_ ;
	wire _w28571_ ;
	wire _w28570_ ;
	wire _w28569_ ;
	wire _w28568_ ;
	wire _w28567_ ;
	wire _w28566_ ;
	wire _w28565_ ;
	wire _w28564_ ;
	wire _w28563_ ;
	wire _w28562_ ;
	wire _w28561_ ;
	wire _w28560_ ;
	wire _w28559_ ;
	wire _w28558_ ;
	wire _w28557_ ;
	wire _w28556_ ;
	wire _w28555_ ;
	wire _w28554_ ;
	wire _w28553_ ;
	wire _w28552_ ;
	wire _w28551_ ;
	wire _w28550_ ;
	wire _w28549_ ;
	wire _w28548_ ;
	wire _w28547_ ;
	wire _w28546_ ;
	wire _w28545_ ;
	wire _w28544_ ;
	wire _w28543_ ;
	wire _w28542_ ;
	wire _w28541_ ;
	wire _w28540_ ;
	wire _w28539_ ;
	wire _w28538_ ;
	wire _w28537_ ;
	wire _w28536_ ;
	wire _w28535_ ;
	wire _w28534_ ;
	wire _w28533_ ;
	wire _w28532_ ;
	wire _w28531_ ;
	wire _w28530_ ;
	wire _w28529_ ;
	wire _w28528_ ;
	wire _w28527_ ;
	wire _w28526_ ;
	wire _w28525_ ;
	wire _w28524_ ;
	wire _w28523_ ;
	wire _w28522_ ;
	wire _w28521_ ;
	wire _w28520_ ;
	wire _w28519_ ;
	wire _w28518_ ;
	wire _w28517_ ;
	wire _w28516_ ;
	wire _w28515_ ;
	wire _w28514_ ;
	wire _w28513_ ;
	wire _w28512_ ;
	wire _w28511_ ;
	wire _w28510_ ;
	wire _w28509_ ;
	wire _w28508_ ;
	wire _w28507_ ;
	wire _w28506_ ;
	wire _w28505_ ;
	wire _w28504_ ;
	wire _w28503_ ;
	wire _w28502_ ;
	wire _w28501_ ;
	wire _w28500_ ;
	wire _w28499_ ;
	wire _w28498_ ;
	wire _w28497_ ;
	wire _w28496_ ;
	wire _w28495_ ;
	wire _w28494_ ;
	wire _w28493_ ;
	wire _w28492_ ;
	wire _w28491_ ;
	wire _w28490_ ;
	wire _w28489_ ;
	wire _w28488_ ;
	wire _w28487_ ;
	wire _w28486_ ;
	wire _w28485_ ;
	wire _w28484_ ;
	wire _w28483_ ;
	wire _w28482_ ;
	wire _w28481_ ;
	wire _w28480_ ;
	wire _w28479_ ;
	wire _w28478_ ;
	wire _w28477_ ;
	wire _w28476_ ;
	wire _w28475_ ;
	wire _w28474_ ;
	wire _w28473_ ;
	wire _w28472_ ;
	wire _w28471_ ;
	wire _w28470_ ;
	wire _w28469_ ;
	wire _w28468_ ;
	wire _w28467_ ;
	wire _w28466_ ;
	wire _w28465_ ;
	wire _w28464_ ;
	wire _w28463_ ;
	wire _w28462_ ;
	wire _w28461_ ;
	wire _w28460_ ;
	wire _w28459_ ;
	wire _w28458_ ;
	wire _w28457_ ;
	wire _w28456_ ;
	wire _w28455_ ;
	wire _w28454_ ;
	wire _w28453_ ;
	wire _w28452_ ;
	wire _w28451_ ;
	wire _w28450_ ;
	wire _w28449_ ;
	wire _w28448_ ;
	wire _w28447_ ;
	wire _w28446_ ;
	wire _w28445_ ;
	wire _w28444_ ;
	wire _w28443_ ;
	wire _w28442_ ;
	wire _w28441_ ;
	wire _w28440_ ;
	wire _w28439_ ;
	wire _w28438_ ;
	wire _w28437_ ;
	wire _w28436_ ;
	wire _w28435_ ;
	wire _w28434_ ;
	wire _w28433_ ;
	wire _w28432_ ;
	wire _w28431_ ;
	wire _w28430_ ;
	wire _w28429_ ;
	wire _w28428_ ;
	wire _w28427_ ;
	wire _w28426_ ;
	wire _w28425_ ;
	wire _w28424_ ;
	wire _w28423_ ;
	wire _w28422_ ;
	wire _w28421_ ;
	wire _w28420_ ;
	wire _w28419_ ;
	wire _w28418_ ;
	wire _w28417_ ;
	wire _w28416_ ;
	wire _w28415_ ;
	wire _w28414_ ;
	wire _w28413_ ;
	wire _w28412_ ;
	wire _w28411_ ;
	wire _w28410_ ;
	wire _w28409_ ;
	wire _w28408_ ;
	wire _w28407_ ;
	wire _w28406_ ;
	wire _w28405_ ;
	wire _w28404_ ;
	wire _w28403_ ;
	wire _w28402_ ;
	wire _w28401_ ;
	wire _w28400_ ;
	wire _w28399_ ;
	wire _w28398_ ;
	wire _w28397_ ;
	wire _w28396_ ;
	wire _w28395_ ;
	wire _w28394_ ;
	wire _w28393_ ;
	wire _w28392_ ;
	wire _w28391_ ;
	wire _w28390_ ;
	wire _w28389_ ;
	wire _w28388_ ;
	wire _w28387_ ;
	wire _w28386_ ;
	wire _w28385_ ;
	wire _w28384_ ;
	wire _w28383_ ;
	wire _w28382_ ;
	wire _w28381_ ;
	wire _w28380_ ;
	wire _w28379_ ;
	wire _w28378_ ;
	wire _w28377_ ;
	wire _w28376_ ;
	wire _w28375_ ;
	wire _w28374_ ;
	wire _w28373_ ;
	wire _w28372_ ;
	wire _w28371_ ;
	wire _w28370_ ;
	wire _w28369_ ;
	wire _w28368_ ;
	wire _w28367_ ;
	wire _w28366_ ;
	wire _w28365_ ;
	wire _w28364_ ;
	wire _w28363_ ;
	wire _w28362_ ;
	wire _w28361_ ;
	wire _w28360_ ;
	wire _w28359_ ;
	wire _w28358_ ;
	wire _w28357_ ;
	wire _w28356_ ;
	wire _w28355_ ;
	wire _w28354_ ;
	wire _w28353_ ;
	wire _w28352_ ;
	wire _w28351_ ;
	wire _w28350_ ;
	wire _w28349_ ;
	wire _w28348_ ;
	wire _w28347_ ;
	wire _w28346_ ;
	wire _w28345_ ;
	wire _w28344_ ;
	wire _w28343_ ;
	wire _w28342_ ;
	wire _w28341_ ;
	wire _w28340_ ;
	wire _w28339_ ;
	wire _w28338_ ;
	wire _w28337_ ;
	wire _w28336_ ;
	wire _w28335_ ;
	wire _w28334_ ;
	wire _w28333_ ;
	wire _w28332_ ;
	wire _w28331_ ;
	wire _w28330_ ;
	wire _w28329_ ;
	wire _w28328_ ;
	wire _w28327_ ;
	wire _w28326_ ;
	wire _w28325_ ;
	wire _w28324_ ;
	wire _w28323_ ;
	wire _w28322_ ;
	wire _w28321_ ;
	wire _w28320_ ;
	wire _w28319_ ;
	wire _w28318_ ;
	wire _w28317_ ;
	wire _w28316_ ;
	wire _w28315_ ;
	wire _w28314_ ;
	wire _w28313_ ;
	wire _w28312_ ;
	wire _w28311_ ;
	wire _w28310_ ;
	wire _w28309_ ;
	wire _w28308_ ;
	wire _w28307_ ;
	wire _w28306_ ;
	wire _w28305_ ;
	wire _w28304_ ;
	wire _w28303_ ;
	wire _w28302_ ;
	wire _w28301_ ;
	wire _w28300_ ;
	wire _w28299_ ;
	wire _w28298_ ;
	wire _w28297_ ;
	wire _w28296_ ;
	wire _w28295_ ;
	wire _w28294_ ;
	wire _w28293_ ;
	wire _w28292_ ;
	wire _w28291_ ;
	wire _w28290_ ;
	wire _w28289_ ;
	wire _w28288_ ;
	wire _w28287_ ;
	wire _w28286_ ;
	wire _w28285_ ;
	wire _w28284_ ;
	wire _w28283_ ;
	wire _w28282_ ;
	wire _w28281_ ;
	wire _w28280_ ;
	wire _w28279_ ;
	wire _w28278_ ;
	wire _w28277_ ;
	wire _w28276_ ;
	wire _w28275_ ;
	wire _w28274_ ;
	wire _w28273_ ;
	wire _w28272_ ;
	wire _w28271_ ;
	wire _w28270_ ;
	wire _w28269_ ;
	wire _w28268_ ;
	wire _w28267_ ;
	wire _w28266_ ;
	wire _w28265_ ;
	wire _w28264_ ;
	wire _w28263_ ;
	wire _w28262_ ;
	wire _w28261_ ;
	wire _w28260_ ;
	wire _w28259_ ;
	wire _w28258_ ;
	wire _w28257_ ;
	wire _w28256_ ;
	wire _w28255_ ;
	wire _w28254_ ;
	wire _w28253_ ;
	wire _w28252_ ;
	wire _w28251_ ;
	wire _w28250_ ;
	wire _w28249_ ;
	wire _w28248_ ;
	wire _w28247_ ;
	wire _w28246_ ;
	wire _w28245_ ;
	wire _w28244_ ;
	wire _w28243_ ;
	wire _w28242_ ;
	wire _w28241_ ;
	wire _w28240_ ;
	wire _w28239_ ;
	wire _w28238_ ;
	wire _w28237_ ;
	wire _w28236_ ;
	wire _w28235_ ;
	wire _w28234_ ;
	wire _w28233_ ;
	wire _w28232_ ;
	wire _w28231_ ;
	wire _w28230_ ;
	wire _w28229_ ;
	wire _w28228_ ;
	wire _w28227_ ;
	wire _w28226_ ;
	wire _w28225_ ;
	wire _w28224_ ;
	wire _w28223_ ;
	wire _w28222_ ;
	wire _w28221_ ;
	wire _w28220_ ;
	wire _w28219_ ;
	wire _w28218_ ;
	wire _w28217_ ;
	wire _w28216_ ;
	wire _w28215_ ;
	wire _w28214_ ;
	wire _w28213_ ;
	wire _w28212_ ;
	wire _w28211_ ;
	wire _w28210_ ;
	wire _w28209_ ;
	wire _w28208_ ;
	wire _w28207_ ;
	wire _w28206_ ;
	wire _w28205_ ;
	wire _w28204_ ;
	wire _w28203_ ;
	wire _w28202_ ;
	wire _w28201_ ;
	wire _w28200_ ;
	wire _w28199_ ;
	wire _w28198_ ;
	wire _w28197_ ;
	wire _w28196_ ;
	wire _w28195_ ;
	wire _w28194_ ;
	wire _w28193_ ;
	wire _w28192_ ;
	wire _w28191_ ;
	wire _w28190_ ;
	wire _w28189_ ;
	wire _w28188_ ;
	wire _w28187_ ;
	wire _w28186_ ;
	wire _w28185_ ;
	wire _w28184_ ;
	wire _w28183_ ;
	wire _w28182_ ;
	wire _w28181_ ;
	wire _w28180_ ;
	wire _w28179_ ;
	wire _w28178_ ;
	wire _w28177_ ;
	wire _w28176_ ;
	wire _w28175_ ;
	wire _w28174_ ;
	wire _w28173_ ;
	wire _w28172_ ;
	wire _w28171_ ;
	wire _w28170_ ;
	wire _w28169_ ;
	wire _w28168_ ;
	wire _w28167_ ;
	wire _w28166_ ;
	wire _w28165_ ;
	wire _w28164_ ;
	wire _w28163_ ;
	wire _w28162_ ;
	wire _w28161_ ;
	wire _w28160_ ;
	wire _w28159_ ;
	wire _w28158_ ;
	wire _w28157_ ;
	wire _w28156_ ;
	wire _w28155_ ;
	wire _w28154_ ;
	wire _w28153_ ;
	wire _w28152_ ;
	wire _w28151_ ;
	wire _w28150_ ;
	wire _w28149_ ;
	wire _w28148_ ;
	wire _w28147_ ;
	wire _w28146_ ;
	wire _w28145_ ;
	wire _w28144_ ;
	wire _w28143_ ;
	wire _w28142_ ;
	wire _w28141_ ;
	wire _w28140_ ;
	wire _w28139_ ;
	wire _w28138_ ;
	wire _w28137_ ;
	wire _w28136_ ;
	wire _w28135_ ;
	wire _w28134_ ;
	wire _w28133_ ;
	wire _w28132_ ;
	wire _w28131_ ;
	wire _w28130_ ;
	wire _w28129_ ;
	wire _w28128_ ;
	wire _w28127_ ;
	wire _w28126_ ;
	wire _w28125_ ;
	wire _w28124_ ;
	wire _w28123_ ;
	wire _w28122_ ;
	wire _w28121_ ;
	wire _w28120_ ;
	wire _w28119_ ;
	wire _w28118_ ;
	wire _w28117_ ;
	wire _w28116_ ;
	wire _w28115_ ;
	wire _w28114_ ;
	wire _w28113_ ;
	wire _w28112_ ;
	wire _w28111_ ;
	wire _w28110_ ;
	wire _w28109_ ;
	wire _w28108_ ;
	wire _w28107_ ;
	wire _w28106_ ;
	wire _w28105_ ;
	wire _w28104_ ;
	wire _w28103_ ;
	wire _w28102_ ;
	wire _w28101_ ;
	wire _w28100_ ;
	wire _w28099_ ;
	wire _w28098_ ;
	wire _w28097_ ;
	wire _w28096_ ;
	wire _w28095_ ;
	wire _w28094_ ;
	wire _w28093_ ;
	wire _w28092_ ;
	wire _w28091_ ;
	wire _w28090_ ;
	wire _w28089_ ;
	wire _w28088_ ;
	wire _w28087_ ;
	wire _w28086_ ;
	wire _w28085_ ;
	wire _w28084_ ;
	wire _w28083_ ;
	wire _w28082_ ;
	wire _w28081_ ;
	wire _w28080_ ;
	wire _w28079_ ;
	wire _w28078_ ;
	wire _w28077_ ;
	wire _w28076_ ;
	wire _w28075_ ;
	wire _w28074_ ;
	wire _w28073_ ;
	wire _w28072_ ;
	wire _w28071_ ;
	wire _w28070_ ;
	wire _w28069_ ;
	wire _w28068_ ;
	wire _w28067_ ;
	wire _w28066_ ;
	wire _w28065_ ;
	wire _w28064_ ;
	wire _w28063_ ;
	wire _w28062_ ;
	wire _w28061_ ;
	wire _w28060_ ;
	wire _w28059_ ;
	wire _w28058_ ;
	wire _w28057_ ;
	wire _w28056_ ;
	wire _w28055_ ;
	wire _w28054_ ;
	wire _w28053_ ;
	wire _w28052_ ;
	wire _w28051_ ;
	wire _w28050_ ;
	wire _w28049_ ;
	wire _w28048_ ;
	wire _w28047_ ;
	wire _w28046_ ;
	wire _w28045_ ;
	wire _w28044_ ;
	wire _w28043_ ;
	wire _w28042_ ;
	wire _w28041_ ;
	wire _w28040_ ;
	wire _w28039_ ;
	wire _w28038_ ;
	wire _w28037_ ;
	wire _w28036_ ;
	wire _w28035_ ;
	wire _w28034_ ;
	wire _w28033_ ;
	wire _w28032_ ;
	wire _w28031_ ;
	wire _w28030_ ;
	wire _w28029_ ;
	wire _w28028_ ;
	wire _w28027_ ;
	wire _w28026_ ;
	wire _w28025_ ;
	wire _w28024_ ;
	wire _w28023_ ;
	wire _w28022_ ;
	wire _w28021_ ;
	wire _w28020_ ;
	wire _w28019_ ;
	wire _w28018_ ;
	wire _w28017_ ;
	wire _w28016_ ;
	wire _w28015_ ;
	wire _w28014_ ;
	wire _w28013_ ;
	wire _w28012_ ;
	wire _w28011_ ;
	wire _w28010_ ;
	wire _w28009_ ;
	wire _w28008_ ;
	wire _w28007_ ;
	wire _w28006_ ;
	wire _w28005_ ;
	wire _w28004_ ;
	wire _w28003_ ;
	wire _w28002_ ;
	wire _w28001_ ;
	wire _w28000_ ;
	wire _w27999_ ;
	wire _w27998_ ;
	wire _w27997_ ;
	wire _w27996_ ;
	wire _w27995_ ;
	wire _w27994_ ;
	wire _w27993_ ;
	wire _w27992_ ;
	wire _w27991_ ;
	wire _w27990_ ;
	wire _w27989_ ;
	wire _w27988_ ;
	wire _w27987_ ;
	wire _w27986_ ;
	wire _w27985_ ;
	wire _w27984_ ;
	wire _w27983_ ;
	wire _w27982_ ;
	wire _w27981_ ;
	wire _w27980_ ;
	wire _w27979_ ;
	wire _w27978_ ;
	wire _w27977_ ;
	wire _w27976_ ;
	wire _w27975_ ;
	wire _w27974_ ;
	wire _w27973_ ;
	wire _w27972_ ;
	wire _w27971_ ;
	wire _w27970_ ;
	wire _w27969_ ;
	wire _w27968_ ;
	wire _w27967_ ;
	wire _w27966_ ;
	wire _w27965_ ;
	wire _w27964_ ;
	wire _w27963_ ;
	wire _w27962_ ;
	wire _w27961_ ;
	wire _w27960_ ;
	wire _w27959_ ;
	wire _w27958_ ;
	wire _w27957_ ;
	wire _w27956_ ;
	wire _w27955_ ;
	wire _w27954_ ;
	wire _w27953_ ;
	wire _w27952_ ;
	wire _w27951_ ;
	wire _w27950_ ;
	wire _w27949_ ;
	wire _w27948_ ;
	wire _w27947_ ;
	wire _w27946_ ;
	wire _w27945_ ;
	wire _w27944_ ;
	wire _w27943_ ;
	wire _w27942_ ;
	wire _w27941_ ;
	wire _w27940_ ;
	wire _w27939_ ;
	wire _w27938_ ;
	wire _w27937_ ;
	wire _w27936_ ;
	wire _w27935_ ;
	wire _w27934_ ;
	wire _w27933_ ;
	wire _w27932_ ;
	wire _w27931_ ;
	wire _w27930_ ;
	wire _w27929_ ;
	wire _w27928_ ;
	wire _w27927_ ;
	wire _w27926_ ;
	wire _w27925_ ;
	wire _w27924_ ;
	wire _w27923_ ;
	wire _w27922_ ;
	wire _w27921_ ;
	wire _w27920_ ;
	wire _w27919_ ;
	wire _w27918_ ;
	wire _w27917_ ;
	wire _w27916_ ;
	wire _w27915_ ;
	wire _w27914_ ;
	wire _w27913_ ;
	wire _w27912_ ;
	wire _w27911_ ;
	wire _w27910_ ;
	wire _w27909_ ;
	wire _w27908_ ;
	wire _w27907_ ;
	wire _w27906_ ;
	wire _w27905_ ;
	wire _w27904_ ;
	wire _w27903_ ;
	wire _w27902_ ;
	wire _w27901_ ;
	wire _w27900_ ;
	wire _w27899_ ;
	wire _w27898_ ;
	wire _w27897_ ;
	wire _w27896_ ;
	wire _w27895_ ;
	wire _w27894_ ;
	wire _w27893_ ;
	wire _w27892_ ;
	wire _w27891_ ;
	wire _w27890_ ;
	wire _w27889_ ;
	wire _w27888_ ;
	wire _w27887_ ;
	wire _w27886_ ;
	wire _w27885_ ;
	wire _w27884_ ;
	wire _w27883_ ;
	wire _w27882_ ;
	wire _w27881_ ;
	wire _w27880_ ;
	wire _w27879_ ;
	wire _w27878_ ;
	wire _w27877_ ;
	wire _w27876_ ;
	wire _w27875_ ;
	wire _w27874_ ;
	wire _w27873_ ;
	wire _w27872_ ;
	wire _w27871_ ;
	wire _w27870_ ;
	wire _w27869_ ;
	wire _w27868_ ;
	wire _w27867_ ;
	wire _w27866_ ;
	wire _w27865_ ;
	wire _w27864_ ;
	wire _w27863_ ;
	wire _w27862_ ;
	wire _w27861_ ;
	wire _w27860_ ;
	wire _w27859_ ;
	wire _w27858_ ;
	wire _w27857_ ;
	wire _w27856_ ;
	wire _w27855_ ;
	wire _w27854_ ;
	wire _w27853_ ;
	wire _w27852_ ;
	wire _w27851_ ;
	wire _w27850_ ;
	wire _w27849_ ;
	wire _w27848_ ;
	wire _w27847_ ;
	wire _w27846_ ;
	wire _w27845_ ;
	wire _w27844_ ;
	wire _w27843_ ;
	wire _w27842_ ;
	wire _w27841_ ;
	wire _w27840_ ;
	wire _w27839_ ;
	wire _w27838_ ;
	wire _w27837_ ;
	wire _w27836_ ;
	wire _w27835_ ;
	wire _w27834_ ;
	wire _w27833_ ;
	wire _w27832_ ;
	wire _w27831_ ;
	wire _w27830_ ;
	wire _w27829_ ;
	wire _w27828_ ;
	wire _w27827_ ;
	wire _w27826_ ;
	wire _w27825_ ;
	wire _w27824_ ;
	wire _w27823_ ;
	wire _w27822_ ;
	wire _w27821_ ;
	wire _w27820_ ;
	wire _w27819_ ;
	wire _w27818_ ;
	wire _w27817_ ;
	wire _w27816_ ;
	wire _w27815_ ;
	wire _w27814_ ;
	wire _w27813_ ;
	wire _w27812_ ;
	wire _w27811_ ;
	wire _w27810_ ;
	wire _w27809_ ;
	wire _w27808_ ;
	wire _w27807_ ;
	wire _w27806_ ;
	wire _w27805_ ;
	wire _w27804_ ;
	wire _w27803_ ;
	wire _w27802_ ;
	wire _w27801_ ;
	wire _w27800_ ;
	wire _w27799_ ;
	wire _w27798_ ;
	wire _w27797_ ;
	wire _w27796_ ;
	wire _w27795_ ;
	wire _w27794_ ;
	wire _w27793_ ;
	wire _w27792_ ;
	wire _w27791_ ;
	wire _w27790_ ;
	wire _w27789_ ;
	wire _w27788_ ;
	wire _w27787_ ;
	wire _w27786_ ;
	wire _w27785_ ;
	wire _w27784_ ;
	wire _w27783_ ;
	wire _w27782_ ;
	wire _w27781_ ;
	wire _w27780_ ;
	wire _w27779_ ;
	wire _w27778_ ;
	wire _w27777_ ;
	wire _w27776_ ;
	wire _w27775_ ;
	wire _w27774_ ;
	wire _w27773_ ;
	wire _w27772_ ;
	wire _w27771_ ;
	wire _w27770_ ;
	wire _w27769_ ;
	wire _w27768_ ;
	wire _w27767_ ;
	wire _w27766_ ;
	wire _w27765_ ;
	wire _w27764_ ;
	wire _w27763_ ;
	wire _w27762_ ;
	wire _w27761_ ;
	wire _w27760_ ;
	wire _w27759_ ;
	wire _w27758_ ;
	wire _w27757_ ;
	wire _w27756_ ;
	wire _w27755_ ;
	wire _w27754_ ;
	wire _w27753_ ;
	wire _w27752_ ;
	wire _w27751_ ;
	wire _w27750_ ;
	wire _w27749_ ;
	wire _w27748_ ;
	wire _w27747_ ;
	wire _w27746_ ;
	wire _w27745_ ;
	wire _w27744_ ;
	wire _w27743_ ;
	wire _w27742_ ;
	wire _w27741_ ;
	wire _w27740_ ;
	wire _w27739_ ;
	wire _w27738_ ;
	wire _w27737_ ;
	wire _w27736_ ;
	wire _w27735_ ;
	wire _w27734_ ;
	wire _w27733_ ;
	wire _w27732_ ;
	wire _w27731_ ;
	wire _w27730_ ;
	wire _w27729_ ;
	wire _w27728_ ;
	wire _w27727_ ;
	wire _w27726_ ;
	wire _w27725_ ;
	wire _w27724_ ;
	wire _w27723_ ;
	wire _w27722_ ;
	wire _w27721_ ;
	wire _w27720_ ;
	wire _w27719_ ;
	wire _w27718_ ;
	wire _w27717_ ;
	wire _w27716_ ;
	wire _w27715_ ;
	wire _w27714_ ;
	wire _w27713_ ;
	wire _w27712_ ;
	wire _w27711_ ;
	wire _w27710_ ;
	wire _w27709_ ;
	wire _w27708_ ;
	wire _w27707_ ;
	wire _w27706_ ;
	wire _w27705_ ;
	wire _w27704_ ;
	wire _w27703_ ;
	wire _w27702_ ;
	wire _w27701_ ;
	wire _w27700_ ;
	wire _w27699_ ;
	wire _w27698_ ;
	wire _w27697_ ;
	wire _w27696_ ;
	wire _w27695_ ;
	wire _w27694_ ;
	wire _w27693_ ;
	wire _w27692_ ;
	wire _w27691_ ;
	wire _w27690_ ;
	wire _w27689_ ;
	wire _w27688_ ;
	wire _w27687_ ;
	wire _w27686_ ;
	wire _w27685_ ;
	wire _w27684_ ;
	wire _w27683_ ;
	wire _w27682_ ;
	wire _w27681_ ;
	wire _w27680_ ;
	wire _w27679_ ;
	wire _w27678_ ;
	wire _w27677_ ;
	wire _w27676_ ;
	wire _w27675_ ;
	wire _w27674_ ;
	wire _w27673_ ;
	wire _w27672_ ;
	wire _w27671_ ;
	wire _w27670_ ;
	wire _w27669_ ;
	wire _w27668_ ;
	wire _w27667_ ;
	wire _w27666_ ;
	wire _w27665_ ;
	wire _w27664_ ;
	wire _w27663_ ;
	wire _w27662_ ;
	wire _w27661_ ;
	wire _w27660_ ;
	wire _w27659_ ;
	wire _w27658_ ;
	wire _w27657_ ;
	wire _w27656_ ;
	wire _w27655_ ;
	wire _w27654_ ;
	wire _w27653_ ;
	wire _w27652_ ;
	wire _w27651_ ;
	wire _w27650_ ;
	wire _w27649_ ;
	wire _w27648_ ;
	wire _w27647_ ;
	wire _w27646_ ;
	wire _w27645_ ;
	wire _w27644_ ;
	wire _w27643_ ;
	wire _w27642_ ;
	wire _w27641_ ;
	wire _w27640_ ;
	wire _w27639_ ;
	wire _w27638_ ;
	wire _w27637_ ;
	wire _w27636_ ;
	wire _w27635_ ;
	wire _w27634_ ;
	wire _w27633_ ;
	wire _w27632_ ;
	wire _w27631_ ;
	wire _w27630_ ;
	wire _w27629_ ;
	wire _w27628_ ;
	wire _w27627_ ;
	wire _w27626_ ;
	wire _w27625_ ;
	wire _w27624_ ;
	wire _w27623_ ;
	wire _w27622_ ;
	wire _w27621_ ;
	wire _w27620_ ;
	wire _w27619_ ;
	wire _w27618_ ;
	wire _w27617_ ;
	wire _w27616_ ;
	wire _w27615_ ;
	wire _w27614_ ;
	wire _w27613_ ;
	wire _w27612_ ;
	wire _w27611_ ;
	wire _w27610_ ;
	wire _w27609_ ;
	wire _w27608_ ;
	wire _w27607_ ;
	wire _w27606_ ;
	wire _w27605_ ;
	wire _w27604_ ;
	wire _w27603_ ;
	wire _w27602_ ;
	wire _w27601_ ;
	wire _w27600_ ;
	wire _w27599_ ;
	wire _w27598_ ;
	wire _w27597_ ;
	wire _w27596_ ;
	wire _w27595_ ;
	wire _w27594_ ;
	wire _w27593_ ;
	wire _w27592_ ;
	wire _w27591_ ;
	wire _w27590_ ;
	wire _w27589_ ;
	wire _w27588_ ;
	wire _w27587_ ;
	wire _w27586_ ;
	wire _w27585_ ;
	wire _w27584_ ;
	wire _w27583_ ;
	wire _w27582_ ;
	wire _w27581_ ;
	wire _w27580_ ;
	wire _w27579_ ;
	wire _w27578_ ;
	wire _w27577_ ;
	wire _w27576_ ;
	wire _w27575_ ;
	wire _w27574_ ;
	wire _w27573_ ;
	wire _w27572_ ;
	wire _w27571_ ;
	wire _w27570_ ;
	wire _w27569_ ;
	wire _w27568_ ;
	wire _w27567_ ;
	wire _w27566_ ;
	wire _w27565_ ;
	wire _w27564_ ;
	wire _w27563_ ;
	wire _w27562_ ;
	wire _w27561_ ;
	wire _w27560_ ;
	wire _w27559_ ;
	wire _w27558_ ;
	wire _w27557_ ;
	wire _w27556_ ;
	wire _w27555_ ;
	wire _w27554_ ;
	wire _w27553_ ;
	wire _w27552_ ;
	wire _w27551_ ;
	wire _w27550_ ;
	wire _w27549_ ;
	wire _w27548_ ;
	wire _w27547_ ;
	wire _w27546_ ;
	wire _w27545_ ;
	wire _w27544_ ;
	wire _w27543_ ;
	wire _w27542_ ;
	wire _w27541_ ;
	wire _w27540_ ;
	wire _w27539_ ;
	wire _w27538_ ;
	wire _w27537_ ;
	wire _w27536_ ;
	wire _w27535_ ;
	wire _w27534_ ;
	wire _w27533_ ;
	wire _w27532_ ;
	wire _w27531_ ;
	wire _w27530_ ;
	wire _w27529_ ;
	wire _w27528_ ;
	wire _w27527_ ;
	wire _w27526_ ;
	wire _w27525_ ;
	wire _w27524_ ;
	wire _w27523_ ;
	wire _w27522_ ;
	wire _w27521_ ;
	wire _w27520_ ;
	wire _w27519_ ;
	wire _w27518_ ;
	wire _w27517_ ;
	wire _w27516_ ;
	wire _w27515_ ;
	wire _w27514_ ;
	wire _w27513_ ;
	wire _w27512_ ;
	wire _w27511_ ;
	wire _w27510_ ;
	wire _w27509_ ;
	wire _w27508_ ;
	wire _w27507_ ;
	wire _w27506_ ;
	wire _w27505_ ;
	wire _w27504_ ;
	wire _w27503_ ;
	wire _w27502_ ;
	wire _w27501_ ;
	wire _w27500_ ;
	wire _w27499_ ;
	wire _w27498_ ;
	wire _w27497_ ;
	wire _w27496_ ;
	wire _w27495_ ;
	wire _w27494_ ;
	wire _w27493_ ;
	wire _w27492_ ;
	wire _w27491_ ;
	wire _w27490_ ;
	wire _w27489_ ;
	wire _w27488_ ;
	wire _w27487_ ;
	wire _w27486_ ;
	wire _w27485_ ;
	wire _w27484_ ;
	wire _w27483_ ;
	wire _w27482_ ;
	wire _w27481_ ;
	wire _w27480_ ;
	wire _w27479_ ;
	wire _w27478_ ;
	wire _w27477_ ;
	wire _w27476_ ;
	wire _w27475_ ;
	wire _w27474_ ;
	wire _w27473_ ;
	wire _w27472_ ;
	wire _w27471_ ;
	wire _w27470_ ;
	wire _w27469_ ;
	wire _w27468_ ;
	wire _w27467_ ;
	wire _w27466_ ;
	wire _w27465_ ;
	wire _w27464_ ;
	wire _w27463_ ;
	wire _w27462_ ;
	wire _w27461_ ;
	wire _w27460_ ;
	wire _w27459_ ;
	wire _w27458_ ;
	wire _w27457_ ;
	wire _w27456_ ;
	wire _w27455_ ;
	wire _w27454_ ;
	wire _w27453_ ;
	wire _w27452_ ;
	wire _w27451_ ;
	wire _w27450_ ;
	wire _w27449_ ;
	wire _w27448_ ;
	wire _w27447_ ;
	wire _w27446_ ;
	wire _w27445_ ;
	wire _w27444_ ;
	wire _w27443_ ;
	wire _w27442_ ;
	wire _w27441_ ;
	wire _w27440_ ;
	wire _w27439_ ;
	wire _w27438_ ;
	wire _w27437_ ;
	wire _w27436_ ;
	wire _w27435_ ;
	wire _w27434_ ;
	wire _w27433_ ;
	wire _w27432_ ;
	wire _w27431_ ;
	wire _w27430_ ;
	wire _w27429_ ;
	wire _w27428_ ;
	wire _w27427_ ;
	wire _w27426_ ;
	wire _w27425_ ;
	wire _w27424_ ;
	wire _w27423_ ;
	wire _w27422_ ;
	wire _w27421_ ;
	wire _w27420_ ;
	wire _w27419_ ;
	wire _w27418_ ;
	wire _w27417_ ;
	wire _w27416_ ;
	wire _w27415_ ;
	wire _w27414_ ;
	wire _w27413_ ;
	wire _w27412_ ;
	wire _w27411_ ;
	wire _w27410_ ;
	wire _w27409_ ;
	wire _w27408_ ;
	wire _w27407_ ;
	wire _w27406_ ;
	wire _w27405_ ;
	wire _w27404_ ;
	wire _w27403_ ;
	wire _w27402_ ;
	wire _w27401_ ;
	wire _w27400_ ;
	wire _w27399_ ;
	wire _w27398_ ;
	wire _w27397_ ;
	wire _w27396_ ;
	wire _w27395_ ;
	wire _w27394_ ;
	wire _w27393_ ;
	wire _w27392_ ;
	wire _w27391_ ;
	wire _w27390_ ;
	wire _w27389_ ;
	wire _w27388_ ;
	wire _w27387_ ;
	wire _w27386_ ;
	wire _w27385_ ;
	wire _w27384_ ;
	wire _w27383_ ;
	wire _w27382_ ;
	wire _w27381_ ;
	wire _w27380_ ;
	wire _w27379_ ;
	wire _w27378_ ;
	wire _w27377_ ;
	wire _w27376_ ;
	wire _w27375_ ;
	wire _w27374_ ;
	wire _w27373_ ;
	wire _w27372_ ;
	wire _w27371_ ;
	wire _w27370_ ;
	wire _w27369_ ;
	wire _w27368_ ;
	wire _w27367_ ;
	wire _w27366_ ;
	wire _w27365_ ;
	wire _w27364_ ;
	wire _w27363_ ;
	wire _w27362_ ;
	wire _w27361_ ;
	wire _w27360_ ;
	wire _w27359_ ;
	wire _w27358_ ;
	wire _w27357_ ;
	wire _w27356_ ;
	wire _w27355_ ;
	wire _w27354_ ;
	wire _w27353_ ;
	wire _w27352_ ;
	wire _w27351_ ;
	wire _w27350_ ;
	wire _w27349_ ;
	wire _w27348_ ;
	wire _w27347_ ;
	wire _w27346_ ;
	wire _w27345_ ;
	wire _w27344_ ;
	wire _w27343_ ;
	wire _w27342_ ;
	wire _w27341_ ;
	wire _w27340_ ;
	wire _w27339_ ;
	wire _w27338_ ;
	wire _w27337_ ;
	wire _w27336_ ;
	wire _w27335_ ;
	wire _w27334_ ;
	wire _w27333_ ;
	wire _w27332_ ;
	wire _w27331_ ;
	wire _w27330_ ;
	wire _w27329_ ;
	wire _w27328_ ;
	wire _w27327_ ;
	wire _w27326_ ;
	wire _w27325_ ;
	wire _w27324_ ;
	wire _w27323_ ;
	wire _w27322_ ;
	wire _w27321_ ;
	wire _w27320_ ;
	wire _w27319_ ;
	wire _w27318_ ;
	wire _w27317_ ;
	wire _w27316_ ;
	wire _w27315_ ;
	wire _w27314_ ;
	wire _w27313_ ;
	wire _w27312_ ;
	wire _w27311_ ;
	wire _w27310_ ;
	wire _w27309_ ;
	wire _w27308_ ;
	wire _w27307_ ;
	wire _w27306_ ;
	wire _w27305_ ;
	wire _w27304_ ;
	wire _w27303_ ;
	wire _w27302_ ;
	wire _w27301_ ;
	wire _w27300_ ;
	wire _w27299_ ;
	wire _w27298_ ;
	wire _w27297_ ;
	wire _w27296_ ;
	wire _w27295_ ;
	wire _w27294_ ;
	wire _w27293_ ;
	wire _w27292_ ;
	wire _w27291_ ;
	wire _w27290_ ;
	wire _w27289_ ;
	wire _w27288_ ;
	wire _w27287_ ;
	wire _w27286_ ;
	wire _w27285_ ;
	wire _w27284_ ;
	wire _w27283_ ;
	wire _w27282_ ;
	wire _w27281_ ;
	wire _w27280_ ;
	wire _w27279_ ;
	wire _w27278_ ;
	wire _w27277_ ;
	wire _w27276_ ;
	wire _w27275_ ;
	wire _w27274_ ;
	wire _w27273_ ;
	wire _w27272_ ;
	wire _w27271_ ;
	wire _w27270_ ;
	wire _w27269_ ;
	wire _w27268_ ;
	wire _w27267_ ;
	wire _w27266_ ;
	wire _w27265_ ;
	wire _w27264_ ;
	wire _w27263_ ;
	wire _w27262_ ;
	wire _w27261_ ;
	wire _w27260_ ;
	wire _w27259_ ;
	wire _w27258_ ;
	wire _w27257_ ;
	wire _w27256_ ;
	wire _w27255_ ;
	wire _w27254_ ;
	wire _w27253_ ;
	wire _w27252_ ;
	wire _w27251_ ;
	wire _w27250_ ;
	wire _w27249_ ;
	wire _w27248_ ;
	wire _w27247_ ;
	wire _w27246_ ;
	wire _w27245_ ;
	wire _w27244_ ;
	wire _w27243_ ;
	wire _w27242_ ;
	wire _w27241_ ;
	wire _w27240_ ;
	wire _w27239_ ;
	wire _w27238_ ;
	wire _w27237_ ;
	wire _w27236_ ;
	wire _w27235_ ;
	wire _w27234_ ;
	wire _w27233_ ;
	wire _w27232_ ;
	wire _w27231_ ;
	wire _w27230_ ;
	wire _w27229_ ;
	wire _w27228_ ;
	wire _w27227_ ;
	wire _w27226_ ;
	wire _w27225_ ;
	wire _w27224_ ;
	wire _w27223_ ;
	wire _w27222_ ;
	wire _w27221_ ;
	wire _w27220_ ;
	wire _w27219_ ;
	wire _w27218_ ;
	wire _w27217_ ;
	wire _w27216_ ;
	wire _w27215_ ;
	wire _w27214_ ;
	wire _w27213_ ;
	wire _w27212_ ;
	wire _w27211_ ;
	wire _w27210_ ;
	wire _w27209_ ;
	wire _w27208_ ;
	wire _w27207_ ;
	wire _w27206_ ;
	wire _w27205_ ;
	wire _w27204_ ;
	wire _w27203_ ;
	wire _w27202_ ;
	wire _w27201_ ;
	wire _w27200_ ;
	wire _w27199_ ;
	wire _w27198_ ;
	wire _w27197_ ;
	wire _w27196_ ;
	wire _w27195_ ;
	wire _w27194_ ;
	wire _w27193_ ;
	wire _w27192_ ;
	wire _w27191_ ;
	wire _w27190_ ;
	wire _w27189_ ;
	wire _w27188_ ;
	wire _w27187_ ;
	wire _w27186_ ;
	wire _w27185_ ;
	wire _w27184_ ;
	wire _w27183_ ;
	wire _w27182_ ;
	wire _w27181_ ;
	wire _w27180_ ;
	wire _w27179_ ;
	wire _w27178_ ;
	wire _w27177_ ;
	wire _w27176_ ;
	wire _w27175_ ;
	wire _w27174_ ;
	wire _w27173_ ;
	wire _w27172_ ;
	wire _w27171_ ;
	wire _w27170_ ;
	wire _w27169_ ;
	wire _w27168_ ;
	wire _w27167_ ;
	wire _w27166_ ;
	wire _w27165_ ;
	wire _w27164_ ;
	wire _w27163_ ;
	wire _w27162_ ;
	wire _w27161_ ;
	wire _w27160_ ;
	wire _w27159_ ;
	wire _w27158_ ;
	wire _w27157_ ;
	wire _w27156_ ;
	wire _w27155_ ;
	wire _w27154_ ;
	wire _w27153_ ;
	wire _w27152_ ;
	wire _w27151_ ;
	wire _w27150_ ;
	wire _w27149_ ;
	wire _w27148_ ;
	wire _w27147_ ;
	wire _w27146_ ;
	wire _w27145_ ;
	wire _w27144_ ;
	wire _w27143_ ;
	wire _w27142_ ;
	wire _w27141_ ;
	wire _w27140_ ;
	wire _w27139_ ;
	wire _w27138_ ;
	wire _w27137_ ;
	wire _w27136_ ;
	wire _w27135_ ;
	wire _w27134_ ;
	wire _w27133_ ;
	wire _w27132_ ;
	wire _w27131_ ;
	wire _w27130_ ;
	wire _w27129_ ;
	wire _w27128_ ;
	wire _w27127_ ;
	wire _w27126_ ;
	wire _w27125_ ;
	wire _w27124_ ;
	wire _w27123_ ;
	wire _w27122_ ;
	wire _w27121_ ;
	wire _w27120_ ;
	wire _w27119_ ;
	wire _w27118_ ;
	wire _w27117_ ;
	wire _w27116_ ;
	wire _w27115_ ;
	wire _w27114_ ;
	wire _w27113_ ;
	wire _w27112_ ;
	wire _w27111_ ;
	wire _w27110_ ;
	wire _w27109_ ;
	wire _w27108_ ;
	wire _w27107_ ;
	wire _w27106_ ;
	wire _w27105_ ;
	wire _w27104_ ;
	wire _w27103_ ;
	wire _w27102_ ;
	wire _w27101_ ;
	wire _w27100_ ;
	wire _w27099_ ;
	wire _w27098_ ;
	wire _w27097_ ;
	wire _w27096_ ;
	wire _w27095_ ;
	wire _w27094_ ;
	wire _w27093_ ;
	wire _w27092_ ;
	wire _w27091_ ;
	wire _w27090_ ;
	wire _w27089_ ;
	wire _w27088_ ;
	wire _w27087_ ;
	wire _w27086_ ;
	wire _w27085_ ;
	wire _w27084_ ;
	wire _w27083_ ;
	wire _w27082_ ;
	wire _w27081_ ;
	wire _w27080_ ;
	wire _w27079_ ;
	wire _w27078_ ;
	wire _w27077_ ;
	wire _w27076_ ;
	wire _w27075_ ;
	wire _w27074_ ;
	wire _w27073_ ;
	wire _w27072_ ;
	wire _w27071_ ;
	wire _w27070_ ;
	wire _w27069_ ;
	wire _w27068_ ;
	wire _w27067_ ;
	wire _w27066_ ;
	wire _w27065_ ;
	wire _w27064_ ;
	wire _w27063_ ;
	wire _w27062_ ;
	wire _w27061_ ;
	wire _w27060_ ;
	wire _w27059_ ;
	wire _w27058_ ;
	wire _w27057_ ;
	wire _w27056_ ;
	wire _w27055_ ;
	wire _w27054_ ;
	wire _w27053_ ;
	wire _w27052_ ;
	wire _w27051_ ;
	wire _w27050_ ;
	wire _w27049_ ;
	wire _w27048_ ;
	wire _w27047_ ;
	wire _w27046_ ;
	wire _w27045_ ;
	wire _w27044_ ;
	wire _w27043_ ;
	wire _w27042_ ;
	wire _w27041_ ;
	wire _w27040_ ;
	wire _w27039_ ;
	wire _w27038_ ;
	wire _w27037_ ;
	wire _w27036_ ;
	wire _w27035_ ;
	wire _w27034_ ;
	wire _w27033_ ;
	wire _w27032_ ;
	wire _w27031_ ;
	wire _w27030_ ;
	wire _w27029_ ;
	wire _w27028_ ;
	wire _w27027_ ;
	wire _w27026_ ;
	wire _w27025_ ;
	wire _w27024_ ;
	wire _w27023_ ;
	wire _w27022_ ;
	wire _w27021_ ;
	wire _w27020_ ;
	wire _w27019_ ;
	wire _w27018_ ;
	wire _w27017_ ;
	wire _w27016_ ;
	wire _w27015_ ;
	wire _w27014_ ;
	wire _w27013_ ;
	wire _w27012_ ;
	wire _w27011_ ;
	wire _w27010_ ;
	wire _w27009_ ;
	wire _w27008_ ;
	wire _w27007_ ;
	wire _w27006_ ;
	wire _w27005_ ;
	wire _w27004_ ;
	wire _w27003_ ;
	wire _w27002_ ;
	wire _w27001_ ;
	wire _w27000_ ;
	wire _w26999_ ;
	wire _w26998_ ;
	wire _w26997_ ;
	wire _w26996_ ;
	wire _w26995_ ;
	wire _w26994_ ;
	wire _w26993_ ;
	wire _w26992_ ;
	wire _w26991_ ;
	wire _w26990_ ;
	wire _w26989_ ;
	wire _w26988_ ;
	wire _w26987_ ;
	wire _w26986_ ;
	wire _w26985_ ;
	wire _w26984_ ;
	wire _w26983_ ;
	wire _w26982_ ;
	wire _w26981_ ;
	wire _w26980_ ;
	wire _w26979_ ;
	wire _w26978_ ;
	wire _w26977_ ;
	wire _w26976_ ;
	wire _w26975_ ;
	wire _w26974_ ;
	wire _w26973_ ;
	wire _w26972_ ;
	wire _w26971_ ;
	wire _w26970_ ;
	wire _w26969_ ;
	wire _w26968_ ;
	wire _w26967_ ;
	wire _w26966_ ;
	wire _w26965_ ;
	wire _w26964_ ;
	wire _w26963_ ;
	wire _w26962_ ;
	wire _w26961_ ;
	wire _w26960_ ;
	wire _w26959_ ;
	wire _w26958_ ;
	wire _w26957_ ;
	wire _w26956_ ;
	wire _w26955_ ;
	wire _w26954_ ;
	wire _w26953_ ;
	wire _w26952_ ;
	wire _w26951_ ;
	wire _w26950_ ;
	wire _w26949_ ;
	wire _w26948_ ;
	wire _w26947_ ;
	wire _w26946_ ;
	wire _w26945_ ;
	wire _w26944_ ;
	wire _w26943_ ;
	wire _w26942_ ;
	wire _w26941_ ;
	wire _w26940_ ;
	wire _w26939_ ;
	wire _w26938_ ;
	wire _w26937_ ;
	wire _w26936_ ;
	wire _w26935_ ;
	wire _w26934_ ;
	wire _w26933_ ;
	wire _w26932_ ;
	wire _w26931_ ;
	wire _w26930_ ;
	wire _w26929_ ;
	wire _w26928_ ;
	wire _w26927_ ;
	wire _w26926_ ;
	wire _w26925_ ;
	wire _w26924_ ;
	wire _w26923_ ;
	wire _w26922_ ;
	wire _w26921_ ;
	wire _w26920_ ;
	wire _w26919_ ;
	wire _w26918_ ;
	wire _w26917_ ;
	wire _w26916_ ;
	wire _w26915_ ;
	wire _w26914_ ;
	wire _w26913_ ;
	wire _w26912_ ;
	wire _w26911_ ;
	wire _w26910_ ;
	wire _w26909_ ;
	wire _w26908_ ;
	wire _w26907_ ;
	wire _w26906_ ;
	wire _w26905_ ;
	wire _w26904_ ;
	wire _w26903_ ;
	wire _w26902_ ;
	wire _w26901_ ;
	wire _w26900_ ;
	wire _w26899_ ;
	wire _w26898_ ;
	wire _w26897_ ;
	wire _w26896_ ;
	wire _w26895_ ;
	wire _w26894_ ;
	wire _w26893_ ;
	wire _w26892_ ;
	wire _w26891_ ;
	wire _w26890_ ;
	wire _w26889_ ;
	wire _w26888_ ;
	wire _w26887_ ;
	wire _w26886_ ;
	wire _w26885_ ;
	wire _w26884_ ;
	wire _w26883_ ;
	wire _w26882_ ;
	wire _w26881_ ;
	wire _w26880_ ;
	wire _w26879_ ;
	wire _w26878_ ;
	wire _w26877_ ;
	wire _w26876_ ;
	wire _w26875_ ;
	wire _w26874_ ;
	wire _w26873_ ;
	wire _w26872_ ;
	wire _w26871_ ;
	wire _w26870_ ;
	wire _w26869_ ;
	wire _w26868_ ;
	wire _w26867_ ;
	wire _w26866_ ;
	wire _w26865_ ;
	wire _w26864_ ;
	wire _w26863_ ;
	wire _w26862_ ;
	wire _w26861_ ;
	wire _w26860_ ;
	wire _w26859_ ;
	wire _w26858_ ;
	wire _w26857_ ;
	wire _w26856_ ;
	wire _w26855_ ;
	wire _w26854_ ;
	wire _w26853_ ;
	wire _w26852_ ;
	wire _w26851_ ;
	wire _w26850_ ;
	wire _w26849_ ;
	wire _w26848_ ;
	wire _w26847_ ;
	wire _w26846_ ;
	wire _w26845_ ;
	wire _w26844_ ;
	wire _w26843_ ;
	wire _w26842_ ;
	wire _w26841_ ;
	wire _w26840_ ;
	wire _w26839_ ;
	wire _w26838_ ;
	wire _w26837_ ;
	wire _w26836_ ;
	wire _w26835_ ;
	wire _w26834_ ;
	wire _w26833_ ;
	wire _w26832_ ;
	wire _w26831_ ;
	wire _w26830_ ;
	wire _w26829_ ;
	wire _w26828_ ;
	wire _w26827_ ;
	wire _w26826_ ;
	wire _w26825_ ;
	wire _w26824_ ;
	wire _w26823_ ;
	wire _w26822_ ;
	wire _w26821_ ;
	wire _w26820_ ;
	wire _w26819_ ;
	wire _w26818_ ;
	wire _w26817_ ;
	wire _w26816_ ;
	wire _w26815_ ;
	wire _w26814_ ;
	wire _w26813_ ;
	wire _w26812_ ;
	wire _w26811_ ;
	wire _w26810_ ;
	wire _w26809_ ;
	wire _w26808_ ;
	wire _w26807_ ;
	wire _w26806_ ;
	wire _w26805_ ;
	wire _w26804_ ;
	wire _w26803_ ;
	wire _w26802_ ;
	wire _w26801_ ;
	wire _w26800_ ;
	wire _w26799_ ;
	wire _w26798_ ;
	wire _w26797_ ;
	wire _w26796_ ;
	wire _w26795_ ;
	wire _w26794_ ;
	wire _w26793_ ;
	wire _w26792_ ;
	wire _w26791_ ;
	wire _w26790_ ;
	wire _w26789_ ;
	wire _w26788_ ;
	wire _w26787_ ;
	wire _w26786_ ;
	wire _w26785_ ;
	wire _w26784_ ;
	wire _w26783_ ;
	wire _w26782_ ;
	wire _w26781_ ;
	wire _w26780_ ;
	wire _w26779_ ;
	wire _w26778_ ;
	wire _w26777_ ;
	wire _w26776_ ;
	wire _w26775_ ;
	wire _w26774_ ;
	wire _w26773_ ;
	wire _w26772_ ;
	wire _w26771_ ;
	wire _w26770_ ;
	wire _w26769_ ;
	wire _w26768_ ;
	wire _w26767_ ;
	wire _w26766_ ;
	wire _w26765_ ;
	wire _w26764_ ;
	wire _w26763_ ;
	wire _w26762_ ;
	wire _w26761_ ;
	wire _w26760_ ;
	wire _w26759_ ;
	wire _w26758_ ;
	wire _w26757_ ;
	wire _w26756_ ;
	wire _w26755_ ;
	wire _w26754_ ;
	wire _w26753_ ;
	wire _w26752_ ;
	wire _w26751_ ;
	wire _w26750_ ;
	wire _w26749_ ;
	wire _w26748_ ;
	wire _w26747_ ;
	wire _w26746_ ;
	wire _w26745_ ;
	wire _w26744_ ;
	wire _w26743_ ;
	wire _w26742_ ;
	wire _w26741_ ;
	wire _w26740_ ;
	wire _w26739_ ;
	wire _w26738_ ;
	wire _w26737_ ;
	wire _w26736_ ;
	wire _w26735_ ;
	wire _w26734_ ;
	wire _w26733_ ;
	wire _w26732_ ;
	wire _w26731_ ;
	wire _w26730_ ;
	wire _w26729_ ;
	wire _w26728_ ;
	wire _w26727_ ;
	wire _w26726_ ;
	wire _w26725_ ;
	wire _w26724_ ;
	wire _w26723_ ;
	wire _w26722_ ;
	wire _w26721_ ;
	wire _w26720_ ;
	wire _w26719_ ;
	wire _w26718_ ;
	wire _w26717_ ;
	wire _w26716_ ;
	wire _w26715_ ;
	wire _w26714_ ;
	wire _w26713_ ;
	wire _w26712_ ;
	wire _w26711_ ;
	wire _w26710_ ;
	wire _w26709_ ;
	wire _w26708_ ;
	wire _w26707_ ;
	wire _w26706_ ;
	wire _w26705_ ;
	wire _w26704_ ;
	wire _w26703_ ;
	wire _w26702_ ;
	wire _w26701_ ;
	wire _w26700_ ;
	wire _w26699_ ;
	wire _w26698_ ;
	wire _w26697_ ;
	wire _w26696_ ;
	wire _w26695_ ;
	wire _w26694_ ;
	wire _w26693_ ;
	wire _w26692_ ;
	wire _w26691_ ;
	wire _w26690_ ;
	wire _w26689_ ;
	wire _w26688_ ;
	wire _w26687_ ;
	wire _w26686_ ;
	wire _w26685_ ;
	wire _w26684_ ;
	wire _w26683_ ;
	wire _w26682_ ;
	wire _w26681_ ;
	wire _w26680_ ;
	wire _w26679_ ;
	wire _w26678_ ;
	wire _w26677_ ;
	wire _w26676_ ;
	wire _w26675_ ;
	wire _w26674_ ;
	wire _w26673_ ;
	wire _w26672_ ;
	wire _w26671_ ;
	wire _w26670_ ;
	wire _w26669_ ;
	wire _w26668_ ;
	wire _w26667_ ;
	wire _w26666_ ;
	wire _w26665_ ;
	wire _w26664_ ;
	wire _w26663_ ;
	wire _w26662_ ;
	wire _w26661_ ;
	wire _w26660_ ;
	wire _w26659_ ;
	wire _w26658_ ;
	wire _w26657_ ;
	wire _w26656_ ;
	wire _w26655_ ;
	wire _w26654_ ;
	wire _w26653_ ;
	wire _w26652_ ;
	wire _w26651_ ;
	wire _w26650_ ;
	wire _w26649_ ;
	wire _w26648_ ;
	wire _w26647_ ;
	wire _w26646_ ;
	wire _w26645_ ;
	wire _w26644_ ;
	wire _w26643_ ;
	wire _w26642_ ;
	wire _w26641_ ;
	wire _w26640_ ;
	wire _w26639_ ;
	wire _w26638_ ;
	wire _w26637_ ;
	wire _w26636_ ;
	wire _w26635_ ;
	wire _w26634_ ;
	wire _w26633_ ;
	wire _w26632_ ;
	wire _w26631_ ;
	wire _w26630_ ;
	wire _w26629_ ;
	wire _w26628_ ;
	wire _w26627_ ;
	wire _w26626_ ;
	wire _w26625_ ;
	wire _w26624_ ;
	wire _w26623_ ;
	wire _w26622_ ;
	wire _w26621_ ;
	wire _w26620_ ;
	wire _w26619_ ;
	wire _w26618_ ;
	wire _w26617_ ;
	wire _w26616_ ;
	wire _w26615_ ;
	wire _w26614_ ;
	wire _w26613_ ;
	wire _w26612_ ;
	wire _w26611_ ;
	wire _w26610_ ;
	wire _w26609_ ;
	wire _w26608_ ;
	wire _w26607_ ;
	wire _w26606_ ;
	wire _w26605_ ;
	wire _w26604_ ;
	wire _w26603_ ;
	wire _w26602_ ;
	wire _w26601_ ;
	wire _w26600_ ;
	wire _w26599_ ;
	wire _w26598_ ;
	wire _w26597_ ;
	wire _w26596_ ;
	wire _w26595_ ;
	wire _w26594_ ;
	wire _w26593_ ;
	wire _w26592_ ;
	wire _w26591_ ;
	wire _w26590_ ;
	wire _w26589_ ;
	wire _w26588_ ;
	wire _w26587_ ;
	wire _w26586_ ;
	wire _w26585_ ;
	wire _w26584_ ;
	wire _w26583_ ;
	wire _w26582_ ;
	wire _w26581_ ;
	wire _w26580_ ;
	wire _w16099_ ;
	wire _w16098_ ;
	wire _w16097_ ;
	wire _w16096_ ;
	wire _w16095_ ;
	wire _w16094_ ;
	wire _w16093_ ;
	wire _w16092_ ;
	wire _w16091_ ;
	wire _w16090_ ;
	wire _w16089_ ;
	wire _w16088_ ;
	wire _w16087_ ;
	wire _w16086_ ;
	wire _w16085_ ;
	wire _w16084_ ;
	wire _w16083_ ;
	wire _w16082_ ;
	wire _w16081_ ;
	wire _w16080_ ;
	wire _w16079_ ;
	wire _w16078_ ;
	wire _w16077_ ;
	wire _w16076_ ;
	wire _w16075_ ;
	wire _w16074_ ;
	wire _w16073_ ;
	wire _w16072_ ;
	wire _w16071_ ;
	wire _w16070_ ;
	wire _w16069_ ;
	wire _w16068_ ;
	wire _w16067_ ;
	wire _w16066_ ;
	wire _w16065_ ;
	wire _w16064_ ;
	wire _w16063_ ;
	wire _w16062_ ;
	wire _w16061_ ;
	wire _w16060_ ;
	wire _w16059_ ;
	wire _w16058_ ;
	wire _w16057_ ;
	wire _w16056_ ;
	wire _w16055_ ;
	wire _w16054_ ;
	wire _w16053_ ;
	wire _w16052_ ;
	wire _w16051_ ;
	wire _w16050_ ;
	wire _w16049_ ;
	wire _w16048_ ;
	wire _w16047_ ;
	wire _w16046_ ;
	wire _w16045_ ;
	wire _w16044_ ;
	wire _w16043_ ;
	wire _w16042_ ;
	wire _w16041_ ;
	wire _w16040_ ;
	wire _w16039_ ;
	wire _w16038_ ;
	wire _w16037_ ;
	wire _w16036_ ;
	wire _w16035_ ;
	wire _w16034_ ;
	wire _w16033_ ;
	wire _w16032_ ;
	wire _w16031_ ;
	wire _w16030_ ;
	wire _w16029_ ;
	wire _w16028_ ;
	wire _w16027_ ;
	wire _w16026_ ;
	wire _w16025_ ;
	wire _w16024_ ;
	wire _w16023_ ;
	wire _w16022_ ;
	wire _w16021_ ;
	wire _w16020_ ;
	wire _w16019_ ;
	wire _w16018_ ;
	wire _w16017_ ;
	wire _w16016_ ;
	wire _w16015_ ;
	wire _w16014_ ;
	wire _w16013_ ;
	wire _w16012_ ;
	wire _w16011_ ;
	wire _w16010_ ;
	wire _w16009_ ;
	wire _w16008_ ;
	wire _w16007_ ;
	wire _w16006_ ;
	wire _w16005_ ;
	wire _w16004_ ;
	wire _w16003_ ;
	wire _w16002_ ;
	wire _w16001_ ;
	wire _w16000_ ;
	wire _w15999_ ;
	wire _w15998_ ;
	wire _w15997_ ;
	wire _w15996_ ;
	wire _w15995_ ;
	wire _w15994_ ;
	wire _w15993_ ;
	wire _w15992_ ;
	wire _w15991_ ;
	wire _w15990_ ;
	wire _w15989_ ;
	wire _w15988_ ;
	wire _w15987_ ;
	wire _w15986_ ;
	wire _w15985_ ;
	wire _w15984_ ;
	wire _w15983_ ;
	wire _w15982_ ;
	wire _w15981_ ;
	wire _w15980_ ;
	wire _w15979_ ;
	wire _w15978_ ;
	wire _w15977_ ;
	wire _w15976_ ;
	wire _w15975_ ;
	wire _w15974_ ;
	wire _w15973_ ;
	wire _w15972_ ;
	wire _w15971_ ;
	wire _w15970_ ;
	wire _w15969_ ;
	wire _w15968_ ;
	wire _w15967_ ;
	wire _w15966_ ;
	wire _w15965_ ;
	wire _w15964_ ;
	wire _w15963_ ;
	wire _w15962_ ;
	wire _w15961_ ;
	wire _w15960_ ;
	wire _w15959_ ;
	wire _w15958_ ;
	wire _w15957_ ;
	wire _w15956_ ;
	wire _w15955_ ;
	wire _w15954_ ;
	wire _w15953_ ;
	wire _w15952_ ;
	wire _w15951_ ;
	wire _w15950_ ;
	wire _w15949_ ;
	wire _w15948_ ;
	wire _w15947_ ;
	wire _w15946_ ;
	wire _w15945_ ;
	wire _w15944_ ;
	wire _w15943_ ;
	wire _w15942_ ;
	wire _w15941_ ;
	wire _w15940_ ;
	wire _w15939_ ;
	wire _w15938_ ;
	wire _w15937_ ;
	wire _w15936_ ;
	wire _w15935_ ;
	wire _w15934_ ;
	wire _w15933_ ;
	wire _w15932_ ;
	wire _w15931_ ;
	wire _w15930_ ;
	wire _w15929_ ;
	wire _w15928_ ;
	wire _w15927_ ;
	wire _w15926_ ;
	wire _w15925_ ;
	wire _w15924_ ;
	wire _w15923_ ;
	wire _w15922_ ;
	wire _w15921_ ;
	wire _w15920_ ;
	wire _w15919_ ;
	wire _w15918_ ;
	wire _w15917_ ;
	wire _w15916_ ;
	wire _w15915_ ;
	wire _w15914_ ;
	wire _w15913_ ;
	wire _w15912_ ;
	wire _w15911_ ;
	wire _w15910_ ;
	wire _w15909_ ;
	wire _w15908_ ;
	wire _w15907_ ;
	wire _w15906_ ;
	wire _w15905_ ;
	wire _w15904_ ;
	wire _w15903_ ;
	wire _w15902_ ;
	wire _w15901_ ;
	wire _w15900_ ;
	wire _w15899_ ;
	wire _w15898_ ;
	wire _w15897_ ;
	wire _w15896_ ;
	wire _w15895_ ;
	wire _w15894_ ;
	wire _w15893_ ;
	wire _w15892_ ;
	wire _w15891_ ;
	wire _w15890_ ;
	wire _w15889_ ;
	wire _w15888_ ;
	wire _w15887_ ;
	wire _w15886_ ;
	wire _w15885_ ;
	wire _w15884_ ;
	wire _w15883_ ;
	wire _w15882_ ;
	wire _w15881_ ;
	wire _w15880_ ;
	wire _w15879_ ;
	wire _w15878_ ;
	wire _w15877_ ;
	wire _w15876_ ;
	wire _w15875_ ;
	wire _w15874_ ;
	wire _w15873_ ;
	wire _w15872_ ;
	wire _w15871_ ;
	wire _w15870_ ;
	wire _w15869_ ;
	wire _w15868_ ;
	wire _w15867_ ;
	wire _w15866_ ;
	wire _w15865_ ;
	wire _w15864_ ;
	wire _w15863_ ;
	wire _w15862_ ;
	wire _w15861_ ;
	wire _w15860_ ;
	wire _w15859_ ;
	wire _w15858_ ;
	wire _w15857_ ;
	wire _w15856_ ;
	wire _w15855_ ;
	wire _w15854_ ;
	wire _w15853_ ;
	wire _w15852_ ;
	wire _w15851_ ;
	wire _w15850_ ;
	wire _w15849_ ;
	wire _w15848_ ;
	wire _w15847_ ;
	wire _w15846_ ;
	wire _w15845_ ;
	wire _w15844_ ;
	wire _w15843_ ;
	wire _w15842_ ;
	wire _w15841_ ;
	wire _w15840_ ;
	wire _w15839_ ;
	wire _w15838_ ;
	wire _w15837_ ;
	wire _w15836_ ;
	wire _w15835_ ;
	wire _w15834_ ;
	wire _w15833_ ;
	wire _w15832_ ;
	wire _w15831_ ;
	wire _w15830_ ;
	wire _w15829_ ;
	wire _w15828_ ;
	wire _w15827_ ;
	wire _w15826_ ;
	wire _w15825_ ;
	wire _w15824_ ;
	wire _w15823_ ;
	wire _w15822_ ;
	wire _w15821_ ;
	wire _w15820_ ;
	wire _w15819_ ;
	wire _w15818_ ;
	wire _w15817_ ;
	wire _w15816_ ;
	wire _w15815_ ;
	wire _w15814_ ;
	wire _w15813_ ;
	wire _w15812_ ;
	wire _w15811_ ;
	wire _w15810_ ;
	wire _w15809_ ;
	wire _w15808_ ;
	wire _w15807_ ;
	wire _w15806_ ;
	wire _w15805_ ;
	wire _w15804_ ;
	wire _w15803_ ;
	wire _w15802_ ;
	wire _w15801_ ;
	wire _w15800_ ;
	wire _w15799_ ;
	wire _w15798_ ;
	wire _w15797_ ;
	wire _w15796_ ;
	wire _w15795_ ;
	wire _w15794_ ;
	wire _w15793_ ;
	wire _w15792_ ;
	wire _w15791_ ;
	wire _w15790_ ;
	wire _w15789_ ;
	wire _w15788_ ;
	wire _w15787_ ;
	wire _w15786_ ;
	wire _w15785_ ;
	wire _w15784_ ;
	wire _w15783_ ;
	wire _w15782_ ;
	wire _w15781_ ;
	wire _w15780_ ;
	wire _w15779_ ;
	wire _w15778_ ;
	wire _w15777_ ;
	wire _w15776_ ;
	wire _w15775_ ;
	wire _w15774_ ;
	wire _w15773_ ;
	wire _w15772_ ;
	wire _w15771_ ;
	wire _w15770_ ;
	wire _w15769_ ;
	wire _w15768_ ;
	wire _w15767_ ;
	wire _w15766_ ;
	wire _w15765_ ;
	wire _w15764_ ;
	wire _w15763_ ;
	wire _w15762_ ;
	wire _w15761_ ;
	wire _w15760_ ;
	wire _w15759_ ;
	wire _w15758_ ;
	wire _w15757_ ;
	wire _w15756_ ;
	wire _w15755_ ;
	wire _w15754_ ;
	wire _w15753_ ;
	wire _w15752_ ;
	wire _w15751_ ;
	wire _w15750_ ;
	wire _w15749_ ;
	wire _w15748_ ;
	wire _w15747_ ;
	wire _w15746_ ;
	wire _w15745_ ;
	wire _w15744_ ;
	wire _w15743_ ;
	wire _w15742_ ;
	wire _w15741_ ;
	wire _w15740_ ;
	wire _w15739_ ;
	wire _w15738_ ;
	wire _w15737_ ;
	wire _w15736_ ;
	wire _w15735_ ;
	wire _w15734_ ;
	wire _w15733_ ;
	wire _w15732_ ;
	wire _w15731_ ;
	wire _w15730_ ;
	wire _w15729_ ;
	wire _w15728_ ;
	wire _w15727_ ;
	wire _w15726_ ;
	wire _w15725_ ;
	wire _w15724_ ;
	wire _w15723_ ;
	wire _w15722_ ;
	wire _w15721_ ;
	wire _w15720_ ;
	wire _w15719_ ;
	wire _w15718_ ;
	wire _w15717_ ;
	wire _w15716_ ;
	wire _w15715_ ;
	wire _w15714_ ;
	wire _w15713_ ;
	wire _w15712_ ;
	wire _w15711_ ;
	wire _w15710_ ;
	wire _w15709_ ;
	wire _w15708_ ;
	wire _w15707_ ;
	wire _w15706_ ;
	wire _w15705_ ;
	wire _w15704_ ;
	wire _w15703_ ;
	wire _w15702_ ;
	wire _w15701_ ;
	wire _w15700_ ;
	wire _w15699_ ;
	wire _w15698_ ;
	wire _w15697_ ;
	wire _w15696_ ;
	wire _w15695_ ;
	wire _w15694_ ;
	wire _w15693_ ;
	wire _w15692_ ;
	wire _w15691_ ;
	wire _w15690_ ;
	wire _w15689_ ;
	wire _w15688_ ;
	wire _w15687_ ;
	wire _w15686_ ;
	wire _w15685_ ;
	wire _w15684_ ;
	wire _w15683_ ;
	wire _w15682_ ;
	wire _w15681_ ;
	wire _w15680_ ;
	wire _w15679_ ;
	wire _w15678_ ;
	wire _w15677_ ;
	wire _w15676_ ;
	wire _w15675_ ;
	wire _w15674_ ;
	wire _w15673_ ;
	wire _w15672_ ;
	wire _w15671_ ;
	wire _w15670_ ;
	wire _w15669_ ;
	wire _w15668_ ;
	wire _w15667_ ;
	wire _w15666_ ;
	wire _w15665_ ;
	wire _w15664_ ;
	wire _w15663_ ;
	wire _w15662_ ;
	wire _w15661_ ;
	wire _w15660_ ;
	wire _w15659_ ;
	wire _w15658_ ;
	wire _w15657_ ;
	wire _w15656_ ;
	wire _w15655_ ;
	wire _w15654_ ;
	wire _w15653_ ;
	wire _w15652_ ;
	wire _w15651_ ;
	wire _w15650_ ;
	wire _w15649_ ;
	wire _w15648_ ;
	wire _w15647_ ;
	wire _w15646_ ;
	wire _w15645_ ;
	wire _w15644_ ;
	wire _w15643_ ;
	wire _w15642_ ;
	wire _w15641_ ;
	wire _w15640_ ;
	wire _w15639_ ;
	wire _w15638_ ;
	wire _w15637_ ;
	wire _w15636_ ;
	wire _w15635_ ;
	wire _w15634_ ;
	wire _w15633_ ;
	wire _w15632_ ;
	wire _w15631_ ;
	wire _w15630_ ;
	wire _w15629_ ;
	wire _w15628_ ;
	wire _w15627_ ;
	wire _w15626_ ;
	wire _w15625_ ;
	wire _w15624_ ;
	wire _w15623_ ;
	wire _w15622_ ;
	wire _w15621_ ;
	wire _w15620_ ;
	wire _w15619_ ;
	wire _w15618_ ;
	wire _w15617_ ;
	wire _w15616_ ;
	wire _w15615_ ;
	wire _w15614_ ;
	wire _w15613_ ;
	wire _w15612_ ;
	wire _w15611_ ;
	wire _w15610_ ;
	wire _w15609_ ;
	wire _w15608_ ;
	wire _w15607_ ;
	wire _w15606_ ;
	wire _w15605_ ;
	wire _w15604_ ;
	wire _w15603_ ;
	wire _w15602_ ;
	wire _w15601_ ;
	wire _w15600_ ;
	wire _w15599_ ;
	wire _w15598_ ;
	wire _w15597_ ;
	wire _w15596_ ;
	wire _w15595_ ;
	wire _w15594_ ;
	wire _w15593_ ;
	wire _w15592_ ;
	wire _w15591_ ;
	wire _w15590_ ;
	wire _w15589_ ;
	wire _w15588_ ;
	wire _w15587_ ;
	wire _w15586_ ;
	wire _w15585_ ;
	wire _w15584_ ;
	wire _w15583_ ;
	wire _w15582_ ;
	wire _w15581_ ;
	wire _w15580_ ;
	wire _w15579_ ;
	wire _w15578_ ;
	wire _w15577_ ;
	wire _w15576_ ;
	wire _w15575_ ;
	wire _w15574_ ;
	wire _w15573_ ;
	wire _w15572_ ;
	wire _w15571_ ;
	wire _w15570_ ;
	wire _w15569_ ;
	wire _w15568_ ;
	wire _w15567_ ;
	wire _w15566_ ;
	wire _w15565_ ;
	wire _w15564_ ;
	wire _w15563_ ;
	wire _w15562_ ;
	wire _w15561_ ;
	wire _w15560_ ;
	wire _w15559_ ;
	wire _w15558_ ;
	wire _w15557_ ;
	wire _w15556_ ;
	wire _w15555_ ;
	wire _w15554_ ;
	wire _w15553_ ;
	wire _w15552_ ;
	wire _w15551_ ;
	wire _w15550_ ;
	wire _w15549_ ;
	wire _w15548_ ;
	wire _w15547_ ;
	wire _w15546_ ;
	wire _w15545_ ;
	wire _w15544_ ;
	wire _w15543_ ;
	wire _w15542_ ;
	wire _w15541_ ;
	wire _w15540_ ;
	wire _w15539_ ;
	wire _w15538_ ;
	wire _w15537_ ;
	wire _w15536_ ;
	wire _w15535_ ;
	wire _w15534_ ;
	wire _w15533_ ;
	wire _w15532_ ;
	wire _w15531_ ;
	wire _w15530_ ;
	wire _w15529_ ;
	wire _w15528_ ;
	wire _w15527_ ;
	wire _w15526_ ;
	wire _w15525_ ;
	wire _w15524_ ;
	wire _w15523_ ;
	wire _w15522_ ;
	wire _w15521_ ;
	wire _w15520_ ;
	wire _w15519_ ;
	wire _w15518_ ;
	wire _w15517_ ;
	wire _w15516_ ;
	wire _w15515_ ;
	wire _w15514_ ;
	wire _w15513_ ;
	wire _w15512_ ;
	wire _w15511_ ;
	wire _w15510_ ;
	wire _w15509_ ;
	wire _w15508_ ;
	wire _w15507_ ;
	wire _w15506_ ;
	wire _w15505_ ;
	wire _w15504_ ;
	wire _w15503_ ;
	wire _w15502_ ;
	wire _w15501_ ;
	wire _w15500_ ;
	wire _w15499_ ;
	wire _w15498_ ;
	wire _w15497_ ;
	wire _w15496_ ;
	wire _w15495_ ;
	wire _w15494_ ;
	wire _w15493_ ;
	wire _w15492_ ;
	wire _w15491_ ;
	wire _w15490_ ;
	wire _w15489_ ;
	wire _w15488_ ;
	wire _w15487_ ;
	wire _w15486_ ;
	wire _w15485_ ;
	wire _w15484_ ;
	wire _w15483_ ;
	wire _w15482_ ;
	wire _w15481_ ;
	wire _w15480_ ;
	wire _w15479_ ;
	wire _w15478_ ;
	wire _w15477_ ;
	wire _w15476_ ;
	wire _w15475_ ;
	wire _w15474_ ;
	wire _w15473_ ;
	wire _w15472_ ;
	wire _w15471_ ;
	wire _w15470_ ;
	wire _w15469_ ;
	wire _w15468_ ;
	wire _w15467_ ;
	wire _w15466_ ;
	wire _w15465_ ;
	wire _w15464_ ;
	wire _w15463_ ;
	wire _w15462_ ;
	wire _w15461_ ;
	wire _w15460_ ;
	wire _w15459_ ;
	wire _w15458_ ;
	wire _w15457_ ;
	wire _w15456_ ;
	wire _w15455_ ;
	wire _w15454_ ;
	wire _w15453_ ;
	wire _w15452_ ;
	wire _w15451_ ;
	wire _w15450_ ;
	wire _w15449_ ;
	wire _w15448_ ;
	wire _w15447_ ;
	wire _w15446_ ;
	wire _w15445_ ;
	wire _w15444_ ;
	wire _w15443_ ;
	wire _w15442_ ;
	wire _w15441_ ;
	wire _w15440_ ;
	wire _w15439_ ;
	wire _w15438_ ;
	wire _w15437_ ;
	wire _w15436_ ;
	wire _w15435_ ;
	wire _w15434_ ;
	wire _w15433_ ;
	wire _w15432_ ;
	wire _w15431_ ;
	wire _w15430_ ;
	wire _w15429_ ;
	wire _w15428_ ;
	wire _w15427_ ;
	wire _w15426_ ;
	wire _w15425_ ;
	wire _w15424_ ;
	wire _w15423_ ;
	wire _w15422_ ;
	wire _w15421_ ;
	wire _w15420_ ;
	wire _w15419_ ;
	wire _w15418_ ;
	wire _w15417_ ;
	wire _w15416_ ;
	wire _w15415_ ;
	wire _w15414_ ;
	wire _w15413_ ;
	wire _w15412_ ;
	wire _w15411_ ;
	wire _w15410_ ;
	wire _w15409_ ;
	wire _w15408_ ;
	wire _w15407_ ;
	wire _w15406_ ;
	wire _w15405_ ;
	wire _w15404_ ;
	wire _w15403_ ;
	wire _w15402_ ;
	wire _w15401_ ;
	wire _w15400_ ;
	wire _w15399_ ;
	wire _w15398_ ;
	wire _w15397_ ;
	wire _w15396_ ;
	wire _w15395_ ;
	wire _w15394_ ;
	wire _w15393_ ;
	wire _w15392_ ;
	wire _w15391_ ;
	wire _w15390_ ;
	wire _w15389_ ;
	wire _w15388_ ;
	wire _w15387_ ;
	wire _w15386_ ;
	wire _w15385_ ;
	wire _w15384_ ;
	wire _w15383_ ;
	wire _w15382_ ;
	wire _w15381_ ;
	wire _w15380_ ;
	wire _w15379_ ;
	wire _w15378_ ;
	wire _w15377_ ;
	wire _w15376_ ;
	wire _w15375_ ;
	wire _w15374_ ;
	wire _w15373_ ;
	wire _w15372_ ;
	wire _w15371_ ;
	wire _w15370_ ;
	wire _w15369_ ;
	wire _w15368_ ;
	wire _w15367_ ;
	wire _w15366_ ;
	wire _w15365_ ;
	wire _w15364_ ;
	wire _w15363_ ;
	wire _w15362_ ;
	wire _w15361_ ;
	wire _w15360_ ;
	wire _w15359_ ;
	wire _w15358_ ;
	wire _w15357_ ;
	wire _w15356_ ;
	wire _w15355_ ;
	wire _w15354_ ;
	wire _w15353_ ;
	wire _w15352_ ;
	wire _w15351_ ;
	wire _w15350_ ;
	wire _w15349_ ;
	wire _w15348_ ;
	wire _w15347_ ;
	wire _w15346_ ;
	wire _w15345_ ;
	wire _w15344_ ;
	wire _w15343_ ;
	wire _w15342_ ;
	wire _w15341_ ;
	wire _w15340_ ;
	wire _w15339_ ;
	wire _w15338_ ;
	wire _w15337_ ;
	wire _w15336_ ;
	wire _w15335_ ;
	wire _w15334_ ;
	wire _w15333_ ;
	wire _w15332_ ;
	wire _w15331_ ;
	wire _w15330_ ;
	wire _w15329_ ;
	wire _w15328_ ;
	wire _w15327_ ;
	wire _w15326_ ;
	wire _w15325_ ;
	wire _w15324_ ;
	wire _w15323_ ;
	wire _w15322_ ;
	wire _w15321_ ;
	wire _w15320_ ;
	wire _w15319_ ;
	wire _w15318_ ;
	wire _w15317_ ;
	wire _w15316_ ;
	wire _w15315_ ;
	wire _w15314_ ;
	wire _w15313_ ;
	wire _w15312_ ;
	wire _w15311_ ;
	wire _w15310_ ;
	wire _w15309_ ;
	wire _w15308_ ;
	wire _w15307_ ;
	wire _w15306_ ;
	wire _w15305_ ;
	wire _w15304_ ;
	wire _w15303_ ;
	wire _w15302_ ;
	wire _w15301_ ;
	wire _w15300_ ;
	wire _w15299_ ;
	wire _w15298_ ;
	wire _w15297_ ;
	wire _w15296_ ;
	wire _w15295_ ;
	wire _w15294_ ;
	wire _w15293_ ;
	wire _w15292_ ;
	wire _w15291_ ;
	wire _w15290_ ;
	wire _w15289_ ;
	wire _w15288_ ;
	wire _w15287_ ;
	wire _w15286_ ;
	wire _w15285_ ;
	wire _w15284_ ;
	wire _w15283_ ;
	wire _w15282_ ;
	wire _w15281_ ;
	wire _w15280_ ;
	wire _w15279_ ;
	wire _w15278_ ;
	wire _w15277_ ;
	wire _w15276_ ;
	wire _w15275_ ;
	wire _w15274_ ;
	wire _w15273_ ;
	wire _w15272_ ;
	wire _w15271_ ;
	wire _w15270_ ;
	wire _w15269_ ;
	wire _w15268_ ;
	wire _w15267_ ;
	wire _w15266_ ;
	wire _w15265_ ;
	wire _w15264_ ;
	wire _w15263_ ;
	wire _w15262_ ;
	wire _w15261_ ;
	wire _w15260_ ;
	wire _w15259_ ;
	wire _w15258_ ;
	wire _w15257_ ;
	wire _w15256_ ;
	wire _w15255_ ;
	wire _w15254_ ;
	wire _w15253_ ;
	wire _w15252_ ;
	wire _w15251_ ;
	wire _w15250_ ;
	wire _w15249_ ;
	wire _w15248_ ;
	wire _w15247_ ;
	wire _w15246_ ;
	wire _w15245_ ;
	wire _w15244_ ;
	wire _w15243_ ;
	wire _w15242_ ;
	wire _w15241_ ;
	wire _w15240_ ;
	wire _w15239_ ;
	wire _w15238_ ;
	wire _w15237_ ;
	wire _w15236_ ;
	wire _w15235_ ;
	wire _w15234_ ;
	wire _w15233_ ;
	wire _w15232_ ;
	wire _w15231_ ;
	wire _w15230_ ;
	wire _w15229_ ;
	wire _w15228_ ;
	wire _w15227_ ;
	wire _w15226_ ;
	wire _w15225_ ;
	wire _w15224_ ;
	wire _w15223_ ;
	wire _w15222_ ;
	wire _w15221_ ;
	wire _w15220_ ;
	wire _w15219_ ;
	wire _w15218_ ;
	wire _w15217_ ;
	wire _w15216_ ;
	wire _w15215_ ;
	wire _w15214_ ;
	wire _w15213_ ;
	wire _w15212_ ;
	wire _w15211_ ;
	wire _w15210_ ;
	wire _w15209_ ;
	wire _w15208_ ;
	wire _w15207_ ;
	wire _w15206_ ;
	wire _w15205_ ;
	wire _w15204_ ;
	wire _w15203_ ;
	wire _w15202_ ;
	wire _w15201_ ;
	wire _w15200_ ;
	wire _w15199_ ;
	wire _w15198_ ;
	wire _w15197_ ;
	wire _w15196_ ;
	wire _w15195_ ;
	wire _w15194_ ;
	wire _w15193_ ;
	wire _w15192_ ;
	wire _w15191_ ;
	wire _w15190_ ;
	wire _w15189_ ;
	wire _w15188_ ;
	wire _w15187_ ;
	wire _w15186_ ;
	wire _w15185_ ;
	wire _w15184_ ;
	wire _w15183_ ;
	wire _w15182_ ;
	wire _w15181_ ;
	wire _w15180_ ;
	wire _w15179_ ;
	wire _w15178_ ;
	wire _w15177_ ;
	wire _w15176_ ;
	wire _w15175_ ;
	wire _w15174_ ;
	wire _w15173_ ;
	wire _w15172_ ;
	wire _w15171_ ;
	wire _w15170_ ;
	wire _w15169_ ;
	wire _w15168_ ;
	wire _w15167_ ;
	wire _w15166_ ;
	wire _w15165_ ;
	wire _w15164_ ;
	wire _w15163_ ;
	wire _w15162_ ;
	wire _w15161_ ;
	wire _w15160_ ;
	wire _w15159_ ;
	wire _w15158_ ;
	wire _w15157_ ;
	wire _w15156_ ;
	wire _w15155_ ;
	wire _w15154_ ;
	wire _w15153_ ;
	wire _w15152_ ;
	wire _w15151_ ;
	wire _w15150_ ;
	wire _w15149_ ;
	wire _w15148_ ;
	wire _w15147_ ;
	wire _w15146_ ;
	wire _w15145_ ;
	wire _w15144_ ;
	wire _w15143_ ;
	wire _w15142_ ;
	wire _w15141_ ;
	wire _w15140_ ;
	wire _w15139_ ;
	wire _w15138_ ;
	wire _w15137_ ;
	wire _w15136_ ;
	wire _w15135_ ;
	wire _w15134_ ;
	wire _w15133_ ;
	wire _w15132_ ;
	wire _w15131_ ;
	wire _w15130_ ;
	wire _w15129_ ;
	wire _w15128_ ;
	wire _w15127_ ;
	wire _w15126_ ;
	wire _w15125_ ;
	wire _w15124_ ;
	wire _w15123_ ;
	wire _w15122_ ;
	wire _w15121_ ;
	wire _w15120_ ;
	wire _w15119_ ;
	wire _w15118_ ;
	wire _w15117_ ;
	wire _w15116_ ;
	wire _w15115_ ;
	wire _w15114_ ;
	wire _w15113_ ;
	wire _w15112_ ;
	wire _w15111_ ;
	wire _w15110_ ;
	wire _w15109_ ;
	wire _w15108_ ;
	wire _w15107_ ;
	wire _w15106_ ;
	wire _w15105_ ;
	wire _w15104_ ;
	wire _w15103_ ;
	wire _w15102_ ;
	wire _w15101_ ;
	wire _w15100_ ;
	wire _w15099_ ;
	wire _w15098_ ;
	wire _w15097_ ;
	wire _w15096_ ;
	wire _w15095_ ;
	wire _w15094_ ;
	wire _w15093_ ;
	wire _w15092_ ;
	wire _w15091_ ;
	wire _w15090_ ;
	wire _w15089_ ;
	wire _w15088_ ;
	wire _w15087_ ;
	wire _w15086_ ;
	wire _w15085_ ;
	wire _w15084_ ;
	wire _w15083_ ;
	wire _w15082_ ;
	wire _w15081_ ;
	wire _w15080_ ;
	wire _w15079_ ;
	wire _w15078_ ;
	wire _w15077_ ;
	wire _w15076_ ;
	wire _w15075_ ;
	wire _w15074_ ;
	wire _w15073_ ;
	wire _w15072_ ;
	wire _w15071_ ;
	wire _w15070_ ;
	wire _w15069_ ;
	wire _w15068_ ;
	wire _w15067_ ;
	wire _w15066_ ;
	wire _w15065_ ;
	wire _w15064_ ;
	wire _w15063_ ;
	wire _w15062_ ;
	wire _w15061_ ;
	wire _w15060_ ;
	wire _w15059_ ;
	wire _w15058_ ;
	wire _w15057_ ;
	wire _w15056_ ;
	wire _w15055_ ;
	wire _w15054_ ;
	wire _w15053_ ;
	wire _w15052_ ;
	wire _w15051_ ;
	wire _w15050_ ;
	wire _w15049_ ;
	wire _w15048_ ;
	wire _w15047_ ;
	wire _w15046_ ;
	wire _w15045_ ;
	wire _w15044_ ;
	wire _w15043_ ;
	wire _w15042_ ;
	wire _w15041_ ;
	wire _w15040_ ;
	wire _w15039_ ;
	wire _w15038_ ;
	wire _w15037_ ;
	wire _w15036_ ;
	wire _w15035_ ;
	wire _w15034_ ;
	wire _w15033_ ;
	wire _w15032_ ;
	wire _w15031_ ;
	wire _w15030_ ;
	wire _w15029_ ;
	wire _w15028_ ;
	wire _w15027_ ;
	wire _w15026_ ;
	wire _w15025_ ;
	wire _w15024_ ;
	wire _w15023_ ;
	wire _w15022_ ;
	wire _w15021_ ;
	wire _w15020_ ;
	wire _w15019_ ;
	wire _w15018_ ;
	wire _w15017_ ;
	wire _w15016_ ;
	wire _w15015_ ;
	wire _w15014_ ;
	wire _w15013_ ;
	wire _w15012_ ;
	wire _w15011_ ;
	wire _w15010_ ;
	wire _w15009_ ;
	wire _w15008_ ;
	wire _w15007_ ;
	wire _w15006_ ;
	wire _w15005_ ;
	wire _w15004_ ;
	wire _w15003_ ;
	wire _w15002_ ;
	wire _w15001_ ;
	wire _w15000_ ;
	wire _w14999_ ;
	wire _w14998_ ;
	wire _w14997_ ;
	wire _w14996_ ;
	wire _w14995_ ;
	wire _w14994_ ;
	wire _w14993_ ;
	wire _w14992_ ;
	wire _w14991_ ;
	wire _w14990_ ;
	wire _w14989_ ;
	wire _w14988_ ;
	wire _w14987_ ;
	wire _w14986_ ;
	wire _w14985_ ;
	wire _w14984_ ;
	wire _w14983_ ;
	wire _w14982_ ;
	wire _w14981_ ;
	wire _w14980_ ;
	wire _w14979_ ;
	wire _w14978_ ;
	wire _w14977_ ;
	wire _w14976_ ;
	wire _w14975_ ;
	wire _w14974_ ;
	wire _w14973_ ;
	wire _w14972_ ;
	wire _w14971_ ;
	wire _w14970_ ;
	wire _w14969_ ;
	wire _w14968_ ;
	wire _w14967_ ;
	wire _w14966_ ;
	wire _w14965_ ;
	wire _w14964_ ;
	wire _w14963_ ;
	wire _w14962_ ;
	wire _w14961_ ;
	wire _w14960_ ;
	wire _w14959_ ;
	wire _w14958_ ;
	wire _w14957_ ;
	wire _w14956_ ;
	wire _w14955_ ;
	wire _w14954_ ;
	wire _w14953_ ;
	wire _w14952_ ;
	wire _w14951_ ;
	wire _w14950_ ;
	wire _w14949_ ;
	wire _w14948_ ;
	wire _w14947_ ;
	wire _w14946_ ;
	wire _w14945_ ;
	wire _w14944_ ;
	wire _w14943_ ;
	wire _w14942_ ;
	wire _w14941_ ;
	wire _w14940_ ;
	wire _w14939_ ;
	wire _w14938_ ;
	wire _w14937_ ;
	wire _w14936_ ;
	wire _w14935_ ;
	wire _w14934_ ;
	wire _w14933_ ;
	wire _w14932_ ;
	wire _w14931_ ;
	wire _w14930_ ;
	wire _w14929_ ;
	wire _w14928_ ;
	wire _w14927_ ;
	wire _w14926_ ;
	wire _w14925_ ;
	wire _w14924_ ;
	wire _w14923_ ;
	wire _w14922_ ;
	wire _w14921_ ;
	wire _w14920_ ;
	wire _w14919_ ;
	wire _w14918_ ;
	wire _w14917_ ;
	wire _w14916_ ;
	wire _w14915_ ;
	wire _w14914_ ;
	wire _w14913_ ;
	wire _w14912_ ;
	wire _w14911_ ;
	wire _w14910_ ;
	wire _w14909_ ;
	wire _w14908_ ;
	wire _w14907_ ;
	wire _w14906_ ;
	wire _w14905_ ;
	wire _w14904_ ;
	wire _w14903_ ;
	wire _w14902_ ;
	wire _w14901_ ;
	wire _w14900_ ;
	wire _w14899_ ;
	wire _w14898_ ;
	wire _w14897_ ;
	wire _w14896_ ;
	wire _w14895_ ;
	wire _w14894_ ;
	wire _w14893_ ;
	wire _w14892_ ;
	wire _w14891_ ;
	wire _w14890_ ;
	wire _w14889_ ;
	wire _w14888_ ;
	wire _w14887_ ;
	wire _w14886_ ;
	wire _w14885_ ;
	wire _w14884_ ;
	wire _w14883_ ;
	wire _w14882_ ;
	wire _w14881_ ;
	wire _w14880_ ;
	wire _w14879_ ;
	wire _w14878_ ;
	wire _w14877_ ;
	wire _w14876_ ;
	wire _w14875_ ;
	wire _w14874_ ;
	wire _w14873_ ;
	wire _w14872_ ;
	wire _w14871_ ;
	wire _w14870_ ;
	wire _w14869_ ;
	wire _w14868_ ;
	wire _w14867_ ;
	wire _w14866_ ;
	wire _w14865_ ;
	wire _w14864_ ;
	wire _w14863_ ;
	wire _w14862_ ;
	wire _w14861_ ;
	wire _w14860_ ;
	wire _w14859_ ;
	wire _w14858_ ;
	wire _w14857_ ;
	wire _w14856_ ;
	wire _w14855_ ;
	wire _w14854_ ;
	wire _w14853_ ;
	wire _w14852_ ;
	wire _w14851_ ;
	wire _w14850_ ;
	wire _w14849_ ;
	wire _w14848_ ;
	wire _w14847_ ;
	wire _w14846_ ;
	wire _w14845_ ;
	wire _w14844_ ;
	wire _w14843_ ;
	wire _w14842_ ;
	wire _w14841_ ;
	wire _w14840_ ;
	wire _w14839_ ;
	wire _w14838_ ;
	wire _w14837_ ;
	wire _w14836_ ;
	wire _w14835_ ;
	wire _w14834_ ;
	wire _w14833_ ;
	wire _w14832_ ;
	wire _w14831_ ;
	wire _w14830_ ;
	wire _w14829_ ;
	wire _w14828_ ;
	wire _w14827_ ;
	wire _w14826_ ;
	wire _w14825_ ;
	wire _w14824_ ;
	wire _w14823_ ;
	wire _w14822_ ;
	wire _w14821_ ;
	wire _w14820_ ;
	wire _w14819_ ;
	wire _w14818_ ;
	wire _w14817_ ;
	wire _w14816_ ;
	wire _w14815_ ;
	wire _w14814_ ;
	wire _w14813_ ;
	wire _w14812_ ;
	wire _w14811_ ;
	wire _w14810_ ;
	wire _w14809_ ;
	wire _w14808_ ;
	wire _w14807_ ;
	wire _w14806_ ;
	wire _w14805_ ;
	wire _w14804_ ;
	wire _w14803_ ;
	wire _w14802_ ;
	wire _w14801_ ;
	wire _w14800_ ;
	wire _w14799_ ;
	wire _w14798_ ;
	wire _w14797_ ;
	wire _w14796_ ;
	wire _w14795_ ;
	wire _w14794_ ;
	wire _w14793_ ;
	wire _w14792_ ;
	wire _w14791_ ;
	wire _w14790_ ;
	wire _w14789_ ;
	wire _w14788_ ;
	wire _w14787_ ;
	wire _w14786_ ;
	wire _w14785_ ;
	wire _w14784_ ;
	wire _w14783_ ;
	wire _w14782_ ;
	wire _w14781_ ;
	wire _w14780_ ;
	wire _w14779_ ;
	wire _w14778_ ;
	wire _w14777_ ;
	wire _w14776_ ;
	wire _w14775_ ;
	wire _w14774_ ;
	wire _w14773_ ;
	wire _w14772_ ;
	wire _w14771_ ;
	wire _w14770_ ;
	wire _w14769_ ;
	wire _w14768_ ;
	wire _w14767_ ;
	wire _w14766_ ;
	wire _w14765_ ;
	wire _w14764_ ;
	wire _w14763_ ;
	wire _w14762_ ;
	wire _w14761_ ;
	wire _w14760_ ;
	wire _w14759_ ;
	wire _w14758_ ;
	wire _w14757_ ;
	wire _w14756_ ;
	wire _w14755_ ;
	wire _w14754_ ;
	wire _w14753_ ;
	wire _w14752_ ;
	wire _w14751_ ;
	wire _w14750_ ;
	wire _w14749_ ;
	wire _w14748_ ;
	wire _w14747_ ;
	wire _w14746_ ;
	wire _w14745_ ;
	wire _w14744_ ;
	wire _w14743_ ;
	wire _w14742_ ;
	wire _w14741_ ;
	wire _w14740_ ;
	wire _w14739_ ;
	wire _w14738_ ;
	wire _w14737_ ;
	wire _w14736_ ;
	wire _w14735_ ;
	wire _w14734_ ;
	wire _w14733_ ;
	wire _w14732_ ;
	wire _w14731_ ;
	wire _w14730_ ;
	wire _w14729_ ;
	wire _w14728_ ;
	wire _w14727_ ;
	wire _w14726_ ;
	wire _w14725_ ;
	wire _w14724_ ;
	wire _w14723_ ;
	wire _w14722_ ;
	wire _w14721_ ;
	wire _w14720_ ;
	wire _w14719_ ;
	wire _w14718_ ;
	wire _w14717_ ;
	wire _w14716_ ;
	wire _w14715_ ;
	wire _w14714_ ;
	wire _w14713_ ;
	wire _w14712_ ;
	wire _w14711_ ;
	wire _w14710_ ;
	wire _w14709_ ;
	wire _w14708_ ;
	wire _w14707_ ;
	wire _w14706_ ;
	wire _w14705_ ;
	wire _w14704_ ;
	wire _w14703_ ;
	wire _w14702_ ;
	wire _w14701_ ;
	wire _w14700_ ;
	wire _w14699_ ;
	wire _w14698_ ;
	wire _w14697_ ;
	wire _w14696_ ;
	wire _w14695_ ;
	wire _w14694_ ;
	wire _w14693_ ;
	wire _w14692_ ;
	wire _w14691_ ;
	wire _w14690_ ;
	wire _w14689_ ;
	wire _w14688_ ;
	wire _w14687_ ;
	wire _w14686_ ;
	wire _w14685_ ;
	wire _w14684_ ;
	wire _w14683_ ;
	wire _w14682_ ;
	wire _w14681_ ;
	wire _w14680_ ;
	wire _w14679_ ;
	wire _w14678_ ;
	wire _w14677_ ;
	wire _w14676_ ;
	wire _w14675_ ;
	wire _w14674_ ;
	wire _w14673_ ;
	wire _w14672_ ;
	wire _w14671_ ;
	wire _w14670_ ;
	wire _w14669_ ;
	wire _w14668_ ;
	wire _w14667_ ;
	wire _w14666_ ;
	wire _w14665_ ;
	wire _w14664_ ;
	wire _w14663_ ;
	wire _w14662_ ;
	wire _w14661_ ;
	wire _w14660_ ;
	wire _w14659_ ;
	wire _w14658_ ;
	wire _w14657_ ;
	wire _w14656_ ;
	wire _w14655_ ;
	wire _w14654_ ;
	wire _w14653_ ;
	wire _w14652_ ;
	wire _w14651_ ;
	wire _w14650_ ;
	wire _w14649_ ;
	wire _w14648_ ;
	wire _w14647_ ;
	wire _w14646_ ;
	wire _w14645_ ;
	wire _w14644_ ;
	wire _w14643_ ;
	wire _w14642_ ;
	wire _w14641_ ;
	wire _w14640_ ;
	wire _w14639_ ;
	wire _w14638_ ;
	wire _w14637_ ;
	wire _w14636_ ;
	wire _w14635_ ;
	wire _w14634_ ;
	wire _w14633_ ;
	wire _w14632_ ;
	wire _w14631_ ;
	wire _w14630_ ;
	wire _w14629_ ;
	wire _w14628_ ;
	wire _w14627_ ;
	wire _w14626_ ;
	wire _w14625_ ;
	wire _w14624_ ;
	wire _w14623_ ;
	wire _w14622_ ;
	wire _w14621_ ;
	wire _w14620_ ;
	wire _w14619_ ;
	wire _w14618_ ;
	wire _w14617_ ;
	wire _w14616_ ;
	wire _w14615_ ;
	wire _w14614_ ;
	wire _w14613_ ;
	wire _w14612_ ;
	wire _w14611_ ;
	wire _w14610_ ;
	wire _w14609_ ;
	wire _w14608_ ;
	wire _w14607_ ;
	wire _w14606_ ;
	wire _w14605_ ;
	wire _w14604_ ;
	wire _w14603_ ;
	wire _w14602_ ;
	wire _w14601_ ;
	wire _w14600_ ;
	wire _w14599_ ;
	wire _w14598_ ;
	wire _w14597_ ;
	wire _w14596_ ;
	wire _w14595_ ;
	wire _w14594_ ;
	wire _w14593_ ;
	wire _w14592_ ;
	wire _w14591_ ;
	wire _w14590_ ;
	wire _w14589_ ;
	wire _w14588_ ;
	wire _w14587_ ;
	wire _w14586_ ;
	wire _w14585_ ;
	wire _w14584_ ;
	wire _w14583_ ;
	wire _w14582_ ;
	wire _w14581_ ;
	wire _w14580_ ;
	wire _w14579_ ;
	wire _w14578_ ;
	wire _w14577_ ;
	wire _w14576_ ;
	wire _w14575_ ;
	wire _w14574_ ;
	wire _w14573_ ;
	wire _w14572_ ;
	wire _w14571_ ;
	wire _w14570_ ;
	wire _w14569_ ;
	wire _w14568_ ;
	wire _w14567_ ;
	wire _w14566_ ;
	wire _w14565_ ;
	wire _w14564_ ;
	wire _w14563_ ;
	wire _w14562_ ;
	wire _w14561_ ;
	wire _w14560_ ;
	wire _w14559_ ;
	wire _w14558_ ;
	wire _w14557_ ;
	wire _w14556_ ;
	wire _w14555_ ;
	wire _w14554_ ;
	wire _w14553_ ;
	wire _w14552_ ;
	wire _w14551_ ;
	wire _w14550_ ;
	wire _w14549_ ;
	wire _w14548_ ;
	wire _w14547_ ;
	wire _w14546_ ;
	wire _w14545_ ;
	wire _w14544_ ;
	wire _w14543_ ;
	wire _w14542_ ;
	wire _w14541_ ;
	wire _w14540_ ;
	wire _w14539_ ;
	wire _w14538_ ;
	wire _w14537_ ;
	wire _w14536_ ;
	wire _w14535_ ;
	wire _w14534_ ;
	wire _w14533_ ;
	wire _w14532_ ;
	wire _w14531_ ;
	wire _w14530_ ;
	wire _w14529_ ;
	wire _w14528_ ;
	wire _w14527_ ;
	wire _w14526_ ;
	wire _w14525_ ;
	wire _w14524_ ;
	wire _w14523_ ;
	wire _w14522_ ;
	wire _w14521_ ;
	wire _w14520_ ;
	wire _w14519_ ;
	wire _w14518_ ;
	wire _w14517_ ;
	wire _w14516_ ;
	wire _w14515_ ;
	wire _w14514_ ;
	wire _w14513_ ;
	wire _w14512_ ;
	wire _w14511_ ;
	wire _w14510_ ;
	wire _w14509_ ;
	wire _w14508_ ;
	wire _w14507_ ;
	wire _w14506_ ;
	wire _w14505_ ;
	wire _w14504_ ;
	wire _w14503_ ;
	wire _w14502_ ;
	wire _w14501_ ;
	wire _w14500_ ;
	wire _w14499_ ;
	wire _w14498_ ;
	wire _w14497_ ;
	wire _w14496_ ;
	wire _w14495_ ;
	wire _w14494_ ;
	wire _w14493_ ;
	wire _w14492_ ;
	wire _w14491_ ;
	wire _w14490_ ;
	wire _w14489_ ;
	wire _w14488_ ;
	wire _w14487_ ;
	wire _w14486_ ;
	wire _w14485_ ;
	wire _w14484_ ;
	wire _w14483_ ;
	wire _w14482_ ;
	wire _w14481_ ;
	wire _w14480_ ;
	wire _w14479_ ;
	wire _w14478_ ;
	wire _w14477_ ;
	wire _w14476_ ;
	wire _w14475_ ;
	wire _w14474_ ;
	wire _w14473_ ;
	wire _w14472_ ;
	wire _w14471_ ;
	wire _w14470_ ;
	wire _w14469_ ;
	wire _w14468_ ;
	wire _w14467_ ;
	wire _w14466_ ;
	wire _w14465_ ;
	wire _w14464_ ;
	wire _w14463_ ;
	wire _w14462_ ;
	wire _w14461_ ;
	wire _w14460_ ;
	wire _w14459_ ;
	wire _w14458_ ;
	wire _w14457_ ;
	wire _w14456_ ;
	wire _w14455_ ;
	wire _w14454_ ;
	wire _w14453_ ;
	wire _w14452_ ;
	wire _w14451_ ;
	wire _w14450_ ;
	wire _w14449_ ;
	wire _w14448_ ;
	wire _w14447_ ;
	wire _w14446_ ;
	wire _w14445_ ;
	wire _w14444_ ;
	wire _w14443_ ;
	wire _w14442_ ;
	wire _w14441_ ;
	wire _w14440_ ;
	wire _w14439_ ;
	wire _w14438_ ;
	wire _w14437_ ;
	wire _w14436_ ;
	wire _w14435_ ;
	wire _w14434_ ;
	wire _w14433_ ;
	wire _w14432_ ;
	wire _w14431_ ;
	wire _w14430_ ;
	wire _w14429_ ;
	wire _w14428_ ;
	wire _w14427_ ;
	wire _w14426_ ;
	wire _w14425_ ;
	wire _w14424_ ;
	wire _w14423_ ;
	wire _w14422_ ;
	wire _w14421_ ;
	wire _w14420_ ;
	wire _w14419_ ;
	wire _w14418_ ;
	wire _w14417_ ;
	wire _w14416_ ;
	wire _w14415_ ;
	wire _w14414_ ;
	wire _w14413_ ;
	wire _w14412_ ;
	wire _w14411_ ;
	wire _w14410_ ;
	wire _w14409_ ;
	wire _w14408_ ;
	wire _w14407_ ;
	wire _w14406_ ;
	wire _w14405_ ;
	wire _w14404_ ;
	wire _w14403_ ;
	wire _w14402_ ;
	wire _w14401_ ;
	wire _w14400_ ;
	wire _w14399_ ;
	wire _w14398_ ;
	wire _w14397_ ;
	wire _w14396_ ;
	wire _w14395_ ;
	wire _w14394_ ;
	wire _w14393_ ;
	wire _w14392_ ;
	wire _w14391_ ;
	wire _w14390_ ;
	wire _w14389_ ;
	wire _w14388_ ;
	wire _w14387_ ;
	wire _w14386_ ;
	wire _w14385_ ;
	wire _w14384_ ;
	wire _w14383_ ;
	wire _w14382_ ;
	wire _w14381_ ;
	wire _w14380_ ;
	wire _w14379_ ;
	wire _w14378_ ;
	wire _w14377_ ;
	wire _w14376_ ;
	wire _w14375_ ;
	wire _w14374_ ;
	wire _w14373_ ;
	wire _w14372_ ;
	wire _w14371_ ;
	wire _w14370_ ;
	wire _w14369_ ;
	wire _w14368_ ;
	wire _w14367_ ;
	wire _w14366_ ;
	wire _w14365_ ;
	wire _w14364_ ;
	wire _w14363_ ;
	wire _w14362_ ;
	wire _w14361_ ;
	wire _w14360_ ;
	wire _w14359_ ;
	wire _w14358_ ;
	wire _w14357_ ;
	wire _w14356_ ;
	wire _w14355_ ;
	wire _w14354_ ;
	wire _w14353_ ;
	wire _w14352_ ;
	wire _w14351_ ;
	wire _w14350_ ;
	wire _w14349_ ;
	wire _w14348_ ;
	wire _w14347_ ;
	wire _w14346_ ;
	wire _w14345_ ;
	wire _w14344_ ;
	wire _w14343_ ;
	wire _w14342_ ;
	wire _w14341_ ;
	wire _w14340_ ;
	wire _w14339_ ;
	wire _w14338_ ;
	wire _w14337_ ;
	wire _w14336_ ;
	wire _w14335_ ;
	wire _w14334_ ;
	wire _w14333_ ;
	wire _w14332_ ;
	wire _w14331_ ;
	wire _w14330_ ;
	wire _w14329_ ;
	wire _w14328_ ;
	wire _w14327_ ;
	wire _w14326_ ;
	wire _w14325_ ;
	wire _w14324_ ;
	wire _w14323_ ;
	wire _w14322_ ;
	wire _w14321_ ;
	wire _w14320_ ;
	wire _w14319_ ;
	wire _w14318_ ;
	wire _w14317_ ;
	wire _w14316_ ;
	wire _w14315_ ;
	wire _w14314_ ;
	wire _w14313_ ;
	wire _w14312_ ;
	wire _w14311_ ;
	wire _w14310_ ;
	wire _w14309_ ;
	wire _w14308_ ;
	wire _w14307_ ;
	wire _w14306_ ;
	wire _w14305_ ;
	wire _w14304_ ;
	wire _w14303_ ;
	wire _w14302_ ;
	wire _w14301_ ;
	wire _w14300_ ;
	wire _w14299_ ;
	wire _w14298_ ;
	wire _w14297_ ;
	wire _w14296_ ;
	wire _w14295_ ;
	wire _w14294_ ;
	wire _w14293_ ;
	wire _w14292_ ;
	wire _w14291_ ;
	wire _w14290_ ;
	wire _w14289_ ;
	wire _w14288_ ;
	wire _w14287_ ;
	wire _w14286_ ;
	wire _w14285_ ;
	wire _w14284_ ;
	wire _w14283_ ;
	wire _w14282_ ;
	wire _w14281_ ;
	wire _w14280_ ;
	wire _w14279_ ;
	wire _w14278_ ;
	wire _w14277_ ;
	wire _w14276_ ;
	wire _w14275_ ;
	wire _w14274_ ;
	wire _w14273_ ;
	wire _w14272_ ;
	wire _w14271_ ;
	wire _w14270_ ;
	wire _w14269_ ;
	wire _w14268_ ;
	wire _w14267_ ;
	wire _w14266_ ;
	wire _w14265_ ;
	wire _w14264_ ;
	wire _w14263_ ;
	wire _w14262_ ;
	wire _w14261_ ;
	wire _w14260_ ;
	wire _w14259_ ;
	wire _w14258_ ;
	wire _w14257_ ;
	wire _w14256_ ;
	wire _w14255_ ;
	wire _w14254_ ;
	wire _w14253_ ;
	wire _w14252_ ;
	wire _w14251_ ;
	wire _w14250_ ;
	wire _w14249_ ;
	wire _w14248_ ;
	wire _w14247_ ;
	wire _w14246_ ;
	wire _w14245_ ;
	wire _w14244_ ;
	wire _w14243_ ;
	wire _w14242_ ;
	wire _w14241_ ;
	wire _w14240_ ;
	wire _w14239_ ;
	wire _w14238_ ;
	wire _w14237_ ;
	wire _w14236_ ;
	wire _w14235_ ;
	wire _w14234_ ;
	wire _w14233_ ;
	wire _w14232_ ;
	wire _w14231_ ;
	wire _w14230_ ;
	wire _w14229_ ;
	wire _w14228_ ;
	wire _w14227_ ;
	wire _w14226_ ;
	wire _w14225_ ;
	wire _w14224_ ;
	wire _w14223_ ;
	wire _w14222_ ;
	wire _w14221_ ;
	wire _w14220_ ;
	wire _w14219_ ;
	wire _w14218_ ;
	wire _w14217_ ;
	wire _w14216_ ;
	wire _w14215_ ;
	wire _w14214_ ;
	wire _w14213_ ;
	wire _w14212_ ;
	wire _w14211_ ;
	wire _w14210_ ;
	wire _w14209_ ;
	wire _w14208_ ;
	wire _w14207_ ;
	wire _w14206_ ;
	wire _w14205_ ;
	wire _w14204_ ;
	wire _w14203_ ;
	wire _w14202_ ;
	wire _w14201_ ;
	wire _w14200_ ;
	wire _w14199_ ;
	wire _w14198_ ;
	wire _w14197_ ;
	wire _w14196_ ;
	wire _w14195_ ;
	wire _w14194_ ;
	wire _w14193_ ;
	wire _w14192_ ;
	wire _w14191_ ;
	wire _w14190_ ;
	wire _w14189_ ;
	wire _w14188_ ;
	wire _w14187_ ;
	wire _w14186_ ;
	wire _w14185_ ;
	wire _w14184_ ;
	wire _w14183_ ;
	wire _w14182_ ;
	wire _w14181_ ;
	wire _w14180_ ;
	wire _w14179_ ;
	wire _w14178_ ;
	wire _w14177_ ;
	wire _w14176_ ;
	wire _w14175_ ;
	wire _w14174_ ;
	wire _w14173_ ;
	wire _w14172_ ;
	wire _w14171_ ;
	wire _w14170_ ;
	wire _w14169_ ;
	wire _w14168_ ;
	wire _w14167_ ;
	wire _w14166_ ;
	wire _w14165_ ;
	wire _w14164_ ;
	wire _w14163_ ;
	wire _w14162_ ;
	wire _w14161_ ;
	wire _w14160_ ;
	wire _w14159_ ;
	wire _w14158_ ;
	wire _w14157_ ;
	wire _w14156_ ;
	wire _w14155_ ;
	wire _w14154_ ;
	wire _w14153_ ;
	wire _w14152_ ;
	wire _w14151_ ;
	wire _w14150_ ;
	wire _w14149_ ;
	wire _w14148_ ;
	wire _w14147_ ;
	wire _w14146_ ;
	wire _w14145_ ;
	wire _w14144_ ;
	wire _w14143_ ;
	wire _w14142_ ;
	wire _w14141_ ;
	wire _w14140_ ;
	wire _w14139_ ;
	wire _w14138_ ;
	wire _w14137_ ;
	wire _w14136_ ;
	wire _w14135_ ;
	wire _w14134_ ;
	wire _w14133_ ;
	wire _w14132_ ;
	wire _w14131_ ;
	wire _w14130_ ;
	wire _w14129_ ;
	wire _w14128_ ;
	wire _w14127_ ;
	wire _w14126_ ;
	wire _w14125_ ;
	wire _w14124_ ;
	wire _w14123_ ;
	wire _w14122_ ;
	wire _w14121_ ;
	wire _w14120_ ;
	wire _w14119_ ;
	wire _w14118_ ;
	wire _w14117_ ;
	wire _w14116_ ;
	wire _w14115_ ;
	wire _w14114_ ;
	wire _w14113_ ;
	wire _w14112_ ;
	wire _w14111_ ;
	wire _w14110_ ;
	wire _w14109_ ;
	wire _w14108_ ;
	wire _w14107_ ;
	wire _w14106_ ;
	wire _w14105_ ;
	wire _w14104_ ;
	wire _w14103_ ;
	wire _w14102_ ;
	wire _w14101_ ;
	wire _w14100_ ;
	wire _w14099_ ;
	wire _w14098_ ;
	wire _w14097_ ;
	wire _w14096_ ;
	wire _w14095_ ;
	wire _w14094_ ;
	wire _w14093_ ;
	wire _w14092_ ;
	wire _w14091_ ;
	wire _w14090_ ;
	wire _w14089_ ;
	wire _w14088_ ;
	wire _w14087_ ;
	wire _w14086_ ;
	wire _w14085_ ;
	wire _w14084_ ;
	wire _w14083_ ;
	wire _w14082_ ;
	wire _w14081_ ;
	wire _w14080_ ;
	wire _w14079_ ;
	wire _w14078_ ;
	wire _w14077_ ;
	wire _w14076_ ;
	wire _w14075_ ;
	wire _w14074_ ;
	wire _w14073_ ;
	wire _w14072_ ;
	wire _w14071_ ;
	wire _w14070_ ;
	wire _w14069_ ;
	wire _w14068_ ;
	wire _w14067_ ;
	wire _w14066_ ;
	wire _w14065_ ;
	wire _w14064_ ;
	wire _w14063_ ;
	wire _w14062_ ;
	wire _w14061_ ;
	wire _w14060_ ;
	wire _w14059_ ;
	wire _w14058_ ;
	wire _w14057_ ;
	wire _w14056_ ;
	wire _w14055_ ;
	wire _w14054_ ;
	wire _w14053_ ;
	wire _w14052_ ;
	wire _w14051_ ;
	wire _w14050_ ;
	wire _w14049_ ;
	wire _w14048_ ;
	wire _w14047_ ;
	wire _w14046_ ;
	wire _w14045_ ;
	wire _w14044_ ;
	wire _w14043_ ;
	wire _w14042_ ;
	wire _w14041_ ;
	wire _w14040_ ;
	wire _w14039_ ;
	wire _w14038_ ;
	wire _w14037_ ;
	wire _w14036_ ;
	wire _w14035_ ;
	wire _w14034_ ;
	wire _w14033_ ;
	wire _w14032_ ;
	wire _w14031_ ;
	wire _w14030_ ;
	wire _w14029_ ;
	wire _w14028_ ;
	wire _w14027_ ;
	wire _w14026_ ;
	wire _w14025_ ;
	wire _w14024_ ;
	wire _w14023_ ;
	wire _w14022_ ;
	wire _w14021_ ;
	wire _w14020_ ;
	wire _w14019_ ;
	wire _w14018_ ;
	wire _w14017_ ;
	wire _w14016_ ;
	wire _w14015_ ;
	wire _w14014_ ;
	wire _w14013_ ;
	wire _w14012_ ;
	wire _w14011_ ;
	wire _w14010_ ;
	wire _w14009_ ;
	wire _w14008_ ;
	wire _w14007_ ;
	wire _w14006_ ;
	wire _w14005_ ;
	wire _w14004_ ;
	wire _w14003_ ;
	wire _w14002_ ;
	wire _w14001_ ;
	wire _w14000_ ;
	wire _w13999_ ;
	wire _w13998_ ;
	wire _w13997_ ;
	wire _w13996_ ;
	wire _w13995_ ;
	wire _w13994_ ;
	wire _w13993_ ;
	wire _w13992_ ;
	wire _w13991_ ;
	wire _w13990_ ;
	wire _w13989_ ;
	wire _w13988_ ;
	wire _w13987_ ;
	wire _w13986_ ;
	wire _w13985_ ;
	wire _w13984_ ;
	wire _w13983_ ;
	wire _w13982_ ;
	wire _w13981_ ;
	wire _w13980_ ;
	wire _w13979_ ;
	wire _w13978_ ;
	wire _w13977_ ;
	wire _w13976_ ;
	wire _w13975_ ;
	wire _w13974_ ;
	wire _w13973_ ;
	wire _w13972_ ;
	wire _w13971_ ;
	wire _w13970_ ;
	wire _w13969_ ;
	wire _w13968_ ;
	wire _w13967_ ;
	wire _w13966_ ;
	wire _w13965_ ;
	wire _w13964_ ;
	wire _w13963_ ;
	wire _w13962_ ;
	wire _w13961_ ;
	wire _w13960_ ;
	wire _w13959_ ;
	wire _w13958_ ;
	wire _w13957_ ;
	wire _w13956_ ;
	wire _w13955_ ;
	wire _w13954_ ;
	wire _w13953_ ;
	wire _w13952_ ;
	wire _w13951_ ;
	wire _w13950_ ;
	wire _w13949_ ;
	wire _w13948_ ;
	wire _w13947_ ;
	wire _w13946_ ;
	wire _w13945_ ;
	wire _w13944_ ;
	wire _w13943_ ;
	wire _w13942_ ;
	wire _w13941_ ;
	wire _w13940_ ;
	wire _w13939_ ;
	wire _w13938_ ;
	wire _w13937_ ;
	wire _w13936_ ;
	wire _w13935_ ;
	wire _w13934_ ;
	wire _w13933_ ;
	wire _w13932_ ;
	wire _w13931_ ;
	wire _w13930_ ;
	wire _w13929_ ;
	wire _w13928_ ;
	wire _w13927_ ;
	wire _w13926_ ;
	wire _w13925_ ;
	wire _w13924_ ;
	wire _w13923_ ;
	wire _w13922_ ;
	wire _w13921_ ;
	wire _w13920_ ;
	wire _w13919_ ;
	wire _w13918_ ;
	wire _w13917_ ;
	wire _w13916_ ;
	wire _w13915_ ;
	wire _w13914_ ;
	wire _w13913_ ;
	wire _w13912_ ;
	wire _w13911_ ;
	wire _w13910_ ;
	wire _w13909_ ;
	wire _w13908_ ;
	wire _w13907_ ;
	wire _w13906_ ;
	wire _w13905_ ;
	wire _w13904_ ;
	wire _w13903_ ;
	wire _w13902_ ;
	wire _w13901_ ;
	wire _w13900_ ;
	wire _w13899_ ;
	wire _w13898_ ;
	wire _w13897_ ;
	wire _w13896_ ;
	wire _w13895_ ;
	wire _w13894_ ;
	wire _w13893_ ;
	wire _w13892_ ;
	wire _w13891_ ;
	wire _w13890_ ;
	wire _w13889_ ;
	wire _w13888_ ;
	wire _w13887_ ;
	wire _w13886_ ;
	wire _w13885_ ;
	wire _w13884_ ;
	wire _w13883_ ;
	wire _w13882_ ;
	wire _w13881_ ;
	wire _w13880_ ;
	wire _w13879_ ;
	wire _w13878_ ;
	wire _w13877_ ;
	wire _w13876_ ;
	wire _w13875_ ;
	wire _w13874_ ;
	wire _w13873_ ;
	wire _w13872_ ;
	wire _w13871_ ;
	wire _w13870_ ;
	wire _w13869_ ;
	wire _w13868_ ;
	wire _w13867_ ;
	wire _w13866_ ;
	wire _w13865_ ;
	wire _w13864_ ;
	wire _w13863_ ;
	wire _w13862_ ;
	wire _w13861_ ;
	wire _w13860_ ;
	wire _w13859_ ;
	wire _w13858_ ;
	wire _w13857_ ;
	wire _w13856_ ;
	wire _w13855_ ;
	wire _w13854_ ;
	wire _w13853_ ;
	wire _w13852_ ;
	wire _w13851_ ;
	wire _w13850_ ;
	wire _w13849_ ;
	wire _w13848_ ;
	wire _w13847_ ;
	wire _w13846_ ;
	wire _w13845_ ;
	wire _w13844_ ;
	wire _w13843_ ;
	wire _w13842_ ;
	wire _w13841_ ;
	wire _w13840_ ;
	wire _w13839_ ;
	wire _w13838_ ;
	wire _w13837_ ;
	wire _w13836_ ;
	wire _w13835_ ;
	wire _w13834_ ;
	wire _w13833_ ;
	wire _w13832_ ;
	wire _w13831_ ;
	wire _w13830_ ;
	wire _w13829_ ;
	wire _w13828_ ;
	wire _w13827_ ;
	wire _w13826_ ;
	wire _w13825_ ;
	wire _w13824_ ;
	wire _w13823_ ;
	wire _w13822_ ;
	wire _w13821_ ;
	wire _w13820_ ;
	wire _w13819_ ;
	wire _w13818_ ;
	wire _w13817_ ;
	wire _w13816_ ;
	wire _w13815_ ;
	wire _w13814_ ;
	wire _w13813_ ;
	wire _w13812_ ;
	wire _w13811_ ;
	wire _w13810_ ;
	wire _w13809_ ;
	wire _w13808_ ;
	wire _w13807_ ;
	wire _w13806_ ;
	wire _w13805_ ;
	wire _w13804_ ;
	wire _w13803_ ;
	wire _w13802_ ;
	wire _w13801_ ;
	wire _w13800_ ;
	wire _w13799_ ;
	wire _w13798_ ;
	wire _w13797_ ;
	wire _w13796_ ;
	wire _w13795_ ;
	wire _w13794_ ;
	wire _w13793_ ;
	wire _w13792_ ;
	wire _w13791_ ;
	wire _w13790_ ;
	wire _w13789_ ;
	wire _w13788_ ;
	wire _w13787_ ;
	wire _w13786_ ;
	wire _w13785_ ;
	wire _w13784_ ;
	wire _w13783_ ;
	wire _w13782_ ;
	wire _w13781_ ;
	wire _w13780_ ;
	wire _w13779_ ;
	wire _w13778_ ;
	wire _w13777_ ;
	wire _w13776_ ;
	wire _w13775_ ;
	wire _w13774_ ;
	wire _w13773_ ;
	wire _w13772_ ;
	wire _w13771_ ;
	wire _w13770_ ;
	wire _w13769_ ;
	wire _w13768_ ;
	wire _w13767_ ;
	wire _w13766_ ;
	wire _w13765_ ;
	wire _w13764_ ;
	wire _w13763_ ;
	wire _w13762_ ;
	wire _w13761_ ;
	wire _w13760_ ;
	wire _w13759_ ;
	wire _w13758_ ;
	wire _w13757_ ;
	wire _w13756_ ;
	wire _w13755_ ;
	wire _w13754_ ;
	wire _w13753_ ;
	wire _w13752_ ;
	wire _w13751_ ;
	wire _w13750_ ;
	wire _w13749_ ;
	wire _w13748_ ;
	wire _w13747_ ;
	wire _w13746_ ;
	wire _w13745_ ;
	wire _w13744_ ;
	wire _w13743_ ;
	wire _w13742_ ;
	wire _w13741_ ;
	wire _w13740_ ;
	wire _w13739_ ;
	wire _w13738_ ;
	wire _w13737_ ;
	wire _w13736_ ;
	wire _w13735_ ;
	wire _w13734_ ;
	wire _w13733_ ;
	wire _w13732_ ;
	wire _w13731_ ;
	wire _w13730_ ;
	wire _w13729_ ;
	wire _w13728_ ;
	wire _w13727_ ;
	wire _w13726_ ;
	wire _w13725_ ;
	wire _w13724_ ;
	wire _w13723_ ;
	wire _w13722_ ;
	wire _w13721_ ;
	wire _w13720_ ;
	wire _w13719_ ;
	wire _w13718_ ;
	wire _w13717_ ;
	wire _w13716_ ;
	wire _w13715_ ;
	wire _w13714_ ;
	wire _w13713_ ;
	wire _w13712_ ;
	wire _w13711_ ;
	wire _w13710_ ;
	wire _w13709_ ;
	wire _w13708_ ;
	wire _w13707_ ;
	wire _w13706_ ;
	wire _w13705_ ;
	wire _w13704_ ;
	wire _w13703_ ;
	wire _w13702_ ;
	wire _w13701_ ;
	wire _w13700_ ;
	wire _w13699_ ;
	wire _w13698_ ;
	wire _w13697_ ;
	wire _w13696_ ;
	wire _w13695_ ;
	wire _w13694_ ;
	wire _w13693_ ;
	wire _w13692_ ;
	wire _w13691_ ;
	wire _w13690_ ;
	wire _w13689_ ;
	wire _w13688_ ;
	wire _w13687_ ;
	wire _w13686_ ;
	wire _w13685_ ;
	wire _w13684_ ;
	wire _w13683_ ;
	wire _w13682_ ;
	wire _w13681_ ;
	wire _w13680_ ;
	wire _w13679_ ;
	wire _w13678_ ;
	wire _w13677_ ;
	wire _w13676_ ;
	wire _w13675_ ;
	wire _w13674_ ;
	wire _w13673_ ;
	wire _w13672_ ;
	wire _w13671_ ;
	wire _w13670_ ;
	wire _w13669_ ;
	wire _w13668_ ;
	wire _w13667_ ;
	wire _w13666_ ;
	wire _w13665_ ;
	wire _w13664_ ;
	wire _w13663_ ;
	wire _w13662_ ;
	wire _w13661_ ;
	wire _w13660_ ;
	wire _w13659_ ;
	wire _w13658_ ;
	wire _w13657_ ;
	wire _w13656_ ;
	wire _w13655_ ;
	wire _w13654_ ;
	wire _w13653_ ;
	wire _w13652_ ;
	wire _w13651_ ;
	wire _w13650_ ;
	wire _w13649_ ;
	wire _w13648_ ;
	wire _w13647_ ;
	wire _w13646_ ;
	wire _w13645_ ;
	wire _w13644_ ;
	wire _w13643_ ;
	wire _w13642_ ;
	wire _w13641_ ;
	wire _w13640_ ;
	wire _w13639_ ;
	wire _w13638_ ;
	wire _w13637_ ;
	wire _w13636_ ;
	wire _w13635_ ;
	wire _w13634_ ;
	wire _w13633_ ;
	wire _w13632_ ;
	wire _w13631_ ;
	wire _w13630_ ;
	wire _w13629_ ;
	wire _w13628_ ;
	wire _w13627_ ;
	wire _w13626_ ;
	wire _w13625_ ;
	wire _w13624_ ;
	wire _w13623_ ;
	wire _w13622_ ;
	wire _w13621_ ;
	wire _w13620_ ;
	wire _w13619_ ;
	wire _w13618_ ;
	wire _w13617_ ;
	wire _w13616_ ;
	wire _w13615_ ;
	wire _w13614_ ;
	wire _w13613_ ;
	wire _w13612_ ;
	wire _w13611_ ;
	wire _w13610_ ;
	wire _w13609_ ;
	wire _w13608_ ;
	wire _w13607_ ;
	wire _w13606_ ;
	wire _w13605_ ;
	wire _w13604_ ;
	wire _w13603_ ;
	wire _w13602_ ;
	wire _w13601_ ;
	wire _w13600_ ;
	wire _w13599_ ;
	wire _w13598_ ;
	wire _w13597_ ;
	wire _w13596_ ;
	wire _w13595_ ;
	wire _w13594_ ;
	wire _w13593_ ;
	wire _w13592_ ;
	wire _w13591_ ;
	wire _w13590_ ;
	wire _w13589_ ;
	wire _w13588_ ;
	wire _w13587_ ;
	wire _w13586_ ;
	wire _w13585_ ;
	wire _w13584_ ;
	wire _w13583_ ;
	wire _w13582_ ;
	wire _w13581_ ;
	wire _w13580_ ;
	wire _w13579_ ;
	wire _w13578_ ;
	wire _w13577_ ;
	wire _w13576_ ;
	wire _w13575_ ;
	wire _w13574_ ;
	wire _w13573_ ;
	wire _w13572_ ;
	wire _w13571_ ;
	wire _w13570_ ;
	wire _w13569_ ;
	wire _w13568_ ;
	wire _w13567_ ;
	wire _w13566_ ;
	wire _w13565_ ;
	wire _w13564_ ;
	wire _w13563_ ;
	wire _w13562_ ;
	wire _w13561_ ;
	wire _w13560_ ;
	wire _w13559_ ;
	wire _w13558_ ;
	wire _w13557_ ;
	wire _w13556_ ;
	wire _w13555_ ;
	wire _w13554_ ;
	wire _w13553_ ;
	wire _w13552_ ;
	wire _w13551_ ;
	wire _w13550_ ;
	wire _w13549_ ;
	wire _w13548_ ;
	wire _w13547_ ;
	wire _w13546_ ;
	wire _w13545_ ;
	wire _w13544_ ;
	wire _w13543_ ;
	wire _w13542_ ;
	wire _w13541_ ;
	wire _w13540_ ;
	wire _w13539_ ;
	wire _w13538_ ;
	wire _w13537_ ;
	wire _w13536_ ;
	wire _w13535_ ;
	wire _w13534_ ;
	wire _w13533_ ;
	wire _w13532_ ;
	wire _w13531_ ;
	wire _w13530_ ;
	wire _w13529_ ;
	wire _w13528_ ;
	wire _w13527_ ;
	wire _w13526_ ;
	wire _w13525_ ;
	wire _w13524_ ;
	wire _w13523_ ;
	wire _w13522_ ;
	wire _w13521_ ;
	wire _w13520_ ;
	wire _w13519_ ;
	wire _w13518_ ;
	wire _w13517_ ;
	wire _w13516_ ;
	wire _w13515_ ;
	wire _w13514_ ;
	wire _w13513_ ;
	wire _w13512_ ;
	wire _w13511_ ;
	wire _w13510_ ;
	wire _w13509_ ;
	wire _w13508_ ;
	wire _w13507_ ;
	wire _w13506_ ;
	wire _w13505_ ;
	wire _w13504_ ;
	wire _w13503_ ;
	wire _w13502_ ;
	wire _w13501_ ;
	wire _w13500_ ;
	wire _w13499_ ;
	wire _w13498_ ;
	wire _w13497_ ;
	wire _w13496_ ;
	wire _w13495_ ;
	wire _w13494_ ;
	wire _w13493_ ;
	wire _w13492_ ;
	wire _w13491_ ;
	wire _w13490_ ;
	wire _w13489_ ;
	wire _w13488_ ;
	wire _w13487_ ;
	wire _w13486_ ;
	wire _w13485_ ;
	wire _w13484_ ;
	wire _w13483_ ;
	wire _w13482_ ;
	wire _w13481_ ;
	wire _w13480_ ;
	wire _w13479_ ;
	wire _w13478_ ;
	wire _w13477_ ;
	wire _w13476_ ;
	wire _w13475_ ;
	wire _w13474_ ;
	wire _w13473_ ;
	wire _w13472_ ;
	wire _w13471_ ;
	wire _w13470_ ;
	wire _w13469_ ;
	wire _w13468_ ;
	wire _w13467_ ;
	wire _w13466_ ;
	wire _w13465_ ;
	wire _w13464_ ;
	wire _w13463_ ;
	wire _w13462_ ;
	wire _w13461_ ;
	wire _w13460_ ;
	wire _w13459_ ;
	wire _w13458_ ;
	wire _w13457_ ;
	wire _w13456_ ;
	wire _w13455_ ;
	wire _w13454_ ;
	wire _w13453_ ;
	wire _w13452_ ;
	wire _w13451_ ;
	wire _w13450_ ;
	wire _w13449_ ;
	wire _w13448_ ;
	wire _w13447_ ;
	wire _w13446_ ;
	wire _w13445_ ;
	wire _w13444_ ;
	wire _w13443_ ;
	wire _w13442_ ;
	wire _w13441_ ;
	wire _w13440_ ;
	wire _w13439_ ;
	wire _w13438_ ;
	wire _w13437_ ;
	wire _w13436_ ;
	wire _w13435_ ;
	wire _w13434_ ;
	wire _w13433_ ;
	wire _w13432_ ;
	wire _w13431_ ;
	wire _w13430_ ;
	wire _w13429_ ;
	wire _w13428_ ;
	wire _w13427_ ;
	wire _w13426_ ;
	wire _w13425_ ;
	wire _w13424_ ;
	wire _w13423_ ;
	wire _w13422_ ;
	wire _w13421_ ;
	wire _w13420_ ;
	wire _w13419_ ;
	wire _w13418_ ;
	wire _w13417_ ;
	wire _w13416_ ;
	wire _w13415_ ;
	wire _w13414_ ;
	wire _w13413_ ;
	wire _w13412_ ;
	wire _w13411_ ;
	wire _w13410_ ;
	wire _w13409_ ;
	wire _w13408_ ;
	wire _w13407_ ;
	wire _w13406_ ;
	wire _w13405_ ;
	wire _w13404_ ;
	wire _w13403_ ;
	wire _w13402_ ;
	wire _w13401_ ;
	wire _w13400_ ;
	wire _w13399_ ;
	wire _w13398_ ;
	wire _w13397_ ;
	wire _w13396_ ;
	wire _w13395_ ;
	wire _w13394_ ;
	wire _w13393_ ;
	wire _w13392_ ;
	wire _w13391_ ;
	wire _w13390_ ;
	wire _w13389_ ;
	wire _w13388_ ;
	wire _w13387_ ;
	wire _w13386_ ;
	wire _w13385_ ;
	wire _w13384_ ;
	wire _w13383_ ;
	wire _w13382_ ;
	wire _w13381_ ;
	wire _w13380_ ;
	wire _w13379_ ;
	wire _w13378_ ;
	wire _w13377_ ;
	wire _w13376_ ;
	wire _w13375_ ;
	wire _w13374_ ;
	wire _w13373_ ;
	wire _w13372_ ;
	wire _w13371_ ;
	wire _w13370_ ;
	wire _w13369_ ;
	wire _w13368_ ;
	wire _w13367_ ;
	wire _w13366_ ;
	wire _w13365_ ;
	wire _w13364_ ;
	wire _w13363_ ;
	wire _w13362_ ;
	wire _w13361_ ;
	wire _w13360_ ;
	wire _w13359_ ;
	wire _w13358_ ;
	wire _w13357_ ;
	wire _w13356_ ;
	wire _w13355_ ;
	wire _w13354_ ;
	wire _w13353_ ;
	wire _w13352_ ;
	wire _w13351_ ;
	wire _w13350_ ;
	wire _w13349_ ;
	wire _w13348_ ;
	wire _w13347_ ;
	wire _w13346_ ;
	wire _w13345_ ;
	wire _w13344_ ;
	wire _w13343_ ;
	wire _w13342_ ;
	wire _w13341_ ;
	wire _w13340_ ;
	wire _w13339_ ;
	wire _w13338_ ;
	wire _w13337_ ;
	wire _w13336_ ;
	wire _w13335_ ;
	wire _w13334_ ;
	wire _w13333_ ;
	wire _w13332_ ;
	wire _w13331_ ;
	wire _w13330_ ;
	wire _w13329_ ;
	wire _w13328_ ;
	wire _w13327_ ;
	wire _w13326_ ;
	wire _w13325_ ;
	wire _w13324_ ;
	wire _w13323_ ;
	wire _w13322_ ;
	wire _w13321_ ;
	wire _w13320_ ;
	wire _w13319_ ;
	wire _w13318_ ;
	wire _w13317_ ;
	wire _w13316_ ;
	wire _w13315_ ;
	wire _w13314_ ;
	wire _w13313_ ;
	wire _w13312_ ;
	wire _w13311_ ;
	wire _w13310_ ;
	wire _w13309_ ;
	wire _w13308_ ;
	wire _w13307_ ;
	wire _w13306_ ;
	wire _w13305_ ;
	wire _w13304_ ;
	wire _w13303_ ;
	wire _w13302_ ;
	wire _w13301_ ;
	wire _w13300_ ;
	wire _w13299_ ;
	wire _w13298_ ;
	wire _w13297_ ;
	wire _w13296_ ;
	wire _w13295_ ;
	wire _w13294_ ;
	wire _w13293_ ;
	wire _w13292_ ;
	wire _w13291_ ;
	wire _w13290_ ;
	wire _w13289_ ;
	wire _w13288_ ;
	wire _w13287_ ;
	wire _w13286_ ;
	wire _w13285_ ;
	wire _w13284_ ;
	wire _w13283_ ;
	wire _w13282_ ;
	wire _w13281_ ;
	wire _w13280_ ;
	wire _w13279_ ;
	wire _w13278_ ;
	wire _w13277_ ;
	wire _w13276_ ;
	wire _w13275_ ;
	wire _w13274_ ;
	wire _w13273_ ;
	wire _w13272_ ;
	wire _w13271_ ;
	wire _w13270_ ;
	wire _w13269_ ;
	wire _w13268_ ;
	wire _w13267_ ;
	wire _w13266_ ;
	wire _w13265_ ;
	wire _w13264_ ;
	wire _w13263_ ;
	wire _w13262_ ;
	wire _w13261_ ;
	wire _w13260_ ;
	wire _w13259_ ;
	wire _w13258_ ;
	wire _w13257_ ;
	wire _w13256_ ;
	wire _w13255_ ;
	wire _w13254_ ;
	wire _w13253_ ;
	wire _w13252_ ;
	wire _w13251_ ;
	wire _w13250_ ;
	wire _w13249_ ;
	wire _w13248_ ;
	wire _w13247_ ;
	wire _w13246_ ;
	wire _w13245_ ;
	wire _w13244_ ;
	wire _w13243_ ;
	wire _w13242_ ;
	wire _w13241_ ;
	wire _w13240_ ;
	wire _w13239_ ;
	wire _w13238_ ;
	wire _w13237_ ;
	wire _w13236_ ;
	wire _w13235_ ;
	wire _w13234_ ;
	wire _w13233_ ;
	wire _w13232_ ;
	wire _w13231_ ;
	wire _w13230_ ;
	wire _w13229_ ;
	wire _w13228_ ;
	wire _w13227_ ;
	wire _w13226_ ;
	wire _w13225_ ;
	wire _w13224_ ;
	wire _w13223_ ;
	wire _w13222_ ;
	wire _w13221_ ;
	wire _w13220_ ;
	wire _w13219_ ;
	wire _w13218_ ;
	wire _w13217_ ;
	wire _w13216_ ;
	wire _w13215_ ;
	wire _w13214_ ;
	wire _w13213_ ;
	wire _w13212_ ;
	wire _w13211_ ;
	wire _w13210_ ;
	wire _w13209_ ;
	wire _w13208_ ;
	wire _w13207_ ;
	wire _w13206_ ;
	wire _w13205_ ;
	wire _w13204_ ;
	wire _w13203_ ;
	wire _w13202_ ;
	wire _w13201_ ;
	wire _w13200_ ;
	wire _w13199_ ;
	wire _w13198_ ;
	wire _w13197_ ;
	wire _w13196_ ;
	wire _w13195_ ;
	wire _w13194_ ;
	wire _w13193_ ;
	wire _w13192_ ;
	wire _w13191_ ;
	wire _w13190_ ;
	wire _w13189_ ;
	wire _w13188_ ;
	wire _w13187_ ;
	wire _w13186_ ;
	wire _w13185_ ;
	wire _w13184_ ;
	wire _w13183_ ;
	wire _w13182_ ;
	wire _w13181_ ;
	wire _w13180_ ;
	wire _w13179_ ;
	wire _w13178_ ;
	wire _w13177_ ;
	wire _w13176_ ;
	wire _w13175_ ;
	wire _w13174_ ;
	wire _w13173_ ;
	wire _w13172_ ;
	wire _w13171_ ;
	wire _w13170_ ;
	wire _w13169_ ;
	wire _w13168_ ;
	wire _w13167_ ;
	wire _w13166_ ;
	wire _w13165_ ;
	wire _w13164_ ;
	wire _w13163_ ;
	wire _w13162_ ;
	wire _w13161_ ;
	wire _w13160_ ;
	wire _w13159_ ;
	wire _w13158_ ;
	wire _w13157_ ;
	wire _w13156_ ;
	wire _w13155_ ;
	wire _w13154_ ;
	wire _w13153_ ;
	wire _w13152_ ;
	wire _w13151_ ;
	wire _w13150_ ;
	wire _w13149_ ;
	wire _w13148_ ;
	wire _w13147_ ;
	wire _w13146_ ;
	wire _w13145_ ;
	wire _w13144_ ;
	wire _w13143_ ;
	wire _w13142_ ;
	wire _w13141_ ;
	wire _w13140_ ;
	wire _w13139_ ;
	wire _w13138_ ;
	wire _w13137_ ;
	wire _w13136_ ;
	wire _w13135_ ;
	wire _w13134_ ;
	wire _w13133_ ;
	wire _w13132_ ;
	wire _w13131_ ;
	wire _w13130_ ;
	wire _w13129_ ;
	wire _w13128_ ;
	wire _w13127_ ;
	wire _w13126_ ;
	wire _w13125_ ;
	wire _w13124_ ;
	wire _w13123_ ;
	wire _w13122_ ;
	wire _w13121_ ;
	wire _w13120_ ;
	wire _w13119_ ;
	wire _w13118_ ;
	wire _w13117_ ;
	wire _w13116_ ;
	wire _w13115_ ;
	wire _w13114_ ;
	wire _w13113_ ;
	wire _w13112_ ;
	wire _w13111_ ;
	wire _w13110_ ;
	wire _w13109_ ;
	wire _w13108_ ;
	wire _w13107_ ;
	wire _w13106_ ;
	wire _w13105_ ;
	wire _w13104_ ;
	wire _w13103_ ;
	wire _w13102_ ;
	wire _w13101_ ;
	wire _w13100_ ;
	wire _w13099_ ;
	wire _w13098_ ;
	wire _w13097_ ;
	wire _w13096_ ;
	wire _w13095_ ;
	wire _w13094_ ;
	wire _w13093_ ;
	wire _w13092_ ;
	wire _w13091_ ;
	wire _w13090_ ;
	wire _w13089_ ;
	wire _w13088_ ;
	wire _w13087_ ;
	wire _w13086_ ;
	wire _w13085_ ;
	wire _w13084_ ;
	wire _w13083_ ;
	wire _w13082_ ;
	wire _w13081_ ;
	wire _w13080_ ;
	wire _w13079_ ;
	wire _w13078_ ;
	wire _w13077_ ;
	wire _w13076_ ;
	wire _w13075_ ;
	wire _w13074_ ;
	wire _w13073_ ;
	wire _w13072_ ;
	wire _w13071_ ;
	wire _w13070_ ;
	wire _w13069_ ;
	wire _w13068_ ;
	wire _w13067_ ;
	wire _w13066_ ;
	wire _w13065_ ;
	wire _w13064_ ;
	wire _w13063_ ;
	wire _w13062_ ;
	wire _w13061_ ;
	wire _w13060_ ;
	wire _w13059_ ;
	wire _w13058_ ;
	wire _w13057_ ;
	wire _w13056_ ;
	wire _w13055_ ;
	wire _w13054_ ;
	wire _w13053_ ;
	wire _w13052_ ;
	wire _w13051_ ;
	wire _w13050_ ;
	wire _w13049_ ;
	wire _w13048_ ;
	wire _w13047_ ;
	wire _w13046_ ;
	wire _w13045_ ;
	wire _w13044_ ;
	wire _w13043_ ;
	wire _w13042_ ;
	wire _w13041_ ;
	wire _w13040_ ;
	wire _w13039_ ;
	wire _w13038_ ;
	wire _w13037_ ;
	wire _w13036_ ;
	wire _w13035_ ;
	wire _w13034_ ;
	wire _w13033_ ;
	wire _w13032_ ;
	wire _w13031_ ;
	wire _w13030_ ;
	wire _w13029_ ;
	wire _w13028_ ;
	wire _w13027_ ;
	wire _w13026_ ;
	wire _w13025_ ;
	wire _w13024_ ;
	wire _w13023_ ;
	wire _w13022_ ;
	wire _w13021_ ;
	wire _w13020_ ;
	wire _w13019_ ;
	wire _w13018_ ;
	wire _w13017_ ;
	wire _w13016_ ;
	wire _w13015_ ;
	wire _w13014_ ;
	wire _w13013_ ;
	wire _w13012_ ;
	wire _w13011_ ;
	wire _w13010_ ;
	wire _w13009_ ;
	wire _w13008_ ;
	wire _w13007_ ;
	wire _w13006_ ;
	wire _w13005_ ;
	wire _w13004_ ;
	wire _w13003_ ;
	wire _w13002_ ;
	wire _w13001_ ;
	wire _w13000_ ;
	wire _w12999_ ;
	wire _w12998_ ;
	wire _w12997_ ;
	wire _w12996_ ;
	wire _w12995_ ;
	wire _w12994_ ;
	wire _w12993_ ;
	wire _w12992_ ;
	wire _w12991_ ;
	wire _w12990_ ;
	wire _w12989_ ;
	wire _w12988_ ;
	wire _w12987_ ;
	wire _w12986_ ;
	wire _w12985_ ;
	wire _w12984_ ;
	wire _w12983_ ;
	wire _w12982_ ;
	wire _w12981_ ;
	wire _w12980_ ;
	wire _w12979_ ;
	wire _w12978_ ;
	wire _w12977_ ;
	wire _w12976_ ;
	wire _w12975_ ;
	wire _w12974_ ;
	wire _w12973_ ;
	wire _w12972_ ;
	wire _w12971_ ;
	wire _w12970_ ;
	wire _w12969_ ;
	wire _w12968_ ;
	wire _w12967_ ;
	wire _w12966_ ;
	wire _w12965_ ;
	wire _w12964_ ;
	wire _w12963_ ;
	wire _w12962_ ;
	wire _w12961_ ;
	wire _w12960_ ;
	wire _w12959_ ;
	wire _w12958_ ;
	wire _w12957_ ;
	wire _w12956_ ;
	wire _w12955_ ;
	wire _w12954_ ;
	wire _w12953_ ;
	wire _w12952_ ;
	wire _w12951_ ;
	wire _w12950_ ;
	wire _w12949_ ;
	wire _w12948_ ;
	wire _w12947_ ;
	wire _w12946_ ;
	wire _w12945_ ;
	wire _w12944_ ;
	wire _w12943_ ;
	wire _w12942_ ;
	wire _w12941_ ;
	wire _w12940_ ;
	wire _w12939_ ;
	wire _w12938_ ;
	wire _w12937_ ;
	wire _w12936_ ;
	wire _w12935_ ;
	wire _w12934_ ;
	wire _w12933_ ;
	wire _w12932_ ;
	wire _w12931_ ;
	wire _w12930_ ;
	wire _w12929_ ;
	wire _w12928_ ;
	wire _w12927_ ;
	wire _w12926_ ;
	wire _w12925_ ;
	wire _w12924_ ;
	wire _w12923_ ;
	wire _w12922_ ;
	wire _w12921_ ;
	wire _w12920_ ;
	wire _w12919_ ;
	wire _w12918_ ;
	wire _w12917_ ;
	wire _w12916_ ;
	wire _w12915_ ;
	wire _w12914_ ;
	wire _w12913_ ;
	wire _w12912_ ;
	wire _w12911_ ;
	wire _w12910_ ;
	wire _w12909_ ;
	wire _w12908_ ;
	wire _w12907_ ;
	wire _w12906_ ;
	wire _w12905_ ;
	wire _w12904_ ;
	wire _w12903_ ;
	wire _w12902_ ;
	wire _w12901_ ;
	wire _w12900_ ;
	wire _w12899_ ;
	wire _w12898_ ;
	wire _w12897_ ;
	wire _w12896_ ;
	wire _w12895_ ;
	wire _w12894_ ;
	wire _w12893_ ;
	wire _w12892_ ;
	wire _w12891_ ;
	wire _w12890_ ;
	wire _w12889_ ;
	wire _w12888_ ;
	wire _w12887_ ;
	wire _w12886_ ;
	wire _w12885_ ;
	wire _w12884_ ;
	wire _w12883_ ;
	wire _w12882_ ;
	wire _w12881_ ;
	wire _w12880_ ;
	wire _w12879_ ;
	wire _w12878_ ;
	wire _w12877_ ;
	wire _w12876_ ;
	wire _w12875_ ;
	wire _w12874_ ;
	wire _w12873_ ;
	wire _w12872_ ;
	wire _w12871_ ;
	wire _w12870_ ;
	wire _w12869_ ;
	wire _w12868_ ;
	wire _w12867_ ;
	wire _w12866_ ;
	wire _w12865_ ;
	wire _w12864_ ;
	wire _w12863_ ;
	wire _w12862_ ;
	wire _w12861_ ;
	wire _w12860_ ;
	wire _w12859_ ;
	wire _w12858_ ;
	wire _w12857_ ;
	wire _w12856_ ;
	wire _w12855_ ;
	wire _w12854_ ;
	wire _w12853_ ;
	wire _w12852_ ;
	wire _w12851_ ;
	wire _w12850_ ;
	wire _w12849_ ;
	wire _w12848_ ;
	wire _w12847_ ;
	wire _w12846_ ;
	wire _w12845_ ;
	wire _w12844_ ;
	wire _w12843_ ;
	wire _w12842_ ;
	wire _w12841_ ;
	wire _w12840_ ;
	wire _w12839_ ;
	wire _w12838_ ;
	wire _w12837_ ;
	wire _w12836_ ;
	wire _w12835_ ;
	wire _w12834_ ;
	wire _w12833_ ;
	wire _w12832_ ;
	wire _w12831_ ;
	wire _w12830_ ;
	wire _w12829_ ;
	wire _w12828_ ;
	wire _w12827_ ;
	wire _w12826_ ;
	wire _w12825_ ;
	wire _w12824_ ;
	wire _w12823_ ;
	wire _w12822_ ;
	wire _w12821_ ;
	wire _w12820_ ;
	wire _w12819_ ;
	wire _w12818_ ;
	wire _w12817_ ;
	wire _w12816_ ;
	wire _w12815_ ;
	wire _w12814_ ;
	wire _w12813_ ;
	wire _w12812_ ;
	wire _w12811_ ;
	wire _w12810_ ;
	wire _w12809_ ;
	wire _w12808_ ;
	wire _w12807_ ;
	wire _w12806_ ;
	wire _w12805_ ;
	wire _w12804_ ;
	wire _w12803_ ;
	wire _w12802_ ;
	wire _w12801_ ;
	wire _w12800_ ;
	wire _w12799_ ;
	wire _w12798_ ;
	wire _w12797_ ;
	wire _w12796_ ;
	wire _w12795_ ;
	wire _w12794_ ;
	wire _w12793_ ;
	wire _w12792_ ;
	wire _w12791_ ;
	wire _w12790_ ;
	wire _w12789_ ;
	wire _w12788_ ;
	wire _w12787_ ;
	wire _w12786_ ;
	wire _w12785_ ;
	wire _w12784_ ;
	wire _w12783_ ;
	wire _w12782_ ;
	wire _w12781_ ;
	wire _w12780_ ;
	wire _w12779_ ;
	wire _w12778_ ;
	wire _w12777_ ;
	wire _w12776_ ;
	wire _w12775_ ;
	wire _w12774_ ;
	wire _w12773_ ;
	wire _w12772_ ;
	wire _w12771_ ;
	wire _w12770_ ;
	wire _w12769_ ;
	wire _w12768_ ;
	wire _w12767_ ;
	wire _w12766_ ;
	wire _w12765_ ;
	wire _w12764_ ;
	wire _w12763_ ;
	wire _w12762_ ;
	wire _w12761_ ;
	wire _w12760_ ;
	wire _w12759_ ;
	wire _w12758_ ;
	wire _w12757_ ;
	wire _w12756_ ;
	wire _w12755_ ;
	wire _w12754_ ;
	wire _w12753_ ;
	wire _w12752_ ;
	wire _w12751_ ;
	wire _w12750_ ;
	wire _w12749_ ;
	wire _w12748_ ;
	wire _w12747_ ;
	wire _w12746_ ;
	wire _w12745_ ;
	wire _w12744_ ;
	wire _w12743_ ;
	wire _w12742_ ;
	wire _w12741_ ;
	wire _w12740_ ;
	wire _w12739_ ;
	wire _w12738_ ;
	wire _w12737_ ;
	wire _w12736_ ;
	wire _w12735_ ;
	wire _w12734_ ;
	wire _w12733_ ;
	wire _w12732_ ;
	wire _w12731_ ;
	wire _w12730_ ;
	wire _w12729_ ;
	wire _w12728_ ;
	wire _w12727_ ;
	wire _w12726_ ;
	wire _w12725_ ;
	wire _w12724_ ;
	wire _w12723_ ;
	wire _w12722_ ;
	wire _w12721_ ;
	wire _w12720_ ;
	wire _w12719_ ;
	wire _w12718_ ;
	wire _w12717_ ;
	wire _w12716_ ;
	wire _w12715_ ;
	wire _w12714_ ;
	wire _w12713_ ;
	wire _w12712_ ;
	wire _w12711_ ;
	wire _w12710_ ;
	wire _w12709_ ;
	wire _w12708_ ;
	wire _w12707_ ;
	wire _w12706_ ;
	wire _w12705_ ;
	wire _w12704_ ;
	wire _w12703_ ;
	wire _w12702_ ;
	wire _w12701_ ;
	wire _w12700_ ;
	wire _w12699_ ;
	wire _w12698_ ;
	wire _w12697_ ;
	wire _w12696_ ;
	wire _w12695_ ;
	wire _w12694_ ;
	wire _w12693_ ;
	wire _w12692_ ;
	wire _w12691_ ;
	wire _w12690_ ;
	wire _w12689_ ;
	wire _w12688_ ;
	wire _w12687_ ;
	wire _w12686_ ;
	wire _w12685_ ;
	wire _w12684_ ;
	wire _w12683_ ;
	wire _w12682_ ;
	wire _w12681_ ;
	wire _w12680_ ;
	wire _w12679_ ;
	wire _w12678_ ;
	wire _w12677_ ;
	wire _w12676_ ;
	wire _w12675_ ;
	wire _w12674_ ;
	wire _w12673_ ;
	wire _w12672_ ;
	wire _w12671_ ;
	wire _w12670_ ;
	wire _w12669_ ;
	wire _w12668_ ;
	wire _w12667_ ;
	wire _w12666_ ;
	wire _w12665_ ;
	wire _w12664_ ;
	wire _w12663_ ;
	wire _w12662_ ;
	wire _w12661_ ;
	wire _w12660_ ;
	wire _w12659_ ;
	wire _w12658_ ;
	wire _w12657_ ;
	wire _w12656_ ;
	wire _w12655_ ;
	wire _w12654_ ;
	wire _w12653_ ;
	wire _w12652_ ;
	wire _w12651_ ;
	wire _w12650_ ;
	wire _w12649_ ;
	wire _w12648_ ;
	wire _w12647_ ;
	wire _w12646_ ;
	wire _w12645_ ;
	wire _w12644_ ;
	wire _w12643_ ;
	wire _w12642_ ;
	wire _w12641_ ;
	wire _w12640_ ;
	wire _w12639_ ;
	wire _w12638_ ;
	wire _w12637_ ;
	wire _w12636_ ;
	wire _w12635_ ;
	wire _w12634_ ;
	wire _w12633_ ;
	wire _w12632_ ;
	wire _w12631_ ;
	wire _w12630_ ;
	wire _w12629_ ;
	wire _w12628_ ;
	wire _w12627_ ;
	wire _w12626_ ;
	wire _w12625_ ;
	wire _w12624_ ;
	wire _w12623_ ;
	wire _w12622_ ;
	wire _w12621_ ;
	wire _w12620_ ;
	wire _w12619_ ;
	wire _w12618_ ;
	wire _w12617_ ;
	wire _w12616_ ;
	wire _w12615_ ;
	wire _w12614_ ;
	wire _w12613_ ;
	wire _w12612_ ;
	wire _w12611_ ;
	wire _w12610_ ;
	wire _w12609_ ;
	wire _w12608_ ;
	wire _w12607_ ;
	wire _w12606_ ;
	wire _w12605_ ;
	wire _w12604_ ;
	wire _w12603_ ;
	wire _w12602_ ;
	wire _w12601_ ;
	wire _w12600_ ;
	wire _w12599_ ;
	wire _w12598_ ;
	wire _w12597_ ;
	wire _w12596_ ;
	wire _w12595_ ;
	wire _w12594_ ;
	wire _w12593_ ;
	wire _w12592_ ;
	wire _w12591_ ;
	wire _w12590_ ;
	wire _w12589_ ;
	wire _w12588_ ;
	wire _w12587_ ;
	wire _w12586_ ;
	wire _w12585_ ;
	wire _w12584_ ;
	wire _w12583_ ;
	wire _w12582_ ;
	wire _w12581_ ;
	wire _w12580_ ;
	wire _w12579_ ;
	wire _w12578_ ;
	wire _w12577_ ;
	wire _w12576_ ;
	wire _w12575_ ;
	wire _w12574_ ;
	wire _w12573_ ;
	wire _w12572_ ;
	wire _w12571_ ;
	wire _w12570_ ;
	wire _w12569_ ;
	wire _w12568_ ;
	wire _w12567_ ;
	wire _w12566_ ;
	wire _w12565_ ;
	wire _w12564_ ;
	wire _w12563_ ;
	wire _w12562_ ;
	wire _w12561_ ;
	wire _w12560_ ;
	wire _w12559_ ;
	wire _w12558_ ;
	wire _w12557_ ;
	wire _w12556_ ;
	wire _w12555_ ;
	wire _w12554_ ;
	wire _w12553_ ;
	wire _w12552_ ;
	wire _w12551_ ;
	wire _w12550_ ;
	wire _w12549_ ;
	wire _w12548_ ;
	wire _w12547_ ;
	wire _w12546_ ;
	wire _w12545_ ;
	wire _w12544_ ;
	wire _w12543_ ;
	wire _w12542_ ;
	wire _w12541_ ;
	wire _w12540_ ;
	wire _w12539_ ;
	wire _w12538_ ;
	wire _w12537_ ;
	wire _w12536_ ;
	wire _w12535_ ;
	wire _w12534_ ;
	wire _w12533_ ;
	wire _w12532_ ;
	wire _w12531_ ;
	wire _w12530_ ;
	wire _w12529_ ;
	wire _w12528_ ;
	wire _w12527_ ;
	wire _w12526_ ;
	wire _w12525_ ;
	wire _w12524_ ;
	wire _w12523_ ;
	wire _w12522_ ;
	wire _w12521_ ;
	wire _w12520_ ;
	wire _w12519_ ;
	wire _w12518_ ;
	wire _w12517_ ;
	wire _w12516_ ;
	wire _w12515_ ;
	wire _w12514_ ;
	wire _w12513_ ;
	wire _w12512_ ;
	wire _w12511_ ;
	wire _w12510_ ;
	wire _w12509_ ;
	wire _w12508_ ;
	wire _w12507_ ;
	wire _w12506_ ;
	wire _w12505_ ;
	wire _w12504_ ;
	wire _w12503_ ;
	wire _w12502_ ;
	wire _w12501_ ;
	wire _w12500_ ;
	wire _w12499_ ;
	wire _w12498_ ;
	wire _w12497_ ;
	wire _w12496_ ;
	wire _w12495_ ;
	wire _w12494_ ;
	wire _w12493_ ;
	wire _w12492_ ;
	wire _w12491_ ;
	wire _w12490_ ;
	wire _w12489_ ;
	wire _w12488_ ;
	wire _w12487_ ;
	wire _w12486_ ;
	wire _w12485_ ;
	wire _w12484_ ;
	wire _w12483_ ;
	wire _w12482_ ;
	wire _w12481_ ;
	wire _w12480_ ;
	wire _w12479_ ;
	wire _w12478_ ;
	wire _w12477_ ;
	wire _w12476_ ;
	wire _w12475_ ;
	wire _w12474_ ;
	wire _w12473_ ;
	wire _w12472_ ;
	wire _w12471_ ;
	wire _w12470_ ;
	wire _w12469_ ;
	wire _w12468_ ;
	wire _w12467_ ;
	wire _w12466_ ;
	wire _w12465_ ;
	wire _w12464_ ;
	wire _w12463_ ;
	wire _w12462_ ;
	wire _w12461_ ;
	wire _w12460_ ;
	wire _w12459_ ;
	wire _w12458_ ;
	wire _w12457_ ;
	wire _w12456_ ;
	wire _w12455_ ;
	wire _w12454_ ;
	wire _w12453_ ;
	wire _w12452_ ;
	wire _w12451_ ;
	wire _w12450_ ;
	wire _w12449_ ;
	wire _w12448_ ;
	wire _w12447_ ;
	wire _w12446_ ;
	wire _w12445_ ;
	wire _w12444_ ;
	wire _w12443_ ;
	wire _w12442_ ;
	wire _w12441_ ;
	wire _w12440_ ;
	wire _w12439_ ;
	wire _w12438_ ;
	wire _w12437_ ;
	wire _w12436_ ;
	wire _w12435_ ;
	wire _w12434_ ;
	wire _w12433_ ;
	wire _w12432_ ;
	wire _w12431_ ;
	wire _w12430_ ;
	wire _w12429_ ;
	wire _w12428_ ;
	wire _w12427_ ;
	wire _w12426_ ;
	wire _w12425_ ;
	wire _w12424_ ;
	wire _w12423_ ;
	wire _w12422_ ;
	wire _w12421_ ;
	wire _w12420_ ;
	wire _w12419_ ;
	wire _w12418_ ;
	wire _w12417_ ;
	wire _w12416_ ;
	wire _w12415_ ;
	wire _w12414_ ;
	wire _w12413_ ;
	wire _w12412_ ;
	wire _w12411_ ;
	wire _w12410_ ;
	wire _w12409_ ;
	wire _w12408_ ;
	wire _w12407_ ;
	wire _w12406_ ;
	wire _w12405_ ;
	wire _w12404_ ;
	wire _w12403_ ;
	wire _w12402_ ;
	wire _w12401_ ;
	wire _w12400_ ;
	wire _w12399_ ;
	wire _w12398_ ;
	wire _w12397_ ;
	wire _w12396_ ;
	wire _w12395_ ;
	wire _w12394_ ;
	wire _w12393_ ;
	wire _w12392_ ;
	wire _w12391_ ;
	wire _w12390_ ;
	wire _w12389_ ;
	wire _w12388_ ;
	wire _w12387_ ;
	wire _w12386_ ;
	wire _w12385_ ;
	wire _w12384_ ;
	wire _w12383_ ;
	wire _w12382_ ;
	wire _w12381_ ;
	wire _w12380_ ;
	wire _w12379_ ;
	wire _w12378_ ;
	wire _w12377_ ;
	wire _w12376_ ;
	wire _w12375_ ;
	wire _w12374_ ;
	wire _w12373_ ;
	wire _w12372_ ;
	wire _w12371_ ;
	wire _w12370_ ;
	wire _w12369_ ;
	wire _w12368_ ;
	wire _w12367_ ;
	wire _w12366_ ;
	wire _w12365_ ;
	wire _w12364_ ;
	wire _w12363_ ;
	wire _w12362_ ;
	wire _w12361_ ;
	wire _w12360_ ;
	wire _w12359_ ;
	wire _w12358_ ;
	wire _w12357_ ;
	wire _w12356_ ;
	wire _w12355_ ;
	wire _w12354_ ;
	wire _w12353_ ;
	wire _w12352_ ;
	wire _w12351_ ;
	wire _w12350_ ;
	wire _w12349_ ;
	wire _w12348_ ;
	wire _w12347_ ;
	wire _w12346_ ;
	wire _w12345_ ;
	wire _w12344_ ;
	wire _w12343_ ;
	wire _w12342_ ;
	wire _w12341_ ;
	wire _w12340_ ;
	wire _w12339_ ;
	wire _w12338_ ;
	wire _w12337_ ;
	wire _w12336_ ;
	wire _w12335_ ;
	wire _w12334_ ;
	wire _w12333_ ;
	wire _w12332_ ;
	wire _w12331_ ;
	wire _w12330_ ;
	wire _w12329_ ;
	wire _w12328_ ;
	wire _w12327_ ;
	wire _w12326_ ;
	wire _w12325_ ;
	wire _w12324_ ;
	wire _w12323_ ;
	wire _w12322_ ;
	wire _w12321_ ;
	wire _w12320_ ;
	wire _w12319_ ;
	wire _w12318_ ;
	wire _w12317_ ;
	wire _w12316_ ;
	wire _w12315_ ;
	wire _w12314_ ;
	wire _w12313_ ;
	wire _w12312_ ;
	wire _w12311_ ;
	wire _w12310_ ;
	wire _w12309_ ;
	wire _w12308_ ;
	wire _w12307_ ;
	wire _w12306_ ;
	wire _w12305_ ;
	wire _w12304_ ;
	wire _w12303_ ;
	wire _w12302_ ;
	wire _w12301_ ;
	wire _w12300_ ;
	wire _w12299_ ;
	wire _w12298_ ;
	wire _w12297_ ;
	wire _w12296_ ;
	wire _w12295_ ;
	wire _w12294_ ;
	wire _w12293_ ;
	wire _w12292_ ;
	wire _w12291_ ;
	wire _w12290_ ;
	wire _w12289_ ;
	wire _w12288_ ;
	wire _w12287_ ;
	wire _w12286_ ;
	wire _w12285_ ;
	wire _w12284_ ;
	wire _w12283_ ;
	wire _w12282_ ;
	wire _w12281_ ;
	wire _w12280_ ;
	wire _w12279_ ;
	wire _w12278_ ;
	wire _w12277_ ;
	wire _w12276_ ;
	wire _w12275_ ;
	wire _w12274_ ;
	wire _w12273_ ;
	wire _w12272_ ;
	wire _w12271_ ;
	wire _w12270_ ;
	wire _w12269_ ;
	wire _w12268_ ;
	wire _w12267_ ;
	wire _w12266_ ;
	wire _w12265_ ;
	wire _w12264_ ;
	wire _w12263_ ;
	wire _w12262_ ;
	wire _w12261_ ;
	wire _w12260_ ;
	wire _w12259_ ;
	wire _w12258_ ;
	wire _w12257_ ;
	wire _w12256_ ;
	wire _w12255_ ;
	wire _w12254_ ;
	wire _w12253_ ;
	wire _w12252_ ;
	wire _w12251_ ;
	wire _w12250_ ;
	wire _w12249_ ;
	wire _w12248_ ;
	wire _w12247_ ;
	wire _w12246_ ;
	wire _w12245_ ;
	wire _w12244_ ;
	wire _w12243_ ;
	wire _w12242_ ;
	wire _w12241_ ;
	wire _w12240_ ;
	wire _w12239_ ;
	wire _w12238_ ;
	wire _w12237_ ;
	wire _w12236_ ;
	wire _w12235_ ;
	wire _w12234_ ;
	wire _w12233_ ;
	wire _w12232_ ;
	wire _w12231_ ;
	wire _w12230_ ;
	wire _w12229_ ;
	wire _w12228_ ;
	wire _w12227_ ;
	wire _w12226_ ;
	wire _w12225_ ;
	wire _w12224_ ;
	wire _w12223_ ;
	wire _w12222_ ;
	wire _w12221_ ;
	wire _w12220_ ;
	wire _w12219_ ;
	wire _w12218_ ;
	wire _w12217_ ;
	wire _w12216_ ;
	wire _w12215_ ;
	wire _w12214_ ;
	wire _w12213_ ;
	wire _w12212_ ;
	wire _w12211_ ;
	wire _w12210_ ;
	wire _w12209_ ;
	wire _w12208_ ;
	wire _w12207_ ;
	wire _w12206_ ;
	wire _w12205_ ;
	wire _w12204_ ;
	wire _w12203_ ;
	wire _w12202_ ;
	wire _w12201_ ;
	wire _w12200_ ;
	wire _w12199_ ;
	wire _w12198_ ;
	wire _w12197_ ;
	wire _w12196_ ;
	wire _w12195_ ;
	wire _w12194_ ;
	wire _w12193_ ;
	wire _w12192_ ;
	wire _w12191_ ;
	wire _w12190_ ;
	wire _w12189_ ;
	wire _w12188_ ;
	wire _w12187_ ;
	wire _w12186_ ;
	wire _w12185_ ;
	wire _w12184_ ;
	wire _w12183_ ;
	wire _w12182_ ;
	wire _w12181_ ;
	wire _w12180_ ;
	wire _w12179_ ;
	wire _w12178_ ;
	wire _w12177_ ;
	wire _w12176_ ;
	wire _w12175_ ;
	wire _w12174_ ;
	wire _w12173_ ;
	wire _w12172_ ;
	wire _w12171_ ;
	wire _w12170_ ;
	wire _w12169_ ;
	wire _w12168_ ;
	wire _w12167_ ;
	wire _w12166_ ;
	wire _w12165_ ;
	wire _w12164_ ;
	wire _w12163_ ;
	wire _w12162_ ;
	wire _w12161_ ;
	wire _w12160_ ;
	wire _w12159_ ;
	wire _w12158_ ;
	wire _w12157_ ;
	wire _w12156_ ;
	wire _w12155_ ;
	wire _w12154_ ;
	wire _w12153_ ;
	wire _w12152_ ;
	wire _w12151_ ;
	wire _w12150_ ;
	wire _w12149_ ;
	wire _w12148_ ;
	wire _w12147_ ;
	wire _w12146_ ;
	wire _w12145_ ;
	wire _w12144_ ;
	wire _w12143_ ;
	wire _w12142_ ;
	wire _w12141_ ;
	wire _w12140_ ;
	wire _w12139_ ;
	wire _w12138_ ;
	wire _w12137_ ;
	wire _w12136_ ;
	wire _w12135_ ;
	wire _w12134_ ;
	wire _w12133_ ;
	wire _w12132_ ;
	wire _w12131_ ;
	wire _w12130_ ;
	wire _w12129_ ;
	wire _w12128_ ;
	wire _w12127_ ;
	wire _w12126_ ;
	wire _w12125_ ;
	wire _w12124_ ;
	wire _w12123_ ;
	wire _w12122_ ;
	wire _w12121_ ;
	wire _w12120_ ;
	wire _w12119_ ;
	wire _w12118_ ;
	wire _w12117_ ;
	wire _w12116_ ;
	wire _w12115_ ;
	wire _w12114_ ;
	wire _w12113_ ;
	wire _w12112_ ;
	wire _w12111_ ;
	wire _w12110_ ;
	wire _w12109_ ;
	wire _w12108_ ;
	wire _w12107_ ;
	wire _w12106_ ;
	wire _w12105_ ;
	wire _w12104_ ;
	wire _w12103_ ;
	wire _w12102_ ;
	wire _w12101_ ;
	wire _w12100_ ;
	wire _w12099_ ;
	wire _w12098_ ;
	wire _w12097_ ;
	wire _w12096_ ;
	wire _w12095_ ;
	wire _w12094_ ;
	wire _w12093_ ;
	wire _w12092_ ;
	wire _w12091_ ;
	wire _w12090_ ;
	wire _w12089_ ;
	wire _w12088_ ;
	wire _w12087_ ;
	wire _w12086_ ;
	wire _w12085_ ;
	wire _w12084_ ;
	wire _w12083_ ;
	wire _w12082_ ;
	wire _w12081_ ;
	wire _w12080_ ;
	wire _w12079_ ;
	wire _w12078_ ;
	wire _w12077_ ;
	wire _w12076_ ;
	wire _w12075_ ;
	wire _w12074_ ;
	wire _w12073_ ;
	wire _w12072_ ;
	wire _w12071_ ;
	wire _w12070_ ;
	wire _w12069_ ;
	wire _w12068_ ;
	wire _w12067_ ;
	wire _w12066_ ;
	wire _w12065_ ;
	wire _w12064_ ;
	wire _w12063_ ;
	wire _w12062_ ;
	wire _w12061_ ;
	wire _w12060_ ;
	wire _w12059_ ;
	wire _w12058_ ;
	wire _w12057_ ;
	wire _w12056_ ;
	wire _w12055_ ;
	wire _w12054_ ;
	wire _w12053_ ;
	wire _w12052_ ;
	wire _w12051_ ;
	wire _w12050_ ;
	wire _w12049_ ;
	wire _w12048_ ;
	wire _w12047_ ;
	wire _w12046_ ;
	wire _w12045_ ;
	wire _w12044_ ;
	wire _w12043_ ;
	wire _w12042_ ;
	wire _w12041_ ;
	wire _w12040_ ;
	wire _w12039_ ;
	wire _w12038_ ;
	wire _w12037_ ;
	wire _w12036_ ;
	wire _w12035_ ;
	wire _w12034_ ;
	wire _w12033_ ;
	wire _w12032_ ;
	wire _w12031_ ;
	wire _w12030_ ;
	wire _w12029_ ;
	wire _w12028_ ;
	wire _w12027_ ;
	wire _w12026_ ;
	wire _w12025_ ;
	wire _w12024_ ;
	wire _w12023_ ;
	wire _w12022_ ;
	wire _w12021_ ;
	wire _w12020_ ;
	wire _w12019_ ;
	wire _w12018_ ;
	wire _w12017_ ;
	wire _w12016_ ;
	wire _w12015_ ;
	wire _w12014_ ;
	wire _w12013_ ;
	wire _w12012_ ;
	wire _w12011_ ;
	wire _w12010_ ;
	wire _w12009_ ;
	wire _w12008_ ;
	wire _w12007_ ;
	wire _w12006_ ;
	wire _w12005_ ;
	wire _w12004_ ;
	wire _w12003_ ;
	wire _w12002_ ;
	wire _w12001_ ;
	wire _w12000_ ;
	wire _w11999_ ;
	wire _w11998_ ;
	wire _w11997_ ;
	wire _w11996_ ;
	wire _w11995_ ;
	wire _w11994_ ;
	wire _w11993_ ;
	wire _w11992_ ;
	wire _w11991_ ;
	wire _w11990_ ;
	wire _w11989_ ;
	wire _w11988_ ;
	wire _w11987_ ;
	wire _w11986_ ;
	wire _w11985_ ;
	wire _w11984_ ;
	wire _w11983_ ;
	wire _w11982_ ;
	wire _w11981_ ;
	wire _w11980_ ;
	wire _w11979_ ;
	wire _w11978_ ;
	wire _w11977_ ;
	wire _w11976_ ;
	wire _w11975_ ;
	wire _w11974_ ;
	wire _w11973_ ;
	wire _w11972_ ;
	wire _w11971_ ;
	wire _w11970_ ;
	wire _w11969_ ;
	wire _w11968_ ;
	wire _w11967_ ;
	wire _w11966_ ;
	wire _w11965_ ;
	wire _w11964_ ;
	wire _w11963_ ;
	wire _w11962_ ;
	wire _w11961_ ;
	wire _w11960_ ;
	wire _w11959_ ;
	wire _w11958_ ;
	wire _w11957_ ;
	wire _w11956_ ;
	wire _w11955_ ;
	wire _w11954_ ;
	wire _w11953_ ;
	wire _w11952_ ;
	wire _w11951_ ;
	wire _w11950_ ;
	wire _w11949_ ;
	wire _w11948_ ;
	wire _w11947_ ;
	wire _w11946_ ;
	wire _w11945_ ;
	wire _w11944_ ;
	wire _w11943_ ;
	wire _w11942_ ;
	wire _w11941_ ;
	wire _w11940_ ;
	wire _w11939_ ;
	wire _w11938_ ;
	wire _w11937_ ;
	wire _w11936_ ;
	wire _w11935_ ;
	wire _w11934_ ;
	wire _w11933_ ;
	wire _w11932_ ;
	wire _w11931_ ;
	wire _w11930_ ;
	wire _w11929_ ;
	wire _w11928_ ;
	wire _w11927_ ;
	wire _w11926_ ;
	wire _w11925_ ;
	wire _w11924_ ;
	wire _w11923_ ;
	wire _w11922_ ;
	wire _w11921_ ;
	wire _w11920_ ;
	wire _w11919_ ;
	wire _w11918_ ;
	wire _w11917_ ;
	wire _w11916_ ;
	wire _w11915_ ;
	wire _w11914_ ;
	wire _w11913_ ;
	wire _w11912_ ;
	wire _w11911_ ;
	wire _w11910_ ;
	wire _w11909_ ;
	wire _w11908_ ;
	wire _w11907_ ;
	wire _w11906_ ;
	wire _w11905_ ;
	wire _w11904_ ;
	wire _w11903_ ;
	wire _w11902_ ;
	wire _w11901_ ;
	wire _w11900_ ;
	wire _w11899_ ;
	wire _w11898_ ;
	wire _w11897_ ;
	wire _w11896_ ;
	wire _w11895_ ;
	wire _w11894_ ;
	wire _w11893_ ;
	wire _w11892_ ;
	wire _w11891_ ;
	wire _w11890_ ;
	wire _w11889_ ;
	wire _w11888_ ;
	wire _w11887_ ;
	wire _w11886_ ;
	wire _w11885_ ;
	wire _w11884_ ;
	wire _w11883_ ;
	wire _w11882_ ;
	wire _w11881_ ;
	wire _w11880_ ;
	wire _w11879_ ;
	wire _w11878_ ;
	wire _w11877_ ;
	wire _w11876_ ;
	wire _w11875_ ;
	wire _w11874_ ;
	wire _w11873_ ;
	wire _w11872_ ;
	wire _w11871_ ;
	wire _w11870_ ;
	wire _w11869_ ;
	wire _w11868_ ;
	wire _w11867_ ;
	wire _w11866_ ;
	wire _w11865_ ;
	wire _w11864_ ;
	wire _w11863_ ;
	wire _w11862_ ;
	wire _w11861_ ;
	wire _w11860_ ;
	wire _w11859_ ;
	wire _w11858_ ;
	wire _w11857_ ;
	wire _w11856_ ;
	wire _w11855_ ;
	wire _w11854_ ;
	wire _w11853_ ;
	wire _w11852_ ;
	wire _w11851_ ;
	wire _w11850_ ;
	wire _w11849_ ;
	wire _w11848_ ;
	wire _w11847_ ;
	wire _w11846_ ;
	wire _w11845_ ;
	wire _w11844_ ;
	wire _w11843_ ;
	wire _w11842_ ;
	wire _w11841_ ;
	wire _w11840_ ;
	wire _w11839_ ;
	wire _w11838_ ;
	wire _w11837_ ;
	wire _w11836_ ;
	wire _w11835_ ;
	wire _w11834_ ;
	wire _w11833_ ;
	wire _w11832_ ;
	wire _w11831_ ;
	wire _w11830_ ;
	wire _w11829_ ;
	wire _w11828_ ;
	wire _w11827_ ;
	wire _w11826_ ;
	wire _w11825_ ;
	wire _w11824_ ;
	wire _w11823_ ;
	wire _w11822_ ;
	wire _w11821_ ;
	wire _w11820_ ;
	wire _w11819_ ;
	wire _w11818_ ;
	wire _w11817_ ;
	wire _w11816_ ;
	wire _w11815_ ;
	wire _w11814_ ;
	wire _w11813_ ;
	wire _w11812_ ;
	wire _w11811_ ;
	wire _w11810_ ;
	wire _w11809_ ;
	wire _w11808_ ;
	wire _w11807_ ;
	wire _w11806_ ;
	wire _w11805_ ;
	wire _w11804_ ;
	wire _w11803_ ;
	wire _w11802_ ;
	wire _w11801_ ;
	wire _w11800_ ;
	wire _w11799_ ;
	wire _w11798_ ;
	wire _w11797_ ;
	wire _w11796_ ;
	wire _w11795_ ;
	wire _w11794_ ;
	wire _w11793_ ;
	wire _w11792_ ;
	wire _w11791_ ;
	wire _w11790_ ;
	wire _w11789_ ;
	wire _w11788_ ;
	wire _w11787_ ;
	wire _w11786_ ;
	wire _w11785_ ;
	wire _w11784_ ;
	wire _w11783_ ;
	wire _w11782_ ;
	wire _w11781_ ;
	wire _w11780_ ;
	wire _w11779_ ;
	wire _w11778_ ;
	wire _w11777_ ;
	wire _w11776_ ;
	wire _w11775_ ;
	wire _w11774_ ;
	wire _w11773_ ;
	wire _w11772_ ;
	wire _w11771_ ;
	wire _w11770_ ;
	wire _w11769_ ;
	wire _w11768_ ;
	wire _w11767_ ;
	wire _w11766_ ;
	wire _w11765_ ;
	wire _w11764_ ;
	wire _w11763_ ;
	wire _w11762_ ;
	wire _w11761_ ;
	wire _w11760_ ;
	wire _w11759_ ;
	wire _w11758_ ;
	wire _w11757_ ;
	wire _w11756_ ;
	wire _w11755_ ;
	wire _w11754_ ;
	wire _w11753_ ;
	wire _w11752_ ;
	wire _w11751_ ;
	wire _w11750_ ;
	wire _w11749_ ;
	wire _w11748_ ;
	wire _w11747_ ;
	wire _w11746_ ;
	wire _w11745_ ;
	wire _w11744_ ;
	wire _w11743_ ;
	wire _w11742_ ;
	wire _w11741_ ;
	wire _w11740_ ;
	wire _w11739_ ;
	wire _w11738_ ;
	wire _w11737_ ;
	wire _w11736_ ;
	wire _w11735_ ;
	wire _w11734_ ;
	wire _w11733_ ;
	wire _w11732_ ;
	wire _w11731_ ;
	wire _w11730_ ;
	wire _w11729_ ;
	wire _w11728_ ;
	wire _w11727_ ;
	wire _w11726_ ;
	wire _w11725_ ;
	wire _w11724_ ;
	wire _w11723_ ;
	wire _w11722_ ;
	wire _w11721_ ;
	wire _w11720_ ;
	wire _w11719_ ;
	wire _w11718_ ;
	wire _w11717_ ;
	wire _w11716_ ;
	wire _w11715_ ;
	wire _w11714_ ;
	wire _w11713_ ;
	wire _w11712_ ;
	wire _w11711_ ;
	wire _w11710_ ;
	wire _w11709_ ;
	wire _w11708_ ;
	wire _w11707_ ;
	wire _w11706_ ;
	wire _w11705_ ;
	wire _w11704_ ;
	wire _w11703_ ;
	wire _w11702_ ;
	wire _w11701_ ;
	wire _w11700_ ;
	wire _w11699_ ;
	wire _w11698_ ;
	wire _w11697_ ;
	wire _w11696_ ;
	wire _w11695_ ;
	wire _w11694_ ;
	wire _w11693_ ;
	wire _w11692_ ;
	wire _w11691_ ;
	wire _w11690_ ;
	wire _w11689_ ;
	wire _w11688_ ;
	wire _w11687_ ;
	wire _w11686_ ;
	wire _w11685_ ;
	wire _w11684_ ;
	wire _w11683_ ;
	wire _w11682_ ;
	wire _w11681_ ;
	wire _w11680_ ;
	wire _w11679_ ;
	wire _w11678_ ;
	wire _w11677_ ;
	wire _w11676_ ;
	wire _w11675_ ;
	wire _w11674_ ;
	wire _w11673_ ;
	wire _w11672_ ;
	wire _w11671_ ;
	wire _w11670_ ;
	wire _w11669_ ;
	wire _w11668_ ;
	wire _w11667_ ;
	wire _w11666_ ;
	wire _w11665_ ;
	wire _w11664_ ;
	wire _w11663_ ;
	wire _w11662_ ;
	wire _w11661_ ;
	wire _w11660_ ;
	wire _w11659_ ;
	wire _w11658_ ;
	wire _w11657_ ;
	wire _w11656_ ;
	wire _w11655_ ;
	wire _w11654_ ;
	wire _w11653_ ;
	wire _w11652_ ;
	wire _w11651_ ;
	wire _w11650_ ;
	wire _w11649_ ;
	wire _w11648_ ;
	wire _w11647_ ;
	wire _w11646_ ;
	wire _w11645_ ;
	wire _w11644_ ;
	wire _w11643_ ;
	wire _w11642_ ;
	wire _w11641_ ;
	wire _w11640_ ;
	wire _w11639_ ;
	wire _w11638_ ;
	wire _w11637_ ;
	wire _w11636_ ;
	wire _w11635_ ;
	wire _w11634_ ;
	wire _w11633_ ;
	wire _w11632_ ;
	wire _w11631_ ;
	wire _w11630_ ;
	wire _w11629_ ;
	wire _w11628_ ;
	wire _w11627_ ;
	wire _w11626_ ;
	wire _w11625_ ;
	wire _w11624_ ;
	wire _w11623_ ;
	wire _w11622_ ;
	wire _w11621_ ;
	wire _w11620_ ;
	wire _w11619_ ;
	wire _w11618_ ;
	wire _w11617_ ;
	wire _w11616_ ;
	wire _w11615_ ;
	wire _w11614_ ;
	wire _w11613_ ;
	wire _w11612_ ;
	wire _w11611_ ;
	wire _w11610_ ;
	wire _w11609_ ;
	wire _w11608_ ;
	wire _w11607_ ;
	wire _w11606_ ;
	wire _w11605_ ;
	wire _w11604_ ;
	wire _w11603_ ;
	wire _w11602_ ;
	wire _w11601_ ;
	wire _w11600_ ;
	wire _w11599_ ;
	wire _w11598_ ;
	wire _w11597_ ;
	wire _w11596_ ;
	wire _w11595_ ;
	wire _w11594_ ;
	wire _w11593_ ;
	wire _w11592_ ;
	wire _w11591_ ;
	wire _w11590_ ;
	wire _w11589_ ;
	wire _w11588_ ;
	wire _w11587_ ;
	wire _w11586_ ;
	wire _w11585_ ;
	wire _w11584_ ;
	wire _w11583_ ;
	wire _w11582_ ;
	wire _w11581_ ;
	wire _w11580_ ;
	wire _w11579_ ;
	wire _w11578_ ;
	wire _w11577_ ;
	wire _w11576_ ;
	wire _w11575_ ;
	wire _w11574_ ;
	wire _w11573_ ;
	wire _w11572_ ;
	wire _w11571_ ;
	wire _w11570_ ;
	wire _w11569_ ;
	wire _w11568_ ;
	wire _w11567_ ;
	wire _w11566_ ;
	wire _w11565_ ;
	wire _w11564_ ;
	wire _w11563_ ;
	wire _w11562_ ;
	wire _w11561_ ;
	wire _w11560_ ;
	wire _w11559_ ;
	wire _w11558_ ;
	wire _w11557_ ;
	wire _w11556_ ;
	wire _w11555_ ;
	wire _w11554_ ;
	wire _w11553_ ;
	wire _w11552_ ;
	wire _w11551_ ;
	wire _w11550_ ;
	wire _w11549_ ;
	wire _w11548_ ;
	wire _w11547_ ;
	wire _w11546_ ;
	wire _w11545_ ;
	wire _w11544_ ;
	wire _w11543_ ;
	wire _w11542_ ;
	wire _w11541_ ;
	wire _w11540_ ;
	wire _w11539_ ;
	wire _w11538_ ;
	wire _w11537_ ;
	wire _w11536_ ;
	wire _w11535_ ;
	wire _w11534_ ;
	wire _w11533_ ;
	wire _w11532_ ;
	wire _w11531_ ;
	wire _w11530_ ;
	wire _w11529_ ;
	wire _w11528_ ;
	wire _w11527_ ;
	wire _w11526_ ;
	wire _w11525_ ;
	wire _w11524_ ;
	wire _w11523_ ;
	wire _w11522_ ;
	wire _w11521_ ;
	wire _w11520_ ;
	wire _w11519_ ;
	wire _w11518_ ;
	wire _w11517_ ;
	wire _w11516_ ;
	wire _w11515_ ;
	wire _w11514_ ;
	wire _w11513_ ;
	wire _w11512_ ;
	wire _w11511_ ;
	wire _w11510_ ;
	wire _w11509_ ;
	wire _w11508_ ;
	wire _w11507_ ;
	wire _w11506_ ;
	wire _w11505_ ;
	wire _w11504_ ;
	wire _w11503_ ;
	wire _w11502_ ;
	wire _w11501_ ;
	wire _w11500_ ;
	wire _w11499_ ;
	wire _w11498_ ;
	wire _w11497_ ;
	wire _w11496_ ;
	wire _w11495_ ;
	wire _w11494_ ;
	wire _w11493_ ;
	wire _w11492_ ;
	wire _w11491_ ;
	wire _w11490_ ;
	wire _w11489_ ;
	wire _w11488_ ;
	wire _w11487_ ;
	wire _w11486_ ;
	wire _w11485_ ;
	wire _w11484_ ;
	wire _w11483_ ;
	wire _w11482_ ;
	wire _w11481_ ;
	wire _w11480_ ;
	wire _w11479_ ;
	wire _w11478_ ;
	wire _w11477_ ;
	wire _w11476_ ;
	wire _w11475_ ;
	wire _w11474_ ;
	wire _w11473_ ;
	wire _w11472_ ;
	wire _w11471_ ;
	wire _w11470_ ;
	wire _w11469_ ;
	wire _w11468_ ;
	wire _w11467_ ;
	wire _w11466_ ;
	wire _w11465_ ;
	wire _w11464_ ;
	wire _w11463_ ;
	wire _w11462_ ;
	wire _w11461_ ;
	wire _w11460_ ;
	wire _w11459_ ;
	wire _w11458_ ;
	wire _w11457_ ;
	wire _w11456_ ;
	wire _w11455_ ;
	wire _w11454_ ;
	wire _w11453_ ;
	wire _w11452_ ;
	wire _w11451_ ;
	wire _w11450_ ;
	wire _w11449_ ;
	wire _w11448_ ;
	wire _w11447_ ;
	wire _w11446_ ;
	wire _w11445_ ;
	wire _w11444_ ;
	wire _w11443_ ;
	wire _w11442_ ;
	wire _w11441_ ;
	wire _w11440_ ;
	wire _w11439_ ;
	wire _w11438_ ;
	wire _w11437_ ;
	wire _w11436_ ;
	wire _w11435_ ;
	wire _w11434_ ;
	wire _w11433_ ;
	wire _w11432_ ;
	wire _w11431_ ;
	wire _w11430_ ;
	wire _w11429_ ;
	wire _w11428_ ;
	wire _w11427_ ;
	wire _w11426_ ;
	wire _w11425_ ;
	wire _w11424_ ;
	wire _w11423_ ;
	wire _w11422_ ;
	wire _w11421_ ;
	wire _w11420_ ;
	wire _w11419_ ;
	wire _w11418_ ;
	wire _w11417_ ;
	wire _w11416_ ;
	wire _w11415_ ;
	wire _w11414_ ;
	wire _w11413_ ;
	wire _w11412_ ;
	wire _w11411_ ;
	wire _w11410_ ;
	wire _w11409_ ;
	wire _w11408_ ;
	wire _w11407_ ;
	wire _w11406_ ;
	wire _w11405_ ;
	wire _w11404_ ;
	wire _w11403_ ;
	wire _w11402_ ;
	wire _w11401_ ;
	wire _w11400_ ;
	wire _w11399_ ;
	wire _w11398_ ;
	wire _w11397_ ;
	wire _w11396_ ;
	wire _w11395_ ;
	wire _w11394_ ;
	wire _w11393_ ;
	wire _w11392_ ;
	wire _w11391_ ;
	wire _w11390_ ;
	wire _w11389_ ;
	wire _w11388_ ;
	wire _w11387_ ;
	wire _w11386_ ;
	wire _w11385_ ;
	wire _w11384_ ;
	wire _w11383_ ;
	wire _w11382_ ;
	wire _w11381_ ;
	wire _w11380_ ;
	wire _w11379_ ;
	wire _w11378_ ;
	wire _w11377_ ;
	wire _w11376_ ;
	wire _w11375_ ;
	wire _w11374_ ;
	wire _w11373_ ;
	wire _w11372_ ;
	wire _w11371_ ;
	wire _w11370_ ;
	wire _w11369_ ;
	wire _w11368_ ;
	wire _w11367_ ;
	wire _w11366_ ;
	wire _w11365_ ;
	wire _w11364_ ;
	wire _w11363_ ;
	wire _w11362_ ;
	wire _w11361_ ;
	wire _w11360_ ;
	wire _w11359_ ;
	wire _w11358_ ;
	wire _w11357_ ;
	wire _w11356_ ;
	wire _w11355_ ;
	wire _w11354_ ;
	wire _w11353_ ;
	wire _w11352_ ;
	wire _w11351_ ;
	wire _w11350_ ;
	wire _w11349_ ;
	wire _w11348_ ;
	wire _w11347_ ;
	wire _w11346_ ;
	wire _w11345_ ;
	wire _w11344_ ;
	wire _w11343_ ;
	wire _w11342_ ;
	wire _w11341_ ;
	wire _w11340_ ;
	wire _w11339_ ;
	wire _w11338_ ;
	wire _w11337_ ;
	wire _w11336_ ;
	wire _w11335_ ;
	wire _w11334_ ;
	wire _w11333_ ;
	wire _w11332_ ;
	wire _w11331_ ;
	wire _w11330_ ;
	wire _w11329_ ;
	wire _w11328_ ;
	wire _w11327_ ;
	wire _w11326_ ;
	wire _w11325_ ;
	wire _w11324_ ;
	wire _w11323_ ;
	wire _w11322_ ;
	wire _w11321_ ;
	wire _w11320_ ;
	wire _w11319_ ;
	wire _w11318_ ;
	wire _w11317_ ;
	wire _w11316_ ;
	wire _w11315_ ;
	wire _w11314_ ;
	wire _w11313_ ;
	wire _w11312_ ;
	wire _w11311_ ;
	wire _w11310_ ;
	wire _w11309_ ;
	wire _w11308_ ;
	wire _w11307_ ;
	wire _w11306_ ;
	wire _w11305_ ;
	wire _w11304_ ;
	wire _w11303_ ;
	wire _w11302_ ;
	wire _w11301_ ;
	wire _w11300_ ;
	wire _w11299_ ;
	wire _w11298_ ;
	wire _w11297_ ;
	wire _w11296_ ;
	wire _w11295_ ;
	wire _w11294_ ;
	wire _w11293_ ;
	wire _w11292_ ;
	wire _w11291_ ;
	wire _w11290_ ;
	wire _w11289_ ;
	wire _w11288_ ;
	wire _w11287_ ;
	wire _w11286_ ;
	wire _w11285_ ;
	wire _w11284_ ;
	wire _w11283_ ;
	wire _w11282_ ;
	wire _w11281_ ;
	wire _w11280_ ;
	wire _w11279_ ;
	wire _w11278_ ;
	wire _w11277_ ;
	wire _w11276_ ;
	wire _w11275_ ;
	wire _w11274_ ;
	wire _w11273_ ;
	wire _w11272_ ;
	wire _w11271_ ;
	wire _w11270_ ;
	wire _w11269_ ;
	wire _w11268_ ;
	wire _w11267_ ;
	wire _w11266_ ;
	wire _w11265_ ;
	wire _w11264_ ;
	wire _w11263_ ;
	wire _w11262_ ;
	wire _w11261_ ;
	wire _w11260_ ;
	wire _w11259_ ;
	wire _w11258_ ;
	wire _w11257_ ;
	wire _w11256_ ;
	wire _w11255_ ;
	wire _w11254_ ;
	wire _w11253_ ;
	wire _w11252_ ;
	wire _w11251_ ;
	wire _w11250_ ;
	wire _w11249_ ;
	wire _w11248_ ;
	wire _w11247_ ;
	wire _w11246_ ;
	wire _w11245_ ;
	wire _w11244_ ;
	wire _w11243_ ;
	wire _w11242_ ;
	wire _w11241_ ;
	wire _w11240_ ;
	wire _w11239_ ;
	wire _w11238_ ;
	wire _w11237_ ;
	wire _w11236_ ;
	wire _w11235_ ;
	wire _w11234_ ;
	wire _w11233_ ;
	wire _w11232_ ;
	wire _w11231_ ;
	wire _w11230_ ;
	wire _w11229_ ;
	wire _w11228_ ;
	wire _w11227_ ;
	wire _w11226_ ;
	wire _w11225_ ;
	wire _w11224_ ;
	wire _w11223_ ;
	wire _w11222_ ;
	wire _w11221_ ;
	wire _w11220_ ;
	wire _w11219_ ;
	wire _w11218_ ;
	wire _w11217_ ;
	wire _w11216_ ;
	wire _w11215_ ;
	wire _w11214_ ;
	wire _w11213_ ;
	wire _w11212_ ;
	wire _w11211_ ;
	wire _w11210_ ;
	wire _w11209_ ;
	wire _w11208_ ;
	wire _w11207_ ;
	wire _w11206_ ;
	wire _w11205_ ;
	wire _w11204_ ;
	wire _w11203_ ;
	wire _w11202_ ;
	wire _w11201_ ;
	wire _w11200_ ;
	wire _w11199_ ;
	wire _w11198_ ;
	wire _w11197_ ;
	wire _w11196_ ;
	wire _w11195_ ;
	wire _w11194_ ;
	wire _w11193_ ;
	wire _w11192_ ;
	wire _w11191_ ;
	wire _w11190_ ;
	wire _w11189_ ;
	wire _w11188_ ;
	wire _w11187_ ;
	wire _w11186_ ;
	wire _w11185_ ;
	wire _w11184_ ;
	wire _w11183_ ;
	wire _w11182_ ;
	wire _w11181_ ;
	wire _w11180_ ;
	wire _w11179_ ;
	wire _w11178_ ;
	wire _w11177_ ;
	wire _w11176_ ;
	wire _w11175_ ;
	wire _w11174_ ;
	wire _w11173_ ;
	wire _w11172_ ;
	wire _w11171_ ;
	wire _w11170_ ;
	wire _w11169_ ;
	wire _w11168_ ;
	wire _w11167_ ;
	wire _w11166_ ;
	wire _w11165_ ;
	wire _w11164_ ;
	wire _w11163_ ;
	wire _w11162_ ;
	wire _w11161_ ;
	wire _w11160_ ;
	wire _w11159_ ;
	wire _w11158_ ;
	wire _w11157_ ;
	wire _w11156_ ;
	wire _w11155_ ;
	wire _w11154_ ;
	wire _w11153_ ;
	wire _w11152_ ;
	wire _w11151_ ;
	wire _w11150_ ;
	wire _w11149_ ;
	wire _w11148_ ;
	wire _w11147_ ;
	wire _w11146_ ;
	wire _w11145_ ;
	wire _w11144_ ;
	wire _w11143_ ;
	wire _w11142_ ;
	wire _w11141_ ;
	wire _w11140_ ;
	wire _w11139_ ;
	wire _w11138_ ;
	wire _w11137_ ;
	wire _w11136_ ;
	wire _w11135_ ;
	wire _w11134_ ;
	wire _w11133_ ;
	wire _w11132_ ;
	wire _w11131_ ;
	wire _w11130_ ;
	wire _w11129_ ;
	wire _w11128_ ;
	wire _w11127_ ;
	wire _w11126_ ;
	wire _w11125_ ;
	wire _w11124_ ;
	wire _w11123_ ;
	wire _w11122_ ;
	wire _w11121_ ;
	wire _w11120_ ;
	wire _w11119_ ;
	wire _w11118_ ;
	wire _w11117_ ;
	wire _w11116_ ;
	wire _w11115_ ;
	wire _w11114_ ;
	wire _w11113_ ;
	wire _w11112_ ;
	wire _w11111_ ;
	wire _w11110_ ;
	wire _w11109_ ;
	wire _w11108_ ;
	wire _w11107_ ;
	wire _w11106_ ;
	wire _w11105_ ;
	wire _w11104_ ;
	wire _w11103_ ;
	wire _w11102_ ;
	wire _w11101_ ;
	wire _w11100_ ;
	wire _w11099_ ;
	wire _w11098_ ;
	wire _w11097_ ;
	wire _w11096_ ;
	wire _w11095_ ;
	wire _w11094_ ;
	wire _w11093_ ;
	wire _w11092_ ;
	wire _w11091_ ;
	wire _w11090_ ;
	wire _w11089_ ;
	wire _w11088_ ;
	wire _w11087_ ;
	wire _w11086_ ;
	wire _w11085_ ;
	wire _w11084_ ;
	wire _w11083_ ;
	wire _w11082_ ;
	wire _w11081_ ;
	wire _w11080_ ;
	wire _w11079_ ;
	wire _w11078_ ;
	wire _w11077_ ;
	wire _w11076_ ;
	wire _w11075_ ;
	wire _w11074_ ;
	wire _w11073_ ;
	wire _w11072_ ;
	wire _w11071_ ;
	wire _w11070_ ;
	wire _w11069_ ;
	wire _w11068_ ;
	wire _w11067_ ;
	wire _w11066_ ;
	wire _w11065_ ;
	wire _w11064_ ;
	wire _w11063_ ;
	wire _w11062_ ;
	wire _w11061_ ;
	wire _w11060_ ;
	wire _w11059_ ;
	wire _w11058_ ;
	wire _w11057_ ;
	wire _w11056_ ;
	wire _w11055_ ;
	wire _w11054_ ;
	wire _w11053_ ;
	wire _w11052_ ;
	wire _w11051_ ;
	wire _w11050_ ;
	wire _w11049_ ;
	wire _w11048_ ;
	wire _w11047_ ;
	wire _w11046_ ;
	wire _w11045_ ;
	wire _w11044_ ;
	wire _w11043_ ;
	wire _w11042_ ;
	wire _w11041_ ;
	wire _w11040_ ;
	wire _w11039_ ;
	wire _w11038_ ;
	wire _w11037_ ;
	wire _w11036_ ;
	wire _w11035_ ;
	wire _w11034_ ;
	wire _w11033_ ;
	wire _w11032_ ;
	wire _w11031_ ;
	wire _w11030_ ;
	wire _w11029_ ;
	wire _w11028_ ;
	wire _w11027_ ;
	wire _w11026_ ;
	wire _w11025_ ;
	wire _w11024_ ;
	wire _w11023_ ;
	wire _w11022_ ;
	wire _w11021_ ;
	wire _w11020_ ;
	wire _w11019_ ;
	wire _w11018_ ;
	wire _w11017_ ;
	wire _w11016_ ;
	wire _w11015_ ;
	wire _w11014_ ;
	wire _w11013_ ;
	wire _w11012_ ;
	wire _w11011_ ;
	wire _w11010_ ;
	wire _w11009_ ;
	wire _w11008_ ;
	wire _w11007_ ;
	wire _w11006_ ;
	wire _w11005_ ;
	wire _w11004_ ;
	wire _w11003_ ;
	wire _w11002_ ;
	wire _w11001_ ;
	wire _w11000_ ;
	wire _w10999_ ;
	wire _w10998_ ;
	wire _w10997_ ;
	wire _w10996_ ;
	wire _w10995_ ;
	wire _w10994_ ;
	wire _w10993_ ;
	wire _w10992_ ;
	wire _w10991_ ;
	wire _w10990_ ;
	wire _w10989_ ;
	wire _w10988_ ;
	wire _w10987_ ;
	wire _w10986_ ;
	wire _w10985_ ;
	wire _w10984_ ;
	wire _w10983_ ;
	wire _w10982_ ;
	wire _w10981_ ;
	wire _w10980_ ;
	wire _w10979_ ;
	wire _w10978_ ;
	wire _w10977_ ;
	wire _w10976_ ;
	wire _w10975_ ;
	wire _w10974_ ;
	wire _w10973_ ;
	wire _w10972_ ;
	wire _w10971_ ;
	wire _w10970_ ;
	wire _w10969_ ;
	wire _w10968_ ;
	wire _w10967_ ;
	wire _w10966_ ;
	wire _w10965_ ;
	wire _w10964_ ;
	wire _w10963_ ;
	wire _w10962_ ;
	wire _w10961_ ;
	wire _w10960_ ;
	wire _w10959_ ;
	wire _w10958_ ;
	wire _w10957_ ;
	wire _w10956_ ;
	wire _w10955_ ;
	wire _w10954_ ;
	wire _w10953_ ;
	wire _w10952_ ;
	wire _w10951_ ;
	wire _w10950_ ;
	wire _w10949_ ;
	wire _w10948_ ;
	wire _w10947_ ;
	wire _w10946_ ;
	wire _w10945_ ;
	wire _w10944_ ;
	wire _w10943_ ;
	wire _w10942_ ;
	wire _w10941_ ;
	wire _w10940_ ;
	wire _w10939_ ;
	wire _w10938_ ;
	wire _w10937_ ;
	wire _w10936_ ;
	wire _w10935_ ;
	wire _w10934_ ;
	wire _w10933_ ;
	wire _w10932_ ;
	wire _w10931_ ;
	wire _w10930_ ;
	wire _w10929_ ;
	wire _w10928_ ;
	wire _w10927_ ;
	wire _w10926_ ;
	wire _w10925_ ;
	wire _w10924_ ;
	wire _w10923_ ;
	wire _w10922_ ;
	wire _w10921_ ;
	wire _w10920_ ;
	wire _w10919_ ;
	wire _w10918_ ;
	wire _w10917_ ;
	wire _w10916_ ;
	wire _w10915_ ;
	wire _w10914_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8038_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w8184_ ;
	wire _w8185_ ;
	wire _w8186_ ;
	wire _w8187_ ;
	wire _w8188_ ;
	wire _w8189_ ;
	wire _w8190_ ;
	wire _w8191_ ;
	wire _w8192_ ;
	wire _w8193_ ;
	wire _w8194_ ;
	wire _w8195_ ;
	wire _w8196_ ;
	wire _w8197_ ;
	wire _w8198_ ;
	wire _w8199_ ;
	wire _w8200_ ;
	wire _w8201_ ;
	wire _w8202_ ;
	wire _w8203_ ;
	wire _w8204_ ;
	wire _w8205_ ;
	wire _w8206_ ;
	wire _w8207_ ;
	wire _w8208_ ;
	wire _w8209_ ;
	wire _w8210_ ;
	wire _w8211_ ;
	wire _w8212_ ;
	wire _w8213_ ;
	wire _w8214_ ;
	wire _w8215_ ;
	wire _w8216_ ;
	wire _w8217_ ;
	wire _w8218_ ;
	wire _w8219_ ;
	wire _w8220_ ;
	wire _w8221_ ;
	wire _w8222_ ;
	wire _w8223_ ;
	wire _w8224_ ;
	wire _w8225_ ;
	wire _w8226_ ;
	wire _w8227_ ;
	wire _w8228_ ;
	wire _w8229_ ;
	wire _w8230_ ;
	wire _w8231_ ;
	wire _w8232_ ;
	wire _w8233_ ;
	wire _w8234_ ;
	wire _w8235_ ;
	wire _w8236_ ;
	wire _w8237_ ;
	wire _w8238_ ;
	wire _w8239_ ;
	wire _w8240_ ;
	wire _w8241_ ;
	wire _w8242_ ;
	wire _w8243_ ;
	wire _w8244_ ;
	wire _w8245_ ;
	wire _w8246_ ;
	wire _w8247_ ;
	wire _w8248_ ;
	wire _w8249_ ;
	wire _w8250_ ;
	wire _w8251_ ;
	wire _w8252_ ;
	wire _w8253_ ;
	wire _w8254_ ;
	wire _w8255_ ;
	wire _w8256_ ;
	wire _w8257_ ;
	wire _w8258_ ;
	wire _w8259_ ;
	wire _w8260_ ;
	wire _w8261_ ;
	wire _w8262_ ;
	wire _w8263_ ;
	wire _w8264_ ;
	wire _w8265_ ;
	wire _w8266_ ;
	wire _w8267_ ;
	wire _w8268_ ;
	wire _w8269_ ;
	wire _w8270_ ;
	wire _w8271_ ;
	wire _w8272_ ;
	wire _w8273_ ;
	wire _w8274_ ;
	wire _w8275_ ;
	wire _w8276_ ;
	wire _w8277_ ;
	wire _w8278_ ;
	wire _w8279_ ;
	wire _w8280_ ;
	wire _w8281_ ;
	wire _w8282_ ;
	wire _w8283_ ;
	wire _w8284_ ;
	wire _w8285_ ;
	wire _w8286_ ;
	wire _w8287_ ;
	wire _w8288_ ;
	wire _w8289_ ;
	wire _w8290_ ;
	wire _w8291_ ;
	wire _w8292_ ;
	wire _w8293_ ;
	wire _w8294_ ;
	wire _w8295_ ;
	wire _w8296_ ;
	wire _w8297_ ;
	wire _w8298_ ;
	wire _w8299_ ;
	wire _w8300_ ;
	wire _w8301_ ;
	wire _w8302_ ;
	wire _w8303_ ;
	wire _w8304_ ;
	wire _w8305_ ;
	wire _w8306_ ;
	wire _w8307_ ;
	wire _w8308_ ;
	wire _w8309_ ;
	wire _w8310_ ;
	wire _w8311_ ;
	wire _w8312_ ;
	wire _w8313_ ;
	wire _w8314_ ;
	wire _w8315_ ;
	wire _w8316_ ;
	wire _w8317_ ;
	wire _w8318_ ;
	wire _w8319_ ;
	wire _w8320_ ;
	wire _w8321_ ;
	wire _w8322_ ;
	wire _w8323_ ;
	wire _w8324_ ;
	wire _w8325_ ;
	wire _w8326_ ;
	wire _w8327_ ;
	wire _w8328_ ;
	wire _w8329_ ;
	wire _w8330_ ;
	wire _w8331_ ;
	wire _w8332_ ;
	wire _w8333_ ;
	wire _w8334_ ;
	wire _w8335_ ;
	wire _w8336_ ;
	wire _w8337_ ;
	wire _w8338_ ;
	wire _w8339_ ;
	wire _w8340_ ;
	wire _w8341_ ;
	wire _w8342_ ;
	wire _w8343_ ;
	wire _w8344_ ;
	wire _w8345_ ;
	wire _w8346_ ;
	wire _w8347_ ;
	wire _w8348_ ;
	wire _w8349_ ;
	wire _w8350_ ;
	wire _w8351_ ;
	wire _w8352_ ;
	wire _w8353_ ;
	wire _w8354_ ;
	wire _w8355_ ;
	wire _w8356_ ;
	wire _w8357_ ;
	wire _w8358_ ;
	wire _w8359_ ;
	wire _w8360_ ;
	wire _w8361_ ;
	wire _w8362_ ;
	wire _w8363_ ;
	wire _w8364_ ;
	wire _w8365_ ;
	wire _w8366_ ;
	wire _w8367_ ;
	wire _w8368_ ;
	wire _w8369_ ;
	wire _w8370_ ;
	wire _w8371_ ;
	wire _w8372_ ;
	wire _w8373_ ;
	wire _w8374_ ;
	wire _w8375_ ;
	wire _w8376_ ;
	wire _w8377_ ;
	wire _w8378_ ;
	wire _w8379_ ;
	wire _w8380_ ;
	wire _w8381_ ;
	wire _w8382_ ;
	wire _w8383_ ;
	wire _w8384_ ;
	wire _w8385_ ;
	wire _w8386_ ;
	wire _w8387_ ;
	wire _w8388_ ;
	wire _w8389_ ;
	wire _w8390_ ;
	wire _w8391_ ;
	wire _w8392_ ;
	wire _w8393_ ;
	wire _w8394_ ;
	wire _w8395_ ;
	wire _w8396_ ;
	wire _w8397_ ;
	wire _w8398_ ;
	wire _w8399_ ;
	wire _w8400_ ;
	wire _w8401_ ;
	wire _w8402_ ;
	wire _w8403_ ;
	wire _w8404_ ;
	wire _w8405_ ;
	wire _w8406_ ;
	wire _w8407_ ;
	wire _w8408_ ;
	wire _w8409_ ;
	wire _w8410_ ;
	wire _w8411_ ;
	wire _w8412_ ;
	wire _w8413_ ;
	wire _w8414_ ;
	wire _w8415_ ;
	wire _w8416_ ;
	wire _w8417_ ;
	wire _w8418_ ;
	wire _w8419_ ;
	wire _w8420_ ;
	wire _w8421_ ;
	wire _w8422_ ;
	wire _w8423_ ;
	wire _w8424_ ;
	wire _w8425_ ;
	wire _w8426_ ;
	wire _w8427_ ;
	wire _w8428_ ;
	wire _w8429_ ;
	wire _w8430_ ;
	wire _w8431_ ;
	wire _w8432_ ;
	wire _w8433_ ;
	wire _w8434_ ;
	wire _w8435_ ;
	wire _w8436_ ;
	wire _w8437_ ;
	wire _w8438_ ;
	wire _w8439_ ;
	wire _w8440_ ;
	wire _w8441_ ;
	wire _w8442_ ;
	wire _w8443_ ;
	wire _w8444_ ;
	wire _w8445_ ;
	wire _w8446_ ;
	wire _w8447_ ;
	wire _w8448_ ;
	wire _w8449_ ;
	wire _w8450_ ;
	wire _w8451_ ;
	wire _w8452_ ;
	wire _w8453_ ;
	wire _w8454_ ;
	wire _w8455_ ;
	wire _w8456_ ;
	wire _w8457_ ;
	wire _w8458_ ;
	wire _w8459_ ;
	wire _w8460_ ;
	wire _w8461_ ;
	wire _w8462_ ;
	wire _w8463_ ;
	wire _w8464_ ;
	wire _w8465_ ;
	wire _w8466_ ;
	wire _w8467_ ;
	wire _w8468_ ;
	wire _w8469_ ;
	wire _w8470_ ;
	wire _w8471_ ;
	wire _w8472_ ;
	wire _w8473_ ;
	wire _w8474_ ;
	wire _w8475_ ;
	wire _w8476_ ;
	wire _w8477_ ;
	wire _w8478_ ;
	wire _w8479_ ;
	wire _w8480_ ;
	wire _w8481_ ;
	wire _w8482_ ;
	wire _w8483_ ;
	wire _w8484_ ;
	wire _w8485_ ;
	wire _w8486_ ;
	wire _w8487_ ;
	wire _w8488_ ;
	wire _w8489_ ;
	wire _w8490_ ;
	wire _w8491_ ;
	wire _w8492_ ;
	wire _w8493_ ;
	wire _w8494_ ;
	wire _w8495_ ;
	wire _w8496_ ;
	wire _w8497_ ;
	wire _w8498_ ;
	wire _w8499_ ;
	wire _w8500_ ;
	wire _w8501_ ;
	wire _w8502_ ;
	wire _w8503_ ;
	wire _w8504_ ;
	wire _w8505_ ;
	wire _w8506_ ;
	wire _w8507_ ;
	wire _w8508_ ;
	wire _w8509_ ;
	wire _w8510_ ;
	wire _w8511_ ;
	wire _w8512_ ;
	wire _w8513_ ;
	wire _w8514_ ;
	wire _w8515_ ;
	wire _w8516_ ;
	wire _w8517_ ;
	wire _w8518_ ;
	wire _w8519_ ;
	wire _w8520_ ;
	wire _w8521_ ;
	wire _w8522_ ;
	wire _w8523_ ;
	wire _w8524_ ;
	wire _w8525_ ;
	wire _w8526_ ;
	wire _w8527_ ;
	wire _w8528_ ;
	wire _w8529_ ;
	wire _w8530_ ;
	wire _w8531_ ;
	wire _w8532_ ;
	wire _w8533_ ;
	wire _w8534_ ;
	wire _w8535_ ;
	wire _w8536_ ;
	wire _w8537_ ;
	wire _w8538_ ;
	wire _w8539_ ;
	wire _w8540_ ;
	wire _w8541_ ;
	wire _w8542_ ;
	wire _w8543_ ;
	wire _w8544_ ;
	wire _w8545_ ;
	wire _w8546_ ;
	wire _w8547_ ;
	wire _w8548_ ;
	wire _w8549_ ;
	wire _w8550_ ;
	wire _w8551_ ;
	wire _w8552_ ;
	wire _w8553_ ;
	wire _w8554_ ;
	wire _w8555_ ;
	wire _w8556_ ;
	wire _w8557_ ;
	wire _w8558_ ;
	wire _w8559_ ;
	wire _w8560_ ;
	wire _w8561_ ;
	wire _w8562_ ;
	wire _w8563_ ;
	wire _w8564_ ;
	wire _w8565_ ;
	wire _w8566_ ;
	wire _w8567_ ;
	wire _w8568_ ;
	wire _w8569_ ;
	wire _w8570_ ;
	wire _w8571_ ;
	wire _w8572_ ;
	wire _w8573_ ;
	wire _w8574_ ;
	wire _w8575_ ;
	wire _w8576_ ;
	wire _w8577_ ;
	wire _w8578_ ;
	wire _w8579_ ;
	wire _w8580_ ;
	wire _w8581_ ;
	wire _w8582_ ;
	wire _w8583_ ;
	wire _w8584_ ;
	wire _w8585_ ;
	wire _w8586_ ;
	wire _w8587_ ;
	wire _w8588_ ;
	wire _w8589_ ;
	wire _w8590_ ;
	wire _w8591_ ;
	wire _w8592_ ;
	wire _w8593_ ;
	wire _w8594_ ;
	wire _w8595_ ;
	wire _w8596_ ;
	wire _w8597_ ;
	wire _w8598_ ;
	wire _w8599_ ;
	wire _w8600_ ;
	wire _w8601_ ;
	wire _w8602_ ;
	wire _w8603_ ;
	wire _w8604_ ;
	wire _w8605_ ;
	wire _w8606_ ;
	wire _w8607_ ;
	wire _w8608_ ;
	wire _w8609_ ;
	wire _w8610_ ;
	wire _w8611_ ;
	wire _w8612_ ;
	wire _w8613_ ;
	wire _w8614_ ;
	wire _w8615_ ;
	wire _w8616_ ;
	wire _w8617_ ;
	wire _w8618_ ;
	wire _w8619_ ;
	wire _w8620_ ;
	wire _w8621_ ;
	wire _w8622_ ;
	wire _w8623_ ;
	wire _w8624_ ;
	wire _w8625_ ;
	wire _w8626_ ;
	wire _w8627_ ;
	wire _w8628_ ;
	wire _w8629_ ;
	wire _w8630_ ;
	wire _w8631_ ;
	wire _w8632_ ;
	wire _w8633_ ;
	wire _w8634_ ;
	wire _w8635_ ;
	wire _w8636_ ;
	wire _w8637_ ;
	wire _w8638_ ;
	wire _w8639_ ;
	wire _w8640_ ;
	wire _w8641_ ;
	wire _w8642_ ;
	wire _w8643_ ;
	wire _w8644_ ;
	wire _w8645_ ;
	wire _w8646_ ;
	wire _w8647_ ;
	wire _w8648_ ;
	wire _w8649_ ;
	wire _w8650_ ;
	wire _w8651_ ;
	wire _w8652_ ;
	wire _w8653_ ;
	wire _w8654_ ;
	wire _w8655_ ;
	wire _w8656_ ;
	wire _w8657_ ;
	wire _w8658_ ;
	wire _w8659_ ;
	wire _w8660_ ;
	wire _w8661_ ;
	wire _w8662_ ;
	wire _w8663_ ;
	wire _w8664_ ;
	wire _w8665_ ;
	wire _w8666_ ;
	wire _w8667_ ;
	wire _w8668_ ;
	wire _w8669_ ;
	wire _w8670_ ;
	wire _w8671_ ;
	wire _w8672_ ;
	wire _w8673_ ;
	wire _w8674_ ;
	wire _w8675_ ;
	wire _w8676_ ;
	wire _w8677_ ;
	wire _w8678_ ;
	wire _w8679_ ;
	wire _w8680_ ;
	wire _w8681_ ;
	wire _w8682_ ;
	wire _w8683_ ;
	wire _w8684_ ;
	wire _w8685_ ;
	wire _w8686_ ;
	wire _w8687_ ;
	wire _w8688_ ;
	wire _w8689_ ;
	wire _w8690_ ;
	wire _w8691_ ;
	wire _w8692_ ;
	wire _w8693_ ;
	wire _w8694_ ;
	wire _w8695_ ;
	wire _w8696_ ;
	wire _w8697_ ;
	wire _w8698_ ;
	wire _w8699_ ;
	wire _w8700_ ;
	wire _w8701_ ;
	wire _w8702_ ;
	wire _w8703_ ;
	wire _w8704_ ;
	wire _w8705_ ;
	wire _w8706_ ;
	wire _w8707_ ;
	wire _w8708_ ;
	wire _w8709_ ;
	wire _w8710_ ;
	wire _w8711_ ;
	wire _w8712_ ;
	wire _w8713_ ;
	wire _w8714_ ;
	wire _w8715_ ;
	wire _w8716_ ;
	wire _w8717_ ;
	wire _w8718_ ;
	wire _w8719_ ;
	wire _w8720_ ;
	wire _w8721_ ;
	wire _w8722_ ;
	wire _w8723_ ;
	wire _w8724_ ;
	wire _w8725_ ;
	wire _w8726_ ;
	wire _w8727_ ;
	wire _w8728_ ;
	wire _w8729_ ;
	wire _w8730_ ;
	wire _w8731_ ;
	wire _w8732_ ;
	wire _w8733_ ;
	wire _w8734_ ;
	wire _w8735_ ;
	wire _w8736_ ;
	wire _w8737_ ;
	wire _w8738_ ;
	wire _w8739_ ;
	wire _w8740_ ;
	wire _w8741_ ;
	wire _w8742_ ;
	wire _w8743_ ;
	wire _w8744_ ;
	wire _w8745_ ;
	wire _w8746_ ;
	wire _w8747_ ;
	wire _w8748_ ;
	wire _w8749_ ;
	wire _w8750_ ;
	wire _w8751_ ;
	wire _w8752_ ;
	wire _w8753_ ;
	wire _w8754_ ;
	wire _w8755_ ;
	wire _w8756_ ;
	wire _w8757_ ;
	wire _w8758_ ;
	wire _w8759_ ;
	wire _w8760_ ;
	wire _w8761_ ;
	wire _w8762_ ;
	wire _w8763_ ;
	wire _w8764_ ;
	wire _w8765_ ;
	wire _w8766_ ;
	wire _w8767_ ;
	wire _w8768_ ;
	wire _w8769_ ;
	wire _w8770_ ;
	wire _w8771_ ;
	wire _w8772_ ;
	wire _w8773_ ;
	wire _w8774_ ;
	wire _w8775_ ;
	wire _w8776_ ;
	wire _w8777_ ;
	wire _w8778_ ;
	wire _w8779_ ;
	wire _w8780_ ;
	wire _w8781_ ;
	wire _w8782_ ;
	wire _w8783_ ;
	wire _w8784_ ;
	wire _w8785_ ;
	wire _w8786_ ;
	wire _w8787_ ;
	wire _w8788_ ;
	wire _w8789_ ;
	wire _w8790_ ;
	wire _w8791_ ;
	wire _w8792_ ;
	wire _w8793_ ;
	wire _w8794_ ;
	wire _w8795_ ;
	wire _w8796_ ;
	wire _w8797_ ;
	wire _w8798_ ;
	wire _w8799_ ;
	wire _w8800_ ;
	wire _w8801_ ;
	wire _w8802_ ;
	wire _w8803_ ;
	wire _w8804_ ;
	wire _w8805_ ;
	wire _w8806_ ;
	wire _w8807_ ;
	wire _w8808_ ;
	wire _w8809_ ;
	wire _w8810_ ;
	wire _w8811_ ;
	wire _w8812_ ;
	wire _w8813_ ;
	wire _w8814_ ;
	wire _w8815_ ;
	wire _w8816_ ;
	wire _w8817_ ;
	wire _w8818_ ;
	wire _w8819_ ;
	wire _w8820_ ;
	wire _w8821_ ;
	wire _w8822_ ;
	wire _w8823_ ;
	wire _w8824_ ;
	wire _w8825_ ;
	wire _w8826_ ;
	wire _w8827_ ;
	wire _w8828_ ;
	wire _w8829_ ;
	wire _w8830_ ;
	wire _w8831_ ;
	wire _w8832_ ;
	wire _w8833_ ;
	wire _w8834_ ;
	wire _w8835_ ;
	wire _w8836_ ;
	wire _w8837_ ;
	wire _w8838_ ;
	wire _w8839_ ;
	wire _w8840_ ;
	wire _w8841_ ;
	wire _w8842_ ;
	wire _w8843_ ;
	wire _w8844_ ;
	wire _w8845_ ;
	wire _w8846_ ;
	wire _w8847_ ;
	wire _w8848_ ;
	wire _w8849_ ;
	wire _w8850_ ;
	wire _w8851_ ;
	wire _w8852_ ;
	wire _w8853_ ;
	wire _w8854_ ;
	wire _w8855_ ;
	wire _w8856_ ;
	wire _w8857_ ;
	wire _w8858_ ;
	wire _w8859_ ;
	wire _w8860_ ;
	wire _w8861_ ;
	wire _w8862_ ;
	wire _w8863_ ;
	wire _w8864_ ;
	wire _w8865_ ;
	wire _w8866_ ;
	wire _w8867_ ;
	wire _w8868_ ;
	wire _w8869_ ;
	wire _w8870_ ;
	wire _w8871_ ;
	wire _w8872_ ;
	wire _w8873_ ;
	wire _w8874_ ;
	wire _w8875_ ;
	wire _w8876_ ;
	wire _w8877_ ;
	wire _w8878_ ;
	wire _w8879_ ;
	wire _w8880_ ;
	wire _w8881_ ;
	wire _w8882_ ;
	wire _w8883_ ;
	wire _w8884_ ;
	wire _w8885_ ;
	wire _w8886_ ;
	wire _w8887_ ;
	wire _w8888_ ;
	wire _w8889_ ;
	wire _w8890_ ;
	wire _w8891_ ;
	wire _w8892_ ;
	wire _w8893_ ;
	wire _w8894_ ;
	wire _w8895_ ;
	wire _w8896_ ;
	wire _w8897_ ;
	wire _w8898_ ;
	wire _w8899_ ;
	wire _w8900_ ;
	wire _w8901_ ;
	wire _w8902_ ;
	wire _w8903_ ;
	wire _w8904_ ;
	wire _w8905_ ;
	wire _w8906_ ;
	wire _w8907_ ;
	wire _w8908_ ;
	wire _w8909_ ;
	wire _w8910_ ;
	wire _w8911_ ;
	wire _w8912_ ;
	wire _w8913_ ;
	wire _w8914_ ;
	wire _w8915_ ;
	wire _w8916_ ;
	wire _w8917_ ;
	wire _w8918_ ;
	wire _w8919_ ;
	wire _w8920_ ;
	wire _w8921_ ;
	wire _w8922_ ;
	wire _w8923_ ;
	wire _w8924_ ;
	wire _w8925_ ;
	wire _w8926_ ;
	wire _w8927_ ;
	wire _w8928_ ;
	wire _w8929_ ;
	wire _w8930_ ;
	wire _w8931_ ;
	wire _w8932_ ;
	wire _w8933_ ;
	wire _w8934_ ;
	wire _w8935_ ;
	wire _w8936_ ;
	wire _w8937_ ;
	wire _w8938_ ;
	wire _w8939_ ;
	wire _w8940_ ;
	wire _w8941_ ;
	wire _w8942_ ;
	wire _w8943_ ;
	wire _w8944_ ;
	wire _w8945_ ;
	wire _w8946_ ;
	wire _w8947_ ;
	wire _w8948_ ;
	wire _w8949_ ;
	wire _w8950_ ;
	wire _w8951_ ;
	wire _w8952_ ;
	wire _w8953_ ;
	wire _w8954_ ;
	wire _w8955_ ;
	wire _w8956_ ;
	wire _w8957_ ;
	wire _w8958_ ;
	wire _w8959_ ;
	wire _w8960_ ;
	wire _w8961_ ;
	wire _w8962_ ;
	wire _w8963_ ;
	wire _w8964_ ;
	wire _w8965_ ;
	wire _w8966_ ;
	wire _w8967_ ;
	wire _w8968_ ;
	wire _w8969_ ;
	wire _w8970_ ;
	wire _w8971_ ;
	wire _w8972_ ;
	wire _w8973_ ;
	wire _w8974_ ;
	wire _w8975_ ;
	wire _w8976_ ;
	wire _w8977_ ;
	wire _w8978_ ;
	wire _w8979_ ;
	wire _w8980_ ;
	wire _w8981_ ;
	wire _w8982_ ;
	wire _w8983_ ;
	wire _w8984_ ;
	wire _w8985_ ;
	wire _w8986_ ;
	wire _w8987_ ;
	wire _w8988_ ;
	wire _w8989_ ;
	wire _w8990_ ;
	wire _w8991_ ;
	wire _w8992_ ;
	wire _w8993_ ;
	wire _w8994_ ;
	wire _w8995_ ;
	wire _w8996_ ;
	wire _w8997_ ;
	wire _w8998_ ;
	wire _w8999_ ;
	wire _w9000_ ;
	wire _w9001_ ;
	wire _w9002_ ;
	wire _w9003_ ;
	wire _w9004_ ;
	wire _w9005_ ;
	wire _w9006_ ;
	wire _w9007_ ;
	wire _w9008_ ;
	wire _w9009_ ;
	wire _w9010_ ;
	wire _w9011_ ;
	wire _w9012_ ;
	wire _w9013_ ;
	wire _w9014_ ;
	wire _w9015_ ;
	wire _w9016_ ;
	wire _w9017_ ;
	wire _w9018_ ;
	wire _w9019_ ;
	wire _w9020_ ;
	wire _w9021_ ;
	wire _w9022_ ;
	wire _w9023_ ;
	wire _w9024_ ;
	wire _w9025_ ;
	wire _w9026_ ;
	wire _w9027_ ;
	wire _w9028_ ;
	wire _w9029_ ;
	wire _w9030_ ;
	wire _w9031_ ;
	wire _w9032_ ;
	wire _w9033_ ;
	wire _w9034_ ;
	wire _w9035_ ;
	wire _w9036_ ;
	wire _w9037_ ;
	wire _w9038_ ;
	wire _w9039_ ;
	wire _w9040_ ;
	wire _w9041_ ;
	wire _w9042_ ;
	wire _w9043_ ;
	wire _w9044_ ;
	wire _w9045_ ;
	wire _w9046_ ;
	wire _w9047_ ;
	wire _w9048_ ;
	wire _w9049_ ;
	wire _w9050_ ;
	wire _w9051_ ;
	wire _w9052_ ;
	wire _w9053_ ;
	wire _w9054_ ;
	wire _w9055_ ;
	wire _w9056_ ;
	wire _w9057_ ;
	wire _w9058_ ;
	wire _w9059_ ;
	wire _w9060_ ;
	wire _w9061_ ;
	wire _w9062_ ;
	wire _w9063_ ;
	wire _w9064_ ;
	wire _w9065_ ;
	wire _w9066_ ;
	wire _w9067_ ;
	wire _w9068_ ;
	wire _w9069_ ;
	wire _w9070_ ;
	wire _w9071_ ;
	wire _w9072_ ;
	wire _w9073_ ;
	wire _w9074_ ;
	wire _w9075_ ;
	wire _w9076_ ;
	wire _w9077_ ;
	wire _w9078_ ;
	wire _w9079_ ;
	wire _w9080_ ;
	wire _w9081_ ;
	wire _w9082_ ;
	wire _w9083_ ;
	wire _w9084_ ;
	wire _w9085_ ;
	wire _w9086_ ;
	wire _w9087_ ;
	wire _w9088_ ;
	wire _w9089_ ;
	wire _w9090_ ;
	wire _w9091_ ;
	wire _w9092_ ;
	wire _w9093_ ;
	wire _w9094_ ;
	wire _w9095_ ;
	wire _w9096_ ;
	wire _w9097_ ;
	wire _w9098_ ;
	wire _w9099_ ;
	wire _w9100_ ;
	wire _w9101_ ;
	wire _w9102_ ;
	wire _w9103_ ;
	wire _w9104_ ;
	wire _w9105_ ;
	wire _w9106_ ;
	wire _w9107_ ;
	wire _w9108_ ;
	wire _w9109_ ;
	wire _w9110_ ;
	wire _w9111_ ;
	wire _w9112_ ;
	wire _w9113_ ;
	wire _w9114_ ;
	wire _w9115_ ;
	wire _w9116_ ;
	wire _w9117_ ;
	wire _w9118_ ;
	wire _w9119_ ;
	wire _w9120_ ;
	wire _w9121_ ;
	wire _w9122_ ;
	wire _w9123_ ;
	wire _w9124_ ;
	wire _w9125_ ;
	wire _w9126_ ;
	wire _w9127_ ;
	wire _w9128_ ;
	wire _w9129_ ;
	wire _w9130_ ;
	wire _w9131_ ;
	wire _w9132_ ;
	wire _w9133_ ;
	wire _w9134_ ;
	wire _w9135_ ;
	wire _w9136_ ;
	wire _w9137_ ;
	wire _w9138_ ;
	wire _w9139_ ;
	wire _w9140_ ;
	wire _w9141_ ;
	wire _w9142_ ;
	wire _w9143_ ;
	wire _w9144_ ;
	wire _w9145_ ;
	wire _w9146_ ;
	wire _w9147_ ;
	wire _w9148_ ;
	wire _w9149_ ;
	wire _w9150_ ;
	wire _w9151_ ;
	wire _w9152_ ;
	wire _w9153_ ;
	wire _w9154_ ;
	wire _w9155_ ;
	wire _w9156_ ;
	wire _w9157_ ;
	wire _w9158_ ;
	wire _w9159_ ;
	wire _w9160_ ;
	wire _w9161_ ;
	wire _w9162_ ;
	wire _w9163_ ;
	wire _w9164_ ;
	wire _w9165_ ;
	wire _w9166_ ;
	wire _w9167_ ;
	wire _w9168_ ;
	wire _w9169_ ;
	wire _w9170_ ;
	wire _w9171_ ;
	wire _w9172_ ;
	wire _w9173_ ;
	wire _w9174_ ;
	wire _w9175_ ;
	wire _w9176_ ;
	wire _w9177_ ;
	wire _w9178_ ;
	wire _w9179_ ;
	wire _w9180_ ;
	wire _w9181_ ;
	wire _w9182_ ;
	wire _w9183_ ;
	wire _w9184_ ;
	wire _w9185_ ;
	wire _w9186_ ;
	wire _w9187_ ;
	wire _w9188_ ;
	wire _w9189_ ;
	wire _w9190_ ;
	wire _w9191_ ;
	wire _w9192_ ;
	wire _w9193_ ;
	wire _w9194_ ;
	wire _w9195_ ;
	wire _w9196_ ;
	wire _w9197_ ;
	wire _w9198_ ;
	wire _w9199_ ;
	wire _w9200_ ;
	wire _w9201_ ;
	wire _w9202_ ;
	wire _w9203_ ;
	wire _w9204_ ;
	wire _w9205_ ;
	wire _w9206_ ;
	wire _w9207_ ;
	wire _w9208_ ;
	wire _w9209_ ;
	wire _w9210_ ;
	wire _w9211_ ;
	wire _w9212_ ;
	wire _w9213_ ;
	wire _w9214_ ;
	wire _w9215_ ;
	wire _w9216_ ;
	wire _w9217_ ;
	wire _w9218_ ;
	wire _w9219_ ;
	wire _w9220_ ;
	wire _w9221_ ;
	wire _w9222_ ;
	wire _w9223_ ;
	wire _w9224_ ;
	wire _w9225_ ;
	wire _w9226_ ;
	wire _w9227_ ;
	wire _w9228_ ;
	wire _w9229_ ;
	wire _w9230_ ;
	wire _w9231_ ;
	wire _w9232_ ;
	wire _w9233_ ;
	wire _w9234_ ;
	wire _w9235_ ;
	wire _w9236_ ;
	wire _w9237_ ;
	wire _w9238_ ;
	wire _w9239_ ;
	wire _w9240_ ;
	wire _w9241_ ;
	wire _w9242_ ;
	wire _w9243_ ;
	wire _w9244_ ;
	wire _w9245_ ;
	wire _w9246_ ;
	wire _w9247_ ;
	wire _w9248_ ;
	wire _w9249_ ;
	wire _w9250_ ;
	wire _w9251_ ;
	wire _w9252_ ;
	wire _w9253_ ;
	wire _w9254_ ;
	wire _w9255_ ;
	wire _w9256_ ;
	wire _w9257_ ;
	wire _w9258_ ;
	wire _w9259_ ;
	wire _w9260_ ;
	wire _w9261_ ;
	wire _w9262_ ;
	wire _w9263_ ;
	wire _w9264_ ;
	wire _w9265_ ;
	wire _w9266_ ;
	wire _w9267_ ;
	wire _w9268_ ;
	wire _w9269_ ;
	wire _w9270_ ;
	wire _w9271_ ;
	wire _w9272_ ;
	wire _w9273_ ;
	wire _w9274_ ;
	wire _w9275_ ;
	wire _w9276_ ;
	wire _w9277_ ;
	wire _w9278_ ;
	wire _w9279_ ;
	wire _w9280_ ;
	wire _w9281_ ;
	wire _w9282_ ;
	wire _w9283_ ;
	wire _w9284_ ;
	wire _w9285_ ;
	wire _w9286_ ;
	wire _w9287_ ;
	wire _w9288_ ;
	wire _w9289_ ;
	wire _w9290_ ;
	wire _w9291_ ;
	wire _w9292_ ;
	wire _w9293_ ;
	wire _w9294_ ;
	wire _w9295_ ;
	wire _w9296_ ;
	wire _w9297_ ;
	wire _w9298_ ;
	wire _w9299_ ;
	wire _w9300_ ;
	wire _w9301_ ;
	wire _w9302_ ;
	wire _w9303_ ;
	wire _w9304_ ;
	wire _w9305_ ;
	wire _w9306_ ;
	wire _w9307_ ;
	wire _w9308_ ;
	wire _w9309_ ;
	wire _w9310_ ;
	wire _w9311_ ;
	wire _w9312_ ;
	wire _w9313_ ;
	wire _w9314_ ;
	wire _w9315_ ;
	wire _w9316_ ;
	wire _w9317_ ;
	wire _w9318_ ;
	wire _w9319_ ;
	wire _w9320_ ;
	wire _w9321_ ;
	wire _w9322_ ;
	wire _w9323_ ;
	wire _w9324_ ;
	wire _w9325_ ;
	wire _w9326_ ;
	wire _w9327_ ;
	wire _w9328_ ;
	wire _w9329_ ;
	wire _w9330_ ;
	wire _w9331_ ;
	wire _w9332_ ;
	wire _w9333_ ;
	wire _w9334_ ;
	wire _w9335_ ;
	wire _w9336_ ;
	wire _w9337_ ;
	wire _w9338_ ;
	wire _w9339_ ;
	wire _w9340_ ;
	wire _w9341_ ;
	wire _w9342_ ;
	wire _w9343_ ;
	wire _w9344_ ;
	wire _w9345_ ;
	wire _w9346_ ;
	wire _w9347_ ;
	wire _w9348_ ;
	wire _w9349_ ;
	wire _w9350_ ;
	wire _w9351_ ;
	wire _w9352_ ;
	wire _w9353_ ;
	wire _w9354_ ;
	wire _w9355_ ;
	wire _w9356_ ;
	wire _w9357_ ;
	wire _w9358_ ;
	wire _w9359_ ;
	wire _w9360_ ;
	wire _w9361_ ;
	wire _w9362_ ;
	wire _w9363_ ;
	wire _w9364_ ;
	wire _w9365_ ;
	wire _w9366_ ;
	wire _w9367_ ;
	wire _w9368_ ;
	wire _w9369_ ;
	wire _w9370_ ;
	wire _w9371_ ;
	wire _w9372_ ;
	wire _w9373_ ;
	wire _w9374_ ;
	wire _w9375_ ;
	wire _w9376_ ;
	wire _w9377_ ;
	wire _w9378_ ;
	wire _w9379_ ;
	wire _w9380_ ;
	wire _w9381_ ;
	wire _w9382_ ;
	wire _w9383_ ;
	wire _w9384_ ;
	wire _w9385_ ;
	wire _w9386_ ;
	wire _w9387_ ;
	wire _w9388_ ;
	wire _w9389_ ;
	wire _w9390_ ;
	wire _w9391_ ;
	wire _w9392_ ;
	wire _w9393_ ;
	wire _w9394_ ;
	wire _w9395_ ;
	wire _w9396_ ;
	wire _w9397_ ;
	wire _w9398_ ;
	wire _w9399_ ;
	wire _w9400_ ;
	wire _w9401_ ;
	wire _w9402_ ;
	wire _w9403_ ;
	wire _w9404_ ;
	wire _w9405_ ;
	wire _w9406_ ;
	wire _w9407_ ;
	wire _w9408_ ;
	wire _w9409_ ;
	wire _w9410_ ;
	wire _w9411_ ;
	wire _w9412_ ;
	wire _w9413_ ;
	wire _w9414_ ;
	wire _w9415_ ;
	wire _w9416_ ;
	wire _w9417_ ;
	wire _w9418_ ;
	wire _w9419_ ;
	wire _w9420_ ;
	wire _w9421_ ;
	wire _w9422_ ;
	wire _w9423_ ;
	wire _w9424_ ;
	wire _w9425_ ;
	wire _w9426_ ;
	wire _w9427_ ;
	wire _w9428_ ;
	wire _w9429_ ;
	wire _w9430_ ;
	wire _w9431_ ;
	wire _w9432_ ;
	wire _w9433_ ;
	wire _w9434_ ;
	wire _w9435_ ;
	wire _w9436_ ;
	wire _w9437_ ;
	wire _w9438_ ;
	wire _w9439_ ;
	wire _w9440_ ;
	wire _w9441_ ;
	wire _w9442_ ;
	wire _w9443_ ;
	wire _w9444_ ;
	wire _w9445_ ;
	wire _w9446_ ;
	wire _w9447_ ;
	wire _w9448_ ;
	wire _w9449_ ;
	wire _w9450_ ;
	wire _w9451_ ;
	wire _w9452_ ;
	wire _w9453_ ;
	wire _w9454_ ;
	wire _w9455_ ;
	wire _w9456_ ;
	wire _w9457_ ;
	wire _w9458_ ;
	wire _w9459_ ;
	wire _w9460_ ;
	wire _w9461_ ;
	wire _w9462_ ;
	wire _w9463_ ;
	wire _w9464_ ;
	wire _w9465_ ;
	wire _w9466_ ;
	wire _w9467_ ;
	wire _w9468_ ;
	wire _w9469_ ;
	wire _w9470_ ;
	wire _w9471_ ;
	wire _w9472_ ;
	wire _w9473_ ;
	wire _w9474_ ;
	wire _w9475_ ;
	wire _w9476_ ;
	wire _w9477_ ;
	wire _w9478_ ;
	wire _w9479_ ;
	wire _w9480_ ;
	wire _w9481_ ;
	wire _w9482_ ;
	wire _w9483_ ;
	wire _w9484_ ;
	wire _w9485_ ;
	wire _w9486_ ;
	wire _w9487_ ;
	wire _w9488_ ;
	wire _w9489_ ;
	wire _w9490_ ;
	wire _w9491_ ;
	wire _w9492_ ;
	wire _w9493_ ;
	wire _w9494_ ;
	wire _w9495_ ;
	wire _w9496_ ;
	wire _w9497_ ;
	wire _w9498_ ;
	wire _w9499_ ;
	wire _w9500_ ;
	wire _w9501_ ;
	wire _w9502_ ;
	wire _w9503_ ;
	wire _w9504_ ;
	wire _w9505_ ;
	wire _w9506_ ;
	wire _w9507_ ;
	wire _w9508_ ;
	wire _w9509_ ;
	wire _w9510_ ;
	wire _w9511_ ;
	wire _w9512_ ;
	wire _w9513_ ;
	wire _w9514_ ;
	wire _w9515_ ;
	wire _w9516_ ;
	wire _w9517_ ;
	wire _w9518_ ;
	wire _w9519_ ;
	wire _w9520_ ;
	wire _w9521_ ;
	wire _w9522_ ;
	wire _w9523_ ;
	wire _w9524_ ;
	wire _w9525_ ;
	wire _w9526_ ;
	wire _w9527_ ;
	wire _w9528_ ;
	wire _w9529_ ;
	wire _w9530_ ;
	wire _w9531_ ;
	wire _w9532_ ;
	wire _w9533_ ;
	wire _w9534_ ;
	wire _w9535_ ;
	wire _w9536_ ;
	wire _w9537_ ;
	wire _w9538_ ;
	wire _w9539_ ;
	wire _w9540_ ;
	wire _w9541_ ;
	wire _w9542_ ;
	wire _w9543_ ;
	wire _w9544_ ;
	wire _w9545_ ;
	wire _w9546_ ;
	wire _w9547_ ;
	wire _w9548_ ;
	wire _w9549_ ;
	wire _w9550_ ;
	wire _w9551_ ;
	wire _w9552_ ;
	wire _w9553_ ;
	wire _w9554_ ;
	wire _w9555_ ;
	wire _w9556_ ;
	wire _w9557_ ;
	wire _w9558_ ;
	wire _w9559_ ;
	wire _w9560_ ;
	wire _w9561_ ;
	wire _w9562_ ;
	wire _w9563_ ;
	wire _w9564_ ;
	wire _w9565_ ;
	wire _w9566_ ;
	wire _w9567_ ;
	wire _w9568_ ;
	wire _w9569_ ;
	wire _w9570_ ;
	wire _w9571_ ;
	wire _w9572_ ;
	wire _w9573_ ;
	wire _w9574_ ;
	wire _w9575_ ;
	wire _w9576_ ;
	wire _w9577_ ;
	wire _w9578_ ;
	wire _w9579_ ;
	wire _w9580_ ;
	wire _w9581_ ;
	wire _w9582_ ;
	wire _w9583_ ;
	wire _w9584_ ;
	wire _w9585_ ;
	wire _w9586_ ;
	wire _w9587_ ;
	wire _w9588_ ;
	wire _w9589_ ;
	wire _w9590_ ;
	wire _w9591_ ;
	wire _w9592_ ;
	wire _w9593_ ;
	wire _w9594_ ;
	wire _w9595_ ;
	wire _w9596_ ;
	wire _w9597_ ;
	wire _w9598_ ;
	wire _w9599_ ;
	wire _w9600_ ;
	wire _w9601_ ;
	wire _w9602_ ;
	wire _w9603_ ;
	wire _w9604_ ;
	wire _w9605_ ;
	wire _w9606_ ;
	wire _w9607_ ;
	wire _w9608_ ;
	wire _w9609_ ;
	wire _w9610_ ;
	wire _w9611_ ;
	wire _w9612_ ;
	wire _w9613_ ;
	wire _w9614_ ;
	wire _w9615_ ;
	wire _w9616_ ;
	wire _w9617_ ;
	wire _w9618_ ;
	wire _w9619_ ;
	wire _w9620_ ;
	wire _w9621_ ;
	wire _w9622_ ;
	wire _w9623_ ;
	wire _w9624_ ;
	wire _w9625_ ;
	wire _w9626_ ;
	wire _w9627_ ;
	wire _w9628_ ;
	wire _w9629_ ;
	wire _w9630_ ;
	wire _w9631_ ;
	wire _w9632_ ;
	wire _w9633_ ;
	wire _w9634_ ;
	wire _w9635_ ;
	wire _w9636_ ;
	wire _w9637_ ;
	wire _w9638_ ;
	wire _w9639_ ;
	wire _w9640_ ;
	wire _w9641_ ;
	wire _w9642_ ;
	wire _w9643_ ;
	wire _w9644_ ;
	wire _w9645_ ;
	wire _w9646_ ;
	wire _w9647_ ;
	wire _w9648_ ;
	wire _w9649_ ;
	wire _w9650_ ;
	wire _w9651_ ;
	wire _w9652_ ;
	wire _w9653_ ;
	wire _w9654_ ;
	wire _w9655_ ;
	wire _w9656_ ;
	wire _w9657_ ;
	wire _w9658_ ;
	wire _w9659_ ;
	wire _w9660_ ;
	wire _w9661_ ;
	wire _w9662_ ;
	wire _w9663_ ;
	wire _w9664_ ;
	wire _w9665_ ;
	wire _w9666_ ;
	wire _w9667_ ;
	wire _w9668_ ;
	wire _w9669_ ;
	wire _w9670_ ;
	wire _w9671_ ;
	wire _w9672_ ;
	wire _w9673_ ;
	wire _w9674_ ;
	wire _w9675_ ;
	wire _w9676_ ;
	wire _w9677_ ;
	wire _w9678_ ;
	wire _w9679_ ;
	wire _w9680_ ;
	wire _w9681_ ;
	wire _w9682_ ;
	wire _w9683_ ;
	wire _w9684_ ;
	wire _w9685_ ;
	wire _w9686_ ;
	wire _w9687_ ;
	wire _w9688_ ;
	wire _w9689_ ;
	wire _w9690_ ;
	wire _w9691_ ;
	wire _w9692_ ;
	wire _w9693_ ;
	wire _w9694_ ;
	wire _w9695_ ;
	wire _w9696_ ;
	wire _w9697_ ;
	wire _w9698_ ;
	wire _w9699_ ;
	wire _w9700_ ;
	wire _w9701_ ;
	wire _w9702_ ;
	wire _w9703_ ;
	wire _w9704_ ;
	wire _w9705_ ;
	wire _w9706_ ;
	wire _w9707_ ;
	wire _w9708_ ;
	wire _w9709_ ;
	wire _w9710_ ;
	wire _w9711_ ;
	wire _w9712_ ;
	wire _w9713_ ;
	wire _w9714_ ;
	wire _w9715_ ;
	wire _w9716_ ;
	wire _w9717_ ;
	wire _w9718_ ;
	wire _w9719_ ;
	wire _w9720_ ;
	wire _w9721_ ;
	wire _w9722_ ;
	wire _w9723_ ;
	wire _w9724_ ;
	wire _w9725_ ;
	wire _w9726_ ;
	wire _w9727_ ;
	wire _w9728_ ;
	wire _w9729_ ;
	wire _w9730_ ;
	wire _w9731_ ;
	wire _w9732_ ;
	wire _w9733_ ;
	wire _w9734_ ;
	wire _w9735_ ;
	wire _w9736_ ;
	wire _w9737_ ;
	wire _w9738_ ;
	wire _w9739_ ;
	wire _w9740_ ;
	wire _w9741_ ;
	wire _w9742_ ;
	wire _w9743_ ;
	wire _w9744_ ;
	wire _w9745_ ;
	wire _w9746_ ;
	wire _w9747_ ;
	wire _w9748_ ;
	wire _w9749_ ;
	wire _w9750_ ;
	wire _w9751_ ;
	wire _w9752_ ;
	wire _w9753_ ;
	wire _w9754_ ;
	wire _w9755_ ;
	wire _w9756_ ;
	wire _w9757_ ;
	wire _w9758_ ;
	wire _w9759_ ;
	wire _w9760_ ;
	wire _w9761_ ;
	wire _w9762_ ;
	wire _w9763_ ;
	wire _w9764_ ;
	wire _w9765_ ;
	wire _w9766_ ;
	wire _w9767_ ;
	wire _w9768_ ;
	wire _w9769_ ;
	wire _w9770_ ;
	wire _w9771_ ;
	wire _w9772_ ;
	wire _w9773_ ;
	wire _w9774_ ;
	wire _w9775_ ;
	wire _w9776_ ;
	wire _w9777_ ;
	wire _w9778_ ;
	wire _w9779_ ;
	wire _w9780_ ;
	wire _w9781_ ;
	wire _w9782_ ;
	wire _w9783_ ;
	wire _w9784_ ;
	wire _w9785_ ;
	wire _w9786_ ;
	wire _w9787_ ;
	wire _w9788_ ;
	wire _w9789_ ;
	wire _w9790_ ;
	wire _w9791_ ;
	wire _w9792_ ;
	wire _w9793_ ;
	wire _w9794_ ;
	wire _w9795_ ;
	wire _w9796_ ;
	wire _w9797_ ;
	wire _w9798_ ;
	wire _w9799_ ;
	wire _w9800_ ;
	wire _w9801_ ;
	wire _w9802_ ;
	wire _w9803_ ;
	wire _w9804_ ;
	wire _w9805_ ;
	wire _w9806_ ;
	wire _w9807_ ;
	wire _w9808_ ;
	wire _w9809_ ;
	wire _w9810_ ;
	wire _w9811_ ;
	wire _w9812_ ;
	wire _w9813_ ;
	wire _w9814_ ;
	wire _w9815_ ;
	wire _w9816_ ;
	wire _w9817_ ;
	wire _w9818_ ;
	wire _w9819_ ;
	wire _w9820_ ;
	wire _w9821_ ;
	wire _w9822_ ;
	wire _w9823_ ;
	wire _w9824_ ;
	wire _w9825_ ;
	wire _w9826_ ;
	wire _w9827_ ;
	wire _w9828_ ;
	wire _w9829_ ;
	wire _w9830_ ;
	wire _w9831_ ;
	wire _w9832_ ;
	wire _w9833_ ;
	wire _w9834_ ;
	wire _w9835_ ;
	wire _w9836_ ;
	wire _w9837_ ;
	wire _w9838_ ;
	wire _w9839_ ;
	wire _w9840_ ;
	wire _w9841_ ;
	wire _w9842_ ;
	wire _w9843_ ;
	wire _w9844_ ;
	wire _w9845_ ;
	wire _w9846_ ;
	wire _w9847_ ;
	wire _w9848_ ;
	wire _w9849_ ;
	wire _w9850_ ;
	wire _w9851_ ;
	wire _w9852_ ;
	wire _w9853_ ;
	wire _w9854_ ;
	wire _w9855_ ;
	wire _w9856_ ;
	wire _w9857_ ;
	wire _w9858_ ;
	wire _w9859_ ;
	wire _w9860_ ;
	wire _w9861_ ;
	wire _w9862_ ;
	wire _w9863_ ;
	wire _w9864_ ;
	wire _w9865_ ;
	wire _w9866_ ;
	wire _w9867_ ;
	wire _w9868_ ;
	wire _w9869_ ;
	wire _w9870_ ;
	wire _w9871_ ;
	wire _w9872_ ;
	wire _w9873_ ;
	wire _w9874_ ;
	wire _w9875_ ;
	wire _w9876_ ;
	wire _w9877_ ;
	wire _w9878_ ;
	wire _w9879_ ;
	wire _w9880_ ;
	wire _w9881_ ;
	wire _w9882_ ;
	wire _w9883_ ;
	wire _w9884_ ;
	wire _w9885_ ;
	wire _w9886_ ;
	wire _w9887_ ;
	wire _w9888_ ;
	wire _w9889_ ;
	wire _w9890_ ;
	wire _w9891_ ;
	wire _w9892_ ;
	wire _w9893_ ;
	wire _w9894_ ;
	wire _w9895_ ;
	wire _w9896_ ;
	wire _w9897_ ;
	wire _w9898_ ;
	wire _w9899_ ;
	wire _w9900_ ;
	wire _w9901_ ;
	wire _w9902_ ;
	wire _w9903_ ;
	wire _w9904_ ;
	wire _w9905_ ;
	wire _w9906_ ;
	wire _w9907_ ;
	wire _w9908_ ;
	wire _w9909_ ;
	wire _w9910_ ;
	wire _w9911_ ;
	wire _w9912_ ;
	wire _w9913_ ;
	wire _w9914_ ;
	wire _w9915_ ;
	wire _w9916_ ;
	wire _w9917_ ;
	wire _w9918_ ;
	wire _w9919_ ;
	wire _w9920_ ;
	wire _w9921_ ;
	wire _w9922_ ;
	wire _w9923_ ;
	wire _w9924_ ;
	wire _w9925_ ;
	wire _w9926_ ;
	wire _w9927_ ;
	wire _w9928_ ;
	wire _w9929_ ;
	wire _w9930_ ;
	wire _w9931_ ;
	wire _w9932_ ;
	wire _w9933_ ;
	wire _w9934_ ;
	wire _w9935_ ;
	wire _w9936_ ;
	wire _w9937_ ;
	wire _w9938_ ;
	wire _w9939_ ;
	wire _w9940_ ;
	wire _w9941_ ;
	wire _w9942_ ;
	wire _w9943_ ;
	wire _w9944_ ;
	wire _w9945_ ;
	wire _w9946_ ;
	wire _w9947_ ;
	wire _w9948_ ;
	wire _w9949_ ;
	wire _w9950_ ;
	wire _w9951_ ;
	wire _w9952_ ;
	wire _w9953_ ;
	wire _w9954_ ;
	wire _w9955_ ;
	wire _w9956_ ;
	wire _w9957_ ;
	wire _w9958_ ;
	wire _w9959_ ;
	wire _w9960_ ;
	wire _w9961_ ;
	wire _w9962_ ;
	wire _w9963_ ;
	wire _w9964_ ;
	wire _w9965_ ;
	wire _w9966_ ;
	wire _w9967_ ;
	wire _w9968_ ;
	wire _w9969_ ;
	wire _w9970_ ;
	wire _w9971_ ;
	wire _w9972_ ;
	wire _w9973_ ;
	wire _w9974_ ;
	wire _w9975_ ;
	wire _w9976_ ;
	wire _w9977_ ;
	wire _w9978_ ;
	wire _w9979_ ;
	wire _w9980_ ;
	wire _w9981_ ;
	wire _w9982_ ;
	wire _w9983_ ;
	wire _w9984_ ;
	wire _w9985_ ;
	wire _w9986_ ;
	wire _w9987_ ;
	wire _w9988_ ;
	wire _w9989_ ;
	wire _w9990_ ;
	wire _w9991_ ;
	wire _w9992_ ;
	wire _w9993_ ;
	wire _w9994_ ;
	wire _w9995_ ;
	wire _w9996_ ;
	wire _w9997_ ;
	wire _w9998_ ;
	wire _w9999_ ;
	wire _w10000_ ;
	wire _w10001_ ;
	wire _w10002_ ;
	wire _w10003_ ;
	wire _w10004_ ;
	wire _w10005_ ;
	wire _w10006_ ;
	wire _w10007_ ;
	wire _w10008_ ;
	wire _w10009_ ;
	wire _w10010_ ;
	wire _w10011_ ;
	wire _w10012_ ;
	wire _w10013_ ;
	wire _w10014_ ;
	wire _w10015_ ;
	wire _w10016_ ;
	wire _w10017_ ;
	wire _w10018_ ;
	wire _w10019_ ;
	wire _w10020_ ;
	wire _w10021_ ;
	wire _w10022_ ;
	wire _w10023_ ;
	wire _w10024_ ;
	wire _w10025_ ;
	wire _w10026_ ;
	wire _w10027_ ;
	wire _w10028_ ;
	wire _w10029_ ;
	wire _w10030_ ;
	wire _w10031_ ;
	wire _w10032_ ;
	wire _w10033_ ;
	wire _w10034_ ;
	wire _w10035_ ;
	wire _w10036_ ;
	wire _w10037_ ;
	wire _w10038_ ;
	wire _w10039_ ;
	wire _w10040_ ;
	wire _w10041_ ;
	wire _w10042_ ;
	wire _w10043_ ;
	wire _w10044_ ;
	wire _w10045_ ;
	wire _w10046_ ;
	wire _w10047_ ;
	wire _w10048_ ;
	wire _w10049_ ;
	wire _w10050_ ;
	wire _w10051_ ;
	wire _w10052_ ;
	wire _w10053_ ;
	wire _w10054_ ;
	wire _w10055_ ;
	wire _w10056_ ;
	wire _w10057_ ;
	wire _w10058_ ;
	wire _w10059_ ;
	wire _w10060_ ;
	wire _w10061_ ;
	wire _w10062_ ;
	wire _w10063_ ;
	wire _w10064_ ;
	wire _w10065_ ;
	wire _w10066_ ;
	wire _w10067_ ;
	wire _w10068_ ;
	wire _w10069_ ;
	wire _w10070_ ;
	wire _w10071_ ;
	wire _w10072_ ;
	wire _w10073_ ;
	wire _w10074_ ;
	wire _w10075_ ;
	wire _w10076_ ;
	wire _w10077_ ;
	wire _w10078_ ;
	wire _w10079_ ;
	wire _w10080_ ;
	wire _w10081_ ;
	wire _w10082_ ;
	wire _w10083_ ;
	wire _w10084_ ;
	wire _w10085_ ;
	wire _w10086_ ;
	wire _w10087_ ;
	wire _w10088_ ;
	wire _w10089_ ;
	wire _w10090_ ;
	wire _w10091_ ;
	wire _w10092_ ;
	wire _w10093_ ;
	wire _w10094_ ;
	wire _w10095_ ;
	wire _w10096_ ;
	wire _w10097_ ;
	wire _w10098_ ;
	wire _w10099_ ;
	wire _w10100_ ;
	wire _w10101_ ;
	wire _w10102_ ;
	wire _w10103_ ;
	wire _w10104_ ;
	wire _w10105_ ;
	wire _w10106_ ;
	wire _w10107_ ;
	wire _w10108_ ;
	wire _w10109_ ;
	wire _w10110_ ;
	wire _w10111_ ;
	wire _w10112_ ;
	wire _w10113_ ;
	wire _w10114_ ;
	wire _w10115_ ;
	wire _w10116_ ;
	wire _w10117_ ;
	wire _w10118_ ;
	wire _w10119_ ;
	wire _w10120_ ;
	wire _w10121_ ;
	wire _w10122_ ;
	wire _w10123_ ;
	wire _w10124_ ;
	wire _w10125_ ;
	wire _w10126_ ;
	wire _w10127_ ;
	wire _w10128_ ;
	wire _w10129_ ;
	wire _w10130_ ;
	wire _w10131_ ;
	wire _w10132_ ;
	wire _w10133_ ;
	wire _w10134_ ;
	wire _w10135_ ;
	wire _w10136_ ;
	wire _w10137_ ;
	wire _w10138_ ;
	wire _w10139_ ;
	wire _w10140_ ;
	wire _w10141_ ;
	wire _w10142_ ;
	wire _w10143_ ;
	wire _w10144_ ;
	wire _w10145_ ;
	wire _w10146_ ;
	wire _w10147_ ;
	wire _w10148_ ;
	wire _w10149_ ;
	wire _w10150_ ;
	wire _w10151_ ;
	wire _w10152_ ;
	wire _w10153_ ;
	wire _w10154_ ;
	wire _w10155_ ;
	wire _w10156_ ;
	wire _w10157_ ;
	wire _w10158_ ;
	wire _w10159_ ;
	wire _w10160_ ;
	wire _w10161_ ;
	wire _w10162_ ;
	wire _w10163_ ;
	wire _w10164_ ;
	wire _w10165_ ;
	wire _w10166_ ;
	wire _w10167_ ;
	wire _w10168_ ;
	wire _w10169_ ;
	wire _w10170_ ;
	wire _w10171_ ;
	wire _w10172_ ;
	wire _w10173_ ;
	wire _w10174_ ;
	wire _w10175_ ;
	wire _w10176_ ;
	wire _w10177_ ;
	wire _w10178_ ;
	wire _w10179_ ;
	wire _w10180_ ;
	wire _w10181_ ;
	wire _w10182_ ;
	wire _w10183_ ;
	wire _w10184_ ;
	wire _w10185_ ;
	wire _w10186_ ;
	wire _w10187_ ;
	wire _w10188_ ;
	wire _w10189_ ;
	wire _w10190_ ;
	wire _w10191_ ;
	wire _w10192_ ;
	wire _w10193_ ;
	wire _w10194_ ;
	wire _w10195_ ;
	wire _w10196_ ;
	wire _w10197_ ;
	wire _w10198_ ;
	wire _w10199_ ;
	wire _w10200_ ;
	wire _w10201_ ;
	wire _w10202_ ;
	wire _w10203_ ;
	wire _w10204_ ;
	wire _w10205_ ;
	wire _w10206_ ;
	wire _w10207_ ;
	wire _w10208_ ;
	wire _w10209_ ;
	wire _w10210_ ;
	wire _w10211_ ;
	wire _w10212_ ;
	wire _w10213_ ;
	wire _w10214_ ;
	wire _w10215_ ;
	wire _w10216_ ;
	wire _w10217_ ;
	wire _w10218_ ;
	wire _w10219_ ;
	wire _w10220_ ;
	wire _w10221_ ;
	wire _w10222_ ;
	wire _w10223_ ;
	wire _w10224_ ;
	wire _w10225_ ;
	wire _w10226_ ;
	wire _w10227_ ;
	wire _w10228_ ;
	wire _w10229_ ;
	wire _w10230_ ;
	wire _w10231_ ;
	wire _w10232_ ;
	wire _w10233_ ;
	wire _w10234_ ;
	wire _w10235_ ;
	wire _w10236_ ;
	wire _w10237_ ;
	wire _w10238_ ;
	wire _w10239_ ;
	wire _w10240_ ;
	wire _w10241_ ;
	wire _w10242_ ;
	wire _w10243_ ;
	wire _w10244_ ;
	wire _w10245_ ;
	wire _w10246_ ;
	wire _w10247_ ;
	wire _w10248_ ;
	wire _w10249_ ;
	wire _w10250_ ;
	wire _w10251_ ;
	wire _w10252_ ;
	wire _w10253_ ;
	wire _w10254_ ;
	wire _w10255_ ;
	wire _w10256_ ;
	wire _w10257_ ;
	wire _w10258_ ;
	wire _w10259_ ;
	wire _w10260_ ;
	wire _w10261_ ;
	wire _w10262_ ;
	wire _w10263_ ;
	wire _w10264_ ;
	wire _w10265_ ;
	wire _w10266_ ;
	wire _w10267_ ;
	wire _w10268_ ;
	wire _w10269_ ;
	wire _w10270_ ;
	wire _w10271_ ;
	wire _w10272_ ;
	wire _w10273_ ;
	wire _w10274_ ;
	wire _w10275_ ;
	wire _w10276_ ;
	wire _w10277_ ;
	wire _w10278_ ;
	wire _w10279_ ;
	wire _w10280_ ;
	wire _w10281_ ;
	wire _w10282_ ;
	wire _w10283_ ;
	wire _w10284_ ;
	wire _w10285_ ;
	wire _w10286_ ;
	wire _w10287_ ;
	wire _w10288_ ;
	wire _w10289_ ;
	wire _w10290_ ;
	wire _w10291_ ;
	wire _w10292_ ;
	wire _w10293_ ;
	wire _w10294_ ;
	wire _w10295_ ;
	wire _w10296_ ;
	wire _w10297_ ;
	wire _w10298_ ;
	wire _w10299_ ;
	wire _w10300_ ;
	wire _w10301_ ;
	wire _w10302_ ;
	wire _w10303_ ;
	wire _w10304_ ;
	wire _w10305_ ;
	wire _w10306_ ;
	wire _w10307_ ;
	wire _w10308_ ;
	wire _w10309_ ;
	wire _w10310_ ;
	wire _w10311_ ;
	wire _w10312_ ;
	wire _w10313_ ;
	wire _w10314_ ;
	wire _w10315_ ;
	wire _w10316_ ;
	wire _w10317_ ;
	wire _w10318_ ;
	wire _w10319_ ;
	wire _w10320_ ;
	wire _w10321_ ;
	wire _w10322_ ;
	wire _w10323_ ;
	wire _w10324_ ;
	wire _w10325_ ;
	wire _w10326_ ;
	wire _w10327_ ;
	wire _w10328_ ;
	wire _w10329_ ;
	wire _w10330_ ;
	wire _w10331_ ;
	wire _w10332_ ;
	wire _w10333_ ;
	wire _w10334_ ;
	wire _w10335_ ;
	wire _w10336_ ;
	wire _w10337_ ;
	wire _w10338_ ;
	wire _w10339_ ;
	wire _w10340_ ;
	wire _w10341_ ;
	wire _w10342_ ;
	wire _w10343_ ;
	wire _w10344_ ;
	wire _w10345_ ;
	wire _w10346_ ;
	wire _w10347_ ;
	wire _w10348_ ;
	wire _w10349_ ;
	wire _w10350_ ;
	wire _w10351_ ;
	wire _w10352_ ;
	wire _w10353_ ;
	wire _w10354_ ;
	wire _w10355_ ;
	wire _w10356_ ;
	wire _w10357_ ;
	wire _w10358_ ;
	wire _w10359_ ;
	wire _w10360_ ;
	wire _w10361_ ;
	wire _w10362_ ;
	wire _w10363_ ;
	wire _w10364_ ;
	wire _w10365_ ;
	wire _w10366_ ;
	wire _w10367_ ;
	wire _w10368_ ;
	wire _w10369_ ;
	wire _w10370_ ;
	wire _w10371_ ;
	wire _w10372_ ;
	wire _w10373_ ;
	wire _w10374_ ;
	wire _w10375_ ;
	wire _w10376_ ;
	wire _w10377_ ;
	wire _w10378_ ;
	wire _w10379_ ;
	wire _w10380_ ;
	wire _w10381_ ;
	wire _w10382_ ;
	wire _w10383_ ;
	wire _w10384_ ;
	wire _w10385_ ;
	wire _w10386_ ;
	wire _w10387_ ;
	wire _w10388_ ;
	wire _w10389_ ;
	wire _w10390_ ;
	wire _w10391_ ;
	wire _w10392_ ;
	wire _w10393_ ;
	wire _w10394_ ;
	wire _w10395_ ;
	wire _w10396_ ;
	wire _w10397_ ;
	wire _w10398_ ;
	wire _w10399_ ;
	wire _w10400_ ;
	wire _w10401_ ;
	wire _w10402_ ;
	wire _w10403_ ;
	wire _w10404_ ;
	wire _w10405_ ;
	wire _w10406_ ;
	wire _w10407_ ;
	wire _w10408_ ;
	wire _w10409_ ;
	wire _w10410_ ;
	wire _w10411_ ;
	wire _w10412_ ;
	wire _w10413_ ;
	wire _w10414_ ;
	wire _w10415_ ;
	wire _w10416_ ;
	wire _w10417_ ;
	wire _w10418_ ;
	wire _w10419_ ;
	wire _w10420_ ;
	wire _w10421_ ;
	wire _w10422_ ;
	wire _w10423_ ;
	wire _w10424_ ;
	wire _w10425_ ;
	wire _w10426_ ;
	wire _w10427_ ;
	wire _w10428_ ;
	wire _w10429_ ;
	wire _w10430_ ;
	wire _w10431_ ;
	wire _w10432_ ;
	wire _w10433_ ;
	wire _w10434_ ;
	wire _w10435_ ;
	wire _w10436_ ;
	wire _w10437_ ;
	wire _w10438_ ;
	wire _w10439_ ;
	wire _w10440_ ;
	wire _w10441_ ;
	wire _w10442_ ;
	wire _w10443_ ;
	wire _w10444_ ;
	wire _w10445_ ;
	wire _w10446_ ;
	wire _w10447_ ;
	wire _w10448_ ;
	wire _w10449_ ;
	wire _w10450_ ;
	wire _w10451_ ;
	wire _w10452_ ;
	wire _w10453_ ;
	wire _w10454_ ;
	wire _w10455_ ;
	wire _w10456_ ;
	wire _w10457_ ;
	wire _w10458_ ;
	wire _w10459_ ;
	wire _w10460_ ;
	wire _w10461_ ;
	wire _w10462_ ;
	wire _w10463_ ;
	wire _w10464_ ;
	wire _w10465_ ;
	wire _w10466_ ;
	wire _w10467_ ;
	wire _w10468_ ;
	wire _w10469_ ;
	wire _w10470_ ;
	wire _w10471_ ;
	wire _w10472_ ;
	wire _w10473_ ;
	wire _w10474_ ;
	wire _w10475_ ;
	wire _w10476_ ;
	wire _w10477_ ;
	wire _w10478_ ;
	wire _w10479_ ;
	wire _w10480_ ;
	wire _w10481_ ;
	wire _w10482_ ;
	wire _w10483_ ;
	wire _w10484_ ;
	wire _w10485_ ;
	wire _w10486_ ;
	wire _w10487_ ;
	wire _w10488_ ;
	wire _w10489_ ;
	wire _w10490_ ;
	wire _w10491_ ;
	wire _w10492_ ;
	wire _w10493_ ;
	wire _w10494_ ;
	wire _w10495_ ;
	wire _w10496_ ;
	wire _w10497_ ;
	wire _w10498_ ;
	wire _w10499_ ;
	wire _w10500_ ;
	wire _w10501_ ;
	wire _w10502_ ;
	wire _w10503_ ;
	wire _w10504_ ;
	wire _w10505_ ;
	wire _w10506_ ;
	wire _w10507_ ;
	wire _w10508_ ;
	wire _w10509_ ;
	wire _w10510_ ;
	wire _w10511_ ;
	wire _w10512_ ;
	wire _w10513_ ;
	wire _w10514_ ;
	wire _w10515_ ;
	wire _w10516_ ;
	wire _w10517_ ;
	wire _w10518_ ;
	wire _w10519_ ;
	wire _w10520_ ;
	wire _w10521_ ;
	wire _w10522_ ;
	wire _w10523_ ;
	wire _w10524_ ;
	wire _w10525_ ;
	wire _w10526_ ;
	wire _w10527_ ;
	wire _w10528_ ;
	wire _w10529_ ;
	wire _w10530_ ;
	wire _w10531_ ;
	wire _w10532_ ;
	wire _w10533_ ;
	wire _w10534_ ;
	wire _w10535_ ;
	wire _w10536_ ;
	wire _w10537_ ;
	wire _w10538_ ;
	wire _w10539_ ;
	wire _w10540_ ;
	wire _w10541_ ;
	wire _w10542_ ;
	wire _w10543_ ;
	wire _w10544_ ;
	wire _w10545_ ;
	wire _w10546_ ;
	wire _w10547_ ;
	wire _w10548_ ;
	wire _w10549_ ;
	wire _w10550_ ;
	wire _w10551_ ;
	wire _w10552_ ;
	wire _w10553_ ;
	wire _w10554_ ;
	wire _w10555_ ;
	wire _w10556_ ;
	wire _w10557_ ;
	wire _w10558_ ;
	wire _w10559_ ;
	wire _w10560_ ;
	wire _w10561_ ;
	wire _w10562_ ;
	wire _w10563_ ;
	wire _w10564_ ;
	wire _w10565_ ;
	wire _w10566_ ;
	wire _w10567_ ;
	wire _w10568_ ;
	wire _w10569_ ;
	wire _w10570_ ;
	wire _w10571_ ;
	wire _w10572_ ;
	wire _w10573_ ;
	wire _w10574_ ;
	wire _w10575_ ;
	wire _w10576_ ;
	wire _w10577_ ;
	wire _w10578_ ;
	wire _w10579_ ;
	wire _w10580_ ;
	wire _w10581_ ;
	wire _w10582_ ;
	wire _w10583_ ;
	wire _w10584_ ;
	wire _w10585_ ;
	wire _w10586_ ;
	wire _w10587_ ;
	wire _w10588_ ;
	wire _w10589_ ;
	wire _w10590_ ;
	wire _w10591_ ;
	wire _w10592_ ;
	wire _w10593_ ;
	wire _w10594_ ;
	wire _w10595_ ;
	wire _w10596_ ;
	wire _w10597_ ;
	wire _w10598_ ;
	wire _w10599_ ;
	wire _w10600_ ;
	wire _w10601_ ;
	wire _w10602_ ;
	wire _w10603_ ;
	wire _w10604_ ;
	wire _w10605_ ;
	wire _w10606_ ;
	wire _w10607_ ;
	wire _w10608_ ;
	wire _w10609_ ;
	wire _w10610_ ;
	wire _w10611_ ;
	wire _w10612_ ;
	wire _w10613_ ;
	wire _w10614_ ;
	wire _w10615_ ;
	wire _w10616_ ;
	wire _w10617_ ;
	wire _w10618_ ;
	wire _w10619_ ;
	wire _w10620_ ;
	wire _w10621_ ;
	wire _w10622_ ;
	wire _w10623_ ;
	wire _w10624_ ;
	wire _w10625_ ;
	wire _w10626_ ;
	wire _w10627_ ;
	wire _w10628_ ;
	wire _w10629_ ;
	wire _w10630_ ;
	wire _w10631_ ;
	wire _w10632_ ;
	wire _w10633_ ;
	wire _w10634_ ;
	wire _w10635_ ;
	wire _w10636_ ;
	wire _w10637_ ;
	wire _w10638_ ;
	wire _w10639_ ;
	wire _w10640_ ;
	wire _w10641_ ;
	wire _w10642_ ;
	wire _w10643_ ;
	wire _w10644_ ;
	wire _w10645_ ;
	wire _w10646_ ;
	wire _w10647_ ;
	wire _w10648_ ;
	wire _w10649_ ;
	wire _w10650_ ;
	wire _w10651_ ;
	wire _w10652_ ;
	wire _w10653_ ;
	wire _w10654_ ;
	wire _w10655_ ;
	wire _w10656_ ;
	wire _w10657_ ;
	wire _w10658_ ;
	wire _w10659_ ;
	wire _w10660_ ;
	wire _w10661_ ;
	wire _w10662_ ;
	wire _w10663_ ;
	wire _w10664_ ;
	wire _w10665_ ;
	wire _w10666_ ;
	wire _w10667_ ;
	wire _w10668_ ;
	wire _w10669_ ;
	wire _w10670_ ;
	wire _w10671_ ;
	wire _w10672_ ;
	wire _w10673_ ;
	wire _w10674_ ;
	wire _w10675_ ;
	wire _w10676_ ;
	wire _w10677_ ;
	wire _w10678_ ;
	wire _w10679_ ;
	wire _w10680_ ;
	wire _w10681_ ;
	wire _w10682_ ;
	wire _w10683_ ;
	wire _w10684_ ;
	wire _w10685_ ;
	wire _w10686_ ;
	wire _w10687_ ;
	wire _w10688_ ;
	wire _w10689_ ;
	wire _w10690_ ;
	wire _w10691_ ;
	wire _w10692_ ;
	wire _w10693_ ;
	wire _w10694_ ;
	wire _w10695_ ;
	wire _w10696_ ;
	wire _w10697_ ;
	wire _w10698_ ;
	wire _w10699_ ;
	wire _w10700_ ;
	wire _w10701_ ;
	wire _w10702_ ;
	wire _w10703_ ;
	wire _w10704_ ;
	wire _w10705_ ;
	wire _w10706_ ;
	wire _w10707_ ;
	wire _w10708_ ;
	wire _w10709_ ;
	wire _w10710_ ;
	wire _w10711_ ;
	wire _w10712_ ;
	wire _w10713_ ;
	wire _w10714_ ;
	wire _w10715_ ;
	wire _w10716_ ;
	wire _w10717_ ;
	wire _w10718_ ;
	wire _w10719_ ;
	wire _w10720_ ;
	wire _w10721_ ;
	wire _w10722_ ;
	wire _w10723_ ;
	wire _w10724_ ;
	wire _w10725_ ;
	wire _w10726_ ;
	wire _w10727_ ;
	wire _w10728_ ;
	wire _w10729_ ;
	wire _w10730_ ;
	wire _w10731_ ;
	wire _w10732_ ;
	wire _w10733_ ;
	wire _w10734_ ;
	wire _w10735_ ;
	wire _w10736_ ;
	wire _w10737_ ;
	wire _w10738_ ;
	wire _w10739_ ;
	wire _w10740_ ;
	wire _w10741_ ;
	wire _w10742_ ;
	wire _w10743_ ;
	wire _w10744_ ;
	wire _w10745_ ;
	wire _w10746_ ;
	wire _w10747_ ;
	wire _w10748_ ;
	wire _w10749_ ;
	wire _w10750_ ;
	wire _w10751_ ;
	wire _w10752_ ;
	wire _w10753_ ;
	wire _w10754_ ;
	wire _w10755_ ;
	wire _w10756_ ;
	wire _w10757_ ;
	wire _w10758_ ;
	wire _w10759_ ;
	wire _w10760_ ;
	wire _w10761_ ;
	wire _w10762_ ;
	wire _w10763_ ;
	wire _w10764_ ;
	wire _w10765_ ;
	wire _w10766_ ;
	wire _w10767_ ;
	wire _w10768_ ;
	wire _w10769_ ;
	wire _w10770_ ;
	wire _w10771_ ;
	wire _w10772_ ;
	wire _w10773_ ;
	wire _w10774_ ;
	wire _w10775_ ;
	wire _w10776_ ;
	wire _w10777_ ;
	wire _w10778_ ;
	wire _w10779_ ;
	wire _w10780_ ;
	wire _w10781_ ;
	wire _w10782_ ;
	wire _w10783_ ;
	wire _w10784_ ;
	wire _w10785_ ;
	wire _w10786_ ;
	wire _w10787_ ;
	wire _w10788_ ;
	wire _w10789_ ;
	wire _w10790_ ;
	wire _w10791_ ;
	wire _w10792_ ;
	wire _w10793_ ;
	wire _w10794_ ;
	wire _w10795_ ;
	wire _w10796_ ;
	wire _w10797_ ;
	wire _w10798_ ;
	wire _w10799_ ;
	wire _w10800_ ;
	wire _w10801_ ;
	wire _w10802_ ;
	wire _w10803_ ;
	wire _w10804_ ;
	wire _w10805_ ;
	wire _w10806_ ;
	wire _w10807_ ;
	wire _w10808_ ;
	wire _w10809_ ;
	wire _w10810_ ;
	wire _w10811_ ;
	wire _w10812_ ;
	wire _w10813_ ;
	wire _w10814_ ;
	wire _w10815_ ;
	wire _w10816_ ;
	wire _w10817_ ;
	wire _w10818_ ;
	wire _w10819_ ;
	wire _w10820_ ;
	wire _w10821_ ;
	wire _w10822_ ;
	wire _w10823_ ;
	wire _w10824_ ;
	wire _w10825_ ;
	wire _w10826_ ;
	wire _w10827_ ;
	wire _w10828_ ;
	wire _w10829_ ;
	wire _w10830_ ;
	wire _w10831_ ;
	wire _w10832_ ;
	wire _w10833_ ;
	wire _w10834_ ;
	wire _w10835_ ;
	wire _w10836_ ;
	wire _w10837_ ;
	wire _w10838_ ;
	wire _w10839_ ;
	wire _w10840_ ;
	wire _w10841_ ;
	wire _w10842_ ;
	wire _w10843_ ;
	wire _w10844_ ;
	wire _w10845_ ;
	wire _w10846_ ;
	wire _w10847_ ;
	wire _w10848_ ;
	wire _w10849_ ;
	wire _w10850_ ;
	wire _w10851_ ;
	wire _w10852_ ;
	wire _w10853_ ;
	wire _w10854_ ;
	wire _w10855_ ;
	wire _w10856_ ;
	wire _w10857_ ;
	wire _w10858_ ;
	wire _w10859_ ;
	wire _w10860_ ;
	wire _w10861_ ;
	wire _w10862_ ;
	wire _w10863_ ;
	wire _w10864_ ;
	wire _w10865_ ;
	wire _w10866_ ;
	wire _w10867_ ;
	wire _w10868_ ;
	wire _w10869_ ;
	wire _w10870_ ;
	wire _w10871_ ;
	wire _w10872_ ;
	wire _w10873_ ;
	wire _w10874_ ;
	wire _w10875_ ;
	wire _w10876_ ;
	wire _w10877_ ;
	wire _w10878_ ;
	wire _w10879_ ;
	wire _w10880_ ;
	wire _w10881_ ;
	wire _w10882_ ;
	wire _w10883_ ;
	wire _w10884_ ;
	wire _w10885_ ;
	wire _w10886_ ;
	wire _w10887_ ;
	wire _w10888_ ;
	wire _w10889_ ;
	wire _w10890_ ;
	wire _w10891_ ;
	wire _w10892_ ;
	wire _w10893_ ;
	wire _w10894_ ;
	wire _w10895_ ;
	wire _w10896_ ;
	wire _w10897_ ;
	wire _w10898_ ;
	wire _w10899_ ;
	wire _w10900_ ;
	wire _w10901_ ;
	wire _w10902_ ;
	wire _w10903_ ;
	wire _w10904_ ;
	wire _w10905_ ;
	wire _w10906_ ;
	wire _w10907_ ;
	wire _w10908_ ;
	wire _w10909_ ;
	wire _w10910_ ;
	wire _w10911_ ;
	wire _w10912_ ;
	wire _w10913_ ;
	wire _w16100_ ;
	wire _w16101_ ;
	wire _w16102_ ;
	wire _w16103_ ;
	wire _w16104_ ;
	wire _w16105_ ;
	wire _w16106_ ;
	wire _w16107_ ;
	wire _w16108_ ;
	wire _w16109_ ;
	wire _w16110_ ;
	wire _w16111_ ;
	wire _w16112_ ;
	wire _w16113_ ;
	wire _w16114_ ;
	wire _w16115_ ;
	wire _w16116_ ;
	wire _w16117_ ;
	wire _w16118_ ;
	wire _w16119_ ;
	wire _w16120_ ;
	wire _w16121_ ;
	wire _w16122_ ;
	wire _w16123_ ;
	wire _w16124_ ;
	wire _w16125_ ;
	wire _w16126_ ;
	wire _w16127_ ;
	wire _w16128_ ;
	wire _w16129_ ;
	wire _w16130_ ;
	wire _w16131_ ;
	wire _w16132_ ;
	wire _w16133_ ;
	wire _w16134_ ;
	wire _w16135_ ;
	wire _w16136_ ;
	wire _w16137_ ;
	wire _w16138_ ;
	wire _w16139_ ;
	wire _w16140_ ;
	wire _w16141_ ;
	wire _w16142_ ;
	wire _w16143_ ;
	wire _w16144_ ;
	wire _w16145_ ;
	wire _w16146_ ;
	wire _w16147_ ;
	wire _w16148_ ;
	wire _w16149_ ;
	wire _w16150_ ;
	wire _w16151_ ;
	wire _w16152_ ;
	wire _w16153_ ;
	wire _w16154_ ;
	wire _w16155_ ;
	wire _w16156_ ;
	wire _w16157_ ;
	wire _w16158_ ;
	wire _w16159_ ;
	wire _w16160_ ;
	wire _w16161_ ;
	wire _w16162_ ;
	wire _w16163_ ;
	wire _w16164_ ;
	wire _w16165_ ;
	wire _w16166_ ;
	wire _w16167_ ;
	wire _w16168_ ;
	wire _w16169_ ;
	wire _w16170_ ;
	wire _w16171_ ;
	wire _w16172_ ;
	wire _w16173_ ;
	wire _w16174_ ;
	wire _w16175_ ;
	wire _w16176_ ;
	wire _w16177_ ;
	wire _w16178_ ;
	wire _w16179_ ;
	wire _w16180_ ;
	wire _w16181_ ;
	wire _w16182_ ;
	wire _w16183_ ;
	wire _w16184_ ;
	wire _w16185_ ;
	wire _w16186_ ;
	wire _w16187_ ;
	wire _w16188_ ;
	wire _w16189_ ;
	wire _w16190_ ;
	wire _w16191_ ;
	wire _w16192_ ;
	wire _w16193_ ;
	wire _w16194_ ;
	wire _w16195_ ;
	wire _w16196_ ;
	wire _w16197_ ;
	wire _w16198_ ;
	wire _w16199_ ;
	wire _w16200_ ;
	wire _w16201_ ;
	wire _w16202_ ;
	wire _w16203_ ;
	wire _w16204_ ;
	wire _w16205_ ;
	wire _w16206_ ;
	wire _w16207_ ;
	wire _w16208_ ;
	wire _w16209_ ;
	wire _w16210_ ;
	wire _w16211_ ;
	wire _w16212_ ;
	wire _w16213_ ;
	wire _w16214_ ;
	wire _w16215_ ;
	wire _w16216_ ;
	wire _w16217_ ;
	wire _w16218_ ;
	wire _w16219_ ;
	wire _w16220_ ;
	wire _w16221_ ;
	wire _w16222_ ;
	wire _w16223_ ;
	wire _w16224_ ;
	wire _w16225_ ;
	wire _w16226_ ;
	wire _w16227_ ;
	wire _w16228_ ;
	wire _w16229_ ;
	wire _w16230_ ;
	wire _w16231_ ;
	wire _w16232_ ;
	wire _w16233_ ;
	wire _w16234_ ;
	wire _w16235_ ;
	wire _w16236_ ;
	wire _w16237_ ;
	wire _w16238_ ;
	wire _w16239_ ;
	wire _w16240_ ;
	wire _w16241_ ;
	wire _w16242_ ;
	wire _w16243_ ;
	wire _w16244_ ;
	wire _w16245_ ;
	wire _w16246_ ;
	wire _w16247_ ;
	wire _w16248_ ;
	wire _w16249_ ;
	wire _w16250_ ;
	wire _w16251_ ;
	wire _w16252_ ;
	wire _w16253_ ;
	wire _w16254_ ;
	wire _w16255_ ;
	wire _w16256_ ;
	wire _w16257_ ;
	wire _w16258_ ;
	wire _w16259_ ;
	wire _w16260_ ;
	wire _w16261_ ;
	wire _w16262_ ;
	wire _w16263_ ;
	wire _w16264_ ;
	wire _w16265_ ;
	wire _w16266_ ;
	wire _w16267_ ;
	wire _w16268_ ;
	wire _w16269_ ;
	wire _w16270_ ;
	wire _w16271_ ;
	wire _w16272_ ;
	wire _w16273_ ;
	wire _w16274_ ;
	wire _w16275_ ;
	wire _w16276_ ;
	wire _w16277_ ;
	wire _w16278_ ;
	wire _w16279_ ;
	wire _w16280_ ;
	wire _w16281_ ;
	wire _w16282_ ;
	wire _w16283_ ;
	wire _w16284_ ;
	wire _w16285_ ;
	wire _w16286_ ;
	wire _w16287_ ;
	wire _w16288_ ;
	wire _w16289_ ;
	wire _w16290_ ;
	wire _w16291_ ;
	wire _w16292_ ;
	wire _w16293_ ;
	wire _w16294_ ;
	wire _w16295_ ;
	wire _w16296_ ;
	wire _w16297_ ;
	wire _w16298_ ;
	wire _w16299_ ;
	wire _w16300_ ;
	wire _w16301_ ;
	wire _w16302_ ;
	wire _w16303_ ;
	wire _w16304_ ;
	wire _w16305_ ;
	wire _w16306_ ;
	wire _w16307_ ;
	wire _w16308_ ;
	wire _w16309_ ;
	wire _w16310_ ;
	wire _w16311_ ;
	wire _w16312_ ;
	wire _w16313_ ;
	wire _w16314_ ;
	wire _w16315_ ;
	wire _w16316_ ;
	wire _w16317_ ;
	wire _w16318_ ;
	wire _w16319_ ;
	wire _w16320_ ;
	wire _w16321_ ;
	wire _w16322_ ;
	wire _w16323_ ;
	wire _w16324_ ;
	wire _w16325_ ;
	wire _w16326_ ;
	wire _w16327_ ;
	wire _w16328_ ;
	wire _w16329_ ;
	wire _w16330_ ;
	wire _w16331_ ;
	wire _w16332_ ;
	wire _w16333_ ;
	wire _w16334_ ;
	wire _w16335_ ;
	wire _w16336_ ;
	wire _w16337_ ;
	wire _w16338_ ;
	wire _w16339_ ;
	wire _w16340_ ;
	wire _w16341_ ;
	wire _w16342_ ;
	wire _w16343_ ;
	wire _w16344_ ;
	wire _w16345_ ;
	wire _w16346_ ;
	wire _w16347_ ;
	wire _w16348_ ;
	wire _w16349_ ;
	wire _w16350_ ;
	wire _w16351_ ;
	wire _w16352_ ;
	wire _w16353_ ;
	wire _w16354_ ;
	wire _w16355_ ;
	wire _w16356_ ;
	wire _w16357_ ;
	wire _w16358_ ;
	wire _w16359_ ;
	wire _w16360_ ;
	wire _w16361_ ;
	wire _w16362_ ;
	wire _w16363_ ;
	wire _w16364_ ;
	wire _w16365_ ;
	wire _w16366_ ;
	wire _w16367_ ;
	wire _w16368_ ;
	wire _w16369_ ;
	wire _w16370_ ;
	wire _w16371_ ;
	wire _w16372_ ;
	wire _w16373_ ;
	wire _w16374_ ;
	wire _w16375_ ;
	wire _w16376_ ;
	wire _w16377_ ;
	wire _w16378_ ;
	wire _w16379_ ;
	wire _w16380_ ;
	wire _w16381_ ;
	wire _w16382_ ;
	wire _w16383_ ;
	wire _w16384_ ;
	wire _w16385_ ;
	wire _w16386_ ;
	wire _w16387_ ;
	wire _w16388_ ;
	wire _w16389_ ;
	wire _w16390_ ;
	wire _w16391_ ;
	wire _w16392_ ;
	wire _w16393_ ;
	wire _w16394_ ;
	wire _w16395_ ;
	wire _w16396_ ;
	wire _w16397_ ;
	wire _w16398_ ;
	wire _w16399_ ;
	wire _w16400_ ;
	wire _w16401_ ;
	wire _w16402_ ;
	wire _w16403_ ;
	wire _w16404_ ;
	wire _w16405_ ;
	wire _w16406_ ;
	wire _w16407_ ;
	wire _w16408_ ;
	wire _w16409_ ;
	wire _w16410_ ;
	wire _w16411_ ;
	wire _w16412_ ;
	wire _w16413_ ;
	wire _w16414_ ;
	wire _w16415_ ;
	wire _w16416_ ;
	wire _w16417_ ;
	wire _w16418_ ;
	wire _w16419_ ;
	wire _w16420_ ;
	wire _w16421_ ;
	wire _w16422_ ;
	wire _w16423_ ;
	wire _w16424_ ;
	wire _w16425_ ;
	wire _w16426_ ;
	wire _w16427_ ;
	wire _w16428_ ;
	wire _w16429_ ;
	wire _w16430_ ;
	wire _w16431_ ;
	wire _w16432_ ;
	wire _w16433_ ;
	wire _w16434_ ;
	wire _w16435_ ;
	wire _w16436_ ;
	wire _w16437_ ;
	wire _w16438_ ;
	wire _w16439_ ;
	wire _w16440_ ;
	wire _w16441_ ;
	wire _w16442_ ;
	wire _w16443_ ;
	wire _w16444_ ;
	wire _w16445_ ;
	wire _w16446_ ;
	wire _w16447_ ;
	wire _w16448_ ;
	wire _w16449_ ;
	wire _w16450_ ;
	wire _w16451_ ;
	wire _w16452_ ;
	wire _w16453_ ;
	wire _w16454_ ;
	wire _w16455_ ;
	wire _w16456_ ;
	wire _w16457_ ;
	wire _w16458_ ;
	wire _w16459_ ;
	wire _w16460_ ;
	wire _w16461_ ;
	wire _w16462_ ;
	wire _w16463_ ;
	wire _w16464_ ;
	wire _w16465_ ;
	wire _w16466_ ;
	wire _w16467_ ;
	wire _w16468_ ;
	wire _w16469_ ;
	wire _w16470_ ;
	wire _w16471_ ;
	wire _w16472_ ;
	wire _w16473_ ;
	wire _w16474_ ;
	wire _w16475_ ;
	wire _w16476_ ;
	wire _w16477_ ;
	wire _w16478_ ;
	wire _w16479_ ;
	wire _w16480_ ;
	wire _w16481_ ;
	wire _w16482_ ;
	wire _w16483_ ;
	wire _w16484_ ;
	wire _w16485_ ;
	wire _w16486_ ;
	wire _w16487_ ;
	wire _w16488_ ;
	wire _w16489_ ;
	wire _w16490_ ;
	wire _w16491_ ;
	wire _w16492_ ;
	wire _w16493_ ;
	wire _w16494_ ;
	wire _w16495_ ;
	wire _w16496_ ;
	wire _w16497_ ;
	wire _w16498_ ;
	wire _w16499_ ;
	wire _w16500_ ;
	wire _w16501_ ;
	wire _w16502_ ;
	wire _w16503_ ;
	wire _w16504_ ;
	wire _w16505_ ;
	wire _w16506_ ;
	wire _w16507_ ;
	wire _w16508_ ;
	wire _w16509_ ;
	wire _w16510_ ;
	wire _w16511_ ;
	wire _w16512_ ;
	wire _w16513_ ;
	wire _w16514_ ;
	wire _w16515_ ;
	wire _w16516_ ;
	wire _w16517_ ;
	wire _w16518_ ;
	wire _w16519_ ;
	wire _w16520_ ;
	wire _w16521_ ;
	wire _w16522_ ;
	wire _w16523_ ;
	wire _w16524_ ;
	wire _w16525_ ;
	wire _w16526_ ;
	wire _w16527_ ;
	wire _w16528_ ;
	wire _w16529_ ;
	wire _w16530_ ;
	wire _w16531_ ;
	wire _w16532_ ;
	wire _w16533_ ;
	wire _w16534_ ;
	wire _w16535_ ;
	wire _w16536_ ;
	wire _w16537_ ;
	wire _w16538_ ;
	wire _w16539_ ;
	wire _w16540_ ;
	wire _w16541_ ;
	wire _w16542_ ;
	wire _w16543_ ;
	wire _w16544_ ;
	wire _w16545_ ;
	wire _w16546_ ;
	wire _w16547_ ;
	wire _w16548_ ;
	wire _w16549_ ;
	wire _w16550_ ;
	wire _w16551_ ;
	wire _w16552_ ;
	wire _w16553_ ;
	wire _w16554_ ;
	wire _w16555_ ;
	wire _w16556_ ;
	wire _w16557_ ;
	wire _w16558_ ;
	wire _w16559_ ;
	wire _w16560_ ;
	wire _w16561_ ;
	wire _w16562_ ;
	wire _w16563_ ;
	wire _w16564_ ;
	wire _w16565_ ;
	wire _w16566_ ;
	wire _w16567_ ;
	wire _w16568_ ;
	wire _w16569_ ;
	wire _w16570_ ;
	wire _w16571_ ;
	wire _w16572_ ;
	wire _w16573_ ;
	wire _w16574_ ;
	wire _w16575_ ;
	wire _w16576_ ;
	wire _w16577_ ;
	wire _w16578_ ;
	wire _w16579_ ;
	wire _w16580_ ;
	wire _w16581_ ;
	wire _w16582_ ;
	wire _w16583_ ;
	wire _w16584_ ;
	wire _w16585_ ;
	wire _w16586_ ;
	wire _w16587_ ;
	wire _w16588_ ;
	wire _w16589_ ;
	wire _w16590_ ;
	wire _w16591_ ;
	wire _w16592_ ;
	wire _w16593_ ;
	wire _w16594_ ;
	wire _w16595_ ;
	wire _w16596_ ;
	wire _w16597_ ;
	wire _w16598_ ;
	wire _w16599_ ;
	wire _w16600_ ;
	wire _w16601_ ;
	wire _w16602_ ;
	wire _w16603_ ;
	wire _w16604_ ;
	wire _w16605_ ;
	wire _w16606_ ;
	wire _w16607_ ;
	wire _w16608_ ;
	wire _w16609_ ;
	wire _w16610_ ;
	wire _w16611_ ;
	wire _w16612_ ;
	wire _w16613_ ;
	wire _w16614_ ;
	wire _w16615_ ;
	wire _w16616_ ;
	wire _w16617_ ;
	wire _w16618_ ;
	wire _w16619_ ;
	wire _w16620_ ;
	wire _w16621_ ;
	wire _w16622_ ;
	wire _w16623_ ;
	wire _w16624_ ;
	wire _w16625_ ;
	wire _w16626_ ;
	wire _w16627_ ;
	wire _w16628_ ;
	wire _w16629_ ;
	wire _w16630_ ;
	wire _w16631_ ;
	wire _w16632_ ;
	wire _w16633_ ;
	wire _w16634_ ;
	wire _w16635_ ;
	wire _w16636_ ;
	wire _w16637_ ;
	wire _w16638_ ;
	wire _w16639_ ;
	wire _w16640_ ;
	wire _w16641_ ;
	wire _w16642_ ;
	wire _w16643_ ;
	wire _w16644_ ;
	wire _w16645_ ;
	wire _w16646_ ;
	wire _w16647_ ;
	wire _w16648_ ;
	wire _w16649_ ;
	wire _w16650_ ;
	wire _w16651_ ;
	wire _w16652_ ;
	wire _w16653_ ;
	wire _w16654_ ;
	wire _w16655_ ;
	wire _w16656_ ;
	wire _w16657_ ;
	wire _w16658_ ;
	wire _w16659_ ;
	wire _w16660_ ;
	wire _w16661_ ;
	wire _w16662_ ;
	wire _w16663_ ;
	wire _w16664_ ;
	wire _w16665_ ;
	wire _w16666_ ;
	wire _w16667_ ;
	wire _w16668_ ;
	wire _w16669_ ;
	wire _w16670_ ;
	wire _w16671_ ;
	wire _w16672_ ;
	wire _w16673_ ;
	wire _w16674_ ;
	wire _w16675_ ;
	wire _w16676_ ;
	wire _w16677_ ;
	wire _w16678_ ;
	wire _w16679_ ;
	wire _w16680_ ;
	wire _w16681_ ;
	wire _w16682_ ;
	wire _w16683_ ;
	wire _w16684_ ;
	wire _w16685_ ;
	wire _w16686_ ;
	wire _w16687_ ;
	wire _w16688_ ;
	wire _w16689_ ;
	wire _w16690_ ;
	wire _w16691_ ;
	wire _w16692_ ;
	wire _w16693_ ;
	wire _w16694_ ;
	wire _w16695_ ;
	wire _w16696_ ;
	wire _w16697_ ;
	wire _w16698_ ;
	wire _w16699_ ;
	wire _w16700_ ;
	wire _w16701_ ;
	wire _w16702_ ;
	wire _w16703_ ;
	wire _w16704_ ;
	wire _w16705_ ;
	wire _w16706_ ;
	wire _w16707_ ;
	wire _w16708_ ;
	wire _w16709_ ;
	wire _w16710_ ;
	wire _w16711_ ;
	wire _w16712_ ;
	wire _w16713_ ;
	wire _w16714_ ;
	wire _w16715_ ;
	wire _w16716_ ;
	wire _w16717_ ;
	wire _w16718_ ;
	wire _w16719_ ;
	wire _w16720_ ;
	wire _w16721_ ;
	wire _w16722_ ;
	wire _w16723_ ;
	wire _w16724_ ;
	wire _w16725_ ;
	wire _w16726_ ;
	wire _w16727_ ;
	wire _w16728_ ;
	wire _w16729_ ;
	wire _w16730_ ;
	wire _w16731_ ;
	wire _w16732_ ;
	wire _w16733_ ;
	wire _w16734_ ;
	wire _w16735_ ;
	wire _w16736_ ;
	wire _w16737_ ;
	wire _w16738_ ;
	wire _w16739_ ;
	wire _w16740_ ;
	wire _w16741_ ;
	wire _w16742_ ;
	wire _w16743_ ;
	wire _w16744_ ;
	wire _w16745_ ;
	wire _w16746_ ;
	wire _w16747_ ;
	wire _w16748_ ;
	wire _w16749_ ;
	wire _w16750_ ;
	wire _w16751_ ;
	wire _w16752_ ;
	wire _w16753_ ;
	wire _w16754_ ;
	wire _w16755_ ;
	wire _w16756_ ;
	wire _w16757_ ;
	wire _w16758_ ;
	wire _w16759_ ;
	wire _w16760_ ;
	wire _w16761_ ;
	wire _w16762_ ;
	wire _w16763_ ;
	wire _w16764_ ;
	wire _w16765_ ;
	wire _w16766_ ;
	wire _w16767_ ;
	wire _w16768_ ;
	wire _w16769_ ;
	wire _w16770_ ;
	wire _w16771_ ;
	wire _w16772_ ;
	wire _w16773_ ;
	wire _w16774_ ;
	wire _w16775_ ;
	wire _w16776_ ;
	wire _w16777_ ;
	wire _w16778_ ;
	wire _w16779_ ;
	wire _w16780_ ;
	wire _w16781_ ;
	wire _w16782_ ;
	wire _w16783_ ;
	wire _w16784_ ;
	wire _w16785_ ;
	wire _w16786_ ;
	wire _w16787_ ;
	wire _w16788_ ;
	wire _w16789_ ;
	wire _w16790_ ;
	wire _w16791_ ;
	wire _w16792_ ;
	wire _w16793_ ;
	wire _w16794_ ;
	wire _w16795_ ;
	wire _w16796_ ;
	wire _w16797_ ;
	wire _w16798_ ;
	wire _w16799_ ;
	wire _w16800_ ;
	wire _w16801_ ;
	wire _w16802_ ;
	wire _w16803_ ;
	wire _w16804_ ;
	wire _w16805_ ;
	wire _w16806_ ;
	wire _w16807_ ;
	wire _w16808_ ;
	wire _w16809_ ;
	wire _w16810_ ;
	wire _w16811_ ;
	wire _w16812_ ;
	wire _w16813_ ;
	wire _w16814_ ;
	wire _w16815_ ;
	wire _w16816_ ;
	wire _w16817_ ;
	wire _w16818_ ;
	wire _w16819_ ;
	wire _w16820_ ;
	wire _w16821_ ;
	wire _w16822_ ;
	wire _w16823_ ;
	wire _w16824_ ;
	wire _w16825_ ;
	wire _w16826_ ;
	wire _w16827_ ;
	wire _w16828_ ;
	wire _w16829_ ;
	wire _w16830_ ;
	wire _w16831_ ;
	wire _w16832_ ;
	wire _w16833_ ;
	wire _w16834_ ;
	wire _w16835_ ;
	wire _w16836_ ;
	wire _w16837_ ;
	wire _w16838_ ;
	wire _w16839_ ;
	wire _w16840_ ;
	wire _w16841_ ;
	wire _w16842_ ;
	wire _w16843_ ;
	wire _w16844_ ;
	wire _w16845_ ;
	wire _w16846_ ;
	wire _w16847_ ;
	wire _w16848_ ;
	wire _w16849_ ;
	wire _w16850_ ;
	wire _w16851_ ;
	wire _w16852_ ;
	wire _w16853_ ;
	wire _w16854_ ;
	wire _w16855_ ;
	wire _w16856_ ;
	wire _w16857_ ;
	wire _w16858_ ;
	wire _w16859_ ;
	wire _w16860_ ;
	wire _w16861_ ;
	wire _w16862_ ;
	wire _w16863_ ;
	wire _w16864_ ;
	wire _w16865_ ;
	wire _w16866_ ;
	wire _w16867_ ;
	wire _w16868_ ;
	wire _w16869_ ;
	wire _w16870_ ;
	wire _w16871_ ;
	wire _w16872_ ;
	wire _w16873_ ;
	wire _w16874_ ;
	wire _w16875_ ;
	wire _w16876_ ;
	wire _w16877_ ;
	wire _w16878_ ;
	wire _w16879_ ;
	wire _w16880_ ;
	wire _w16881_ ;
	wire _w16882_ ;
	wire _w16883_ ;
	wire _w16884_ ;
	wire _w16885_ ;
	wire _w16886_ ;
	wire _w16887_ ;
	wire _w16888_ ;
	wire _w16889_ ;
	wire _w16890_ ;
	wire _w16891_ ;
	wire _w16892_ ;
	wire _w16893_ ;
	wire _w16894_ ;
	wire _w16895_ ;
	wire _w16896_ ;
	wire _w16897_ ;
	wire _w16898_ ;
	wire _w16899_ ;
	wire _w16900_ ;
	wire _w16901_ ;
	wire _w16902_ ;
	wire _w16903_ ;
	wire _w16904_ ;
	wire _w16905_ ;
	wire _w16906_ ;
	wire _w16907_ ;
	wire _w16908_ ;
	wire _w16909_ ;
	wire _w16910_ ;
	wire _w16911_ ;
	wire _w16912_ ;
	wire _w16913_ ;
	wire _w16914_ ;
	wire _w16915_ ;
	wire _w16916_ ;
	wire _w16917_ ;
	wire _w16918_ ;
	wire _w16919_ ;
	wire _w16920_ ;
	wire _w16921_ ;
	wire _w16922_ ;
	wire _w16923_ ;
	wire _w16924_ ;
	wire _w16925_ ;
	wire _w16926_ ;
	wire _w16927_ ;
	wire _w16928_ ;
	wire _w16929_ ;
	wire _w16930_ ;
	wire _w16931_ ;
	wire _w16932_ ;
	wire _w16933_ ;
	wire _w16934_ ;
	wire _w16935_ ;
	wire _w16936_ ;
	wire _w16937_ ;
	wire _w16938_ ;
	wire _w16939_ ;
	wire _w16940_ ;
	wire _w16941_ ;
	wire _w16942_ ;
	wire _w16943_ ;
	wire _w16944_ ;
	wire _w16945_ ;
	wire _w16946_ ;
	wire _w16947_ ;
	wire _w16948_ ;
	wire _w16949_ ;
	wire _w16950_ ;
	wire _w16951_ ;
	wire _w16952_ ;
	wire _w16953_ ;
	wire _w16954_ ;
	wire _w16955_ ;
	wire _w16956_ ;
	wire _w16957_ ;
	wire _w16958_ ;
	wire _w16959_ ;
	wire _w16960_ ;
	wire _w16961_ ;
	wire _w16962_ ;
	wire _w16963_ ;
	wire _w16964_ ;
	wire _w16965_ ;
	wire _w16966_ ;
	wire _w16967_ ;
	wire _w16968_ ;
	wire _w16969_ ;
	wire _w16970_ ;
	wire _w16971_ ;
	wire _w16972_ ;
	wire _w16973_ ;
	wire _w16974_ ;
	wire _w16975_ ;
	wire _w16976_ ;
	wire _w16977_ ;
	wire _w16978_ ;
	wire _w16979_ ;
	wire _w16980_ ;
	wire _w16981_ ;
	wire _w16982_ ;
	wire _w16983_ ;
	wire _w16984_ ;
	wire _w16985_ ;
	wire _w16986_ ;
	wire _w16987_ ;
	wire _w16988_ ;
	wire _w16989_ ;
	wire _w16990_ ;
	wire _w16991_ ;
	wire _w16992_ ;
	wire _w16993_ ;
	wire _w16994_ ;
	wire _w16995_ ;
	wire _w16996_ ;
	wire _w16997_ ;
	wire _w16998_ ;
	wire _w16999_ ;
	wire _w17000_ ;
	wire _w17001_ ;
	wire _w17002_ ;
	wire _w17003_ ;
	wire _w17004_ ;
	wire _w17005_ ;
	wire _w17006_ ;
	wire _w17007_ ;
	wire _w17008_ ;
	wire _w17009_ ;
	wire _w17010_ ;
	wire _w17011_ ;
	wire _w17012_ ;
	wire _w17013_ ;
	wire _w17014_ ;
	wire _w17015_ ;
	wire _w17016_ ;
	wire _w17017_ ;
	wire _w17018_ ;
	wire _w17019_ ;
	wire _w17020_ ;
	wire _w17021_ ;
	wire _w17022_ ;
	wire _w17023_ ;
	wire _w17024_ ;
	wire _w17025_ ;
	wire _w17026_ ;
	wire _w17027_ ;
	wire _w17028_ ;
	wire _w17029_ ;
	wire _w17030_ ;
	wire _w17031_ ;
	wire _w17032_ ;
	wire _w17033_ ;
	wire _w17034_ ;
	wire _w17035_ ;
	wire _w17036_ ;
	wire _w17037_ ;
	wire _w17038_ ;
	wire _w17039_ ;
	wire _w17040_ ;
	wire _w17041_ ;
	wire _w17042_ ;
	wire _w17043_ ;
	wire _w17044_ ;
	wire _w17045_ ;
	wire _w17046_ ;
	wire _w17047_ ;
	wire _w17048_ ;
	wire _w17049_ ;
	wire _w17050_ ;
	wire _w17051_ ;
	wire _w17052_ ;
	wire _w17053_ ;
	wire _w17054_ ;
	wire _w17055_ ;
	wire _w17056_ ;
	wire _w17057_ ;
	wire _w17058_ ;
	wire _w17059_ ;
	wire _w17060_ ;
	wire _w17061_ ;
	wire _w17062_ ;
	wire _w17063_ ;
	wire _w17064_ ;
	wire _w17065_ ;
	wire _w17066_ ;
	wire _w17067_ ;
	wire _w17068_ ;
	wire _w17069_ ;
	wire _w17070_ ;
	wire _w17071_ ;
	wire _w17072_ ;
	wire _w17073_ ;
	wire _w17074_ ;
	wire _w17075_ ;
	wire _w17076_ ;
	wire _w17077_ ;
	wire _w17078_ ;
	wire _w17079_ ;
	wire _w17080_ ;
	wire _w17081_ ;
	wire _w17082_ ;
	wire _w17083_ ;
	wire _w17084_ ;
	wire _w17085_ ;
	wire _w17086_ ;
	wire _w17087_ ;
	wire _w17088_ ;
	wire _w17089_ ;
	wire _w17090_ ;
	wire _w17091_ ;
	wire _w17092_ ;
	wire _w17093_ ;
	wire _w17094_ ;
	wire _w17095_ ;
	wire _w17096_ ;
	wire _w17097_ ;
	wire _w17098_ ;
	wire _w17099_ ;
	wire _w17100_ ;
	wire _w17101_ ;
	wire _w17102_ ;
	wire _w17103_ ;
	wire _w17104_ ;
	wire _w17105_ ;
	wire _w17106_ ;
	wire _w17107_ ;
	wire _w17108_ ;
	wire _w17109_ ;
	wire _w17110_ ;
	wire _w17111_ ;
	wire _w17112_ ;
	wire _w17113_ ;
	wire _w17114_ ;
	wire _w17115_ ;
	wire _w17116_ ;
	wire _w17117_ ;
	wire _w17118_ ;
	wire _w17119_ ;
	wire _w17120_ ;
	wire _w17121_ ;
	wire _w17122_ ;
	wire _w17123_ ;
	wire _w17124_ ;
	wire _w17125_ ;
	wire _w17126_ ;
	wire _w17127_ ;
	wire _w17128_ ;
	wire _w17129_ ;
	wire _w17130_ ;
	wire _w17131_ ;
	wire _w17132_ ;
	wire _w17133_ ;
	wire _w17134_ ;
	wire _w17135_ ;
	wire _w17136_ ;
	wire _w17137_ ;
	wire _w17138_ ;
	wire _w17139_ ;
	wire _w17140_ ;
	wire _w17141_ ;
	wire _w17142_ ;
	wire _w17143_ ;
	wire _w17144_ ;
	wire _w17145_ ;
	wire _w17146_ ;
	wire _w17147_ ;
	wire _w17148_ ;
	wire _w17149_ ;
	wire _w17150_ ;
	wire _w17151_ ;
	wire _w17152_ ;
	wire _w17153_ ;
	wire _w17154_ ;
	wire _w17155_ ;
	wire _w17156_ ;
	wire _w17157_ ;
	wire _w17158_ ;
	wire _w17159_ ;
	wire _w17160_ ;
	wire _w17161_ ;
	wire _w17162_ ;
	wire _w17163_ ;
	wire _w17164_ ;
	wire _w17165_ ;
	wire _w17166_ ;
	wire _w17167_ ;
	wire _w17168_ ;
	wire _w17169_ ;
	wire _w17170_ ;
	wire _w17171_ ;
	wire _w17172_ ;
	wire _w17173_ ;
	wire _w17174_ ;
	wire _w17175_ ;
	wire _w17176_ ;
	wire _w17177_ ;
	wire _w17178_ ;
	wire _w17179_ ;
	wire _w17180_ ;
	wire _w17181_ ;
	wire _w17182_ ;
	wire _w17183_ ;
	wire _w17184_ ;
	wire _w17185_ ;
	wire _w17186_ ;
	wire _w17187_ ;
	wire _w17188_ ;
	wire _w17189_ ;
	wire _w17190_ ;
	wire _w17191_ ;
	wire _w17192_ ;
	wire _w17193_ ;
	wire _w17194_ ;
	wire _w17195_ ;
	wire _w17196_ ;
	wire _w17197_ ;
	wire _w17198_ ;
	wire _w17199_ ;
	wire _w17200_ ;
	wire _w17201_ ;
	wire _w17202_ ;
	wire _w17203_ ;
	wire _w17204_ ;
	wire _w17205_ ;
	wire _w17206_ ;
	wire _w17207_ ;
	wire _w17208_ ;
	wire _w17209_ ;
	wire _w17210_ ;
	wire _w17211_ ;
	wire _w17212_ ;
	wire _w17213_ ;
	wire _w17214_ ;
	wire _w17215_ ;
	wire _w17216_ ;
	wire _w17217_ ;
	wire _w17218_ ;
	wire _w17219_ ;
	wire _w17220_ ;
	wire _w17221_ ;
	wire _w17222_ ;
	wire _w17223_ ;
	wire _w17224_ ;
	wire _w17225_ ;
	wire _w17226_ ;
	wire _w17227_ ;
	wire _w17228_ ;
	wire _w17229_ ;
	wire _w17230_ ;
	wire _w17231_ ;
	wire _w17232_ ;
	wire _w17233_ ;
	wire _w17234_ ;
	wire _w17235_ ;
	wire _w17236_ ;
	wire _w17237_ ;
	wire _w17238_ ;
	wire _w17239_ ;
	wire _w17240_ ;
	wire _w17241_ ;
	wire _w17242_ ;
	wire _w17243_ ;
	wire _w17244_ ;
	wire _w17245_ ;
	wire _w17246_ ;
	wire _w17247_ ;
	wire _w17248_ ;
	wire _w17249_ ;
	wire _w17250_ ;
	wire _w17251_ ;
	wire _w17252_ ;
	wire _w17253_ ;
	wire _w17254_ ;
	wire _w17255_ ;
	wire _w17256_ ;
	wire _w17257_ ;
	wire _w17258_ ;
	wire _w17259_ ;
	wire _w17260_ ;
	wire _w17261_ ;
	wire _w17262_ ;
	wire _w17263_ ;
	wire _w17264_ ;
	wire _w17265_ ;
	wire _w17266_ ;
	wire _w17267_ ;
	wire _w17268_ ;
	wire _w17269_ ;
	wire _w17270_ ;
	wire _w17271_ ;
	wire _w17272_ ;
	wire _w17273_ ;
	wire _w17274_ ;
	wire _w17275_ ;
	wire _w17276_ ;
	wire _w17277_ ;
	wire _w17278_ ;
	wire _w17279_ ;
	wire _w17280_ ;
	wire _w17281_ ;
	wire _w17282_ ;
	wire _w17283_ ;
	wire _w17284_ ;
	wire _w17285_ ;
	wire _w17286_ ;
	wire _w17287_ ;
	wire _w17288_ ;
	wire _w17289_ ;
	wire _w17290_ ;
	wire _w17291_ ;
	wire _w17292_ ;
	wire _w17293_ ;
	wire _w17294_ ;
	wire _w17295_ ;
	wire _w17296_ ;
	wire _w17297_ ;
	wire _w17298_ ;
	wire _w17299_ ;
	wire _w17300_ ;
	wire _w17301_ ;
	wire _w17302_ ;
	wire _w17303_ ;
	wire _w17304_ ;
	wire _w17305_ ;
	wire _w17306_ ;
	wire _w17307_ ;
	wire _w17308_ ;
	wire _w17309_ ;
	wire _w17310_ ;
	wire _w17311_ ;
	wire _w17312_ ;
	wire _w17313_ ;
	wire _w17314_ ;
	wire _w17315_ ;
	wire _w17316_ ;
	wire _w17317_ ;
	wire _w17318_ ;
	wire _w17319_ ;
	wire _w17320_ ;
	wire _w17321_ ;
	wire _w17322_ ;
	wire _w17323_ ;
	wire _w17324_ ;
	wire _w17325_ ;
	wire _w17326_ ;
	wire _w17327_ ;
	wire _w17328_ ;
	wire _w17329_ ;
	wire _w17330_ ;
	wire _w17331_ ;
	wire _w17332_ ;
	wire _w17333_ ;
	wire _w17334_ ;
	wire _w17335_ ;
	wire _w17336_ ;
	wire _w17337_ ;
	wire _w17338_ ;
	wire _w17339_ ;
	wire _w17340_ ;
	wire _w17341_ ;
	wire _w17342_ ;
	wire _w17343_ ;
	wire _w17344_ ;
	wire _w17345_ ;
	wire _w17346_ ;
	wire _w17347_ ;
	wire _w17348_ ;
	wire _w17349_ ;
	wire _w17350_ ;
	wire _w17351_ ;
	wire _w17352_ ;
	wire _w17353_ ;
	wire _w17354_ ;
	wire _w17355_ ;
	wire _w17356_ ;
	wire _w17357_ ;
	wire _w17358_ ;
	wire _w17359_ ;
	wire _w17360_ ;
	wire _w17361_ ;
	wire _w17362_ ;
	wire _w17363_ ;
	wire _w17364_ ;
	wire _w17365_ ;
	wire _w17366_ ;
	wire _w17367_ ;
	wire _w17368_ ;
	wire _w17369_ ;
	wire _w17370_ ;
	wire _w17371_ ;
	wire _w17372_ ;
	wire _w17373_ ;
	wire _w17374_ ;
	wire _w17375_ ;
	wire _w17376_ ;
	wire _w17377_ ;
	wire _w17378_ ;
	wire _w17379_ ;
	wire _w17380_ ;
	wire _w17381_ ;
	wire _w17382_ ;
	wire _w17383_ ;
	wire _w17384_ ;
	wire _w17385_ ;
	wire _w17386_ ;
	wire _w17387_ ;
	wire _w17388_ ;
	wire _w17389_ ;
	wire _w17390_ ;
	wire _w17391_ ;
	wire _w17392_ ;
	wire _w17393_ ;
	wire _w17394_ ;
	wire _w17395_ ;
	wire _w17396_ ;
	wire _w17397_ ;
	wire _w17398_ ;
	wire _w17399_ ;
	wire _w17400_ ;
	wire _w17401_ ;
	wire _w17402_ ;
	wire _w17403_ ;
	wire _w17404_ ;
	wire _w17405_ ;
	wire _w17406_ ;
	wire _w17407_ ;
	wire _w17408_ ;
	wire _w17409_ ;
	wire _w17410_ ;
	wire _w17411_ ;
	wire _w17412_ ;
	wire _w17413_ ;
	wire _w17414_ ;
	wire _w17415_ ;
	wire _w17416_ ;
	wire _w17417_ ;
	wire _w17418_ ;
	wire _w17419_ ;
	wire _w17420_ ;
	wire _w17421_ ;
	wire _w17422_ ;
	wire _w17423_ ;
	wire _w17424_ ;
	wire _w17425_ ;
	wire _w17426_ ;
	wire _w17427_ ;
	wire _w17428_ ;
	wire _w17429_ ;
	wire _w17430_ ;
	wire _w17431_ ;
	wire _w17432_ ;
	wire _w17433_ ;
	wire _w17434_ ;
	wire _w17435_ ;
	wire _w17436_ ;
	wire _w17437_ ;
	wire _w17438_ ;
	wire _w17439_ ;
	wire _w17440_ ;
	wire _w17441_ ;
	wire _w17442_ ;
	wire _w17443_ ;
	wire _w17444_ ;
	wire _w17445_ ;
	wire _w17446_ ;
	wire _w17447_ ;
	wire _w17448_ ;
	wire _w17449_ ;
	wire _w17450_ ;
	wire _w17451_ ;
	wire _w17452_ ;
	wire _w17453_ ;
	wire _w17454_ ;
	wire _w17455_ ;
	wire _w17456_ ;
	wire _w17457_ ;
	wire _w17458_ ;
	wire _w17459_ ;
	wire _w17460_ ;
	wire _w17461_ ;
	wire _w17462_ ;
	wire _w17463_ ;
	wire _w17464_ ;
	wire _w17465_ ;
	wire _w17466_ ;
	wire _w17467_ ;
	wire _w17468_ ;
	wire _w17469_ ;
	wire _w17470_ ;
	wire _w17471_ ;
	wire _w17472_ ;
	wire _w17473_ ;
	wire _w17474_ ;
	wire _w17475_ ;
	wire _w17476_ ;
	wire _w17477_ ;
	wire _w17478_ ;
	wire _w17479_ ;
	wire _w17480_ ;
	wire _w17481_ ;
	wire _w17482_ ;
	wire _w17483_ ;
	wire _w17484_ ;
	wire _w17485_ ;
	wire _w17486_ ;
	wire _w17487_ ;
	wire _w17488_ ;
	wire _w17489_ ;
	wire _w17490_ ;
	wire _w17491_ ;
	wire _w17492_ ;
	wire _w17493_ ;
	wire _w17494_ ;
	wire _w17495_ ;
	wire _w17496_ ;
	wire _w17497_ ;
	wire _w17498_ ;
	wire _w17499_ ;
	wire _w17500_ ;
	wire _w17501_ ;
	wire _w17502_ ;
	wire _w17503_ ;
	wire _w17504_ ;
	wire _w17505_ ;
	wire _w17506_ ;
	wire _w17507_ ;
	wire _w17508_ ;
	wire _w17509_ ;
	wire _w17510_ ;
	wire _w17511_ ;
	wire _w17512_ ;
	wire _w17513_ ;
	wire _w17514_ ;
	wire _w17515_ ;
	wire _w17516_ ;
	wire _w17517_ ;
	wire _w17518_ ;
	wire _w17519_ ;
	wire _w17520_ ;
	wire _w17521_ ;
	wire _w17522_ ;
	wire _w17523_ ;
	wire _w17524_ ;
	wire _w17525_ ;
	wire _w17526_ ;
	wire _w17527_ ;
	wire _w17528_ ;
	wire _w17529_ ;
	wire _w17530_ ;
	wire _w17531_ ;
	wire _w17532_ ;
	wire _w17533_ ;
	wire _w17534_ ;
	wire _w17535_ ;
	wire _w17536_ ;
	wire _w17537_ ;
	wire _w17538_ ;
	wire _w17539_ ;
	wire _w17540_ ;
	wire _w17541_ ;
	wire _w17542_ ;
	wire _w17543_ ;
	wire _w17544_ ;
	wire _w17545_ ;
	wire _w17546_ ;
	wire _w17547_ ;
	wire _w17548_ ;
	wire _w17549_ ;
	wire _w17550_ ;
	wire _w17551_ ;
	wire _w17552_ ;
	wire _w17553_ ;
	wire _w17554_ ;
	wire _w17555_ ;
	wire _w17556_ ;
	wire _w17557_ ;
	wire _w17558_ ;
	wire _w17559_ ;
	wire _w17560_ ;
	wire _w17561_ ;
	wire _w17562_ ;
	wire _w17563_ ;
	wire _w17564_ ;
	wire _w17565_ ;
	wire _w17566_ ;
	wire _w17567_ ;
	wire _w17568_ ;
	wire _w17569_ ;
	wire _w17570_ ;
	wire _w17571_ ;
	wire _w17572_ ;
	wire _w17573_ ;
	wire _w17574_ ;
	wire _w17575_ ;
	wire _w17576_ ;
	wire _w17577_ ;
	wire _w17578_ ;
	wire _w17579_ ;
	wire _w17580_ ;
	wire _w17581_ ;
	wire _w17582_ ;
	wire _w17583_ ;
	wire _w17584_ ;
	wire _w17585_ ;
	wire _w17586_ ;
	wire _w17587_ ;
	wire _w17588_ ;
	wire _w17589_ ;
	wire _w17590_ ;
	wire _w17591_ ;
	wire _w17592_ ;
	wire _w17593_ ;
	wire _w17594_ ;
	wire _w17595_ ;
	wire _w17596_ ;
	wire _w17597_ ;
	wire _w17598_ ;
	wire _w17599_ ;
	wire _w17600_ ;
	wire _w17601_ ;
	wire _w17602_ ;
	wire _w17603_ ;
	wire _w17604_ ;
	wire _w17605_ ;
	wire _w17606_ ;
	wire _w17607_ ;
	wire _w17608_ ;
	wire _w17609_ ;
	wire _w17610_ ;
	wire _w17611_ ;
	wire _w17612_ ;
	wire _w17613_ ;
	wire _w17614_ ;
	wire _w17615_ ;
	wire _w17616_ ;
	wire _w17617_ ;
	wire _w17618_ ;
	wire _w17619_ ;
	wire _w17620_ ;
	wire _w17621_ ;
	wire _w17622_ ;
	wire _w17623_ ;
	wire _w17624_ ;
	wire _w17625_ ;
	wire _w17626_ ;
	wire _w17627_ ;
	wire _w17628_ ;
	wire _w17629_ ;
	wire _w17630_ ;
	wire _w17631_ ;
	wire _w17632_ ;
	wire _w17633_ ;
	wire _w17634_ ;
	wire _w17635_ ;
	wire _w17636_ ;
	wire _w17637_ ;
	wire _w17638_ ;
	wire _w17639_ ;
	wire _w17640_ ;
	wire _w17641_ ;
	wire _w17642_ ;
	wire _w17643_ ;
	wire _w17644_ ;
	wire _w17645_ ;
	wire _w17646_ ;
	wire _w17647_ ;
	wire _w17648_ ;
	wire _w17649_ ;
	wire _w17650_ ;
	wire _w17651_ ;
	wire _w17652_ ;
	wire _w17653_ ;
	wire _w17654_ ;
	wire _w17655_ ;
	wire _w17656_ ;
	wire _w17657_ ;
	wire _w17658_ ;
	wire _w17659_ ;
	wire _w17660_ ;
	wire _w17661_ ;
	wire _w17662_ ;
	wire _w17663_ ;
	wire _w17664_ ;
	wire _w17665_ ;
	wire _w17666_ ;
	wire _w17667_ ;
	wire _w17668_ ;
	wire _w17669_ ;
	wire _w17670_ ;
	wire _w17671_ ;
	wire _w17672_ ;
	wire _w17673_ ;
	wire _w17674_ ;
	wire _w17675_ ;
	wire _w17676_ ;
	wire _w17677_ ;
	wire _w17678_ ;
	wire _w17679_ ;
	wire _w17680_ ;
	wire _w17681_ ;
	wire _w17682_ ;
	wire _w17683_ ;
	wire _w17684_ ;
	wire _w17685_ ;
	wire _w17686_ ;
	wire _w17687_ ;
	wire _w17688_ ;
	wire _w17689_ ;
	wire _w17690_ ;
	wire _w17691_ ;
	wire _w17692_ ;
	wire _w17693_ ;
	wire _w17694_ ;
	wire _w17695_ ;
	wire _w17696_ ;
	wire _w17697_ ;
	wire _w17698_ ;
	wire _w17699_ ;
	wire _w17700_ ;
	wire _w17701_ ;
	wire _w17702_ ;
	wire _w17703_ ;
	wire _w17704_ ;
	wire _w17705_ ;
	wire _w17706_ ;
	wire _w17707_ ;
	wire _w17708_ ;
	wire _w17709_ ;
	wire _w17710_ ;
	wire _w17711_ ;
	wire _w17712_ ;
	wire _w17713_ ;
	wire _w17714_ ;
	wire _w17715_ ;
	wire _w17716_ ;
	wire _w17717_ ;
	wire _w17718_ ;
	wire _w17719_ ;
	wire _w17720_ ;
	wire _w17721_ ;
	wire _w17722_ ;
	wire _w17723_ ;
	wire _w17724_ ;
	wire _w17725_ ;
	wire _w17726_ ;
	wire _w17727_ ;
	wire _w17728_ ;
	wire _w17729_ ;
	wire _w17730_ ;
	wire _w17731_ ;
	wire _w17732_ ;
	wire _w17733_ ;
	wire _w17734_ ;
	wire _w17735_ ;
	wire _w17736_ ;
	wire _w17737_ ;
	wire _w17738_ ;
	wire _w17739_ ;
	wire _w17740_ ;
	wire _w17741_ ;
	wire _w17742_ ;
	wire _w17743_ ;
	wire _w17744_ ;
	wire _w17745_ ;
	wire _w17746_ ;
	wire _w17747_ ;
	wire _w17748_ ;
	wire _w17749_ ;
	wire _w17750_ ;
	wire _w17751_ ;
	wire _w17752_ ;
	wire _w17753_ ;
	wire _w17754_ ;
	wire _w17755_ ;
	wire _w17756_ ;
	wire _w17757_ ;
	wire _w17758_ ;
	wire _w17759_ ;
	wire _w17760_ ;
	wire _w17761_ ;
	wire _w17762_ ;
	wire _w17763_ ;
	wire _w17764_ ;
	wire _w17765_ ;
	wire _w17766_ ;
	wire _w17767_ ;
	wire _w17768_ ;
	wire _w17769_ ;
	wire _w17770_ ;
	wire _w17771_ ;
	wire _w17772_ ;
	wire _w17773_ ;
	wire _w17774_ ;
	wire _w17775_ ;
	wire _w17776_ ;
	wire _w17777_ ;
	wire _w17778_ ;
	wire _w17779_ ;
	wire _w17780_ ;
	wire _w17781_ ;
	wire _w17782_ ;
	wire _w17783_ ;
	wire _w17784_ ;
	wire _w17785_ ;
	wire _w17786_ ;
	wire _w17787_ ;
	wire _w17788_ ;
	wire _w17789_ ;
	wire _w17790_ ;
	wire _w17791_ ;
	wire _w17792_ ;
	wire _w17793_ ;
	wire _w17794_ ;
	wire _w17795_ ;
	wire _w17796_ ;
	wire _w17797_ ;
	wire _w17798_ ;
	wire _w17799_ ;
	wire _w17800_ ;
	wire _w17801_ ;
	wire _w17802_ ;
	wire _w17803_ ;
	wire _w17804_ ;
	wire _w17805_ ;
	wire _w17806_ ;
	wire _w17807_ ;
	wire _w17808_ ;
	wire _w17809_ ;
	wire _w17810_ ;
	wire _w17811_ ;
	wire _w17812_ ;
	wire _w17813_ ;
	wire _w17814_ ;
	wire _w17815_ ;
	wire _w17816_ ;
	wire _w17817_ ;
	wire _w17818_ ;
	wire _w17819_ ;
	wire _w17820_ ;
	wire _w17821_ ;
	wire _w17822_ ;
	wire _w17823_ ;
	wire _w17824_ ;
	wire _w17825_ ;
	wire _w17826_ ;
	wire _w17827_ ;
	wire _w17828_ ;
	wire _w17829_ ;
	wire _w17830_ ;
	wire _w17831_ ;
	wire _w17832_ ;
	wire _w17833_ ;
	wire _w17834_ ;
	wire _w17835_ ;
	wire _w17836_ ;
	wire _w17837_ ;
	wire _w17838_ ;
	wire _w17839_ ;
	wire _w17840_ ;
	wire _w17841_ ;
	wire _w17842_ ;
	wire _w17843_ ;
	wire _w17844_ ;
	wire _w17845_ ;
	wire _w17846_ ;
	wire _w17847_ ;
	wire _w17848_ ;
	wire _w17849_ ;
	wire _w17850_ ;
	wire _w17851_ ;
	wire _w17852_ ;
	wire _w17853_ ;
	wire _w17854_ ;
	wire _w17855_ ;
	wire _w17856_ ;
	wire _w17857_ ;
	wire _w17858_ ;
	wire _w17859_ ;
	wire _w17860_ ;
	wire _w17861_ ;
	wire _w17862_ ;
	wire _w17863_ ;
	wire _w17864_ ;
	wire _w17865_ ;
	wire _w17866_ ;
	wire _w17867_ ;
	wire _w17868_ ;
	wire _w17869_ ;
	wire _w17870_ ;
	wire _w17871_ ;
	wire _w17872_ ;
	wire _w17873_ ;
	wire _w17874_ ;
	wire _w17875_ ;
	wire _w17876_ ;
	wire _w17877_ ;
	wire _w17878_ ;
	wire _w17879_ ;
	wire _w17880_ ;
	wire _w17881_ ;
	wire _w17882_ ;
	wire _w17883_ ;
	wire _w17884_ ;
	wire _w17885_ ;
	wire _w17886_ ;
	wire _w17887_ ;
	wire _w17888_ ;
	wire _w17889_ ;
	wire _w17890_ ;
	wire _w17891_ ;
	wire _w17892_ ;
	wire _w17893_ ;
	wire _w17894_ ;
	wire _w17895_ ;
	wire _w17896_ ;
	wire _w17897_ ;
	wire _w17898_ ;
	wire _w17899_ ;
	wire _w17900_ ;
	wire _w17901_ ;
	wire _w17902_ ;
	wire _w17903_ ;
	wire _w17904_ ;
	wire _w17905_ ;
	wire _w17906_ ;
	wire _w17907_ ;
	wire _w17908_ ;
	wire _w17909_ ;
	wire _w17910_ ;
	wire _w17911_ ;
	wire _w17912_ ;
	wire _w17913_ ;
	wire _w17914_ ;
	wire _w17915_ ;
	wire _w17916_ ;
	wire _w17917_ ;
	wire _w17918_ ;
	wire _w17919_ ;
	wire _w17920_ ;
	wire _w17921_ ;
	wire _w17922_ ;
	wire _w17923_ ;
	wire _w17924_ ;
	wire _w17925_ ;
	wire _w17926_ ;
	wire _w17927_ ;
	wire _w17928_ ;
	wire _w17929_ ;
	wire _w17930_ ;
	wire _w17931_ ;
	wire _w17932_ ;
	wire _w17933_ ;
	wire _w17934_ ;
	wire _w17935_ ;
	wire _w17936_ ;
	wire _w17937_ ;
	wire _w17938_ ;
	wire _w17939_ ;
	wire _w17940_ ;
	wire _w17941_ ;
	wire _w17942_ ;
	wire _w17943_ ;
	wire _w17944_ ;
	wire _w17945_ ;
	wire _w17946_ ;
	wire _w17947_ ;
	wire _w17948_ ;
	wire _w17949_ ;
	wire _w17950_ ;
	wire _w17951_ ;
	wire _w17952_ ;
	wire _w17953_ ;
	wire _w17954_ ;
	wire _w17955_ ;
	wire _w17956_ ;
	wire _w17957_ ;
	wire _w17958_ ;
	wire _w17959_ ;
	wire _w17960_ ;
	wire _w17961_ ;
	wire _w17962_ ;
	wire _w17963_ ;
	wire _w17964_ ;
	wire _w17965_ ;
	wire _w17966_ ;
	wire _w17967_ ;
	wire _w17968_ ;
	wire _w17969_ ;
	wire _w17970_ ;
	wire _w17971_ ;
	wire _w17972_ ;
	wire _w17973_ ;
	wire _w17974_ ;
	wire _w17975_ ;
	wire _w17976_ ;
	wire _w17977_ ;
	wire _w17978_ ;
	wire _w17979_ ;
	wire _w17980_ ;
	wire _w17981_ ;
	wire _w17982_ ;
	wire _w17983_ ;
	wire _w17984_ ;
	wire _w17985_ ;
	wire _w17986_ ;
	wire _w17987_ ;
	wire _w17988_ ;
	wire _w17989_ ;
	wire _w17990_ ;
	wire _w17991_ ;
	wire _w17992_ ;
	wire _w17993_ ;
	wire _w17994_ ;
	wire _w17995_ ;
	wire _w17996_ ;
	wire _w17997_ ;
	wire _w17998_ ;
	wire _w17999_ ;
	wire _w18000_ ;
	wire _w18001_ ;
	wire _w18002_ ;
	wire _w18003_ ;
	wire _w18004_ ;
	wire _w18005_ ;
	wire _w18006_ ;
	wire _w18007_ ;
	wire _w18008_ ;
	wire _w18009_ ;
	wire _w18010_ ;
	wire _w18011_ ;
	wire _w18012_ ;
	wire _w18013_ ;
	wire _w18014_ ;
	wire _w18015_ ;
	wire _w18016_ ;
	wire _w18017_ ;
	wire _w18018_ ;
	wire _w18019_ ;
	wire _w18020_ ;
	wire _w18021_ ;
	wire _w18022_ ;
	wire _w18023_ ;
	wire _w18024_ ;
	wire _w18025_ ;
	wire _w18026_ ;
	wire _w18027_ ;
	wire _w18028_ ;
	wire _w18029_ ;
	wire _w18030_ ;
	wire _w18031_ ;
	wire _w18032_ ;
	wire _w18033_ ;
	wire _w18034_ ;
	wire _w18035_ ;
	wire _w18036_ ;
	wire _w18037_ ;
	wire _w18038_ ;
	wire _w18039_ ;
	wire _w18040_ ;
	wire _w18041_ ;
	wire _w18042_ ;
	wire _w18043_ ;
	wire _w18044_ ;
	wire _w18045_ ;
	wire _w18046_ ;
	wire _w18047_ ;
	wire _w18048_ ;
	wire _w18049_ ;
	wire _w18050_ ;
	wire _w18051_ ;
	wire _w18052_ ;
	wire _w18053_ ;
	wire _w18054_ ;
	wire _w18055_ ;
	wire _w18056_ ;
	wire _w18057_ ;
	wire _w18058_ ;
	wire _w18059_ ;
	wire _w18060_ ;
	wire _w18061_ ;
	wire _w18062_ ;
	wire _w18063_ ;
	wire _w18064_ ;
	wire _w18065_ ;
	wire _w18066_ ;
	wire _w18067_ ;
	wire _w18068_ ;
	wire _w18069_ ;
	wire _w18070_ ;
	wire _w18071_ ;
	wire _w18072_ ;
	wire _w18073_ ;
	wire _w18074_ ;
	wire _w18075_ ;
	wire _w18076_ ;
	wire _w18077_ ;
	wire _w18078_ ;
	wire _w18079_ ;
	wire _w18080_ ;
	wire _w18081_ ;
	wire _w18082_ ;
	wire _w18083_ ;
	wire _w18084_ ;
	wire _w18085_ ;
	wire _w18086_ ;
	wire _w18087_ ;
	wire _w18088_ ;
	wire _w18089_ ;
	wire _w18090_ ;
	wire _w18091_ ;
	wire _w18092_ ;
	wire _w18093_ ;
	wire _w18094_ ;
	wire _w18095_ ;
	wire _w18096_ ;
	wire _w18097_ ;
	wire _w18098_ ;
	wire _w18099_ ;
	wire _w18100_ ;
	wire _w18101_ ;
	wire _w18102_ ;
	wire _w18103_ ;
	wire _w18104_ ;
	wire _w18105_ ;
	wire _w18106_ ;
	wire _w18107_ ;
	wire _w18108_ ;
	wire _w18109_ ;
	wire _w18110_ ;
	wire _w18111_ ;
	wire _w18112_ ;
	wire _w18113_ ;
	wire _w18114_ ;
	wire _w18115_ ;
	wire _w18116_ ;
	wire _w18117_ ;
	wire _w18118_ ;
	wire _w18119_ ;
	wire _w18120_ ;
	wire _w18121_ ;
	wire _w18122_ ;
	wire _w18123_ ;
	wire _w18124_ ;
	wire _w18125_ ;
	wire _w18126_ ;
	wire _w18127_ ;
	wire _w18128_ ;
	wire _w18129_ ;
	wire _w18130_ ;
	wire _w18131_ ;
	wire _w18132_ ;
	wire _w18133_ ;
	wire _w18134_ ;
	wire _w18135_ ;
	wire _w18136_ ;
	wire _w18137_ ;
	wire _w18138_ ;
	wire _w18139_ ;
	wire _w18140_ ;
	wire _w18141_ ;
	wire _w18142_ ;
	wire _w18143_ ;
	wire _w18144_ ;
	wire _w18145_ ;
	wire _w18146_ ;
	wire _w18147_ ;
	wire _w18148_ ;
	wire _w18149_ ;
	wire _w18150_ ;
	wire _w18151_ ;
	wire _w18152_ ;
	wire _w18153_ ;
	wire _w18154_ ;
	wire _w18155_ ;
	wire _w18156_ ;
	wire _w18157_ ;
	wire _w18158_ ;
	wire _w18159_ ;
	wire _w18160_ ;
	wire _w18161_ ;
	wire _w18162_ ;
	wire _w18163_ ;
	wire _w18164_ ;
	wire _w18165_ ;
	wire _w18166_ ;
	wire _w18167_ ;
	wire _w18168_ ;
	wire _w18169_ ;
	wire _w18170_ ;
	wire _w18171_ ;
	wire _w18172_ ;
	wire _w18173_ ;
	wire _w18174_ ;
	wire _w18175_ ;
	wire _w18176_ ;
	wire _w18177_ ;
	wire _w18178_ ;
	wire _w18179_ ;
	wire _w18180_ ;
	wire _w18181_ ;
	wire _w18182_ ;
	wire _w18183_ ;
	wire _w18184_ ;
	wire _w18185_ ;
	wire _w18186_ ;
	wire _w18187_ ;
	wire _w18188_ ;
	wire _w18189_ ;
	wire _w18190_ ;
	wire _w18191_ ;
	wire _w18192_ ;
	wire _w18193_ ;
	wire _w18194_ ;
	wire _w18195_ ;
	wire _w18196_ ;
	wire _w18197_ ;
	wire _w18198_ ;
	wire _w18199_ ;
	wire _w18200_ ;
	wire _w18201_ ;
	wire _w18202_ ;
	wire _w18203_ ;
	wire _w18204_ ;
	wire _w18205_ ;
	wire _w18206_ ;
	wire _w18207_ ;
	wire _w18208_ ;
	wire _w18209_ ;
	wire _w18210_ ;
	wire _w18211_ ;
	wire _w18212_ ;
	wire _w18213_ ;
	wire _w18214_ ;
	wire _w18215_ ;
	wire _w18216_ ;
	wire _w18217_ ;
	wire _w18218_ ;
	wire _w18219_ ;
	wire _w18220_ ;
	wire _w18221_ ;
	wire _w18222_ ;
	wire _w18223_ ;
	wire _w18224_ ;
	wire _w18225_ ;
	wire _w18226_ ;
	wire _w18227_ ;
	wire _w18228_ ;
	wire _w18229_ ;
	wire _w18230_ ;
	wire _w18231_ ;
	wire _w18232_ ;
	wire _w18233_ ;
	wire _w18234_ ;
	wire _w18235_ ;
	wire _w18236_ ;
	wire _w18237_ ;
	wire _w18238_ ;
	wire _w18239_ ;
	wire _w18240_ ;
	wire _w18241_ ;
	wire _w18242_ ;
	wire _w18243_ ;
	wire _w18244_ ;
	wire _w18245_ ;
	wire _w18246_ ;
	wire _w18247_ ;
	wire _w18248_ ;
	wire _w18249_ ;
	wire _w18250_ ;
	wire _w18251_ ;
	wire _w18252_ ;
	wire _w18253_ ;
	wire _w18254_ ;
	wire _w18255_ ;
	wire _w18256_ ;
	wire _w18257_ ;
	wire _w18258_ ;
	wire _w18259_ ;
	wire _w18260_ ;
	wire _w18261_ ;
	wire _w18262_ ;
	wire _w18263_ ;
	wire _w18264_ ;
	wire _w18265_ ;
	wire _w18266_ ;
	wire _w18267_ ;
	wire _w18268_ ;
	wire _w18269_ ;
	wire _w18270_ ;
	wire _w18271_ ;
	wire _w18272_ ;
	wire _w18273_ ;
	wire _w18274_ ;
	wire _w18275_ ;
	wire _w18276_ ;
	wire _w18277_ ;
	wire _w18278_ ;
	wire _w18279_ ;
	wire _w18280_ ;
	wire _w18281_ ;
	wire _w18282_ ;
	wire _w18283_ ;
	wire _w18284_ ;
	wire _w18285_ ;
	wire _w18286_ ;
	wire _w18287_ ;
	wire _w18288_ ;
	wire _w18289_ ;
	wire _w18290_ ;
	wire _w18291_ ;
	wire _w18292_ ;
	wire _w18293_ ;
	wire _w18294_ ;
	wire _w18295_ ;
	wire _w18296_ ;
	wire _w18297_ ;
	wire _w18298_ ;
	wire _w18299_ ;
	wire _w18300_ ;
	wire _w18301_ ;
	wire _w18302_ ;
	wire _w18303_ ;
	wire _w18304_ ;
	wire _w18305_ ;
	wire _w18306_ ;
	wire _w18307_ ;
	wire _w18308_ ;
	wire _w18309_ ;
	wire _w18310_ ;
	wire _w18311_ ;
	wire _w18312_ ;
	wire _w18313_ ;
	wire _w18314_ ;
	wire _w18315_ ;
	wire _w18316_ ;
	wire _w18317_ ;
	wire _w18318_ ;
	wire _w18319_ ;
	wire _w18320_ ;
	wire _w18321_ ;
	wire _w18322_ ;
	wire _w18323_ ;
	wire _w18324_ ;
	wire _w18325_ ;
	wire _w18326_ ;
	wire _w18327_ ;
	wire _w18328_ ;
	wire _w18329_ ;
	wire _w18330_ ;
	wire _w18331_ ;
	wire _w18332_ ;
	wire _w18333_ ;
	wire _w18334_ ;
	wire _w18335_ ;
	wire _w18336_ ;
	wire _w18337_ ;
	wire _w18338_ ;
	wire _w18339_ ;
	wire _w18340_ ;
	wire _w18341_ ;
	wire _w18342_ ;
	wire _w18343_ ;
	wire _w18344_ ;
	wire _w18345_ ;
	wire _w18346_ ;
	wire _w18347_ ;
	wire _w18348_ ;
	wire _w18349_ ;
	wire _w18350_ ;
	wire _w18351_ ;
	wire _w18352_ ;
	wire _w18353_ ;
	wire _w18354_ ;
	wire _w18355_ ;
	wire _w18356_ ;
	wire _w18357_ ;
	wire _w18358_ ;
	wire _w18359_ ;
	wire _w18360_ ;
	wire _w18361_ ;
	wire _w18362_ ;
	wire _w18363_ ;
	wire _w18364_ ;
	wire _w18365_ ;
	wire _w18366_ ;
	wire _w18367_ ;
	wire _w18368_ ;
	wire _w18369_ ;
	wire _w18370_ ;
	wire _w18371_ ;
	wire _w18372_ ;
	wire _w18373_ ;
	wire _w18374_ ;
	wire _w18375_ ;
	wire _w18376_ ;
	wire _w18377_ ;
	wire _w18378_ ;
	wire _w18379_ ;
	wire _w18380_ ;
	wire _w18381_ ;
	wire _w18382_ ;
	wire _w18383_ ;
	wire _w18384_ ;
	wire _w18385_ ;
	wire _w18386_ ;
	wire _w18387_ ;
	wire _w18388_ ;
	wire _w18389_ ;
	wire _w18390_ ;
	wire _w18391_ ;
	wire _w18392_ ;
	wire _w18393_ ;
	wire _w18394_ ;
	wire _w18395_ ;
	wire _w18396_ ;
	wire _w18397_ ;
	wire _w18398_ ;
	wire _w18399_ ;
	wire _w18400_ ;
	wire _w18401_ ;
	wire _w18402_ ;
	wire _w18403_ ;
	wire _w18404_ ;
	wire _w18405_ ;
	wire _w18406_ ;
	wire _w18407_ ;
	wire _w18408_ ;
	wire _w18409_ ;
	wire _w18410_ ;
	wire _w18411_ ;
	wire _w18412_ ;
	wire _w18413_ ;
	wire _w18414_ ;
	wire _w18415_ ;
	wire _w18416_ ;
	wire _w18417_ ;
	wire _w18418_ ;
	wire _w18419_ ;
	wire _w18420_ ;
	wire _w18421_ ;
	wire _w18422_ ;
	wire _w18423_ ;
	wire _w18424_ ;
	wire _w18425_ ;
	wire _w18426_ ;
	wire _w18427_ ;
	wire _w18428_ ;
	wire _w18429_ ;
	wire _w18430_ ;
	wire _w18431_ ;
	wire _w18432_ ;
	wire _w18433_ ;
	wire _w18434_ ;
	wire _w18435_ ;
	wire _w18436_ ;
	wire _w18437_ ;
	wire _w18438_ ;
	wire _w18439_ ;
	wire _w18440_ ;
	wire _w18441_ ;
	wire _w18442_ ;
	wire _w18443_ ;
	wire _w18444_ ;
	wire _w18445_ ;
	wire _w18446_ ;
	wire _w18447_ ;
	wire _w18448_ ;
	wire _w18449_ ;
	wire _w18450_ ;
	wire _w18451_ ;
	wire _w18452_ ;
	wire _w18453_ ;
	wire _w18454_ ;
	wire _w18455_ ;
	wire _w18456_ ;
	wire _w18457_ ;
	wire _w18458_ ;
	wire _w18459_ ;
	wire _w18460_ ;
	wire _w18461_ ;
	wire _w18462_ ;
	wire _w18463_ ;
	wire _w18464_ ;
	wire _w18465_ ;
	wire _w18466_ ;
	wire _w18467_ ;
	wire _w18468_ ;
	wire _w18469_ ;
	wire _w18470_ ;
	wire _w18471_ ;
	wire _w18472_ ;
	wire _w18473_ ;
	wire _w18474_ ;
	wire _w18475_ ;
	wire _w18476_ ;
	wire _w18477_ ;
	wire _w18478_ ;
	wire _w18479_ ;
	wire _w18480_ ;
	wire _w18481_ ;
	wire _w18482_ ;
	wire _w18483_ ;
	wire _w18484_ ;
	wire _w18485_ ;
	wire _w18486_ ;
	wire _w18487_ ;
	wire _w18488_ ;
	wire _w18489_ ;
	wire _w18490_ ;
	wire _w18491_ ;
	wire _w18492_ ;
	wire _w18493_ ;
	wire _w18494_ ;
	wire _w18495_ ;
	wire _w18496_ ;
	wire _w18497_ ;
	wire _w18498_ ;
	wire _w18499_ ;
	wire _w18500_ ;
	wire _w18501_ ;
	wire _w18502_ ;
	wire _w18503_ ;
	wire _w18504_ ;
	wire _w18505_ ;
	wire _w18506_ ;
	wire _w18507_ ;
	wire _w18508_ ;
	wire _w18509_ ;
	wire _w18510_ ;
	wire _w18511_ ;
	wire _w18512_ ;
	wire _w18513_ ;
	wire _w18514_ ;
	wire _w18515_ ;
	wire _w18516_ ;
	wire _w18517_ ;
	wire _w18518_ ;
	wire _w18519_ ;
	wire _w18520_ ;
	wire _w18521_ ;
	wire _w18522_ ;
	wire _w18523_ ;
	wire _w18524_ ;
	wire _w18525_ ;
	wire _w18526_ ;
	wire _w18527_ ;
	wire _w18528_ ;
	wire _w18529_ ;
	wire _w18530_ ;
	wire _w18531_ ;
	wire _w18532_ ;
	wire _w18533_ ;
	wire _w18534_ ;
	wire _w18535_ ;
	wire _w18536_ ;
	wire _w18537_ ;
	wire _w18538_ ;
	wire _w18539_ ;
	wire _w18540_ ;
	wire _w18541_ ;
	wire _w18542_ ;
	wire _w18543_ ;
	wire _w18544_ ;
	wire _w18545_ ;
	wire _w18546_ ;
	wire _w18547_ ;
	wire _w18548_ ;
	wire _w18549_ ;
	wire _w18550_ ;
	wire _w18551_ ;
	wire _w18552_ ;
	wire _w18553_ ;
	wire _w18554_ ;
	wire _w18555_ ;
	wire _w18556_ ;
	wire _w18557_ ;
	wire _w18558_ ;
	wire _w18559_ ;
	wire _w18560_ ;
	wire _w18561_ ;
	wire _w18562_ ;
	wire _w18563_ ;
	wire _w18564_ ;
	wire _w18565_ ;
	wire _w18566_ ;
	wire _w18567_ ;
	wire _w18568_ ;
	wire _w18569_ ;
	wire _w18570_ ;
	wire _w18571_ ;
	wire _w18572_ ;
	wire _w18573_ ;
	wire _w18574_ ;
	wire _w18575_ ;
	wire _w18576_ ;
	wire _w18577_ ;
	wire _w18578_ ;
	wire _w18579_ ;
	wire _w18580_ ;
	wire _w18581_ ;
	wire _w18582_ ;
	wire _w18583_ ;
	wire _w18584_ ;
	wire _w18585_ ;
	wire _w18586_ ;
	wire _w18587_ ;
	wire _w18588_ ;
	wire _w18589_ ;
	wire _w18590_ ;
	wire _w18591_ ;
	wire _w18592_ ;
	wire _w18593_ ;
	wire _w18594_ ;
	wire _w18595_ ;
	wire _w18596_ ;
	wire _w18597_ ;
	wire _w18598_ ;
	wire _w18599_ ;
	wire _w18600_ ;
	wire _w18601_ ;
	wire _w18602_ ;
	wire _w18603_ ;
	wire _w18604_ ;
	wire _w18605_ ;
	wire _w18606_ ;
	wire _w18607_ ;
	wire _w18608_ ;
	wire _w18609_ ;
	wire _w18610_ ;
	wire _w18611_ ;
	wire _w18612_ ;
	wire _w18613_ ;
	wire _w18614_ ;
	wire _w18615_ ;
	wire _w18616_ ;
	wire _w18617_ ;
	wire _w18618_ ;
	wire _w18619_ ;
	wire _w18620_ ;
	wire _w18621_ ;
	wire _w18622_ ;
	wire _w18623_ ;
	wire _w18624_ ;
	wire _w18625_ ;
	wire _w18626_ ;
	wire _w18627_ ;
	wire _w18628_ ;
	wire _w18629_ ;
	wire _w18630_ ;
	wire _w18631_ ;
	wire _w18632_ ;
	wire _w18633_ ;
	wire _w18634_ ;
	wire _w18635_ ;
	wire _w18636_ ;
	wire _w18637_ ;
	wire _w18638_ ;
	wire _w18639_ ;
	wire _w18640_ ;
	wire _w18641_ ;
	wire _w18642_ ;
	wire _w18643_ ;
	wire _w18644_ ;
	wire _w18645_ ;
	wire _w18646_ ;
	wire _w18647_ ;
	wire _w18648_ ;
	wire _w18649_ ;
	wire _w18650_ ;
	wire _w18651_ ;
	wire _w18652_ ;
	wire _w18653_ ;
	wire _w18654_ ;
	wire _w18655_ ;
	wire _w18656_ ;
	wire _w18657_ ;
	wire _w18658_ ;
	wire _w18659_ ;
	wire _w18660_ ;
	wire _w18661_ ;
	wire _w18662_ ;
	wire _w18663_ ;
	wire _w18664_ ;
	wire _w18665_ ;
	wire _w18666_ ;
	wire _w18667_ ;
	wire _w18668_ ;
	wire _w18669_ ;
	wire _w18670_ ;
	wire _w18671_ ;
	wire _w18672_ ;
	wire _w18673_ ;
	wire _w18674_ ;
	wire _w18675_ ;
	wire _w18676_ ;
	wire _w18677_ ;
	wire _w18678_ ;
	wire _w18679_ ;
	wire _w18680_ ;
	wire _w18681_ ;
	wire _w18682_ ;
	wire _w18683_ ;
	wire _w18684_ ;
	wire _w18685_ ;
	wire _w18686_ ;
	wire _w18687_ ;
	wire _w18688_ ;
	wire _w18689_ ;
	wire _w18690_ ;
	wire _w18691_ ;
	wire _w18692_ ;
	wire _w18693_ ;
	wire _w18694_ ;
	wire _w18695_ ;
	wire _w18696_ ;
	wire _w18697_ ;
	wire _w18698_ ;
	wire _w18699_ ;
	wire _w18700_ ;
	wire _w18701_ ;
	wire _w18702_ ;
	wire _w18703_ ;
	wire _w18704_ ;
	wire _w18705_ ;
	wire _w18706_ ;
	wire _w18707_ ;
	wire _w18708_ ;
	wire _w18709_ ;
	wire _w18710_ ;
	wire _w18711_ ;
	wire _w18712_ ;
	wire _w18713_ ;
	wire _w18714_ ;
	wire _w18715_ ;
	wire _w18716_ ;
	wire _w18717_ ;
	wire _w18718_ ;
	wire _w18719_ ;
	wire _w18720_ ;
	wire _w18721_ ;
	wire _w18722_ ;
	wire _w18723_ ;
	wire _w18724_ ;
	wire _w18725_ ;
	wire _w18726_ ;
	wire _w18727_ ;
	wire _w18728_ ;
	wire _w18729_ ;
	wire _w18730_ ;
	wire _w18731_ ;
	wire _w18732_ ;
	wire _w18733_ ;
	wire _w18734_ ;
	wire _w18735_ ;
	wire _w18736_ ;
	wire _w18737_ ;
	wire _w18738_ ;
	wire _w18739_ ;
	wire _w18740_ ;
	wire _w18741_ ;
	wire _w18742_ ;
	wire _w18743_ ;
	wire _w18744_ ;
	wire _w18745_ ;
	wire _w18746_ ;
	wire _w18747_ ;
	wire _w18748_ ;
	wire _w18749_ ;
	wire _w18750_ ;
	wire _w18751_ ;
	wire _w18752_ ;
	wire _w18753_ ;
	wire _w18754_ ;
	wire _w18755_ ;
	wire _w18756_ ;
	wire _w18757_ ;
	wire _w18758_ ;
	wire _w18759_ ;
	wire _w18760_ ;
	wire _w18761_ ;
	wire _w18762_ ;
	wire _w18763_ ;
	wire _w18764_ ;
	wire _w18765_ ;
	wire _w18766_ ;
	wire _w18767_ ;
	wire _w18768_ ;
	wire _w18769_ ;
	wire _w18770_ ;
	wire _w18771_ ;
	wire _w18772_ ;
	wire _w18773_ ;
	wire _w18774_ ;
	wire _w18775_ ;
	wire _w18776_ ;
	wire _w18777_ ;
	wire _w18778_ ;
	wire _w18779_ ;
	wire _w18780_ ;
	wire _w18781_ ;
	wire _w18782_ ;
	wire _w18783_ ;
	wire _w18784_ ;
	wire _w18785_ ;
	wire _w18786_ ;
	wire _w18787_ ;
	wire _w18788_ ;
	wire _w18789_ ;
	wire _w18790_ ;
	wire _w18791_ ;
	wire _w18792_ ;
	wire _w18793_ ;
	wire _w18794_ ;
	wire _w18795_ ;
	wire _w18796_ ;
	wire _w18797_ ;
	wire _w18798_ ;
	wire _w18799_ ;
	wire _w18800_ ;
	wire _w18801_ ;
	wire _w18802_ ;
	wire _w18803_ ;
	wire _w18804_ ;
	wire _w18805_ ;
	wire _w18806_ ;
	wire _w18807_ ;
	wire _w18808_ ;
	wire _w18809_ ;
	wire _w18810_ ;
	wire _w18811_ ;
	wire _w18812_ ;
	wire _w18813_ ;
	wire _w18814_ ;
	wire _w18815_ ;
	wire _w18816_ ;
	wire _w18817_ ;
	wire _w18818_ ;
	wire _w18819_ ;
	wire _w18820_ ;
	wire _w18821_ ;
	wire _w18822_ ;
	wire _w18823_ ;
	wire _w18824_ ;
	wire _w18825_ ;
	wire _w18826_ ;
	wire _w18827_ ;
	wire _w18828_ ;
	wire _w18829_ ;
	wire _w18830_ ;
	wire _w18831_ ;
	wire _w18832_ ;
	wire _w18833_ ;
	wire _w18834_ ;
	wire _w18835_ ;
	wire _w18836_ ;
	wire _w18837_ ;
	wire _w18838_ ;
	wire _w18839_ ;
	wire _w18840_ ;
	wire _w18841_ ;
	wire _w18842_ ;
	wire _w18843_ ;
	wire _w18844_ ;
	wire _w18845_ ;
	wire _w18846_ ;
	wire _w18847_ ;
	wire _w18848_ ;
	wire _w18849_ ;
	wire _w18850_ ;
	wire _w18851_ ;
	wire _w18852_ ;
	wire _w18853_ ;
	wire _w18854_ ;
	wire _w18855_ ;
	wire _w18856_ ;
	wire _w18857_ ;
	wire _w18858_ ;
	wire _w18859_ ;
	wire _w18860_ ;
	wire _w18861_ ;
	wire _w18862_ ;
	wire _w18863_ ;
	wire _w18864_ ;
	wire _w18865_ ;
	wire _w18866_ ;
	wire _w18867_ ;
	wire _w18868_ ;
	wire _w18869_ ;
	wire _w18870_ ;
	wire _w18871_ ;
	wire _w18872_ ;
	wire _w18873_ ;
	wire _w18874_ ;
	wire _w18875_ ;
	wire _w18876_ ;
	wire _w18877_ ;
	wire _w18878_ ;
	wire _w18879_ ;
	wire _w18880_ ;
	wire _w18881_ ;
	wire _w18882_ ;
	wire _w18883_ ;
	wire _w18884_ ;
	wire _w18885_ ;
	wire _w18886_ ;
	wire _w18887_ ;
	wire _w18888_ ;
	wire _w18889_ ;
	wire _w18890_ ;
	wire _w18891_ ;
	wire _w18892_ ;
	wire _w18893_ ;
	wire _w18894_ ;
	wire _w18895_ ;
	wire _w18896_ ;
	wire _w18897_ ;
	wire _w18898_ ;
	wire _w18899_ ;
	wire _w18900_ ;
	wire _w18901_ ;
	wire _w18902_ ;
	wire _w18903_ ;
	wire _w18904_ ;
	wire _w18905_ ;
	wire _w18906_ ;
	wire _w18907_ ;
	wire _w18908_ ;
	wire _w18909_ ;
	wire _w18910_ ;
	wire _w18911_ ;
	wire _w18912_ ;
	wire _w18913_ ;
	wire _w18914_ ;
	wire _w18915_ ;
	wire _w18916_ ;
	wire _w18917_ ;
	wire _w18918_ ;
	wire _w18919_ ;
	wire _w18920_ ;
	wire _w18921_ ;
	wire _w18922_ ;
	wire _w18923_ ;
	wire _w18924_ ;
	wire _w18925_ ;
	wire _w18926_ ;
	wire _w18927_ ;
	wire _w18928_ ;
	wire _w18929_ ;
	wire _w18930_ ;
	wire _w18931_ ;
	wire _w18932_ ;
	wire _w18933_ ;
	wire _w18934_ ;
	wire _w18935_ ;
	wire _w18936_ ;
	wire _w18937_ ;
	wire _w18938_ ;
	wire _w18939_ ;
	wire _w18940_ ;
	wire _w18941_ ;
	wire _w18942_ ;
	wire _w18943_ ;
	wire _w18944_ ;
	wire _w18945_ ;
	wire _w18946_ ;
	wire _w18947_ ;
	wire _w18948_ ;
	wire _w18949_ ;
	wire _w18950_ ;
	wire _w18951_ ;
	wire _w18952_ ;
	wire _w18953_ ;
	wire _w18954_ ;
	wire _w18955_ ;
	wire _w18956_ ;
	wire _w18957_ ;
	wire _w18958_ ;
	wire _w18959_ ;
	wire _w18960_ ;
	wire _w18961_ ;
	wire _w18962_ ;
	wire _w18963_ ;
	wire _w18964_ ;
	wire _w18965_ ;
	wire _w18966_ ;
	wire _w18967_ ;
	wire _w18968_ ;
	wire _w18969_ ;
	wire _w18970_ ;
	wire _w18971_ ;
	wire _w18972_ ;
	wire _w18973_ ;
	wire _w18974_ ;
	wire _w18975_ ;
	wire _w18976_ ;
	wire _w18977_ ;
	wire _w18978_ ;
	wire _w18979_ ;
	wire _w18980_ ;
	wire _w18981_ ;
	wire _w18982_ ;
	wire _w18983_ ;
	wire _w18984_ ;
	wire _w18985_ ;
	wire _w18986_ ;
	wire _w18987_ ;
	wire _w18988_ ;
	wire _w18989_ ;
	wire _w18990_ ;
	wire _w18991_ ;
	wire _w18992_ ;
	wire _w18993_ ;
	wire _w18994_ ;
	wire _w18995_ ;
	wire _w18996_ ;
	wire _w18997_ ;
	wire _w18998_ ;
	wire _w18999_ ;
	wire _w19000_ ;
	wire _w19001_ ;
	wire _w19002_ ;
	wire _w19003_ ;
	wire _w19004_ ;
	wire _w19005_ ;
	wire _w19006_ ;
	wire _w19007_ ;
	wire _w19008_ ;
	wire _w19009_ ;
	wire _w19010_ ;
	wire _w19011_ ;
	wire _w19012_ ;
	wire _w19013_ ;
	wire _w19014_ ;
	wire _w19015_ ;
	wire _w19016_ ;
	wire _w19017_ ;
	wire _w19018_ ;
	wire _w19019_ ;
	wire _w19020_ ;
	wire _w19021_ ;
	wire _w19022_ ;
	wire _w19023_ ;
	wire _w19024_ ;
	wire _w19025_ ;
	wire _w19026_ ;
	wire _w19027_ ;
	wire _w19028_ ;
	wire _w19029_ ;
	wire _w19030_ ;
	wire _w19031_ ;
	wire _w19032_ ;
	wire _w19033_ ;
	wire _w19034_ ;
	wire _w19035_ ;
	wire _w19036_ ;
	wire _w19037_ ;
	wire _w19038_ ;
	wire _w19039_ ;
	wire _w19040_ ;
	wire _w19041_ ;
	wire _w19042_ ;
	wire _w19043_ ;
	wire _w19044_ ;
	wire _w19045_ ;
	wire _w19046_ ;
	wire _w19047_ ;
	wire _w19048_ ;
	wire _w19049_ ;
	wire _w19050_ ;
	wire _w19051_ ;
	wire _w19052_ ;
	wire _w19053_ ;
	wire _w19054_ ;
	wire _w19055_ ;
	wire _w19056_ ;
	wire _w19057_ ;
	wire _w19058_ ;
	wire _w19059_ ;
	wire _w19060_ ;
	wire _w19061_ ;
	wire _w19062_ ;
	wire _w19063_ ;
	wire _w19064_ ;
	wire _w19065_ ;
	wire _w19066_ ;
	wire _w19067_ ;
	wire _w19068_ ;
	wire _w19069_ ;
	wire _w19070_ ;
	wire _w19071_ ;
	wire _w19072_ ;
	wire _w19073_ ;
	wire _w19074_ ;
	wire _w19075_ ;
	wire _w19076_ ;
	wire _w19077_ ;
	wire _w19078_ ;
	wire _w19079_ ;
	wire _w19080_ ;
	wire _w19081_ ;
	wire _w19082_ ;
	wire _w19083_ ;
	wire _w19084_ ;
	wire _w19085_ ;
	wire _w19086_ ;
	wire _w19087_ ;
	wire _w19088_ ;
	wire _w19089_ ;
	wire _w19090_ ;
	wire _w19091_ ;
	wire _w19092_ ;
	wire _w19093_ ;
	wire _w19094_ ;
	wire _w19095_ ;
	wire _w19096_ ;
	wire _w19097_ ;
	wire _w19098_ ;
	wire _w19099_ ;
	wire _w19100_ ;
	wire _w19101_ ;
	wire _w19102_ ;
	wire _w19103_ ;
	wire _w19104_ ;
	wire _w19105_ ;
	wire _w19106_ ;
	wire _w19107_ ;
	wire _w19108_ ;
	wire _w19109_ ;
	wire _w19110_ ;
	wire _w19111_ ;
	wire _w19112_ ;
	wire _w19113_ ;
	wire _w19114_ ;
	wire _w19115_ ;
	wire _w19116_ ;
	wire _w19117_ ;
	wire _w19118_ ;
	wire _w19119_ ;
	wire _w19120_ ;
	wire _w19121_ ;
	wire _w19122_ ;
	wire _w19123_ ;
	wire _w19124_ ;
	wire _w19125_ ;
	wire _w19126_ ;
	wire _w19127_ ;
	wire _w19128_ ;
	wire _w19129_ ;
	wire _w19130_ ;
	wire _w19131_ ;
	wire _w19132_ ;
	wire _w19133_ ;
	wire _w19134_ ;
	wire _w19135_ ;
	wire _w19136_ ;
	wire _w19137_ ;
	wire _w19138_ ;
	wire _w19139_ ;
	wire _w19140_ ;
	wire _w19141_ ;
	wire _w19142_ ;
	wire _w19143_ ;
	wire _w19144_ ;
	wire _w19145_ ;
	wire _w19146_ ;
	wire _w19147_ ;
	wire _w19148_ ;
	wire _w19149_ ;
	wire _w19150_ ;
	wire _w19151_ ;
	wire _w19152_ ;
	wire _w19153_ ;
	wire _w19154_ ;
	wire _w19155_ ;
	wire _w19156_ ;
	wire _w19157_ ;
	wire _w19158_ ;
	wire _w19159_ ;
	wire _w19160_ ;
	wire _w19161_ ;
	wire _w19162_ ;
	wire _w19163_ ;
	wire _w19164_ ;
	wire _w19165_ ;
	wire _w19166_ ;
	wire _w19167_ ;
	wire _w19168_ ;
	wire _w19169_ ;
	wire _w19170_ ;
	wire _w19171_ ;
	wire _w19172_ ;
	wire _w19173_ ;
	wire _w19174_ ;
	wire _w19175_ ;
	wire _w19176_ ;
	wire _w19177_ ;
	wire _w19178_ ;
	wire _w19179_ ;
	wire _w19180_ ;
	wire _w19181_ ;
	wire _w19182_ ;
	wire _w19183_ ;
	wire _w19184_ ;
	wire _w19185_ ;
	wire _w19186_ ;
	wire _w19187_ ;
	wire _w19188_ ;
	wire _w19189_ ;
	wire _w19190_ ;
	wire _w19191_ ;
	wire _w19192_ ;
	wire _w19193_ ;
	wire _w19194_ ;
	wire _w19195_ ;
	wire _w19196_ ;
	wire _w19197_ ;
	wire _w19198_ ;
	wire _w19199_ ;
	wire _w19200_ ;
	wire _w19201_ ;
	wire _w19202_ ;
	wire _w19203_ ;
	wire _w19204_ ;
	wire _w19205_ ;
	wire _w19206_ ;
	wire _w19207_ ;
	wire _w19208_ ;
	wire _w19209_ ;
	wire _w19210_ ;
	wire _w19211_ ;
	wire _w19212_ ;
	wire _w19213_ ;
	wire _w19214_ ;
	wire _w19215_ ;
	wire _w19216_ ;
	wire _w19217_ ;
	wire _w19218_ ;
	wire _w19219_ ;
	wire _w19220_ ;
	wire _w19221_ ;
	wire _w19222_ ;
	wire _w19223_ ;
	wire _w19224_ ;
	wire _w19225_ ;
	wire _w19226_ ;
	wire _w19227_ ;
	wire _w19228_ ;
	wire _w19229_ ;
	wire _w19230_ ;
	wire _w19231_ ;
	wire _w19232_ ;
	wire _w19233_ ;
	wire _w19234_ ;
	wire _w19235_ ;
	wire _w19236_ ;
	wire _w19237_ ;
	wire _w19238_ ;
	wire _w19239_ ;
	wire _w19240_ ;
	wire _w19241_ ;
	wire _w19242_ ;
	wire _w19243_ ;
	wire _w19244_ ;
	wire _w19245_ ;
	wire _w19246_ ;
	wire _w19247_ ;
	wire _w19248_ ;
	wire _w19249_ ;
	wire _w19250_ ;
	wire _w19251_ ;
	wire _w19252_ ;
	wire _w19253_ ;
	wire _w19254_ ;
	wire _w19255_ ;
	wire _w19256_ ;
	wire _w19257_ ;
	wire _w19258_ ;
	wire _w19259_ ;
	wire _w19260_ ;
	wire _w19261_ ;
	wire _w19262_ ;
	wire _w19263_ ;
	wire _w19264_ ;
	wire _w19265_ ;
	wire _w19266_ ;
	wire _w19267_ ;
	wire _w19268_ ;
	wire _w19269_ ;
	wire _w19270_ ;
	wire _w19271_ ;
	wire _w19272_ ;
	wire _w19273_ ;
	wire _w19274_ ;
	wire _w19275_ ;
	wire _w19276_ ;
	wire _w19277_ ;
	wire _w19278_ ;
	wire _w19279_ ;
	wire _w19280_ ;
	wire _w19281_ ;
	wire _w19282_ ;
	wire _w19283_ ;
	wire _w19284_ ;
	wire _w19285_ ;
	wire _w19286_ ;
	wire _w19287_ ;
	wire _w19288_ ;
	wire _w19289_ ;
	wire _w19290_ ;
	wire _w19291_ ;
	wire _w19292_ ;
	wire _w19293_ ;
	wire _w19294_ ;
	wire _w19295_ ;
	wire _w19296_ ;
	wire _w19297_ ;
	wire _w19298_ ;
	wire _w19299_ ;
	wire _w19300_ ;
	wire _w19301_ ;
	wire _w19302_ ;
	wire _w19303_ ;
	wire _w19304_ ;
	wire _w19305_ ;
	wire _w19306_ ;
	wire _w19307_ ;
	wire _w19308_ ;
	wire _w19309_ ;
	wire _w19310_ ;
	wire _w19311_ ;
	wire _w19312_ ;
	wire _w19313_ ;
	wire _w19314_ ;
	wire _w19315_ ;
	wire _w19316_ ;
	wire _w19317_ ;
	wire _w19318_ ;
	wire _w19319_ ;
	wire _w19320_ ;
	wire _w19321_ ;
	wire _w19322_ ;
	wire _w19323_ ;
	wire _w19324_ ;
	wire _w19325_ ;
	wire _w19326_ ;
	wire _w19327_ ;
	wire _w19328_ ;
	wire _w19329_ ;
	wire _w19330_ ;
	wire _w19331_ ;
	wire _w19332_ ;
	wire _w19333_ ;
	wire _w19334_ ;
	wire _w19335_ ;
	wire _w19336_ ;
	wire _w19337_ ;
	wire _w19338_ ;
	wire _w19339_ ;
	wire _w19340_ ;
	wire _w19341_ ;
	wire _w19342_ ;
	wire _w19343_ ;
	wire _w19344_ ;
	wire _w19345_ ;
	wire _w19346_ ;
	wire _w19347_ ;
	wire _w19348_ ;
	wire _w19349_ ;
	wire _w19350_ ;
	wire _w19351_ ;
	wire _w19352_ ;
	wire _w19353_ ;
	wire _w19354_ ;
	wire _w19355_ ;
	wire _w19356_ ;
	wire _w19357_ ;
	wire _w19358_ ;
	wire _w19359_ ;
	wire _w19360_ ;
	wire _w19361_ ;
	wire _w19362_ ;
	wire _w19363_ ;
	wire _w19364_ ;
	wire _w19365_ ;
	wire _w19366_ ;
	wire _w19367_ ;
	wire _w19368_ ;
	wire _w19369_ ;
	wire _w19370_ ;
	wire _w19371_ ;
	wire _w19372_ ;
	wire _w19373_ ;
	wire _w19374_ ;
	wire _w19375_ ;
	wire _w19376_ ;
	wire _w19377_ ;
	wire _w19378_ ;
	wire _w19379_ ;
	wire _w19380_ ;
	wire _w19381_ ;
	wire _w19382_ ;
	wire _w19383_ ;
	wire _w19384_ ;
	wire _w19385_ ;
	wire _w19386_ ;
	wire _w19387_ ;
	wire _w19388_ ;
	wire _w19389_ ;
	wire _w19390_ ;
	wire _w19391_ ;
	wire _w19392_ ;
	wire _w19393_ ;
	wire _w19394_ ;
	wire _w19395_ ;
	wire _w19396_ ;
	wire _w19397_ ;
	wire _w19398_ ;
	wire _w19399_ ;
	wire _w19400_ ;
	wire _w19401_ ;
	wire _w19402_ ;
	wire _w19403_ ;
	wire _w19404_ ;
	wire _w19405_ ;
	wire _w19406_ ;
	wire _w19407_ ;
	wire _w19408_ ;
	wire _w19409_ ;
	wire _w19410_ ;
	wire _w19411_ ;
	wire _w19412_ ;
	wire _w19413_ ;
	wire _w19414_ ;
	wire _w19415_ ;
	wire _w19416_ ;
	wire _w19417_ ;
	wire _w19418_ ;
	wire _w19419_ ;
	wire _w19420_ ;
	wire _w19421_ ;
	wire _w19422_ ;
	wire _w19423_ ;
	wire _w19424_ ;
	wire _w19425_ ;
	wire _w19426_ ;
	wire _w19427_ ;
	wire _w19428_ ;
	wire _w19429_ ;
	wire _w19430_ ;
	wire _w19431_ ;
	wire _w19432_ ;
	wire _w19433_ ;
	wire _w19434_ ;
	wire _w19435_ ;
	wire _w19436_ ;
	wire _w19437_ ;
	wire _w19438_ ;
	wire _w19439_ ;
	wire _w19440_ ;
	wire _w19441_ ;
	wire _w19442_ ;
	wire _w19443_ ;
	wire _w19444_ ;
	wire _w19445_ ;
	wire _w19446_ ;
	wire _w19447_ ;
	wire _w19448_ ;
	wire _w19449_ ;
	wire _w19450_ ;
	wire _w19451_ ;
	wire _w19452_ ;
	wire _w19453_ ;
	wire _w19454_ ;
	wire _w19455_ ;
	wire _w19456_ ;
	wire _w19457_ ;
	wire _w19458_ ;
	wire _w19459_ ;
	wire _w19460_ ;
	wire _w19461_ ;
	wire _w19462_ ;
	wire _w19463_ ;
	wire _w19464_ ;
	wire _w19465_ ;
	wire _w19466_ ;
	wire _w19467_ ;
	wire _w19468_ ;
	wire _w19469_ ;
	wire _w19470_ ;
	wire _w19471_ ;
	wire _w19472_ ;
	wire _w19473_ ;
	wire _w19474_ ;
	wire _w19475_ ;
	wire _w19476_ ;
	wire _w19477_ ;
	wire _w19478_ ;
	wire _w19479_ ;
	wire _w19480_ ;
	wire _w19481_ ;
	wire _w19482_ ;
	wire _w19483_ ;
	wire _w19484_ ;
	wire _w19485_ ;
	wire _w19486_ ;
	wire _w19487_ ;
	wire _w19488_ ;
	wire _w19489_ ;
	wire _w19490_ ;
	wire _w19491_ ;
	wire _w19492_ ;
	wire _w19493_ ;
	wire _w19494_ ;
	wire _w19495_ ;
	wire _w19496_ ;
	wire _w19497_ ;
	wire _w19498_ ;
	wire _w19499_ ;
	wire _w19500_ ;
	wire _w19501_ ;
	wire _w19502_ ;
	wire _w19503_ ;
	wire _w19504_ ;
	wire _w19505_ ;
	wire _w19506_ ;
	wire _w19507_ ;
	wire _w19508_ ;
	wire _w19509_ ;
	wire _w19510_ ;
	wire _w19511_ ;
	wire _w19512_ ;
	wire _w19513_ ;
	wire _w19514_ ;
	wire _w19515_ ;
	wire _w19516_ ;
	wire _w19517_ ;
	wire _w19518_ ;
	wire _w19519_ ;
	wire _w19520_ ;
	wire _w19521_ ;
	wire _w19522_ ;
	wire _w19523_ ;
	wire _w19524_ ;
	wire _w19525_ ;
	wire _w19526_ ;
	wire _w19527_ ;
	wire _w19528_ ;
	wire _w19529_ ;
	wire _w19530_ ;
	wire _w19531_ ;
	wire _w19532_ ;
	wire _w19533_ ;
	wire _w19534_ ;
	wire _w19535_ ;
	wire _w19536_ ;
	wire _w19537_ ;
	wire _w19538_ ;
	wire _w19539_ ;
	wire _w19540_ ;
	wire _w19541_ ;
	wire _w19542_ ;
	wire _w19543_ ;
	wire _w19544_ ;
	wire _w19545_ ;
	wire _w19546_ ;
	wire _w19547_ ;
	wire _w19548_ ;
	wire _w19549_ ;
	wire _w19550_ ;
	wire _w19551_ ;
	wire _w19552_ ;
	wire _w19553_ ;
	wire _w19554_ ;
	wire _w19555_ ;
	wire _w19556_ ;
	wire _w19557_ ;
	wire _w19558_ ;
	wire _w19559_ ;
	wire _w19560_ ;
	wire _w19561_ ;
	wire _w19562_ ;
	wire _w19563_ ;
	wire _w19564_ ;
	wire _w19565_ ;
	wire _w19566_ ;
	wire _w19567_ ;
	wire _w19568_ ;
	wire _w19569_ ;
	wire _w19570_ ;
	wire _w19571_ ;
	wire _w19572_ ;
	wire _w19573_ ;
	wire _w19574_ ;
	wire _w19575_ ;
	wire _w19576_ ;
	wire _w19577_ ;
	wire _w19578_ ;
	wire _w19579_ ;
	wire _w19580_ ;
	wire _w19581_ ;
	wire _w19582_ ;
	wire _w19583_ ;
	wire _w19584_ ;
	wire _w19585_ ;
	wire _w19586_ ;
	wire _w19587_ ;
	wire _w19588_ ;
	wire _w19589_ ;
	wire _w19590_ ;
	wire _w19591_ ;
	wire _w19592_ ;
	wire _w19593_ ;
	wire _w19594_ ;
	wire _w19595_ ;
	wire _w19596_ ;
	wire _w19597_ ;
	wire _w19598_ ;
	wire _w19599_ ;
	wire _w19600_ ;
	wire _w19601_ ;
	wire _w19602_ ;
	wire _w19603_ ;
	wire _w19604_ ;
	wire _w19605_ ;
	wire _w19606_ ;
	wire _w19607_ ;
	wire _w19608_ ;
	wire _w19609_ ;
	wire _w19610_ ;
	wire _w19611_ ;
	wire _w19612_ ;
	wire _w19613_ ;
	wire _w19614_ ;
	wire _w19615_ ;
	wire _w19616_ ;
	wire _w19617_ ;
	wire _w19618_ ;
	wire _w19619_ ;
	wire _w19620_ ;
	wire _w19621_ ;
	wire _w19622_ ;
	wire _w19623_ ;
	wire _w19624_ ;
	wire _w19625_ ;
	wire _w19626_ ;
	wire _w19627_ ;
	wire _w19628_ ;
	wire _w19629_ ;
	wire _w19630_ ;
	wire _w19631_ ;
	wire _w19632_ ;
	wire _w19633_ ;
	wire _w19634_ ;
	wire _w19635_ ;
	wire _w19636_ ;
	wire _w19637_ ;
	wire _w19638_ ;
	wire _w19639_ ;
	wire _w19640_ ;
	wire _w19641_ ;
	wire _w19642_ ;
	wire _w19643_ ;
	wire _w19644_ ;
	wire _w19645_ ;
	wire _w19646_ ;
	wire _w19647_ ;
	wire _w19648_ ;
	wire _w19649_ ;
	wire _w19650_ ;
	wire _w19651_ ;
	wire _w19652_ ;
	wire _w19653_ ;
	wire _w19654_ ;
	wire _w19655_ ;
	wire _w19656_ ;
	wire _w19657_ ;
	wire _w19658_ ;
	wire _w19659_ ;
	wire _w19660_ ;
	wire _w19661_ ;
	wire _w19662_ ;
	wire _w19663_ ;
	wire _w19664_ ;
	wire _w19665_ ;
	wire _w19666_ ;
	wire _w19667_ ;
	wire _w19668_ ;
	wire _w19669_ ;
	wire _w19670_ ;
	wire _w19671_ ;
	wire _w19672_ ;
	wire _w19673_ ;
	wire _w19674_ ;
	wire _w19675_ ;
	wire _w19676_ ;
	wire _w19677_ ;
	wire _w19678_ ;
	wire _w19679_ ;
	wire _w19680_ ;
	wire _w19681_ ;
	wire _w19682_ ;
	wire _w19683_ ;
	wire _w19684_ ;
	wire _w19685_ ;
	wire _w19686_ ;
	wire _w19687_ ;
	wire _w19688_ ;
	wire _w19689_ ;
	wire _w19690_ ;
	wire _w19691_ ;
	wire _w19692_ ;
	wire _w19693_ ;
	wire _w19694_ ;
	wire _w19695_ ;
	wire _w19696_ ;
	wire _w19697_ ;
	wire _w19698_ ;
	wire _w19699_ ;
	wire _w19700_ ;
	wire _w19701_ ;
	wire _w19702_ ;
	wire _w19703_ ;
	wire _w19704_ ;
	wire _w19705_ ;
	wire _w19706_ ;
	wire _w19707_ ;
	wire _w19708_ ;
	wire _w19709_ ;
	wire _w19710_ ;
	wire _w19711_ ;
	wire _w19712_ ;
	wire _w19713_ ;
	wire _w19714_ ;
	wire _w19715_ ;
	wire _w19716_ ;
	wire _w19717_ ;
	wire _w19718_ ;
	wire _w19719_ ;
	wire _w19720_ ;
	wire _w19721_ ;
	wire _w19722_ ;
	wire _w19723_ ;
	wire _w19724_ ;
	wire _w19725_ ;
	wire _w19726_ ;
	wire _w19727_ ;
	wire _w19728_ ;
	wire _w19729_ ;
	wire _w19730_ ;
	wire _w19731_ ;
	wire _w19732_ ;
	wire _w19733_ ;
	wire _w19734_ ;
	wire _w19735_ ;
	wire _w19736_ ;
	wire _w19737_ ;
	wire _w19738_ ;
	wire _w19739_ ;
	wire _w19740_ ;
	wire _w19741_ ;
	wire _w19742_ ;
	wire _w19743_ ;
	wire _w19744_ ;
	wire _w19745_ ;
	wire _w19746_ ;
	wire _w19747_ ;
	wire _w19748_ ;
	wire _w19749_ ;
	wire _w19750_ ;
	wire _w19751_ ;
	wire _w19752_ ;
	wire _w19753_ ;
	wire _w19754_ ;
	wire _w19755_ ;
	wire _w19756_ ;
	wire _w19757_ ;
	wire _w19758_ ;
	wire _w19759_ ;
	wire _w19760_ ;
	wire _w19761_ ;
	wire _w19762_ ;
	wire _w19763_ ;
	wire _w19764_ ;
	wire _w19765_ ;
	wire _w19766_ ;
	wire _w19767_ ;
	wire _w19768_ ;
	wire _w19769_ ;
	wire _w19770_ ;
	wire _w19771_ ;
	wire _w19772_ ;
	wire _w19773_ ;
	wire _w19774_ ;
	wire _w19775_ ;
	wire _w19776_ ;
	wire _w19777_ ;
	wire _w19778_ ;
	wire _w19779_ ;
	wire _w19780_ ;
	wire _w19781_ ;
	wire _w19782_ ;
	wire _w19783_ ;
	wire _w19784_ ;
	wire _w19785_ ;
	wire _w19786_ ;
	wire _w19787_ ;
	wire _w19788_ ;
	wire _w19789_ ;
	wire _w19790_ ;
	wire _w19791_ ;
	wire _w19792_ ;
	wire _w19793_ ;
	wire _w19794_ ;
	wire _w19795_ ;
	wire _w19796_ ;
	wire _w19797_ ;
	wire _w19798_ ;
	wire _w19799_ ;
	wire _w19800_ ;
	wire _w19801_ ;
	wire _w19802_ ;
	wire _w19803_ ;
	wire _w19804_ ;
	wire _w19805_ ;
	wire _w19806_ ;
	wire _w19807_ ;
	wire _w19808_ ;
	wire _w19809_ ;
	wire _w19810_ ;
	wire _w19811_ ;
	wire _w19812_ ;
	wire _w19813_ ;
	wire _w19814_ ;
	wire _w19815_ ;
	wire _w19816_ ;
	wire _w19817_ ;
	wire _w19818_ ;
	wire _w19819_ ;
	wire _w19820_ ;
	wire _w19821_ ;
	wire _w19822_ ;
	wire _w19823_ ;
	wire _w19824_ ;
	wire _w19825_ ;
	wire _w19826_ ;
	wire _w19827_ ;
	wire _w19828_ ;
	wire _w19829_ ;
	wire _w19830_ ;
	wire _w19831_ ;
	wire _w19832_ ;
	wire _w19833_ ;
	wire _w19834_ ;
	wire _w19835_ ;
	wire _w19836_ ;
	wire _w19837_ ;
	wire _w19838_ ;
	wire _w19839_ ;
	wire _w19840_ ;
	wire _w19841_ ;
	wire _w19842_ ;
	wire _w19843_ ;
	wire _w19844_ ;
	wire _w19845_ ;
	wire _w19846_ ;
	wire _w19847_ ;
	wire _w19848_ ;
	wire _w19849_ ;
	wire _w19850_ ;
	wire _w19851_ ;
	wire _w19852_ ;
	wire _w19853_ ;
	wire _w19854_ ;
	wire _w19855_ ;
	wire _w19856_ ;
	wire _w19857_ ;
	wire _w19858_ ;
	wire _w19859_ ;
	wire _w19860_ ;
	wire _w19861_ ;
	wire _w19862_ ;
	wire _w19863_ ;
	wire _w19864_ ;
	wire _w19865_ ;
	wire _w19866_ ;
	wire _w19867_ ;
	wire _w19868_ ;
	wire _w19869_ ;
	wire _w19870_ ;
	wire _w19871_ ;
	wire _w19872_ ;
	wire _w19873_ ;
	wire _w19874_ ;
	wire _w19875_ ;
	wire _w19876_ ;
	wire _w19877_ ;
	wire _w19878_ ;
	wire _w19879_ ;
	wire _w19880_ ;
	wire _w19881_ ;
	wire _w19882_ ;
	wire _w19883_ ;
	wire _w19884_ ;
	wire _w19885_ ;
	wire _w19886_ ;
	wire _w19887_ ;
	wire _w19888_ ;
	wire _w19889_ ;
	wire _w19890_ ;
	wire _w19891_ ;
	wire _w19892_ ;
	wire _w19893_ ;
	wire _w19894_ ;
	wire _w19895_ ;
	wire _w19896_ ;
	wire _w19897_ ;
	wire _w19898_ ;
	wire _w19899_ ;
	wire _w19900_ ;
	wire _w19901_ ;
	wire _w19902_ ;
	wire _w19903_ ;
	wire _w19904_ ;
	wire _w19905_ ;
	wire _w19906_ ;
	wire _w19907_ ;
	wire _w19908_ ;
	wire _w19909_ ;
	wire _w19910_ ;
	wire _w19911_ ;
	wire _w19912_ ;
	wire _w19913_ ;
	wire _w19914_ ;
	wire _w19915_ ;
	wire _w19916_ ;
	wire _w19917_ ;
	wire _w19918_ ;
	wire _w19919_ ;
	wire _w19920_ ;
	wire _w19921_ ;
	wire _w19922_ ;
	wire _w19923_ ;
	wire _w19924_ ;
	wire _w19925_ ;
	wire _w19926_ ;
	wire _w19927_ ;
	wire _w19928_ ;
	wire _w19929_ ;
	wire _w19930_ ;
	wire _w19931_ ;
	wire _w19932_ ;
	wire _w19933_ ;
	wire _w19934_ ;
	wire _w19935_ ;
	wire _w19936_ ;
	wire _w19937_ ;
	wire _w19938_ ;
	wire _w19939_ ;
	wire _w19940_ ;
	wire _w19941_ ;
	wire _w19942_ ;
	wire _w19943_ ;
	wire _w19944_ ;
	wire _w19945_ ;
	wire _w19946_ ;
	wire _w19947_ ;
	wire _w19948_ ;
	wire _w19949_ ;
	wire _w19950_ ;
	wire _w19951_ ;
	wire _w19952_ ;
	wire _w19953_ ;
	wire _w19954_ ;
	wire _w19955_ ;
	wire _w19956_ ;
	wire _w19957_ ;
	wire _w19958_ ;
	wire _w19959_ ;
	wire _w19960_ ;
	wire _w19961_ ;
	wire _w19962_ ;
	wire _w19963_ ;
	wire _w19964_ ;
	wire _w19965_ ;
	wire _w19966_ ;
	wire _w19967_ ;
	wire _w19968_ ;
	wire _w19969_ ;
	wire _w19970_ ;
	wire _w19971_ ;
	wire _w19972_ ;
	wire _w19973_ ;
	wire _w19974_ ;
	wire _w19975_ ;
	wire _w19976_ ;
	wire _w19977_ ;
	wire _w19978_ ;
	wire _w19979_ ;
	wire _w19980_ ;
	wire _w19981_ ;
	wire _w19982_ ;
	wire _w19983_ ;
	wire _w19984_ ;
	wire _w19985_ ;
	wire _w19986_ ;
	wire _w19987_ ;
	wire _w19988_ ;
	wire _w19989_ ;
	wire _w19990_ ;
	wire _w19991_ ;
	wire _w19992_ ;
	wire _w19993_ ;
	wire _w19994_ ;
	wire _w19995_ ;
	wire _w19996_ ;
	wire _w19997_ ;
	wire _w19998_ ;
	wire _w19999_ ;
	wire _w20000_ ;
	wire _w20001_ ;
	wire _w20002_ ;
	wire _w20003_ ;
	wire _w20004_ ;
	wire _w20005_ ;
	wire _w20006_ ;
	wire _w20007_ ;
	wire _w20008_ ;
	wire _w20009_ ;
	wire _w20010_ ;
	wire _w20011_ ;
	wire _w20012_ ;
	wire _w20013_ ;
	wire _w20014_ ;
	wire _w20015_ ;
	wire _w20016_ ;
	wire _w20017_ ;
	wire _w20018_ ;
	wire _w20019_ ;
	wire _w20020_ ;
	wire _w20021_ ;
	wire _w20022_ ;
	wire _w20023_ ;
	wire _w20024_ ;
	wire _w20025_ ;
	wire _w20026_ ;
	wire _w20027_ ;
	wire _w20028_ ;
	wire _w20029_ ;
	wire _w20030_ ;
	wire _w20031_ ;
	wire _w20032_ ;
	wire _w20033_ ;
	wire _w20034_ ;
	wire _w20035_ ;
	wire _w20036_ ;
	wire _w20037_ ;
	wire _w20038_ ;
	wire _w20039_ ;
	wire _w20040_ ;
	wire _w20041_ ;
	wire _w20042_ ;
	wire _w20043_ ;
	wire _w20044_ ;
	wire _w20045_ ;
	wire _w20046_ ;
	wire _w20047_ ;
	wire _w20048_ ;
	wire _w20049_ ;
	wire _w20050_ ;
	wire _w20051_ ;
	wire _w20052_ ;
	wire _w20053_ ;
	wire _w20054_ ;
	wire _w20055_ ;
	wire _w20056_ ;
	wire _w20057_ ;
	wire _w20058_ ;
	wire _w20059_ ;
	wire _w20060_ ;
	wire _w20061_ ;
	wire _w20062_ ;
	wire _w20063_ ;
	wire _w20064_ ;
	wire _w20065_ ;
	wire _w20066_ ;
	wire _w20067_ ;
	wire _w20068_ ;
	wire _w20069_ ;
	wire _w20070_ ;
	wire _w20071_ ;
	wire _w20072_ ;
	wire _w20073_ ;
	wire _w20074_ ;
	wire _w20075_ ;
	wire _w20076_ ;
	wire _w20077_ ;
	wire _w20078_ ;
	wire _w20079_ ;
	wire _w20080_ ;
	wire _w20081_ ;
	wire _w20082_ ;
	wire _w20083_ ;
	wire _w20084_ ;
	wire _w20085_ ;
	wire _w20086_ ;
	wire _w20087_ ;
	wire _w20088_ ;
	wire _w20089_ ;
	wire _w20090_ ;
	wire _w20091_ ;
	wire _w20092_ ;
	wire _w20093_ ;
	wire _w20094_ ;
	wire _w20095_ ;
	wire _w20096_ ;
	wire _w20097_ ;
	wire _w20098_ ;
	wire _w20099_ ;
	wire _w20100_ ;
	wire _w20101_ ;
	wire _w20102_ ;
	wire _w20103_ ;
	wire _w20104_ ;
	wire _w20105_ ;
	wire _w20106_ ;
	wire _w20107_ ;
	wire _w20108_ ;
	wire _w20109_ ;
	wire _w20110_ ;
	wire _w20111_ ;
	wire _w20112_ ;
	wire _w20113_ ;
	wire _w20114_ ;
	wire _w20115_ ;
	wire _w20116_ ;
	wire _w20117_ ;
	wire _w20118_ ;
	wire _w20119_ ;
	wire _w20120_ ;
	wire _w20121_ ;
	wire _w20122_ ;
	wire _w20123_ ;
	wire _w20124_ ;
	wire _w20125_ ;
	wire _w20126_ ;
	wire _w20127_ ;
	wire _w20128_ ;
	wire _w20129_ ;
	wire _w20130_ ;
	wire _w20131_ ;
	wire _w20132_ ;
	wire _w20133_ ;
	wire _w20134_ ;
	wire _w20135_ ;
	wire _w20136_ ;
	wire _w20137_ ;
	wire _w20138_ ;
	wire _w20139_ ;
	wire _w20140_ ;
	wire _w20141_ ;
	wire _w20142_ ;
	wire _w20143_ ;
	wire _w20144_ ;
	wire _w20145_ ;
	wire _w20146_ ;
	wire _w20147_ ;
	wire _w20148_ ;
	wire _w20149_ ;
	wire _w20150_ ;
	wire _w20151_ ;
	wire _w20152_ ;
	wire _w20153_ ;
	wire _w20154_ ;
	wire _w20155_ ;
	wire _w20156_ ;
	wire _w20157_ ;
	wire _w20158_ ;
	wire _w20159_ ;
	wire _w20160_ ;
	wire _w20161_ ;
	wire _w20162_ ;
	wire _w20163_ ;
	wire _w20164_ ;
	wire _w20165_ ;
	wire _w20166_ ;
	wire _w20167_ ;
	wire _w20168_ ;
	wire _w20169_ ;
	wire _w20170_ ;
	wire _w20171_ ;
	wire _w20172_ ;
	wire _w20173_ ;
	wire _w20174_ ;
	wire _w20175_ ;
	wire _w20176_ ;
	wire _w20177_ ;
	wire _w20178_ ;
	wire _w20179_ ;
	wire _w20180_ ;
	wire _w20181_ ;
	wire _w20182_ ;
	wire _w20183_ ;
	wire _w20184_ ;
	wire _w20185_ ;
	wire _w20186_ ;
	wire _w20187_ ;
	wire _w20188_ ;
	wire _w20189_ ;
	wire _w20190_ ;
	wire _w20191_ ;
	wire _w20192_ ;
	wire _w20193_ ;
	wire _w20194_ ;
	wire _w20195_ ;
	wire _w20196_ ;
	wire _w20197_ ;
	wire _w20198_ ;
	wire _w20199_ ;
	wire _w20200_ ;
	wire _w20201_ ;
	wire _w20202_ ;
	wire _w20203_ ;
	wire _w20204_ ;
	wire _w20205_ ;
	wire _w20206_ ;
	wire _w20207_ ;
	wire _w20208_ ;
	wire _w20209_ ;
	wire _w20210_ ;
	wire _w20211_ ;
	wire _w20212_ ;
	wire _w20213_ ;
	wire _w20214_ ;
	wire _w20215_ ;
	wire _w20216_ ;
	wire _w20217_ ;
	wire _w20218_ ;
	wire _w20219_ ;
	wire _w20220_ ;
	wire _w20221_ ;
	wire _w20222_ ;
	wire _w20223_ ;
	wire _w20224_ ;
	wire _w20225_ ;
	wire _w20226_ ;
	wire _w20227_ ;
	wire _w20228_ ;
	wire _w20229_ ;
	wire _w20230_ ;
	wire _w20231_ ;
	wire _w20232_ ;
	wire _w20233_ ;
	wire _w20234_ ;
	wire _w20235_ ;
	wire _w20236_ ;
	wire _w20237_ ;
	wire _w20238_ ;
	wire _w20239_ ;
	wire _w20240_ ;
	wire _w20241_ ;
	wire _w20242_ ;
	wire _w20243_ ;
	wire _w20244_ ;
	wire _w20245_ ;
	wire _w20246_ ;
	wire _w20247_ ;
	wire _w20248_ ;
	wire _w20249_ ;
	wire _w20250_ ;
	wire _w20251_ ;
	wire _w20252_ ;
	wire _w20253_ ;
	wire _w20254_ ;
	wire _w20255_ ;
	wire _w20256_ ;
	wire _w20257_ ;
	wire _w20258_ ;
	wire _w20259_ ;
	wire _w20260_ ;
	wire _w20261_ ;
	wire _w20262_ ;
	wire _w20263_ ;
	wire _w20264_ ;
	wire _w20265_ ;
	wire _w20266_ ;
	wire _w20267_ ;
	wire _w20268_ ;
	wire _w20269_ ;
	wire _w20270_ ;
	wire _w20271_ ;
	wire _w20272_ ;
	wire _w20273_ ;
	wire _w20274_ ;
	wire _w20275_ ;
	wire _w20276_ ;
	wire _w20277_ ;
	wire _w20278_ ;
	wire _w20279_ ;
	wire _w20280_ ;
	wire _w20281_ ;
	wire _w20282_ ;
	wire _w20283_ ;
	wire _w20284_ ;
	wire _w20285_ ;
	wire _w20286_ ;
	wire _w20287_ ;
	wire _w20288_ ;
	wire _w20289_ ;
	wire _w20290_ ;
	wire _w20291_ ;
	wire _w20292_ ;
	wire _w20293_ ;
	wire _w20294_ ;
	wire _w20295_ ;
	wire _w20296_ ;
	wire _w20297_ ;
	wire _w20298_ ;
	wire _w20299_ ;
	wire _w20300_ ;
	wire _w20301_ ;
	wire _w20302_ ;
	wire _w20303_ ;
	wire _w20304_ ;
	wire _w20305_ ;
	wire _w20306_ ;
	wire _w20307_ ;
	wire _w20308_ ;
	wire _w20309_ ;
	wire _w20310_ ;
	wire _w20311_ ;
	wire _w20312_ ;
	wire _w20313_ ;
	wire _w20314_ ;
	wire _w20315_ ;
	wire _w20316_ ;
	wire _w20317_ ;
	wire _w20318_ ;
	wire _w20319_ ;
	wire _w20320_ ;
	wire _w20321_ ;
	wire _w20322_ ;
	wire _w20323_ ;
	wire _w20324_ ;
	wire _w20325_ ;
	wire _w20326_ ;
	wire _w20327_ ;
	wire _w20328_ ;
	wire _w20329_ ;
	wire _w20330_ ;
	wire _w20331_ ;
	wire _w20332_ ;
	wire _w20333_ ;
	wire _w20334_ ;
	wire _w20335_ ;
	wire _w20336_ ;
	wire _w20337_ ;
	wire _w20338_ ;
	wire _w20339_ ;
	wire _w20340_ ;
	wire _w20341_ ;
	wire _w20342_ ;
	wire _w20343_ ;
	wire _w20344_ ;
	wire _w20345_ ;
	wire _w20346_ ;
	wire _w20347_ ;
	wire _w20348_ ;
	wire _w20349_ ;
	wire _w20350_ ;
	wire _w20351_ ;
	wire _w20352_ ;
	wire _w20353_ ;
	wire _w20354_ ;
	wire _w20355_ ;
	wire _w20356_ ;
	wire _w20357_ ;
	wire _w20358_ ;
	wire _w20359_ ;
	wire _w20360_ ;
	wire _w20361_ ;
	wire _w20362_ ;
	wire _w20363_ ;
	wire _w20364_ ;
	wire _w20365_ ;
	wire _w20366_ ;
	wire _w20367_ ;
	wire _w20368_ ;
	wire _w20369_ ;
	wire _w20370_ ;
	wire _w20371_ ;
	wire _w20372_ ;
	wire _w20373_ ;
	wire _w20374_ ;
	wire _w20375_ ;
	wire _w20376_ ;
	wire _w20377_ ;
	wire _w20378_ ;
	wire _w20379_ ;
	wire _w20380_ ;
	wire _w20381_ ;
	wire _w20382_ ;
	wire _w20383_ ;
	wire _w20384_ ;
	wire _w20385_ ;
	wire _w20386_ ;
	wire _w20387_ ;
	wire _w20388_ ;
	wire _w20389_ ;
	wire _w20390_ ;
	wire _w20391_ ;
	wire _w20392_ ;
	wire _w20393_ ;
	wire _w20394_ ;
	wire _w20395_ ;
	wire _w20396_ ;
	wire _w20397_ ;
	wire _w20398_ ;
	wire _w20399_ ;
	wire _w20400_ ;
	wire _w20401_ ;
	wire _w20402_ ;
	wire _w20403_ ;
	wire _w20404_ ;
	wire _w20405_ ;
	wire _w20406_ ;
	wire _w20407_ ;
	wire _w20408_ ;
	wire _w20409_ ;
	wire _w20410_ ;
	wire _w20411_ ;
	wire _w20412_ ;
	wire _w20413_ ;
	wire _w20414_ ;
	wire _w20415_ ;
	wire _w20416_ ;
	wire _w20417_ ;
	wire _w20418_ ;
	wire _w20419_ ;
	wire _w20420_ ;
	wire _w20421_ ;
	wire _w20422_ ;
	wire _w20423_ ;
	wire _w20424_ ;
	wire _w20425_ ;
	wire _w20426_ ;
	wire _w20427_ ;
	wire _w20428_ ;
	wire _w20429_ ;
	wire _w20430_ ;
	wire _w20431_ ;
	wire _w20432_ ;
	wire _w20433_ ;
	wire _w20434_ ;
	wire _w20435_ ;
	wire _w20436_ ;
	wire _w20437_ ;
	wire _w20438_ ;
	wire _w20439_ ;
	wire _w20440_ ;
	wire _w20441_ ;
	wire _w20442_ ;
	wire _w20443_ ;
	wire _w20444_ ;
	wire _w20445_ ;
	wire _w20446_ ;
	wire _w20447_ ;
	wire _w20448_ ;
	wire _w20449_ ;
	wire _w20450_ ;
	wire _w20451_ ;
	wire _w20452_ ;
	wire _w20453_ ;
	wire _w20454_ ;
	wire _w20455_ ;
	wire _w20456_ ;
	wire _w20457_ ;
	wire _w20458_ ;
	wire _w20459_ ;
	wire _w20460_ ;
	wire _w20461_ ;
	wire _w20462_ ;
	wire _w20463_ ;
	wire _w20464_ ;
	wire _w20465_ ;
	wire _w20466_ ;
	wire _w20467_ ;
	wire _w20468_ ;
	wire _w20469_ ;
	wire _w20470_ ;
	wire _w20471_ ;
	wire _w20472_ ;
	wire _w20473_ ;
	wire _w20474_ ;
	wire _w20475_ ;
	wire _w20476_ ;
	wire _w20477_ ;
	wire _w20478_ ;
	wire _w20479_ ;
	wire _w20480_ ;
	wire _w20481_ ;
	wire _w20482_ ;
	wire _w20483_ ;
	wire _w20484_ ;
	wire _w20485_ ;
	wire _w20486_ ;
	wire _w20487_ ;
	wire _w20488_ ;
	wire _w20489_ ;
	wire _w20490_ ;
	wire _w20491_ ;
	wire _w20492_ ;
	wire _w20493_ ;
	wire _w20494_ ;
	wire _w20495_ ;
	wire _w20496_ ;
	wire _w20497_ ;
	wire _w20498_ ;
	wire _w20499_ ;
	wire _w20500_ ;
	wire _w20501_ ;
	wire _w20502_ ;
	wire _w20503_ ;
	wire _w20504_ ;
	wire _w20505_ ;
	wire _w20506_ ;
	wire _w20507_ ;
	wire _w20508_ ;
	wire _w20509_ ;
	wire _w20510_ ;
	wire _w20511_ ;
	wire _w20512_ ;
	wire _w20513_ ;
	wire _w20514_ ;
	wire _w20515_ ;
	wire _w20516_ ;
	wire _w20517_ ;
	wire _w20518_ ;
	wire _w20519_ ;
	wire _w20520_ ;
	wire _w20521_ ;
	wire _w20522_ ;
	wire _w20523_ ;
	wire _w20524_ ;
	wire _w20525_ ;
	wire _w20526_ ;
	wire _w20527_ ;
	wire _w20528_ ;
	wire _w20529_ ;
	wire _w20530_ ;
	wire _w20531_ ;
	wire _w20532_ ;
	wire _w20533_ ;
	wire _w20534_ ;
	wire _w20535_ ;
	wire _w20536_ ;
	wire _w20537_ ;
	wire _w20538_ ;
	wire _w20539_ ;
	wire _w20540_ ;
	wire _w20541_ ;
	wire _w20542_ ;
	wire _w20543_ ;
	wire _w20544_ ;
	wire _w20545_ ;
	wire _w20546_ ;
	wire _w20547_ ;
	wire _w20548_ ;
	wire _w20549_ ;
	wire _w20550_ ;
	wire _w20551_ ;
	wire _w20552_ ;
	wire _w20553_ ;
	wire _w20554_ ;
	wire _w20555_ ;
	wire _w20556_ ;
	wire _w20557_ ;
	wire _w20558_ ;
	wire _w20559_ ;
	wire _w20560_ ;
	wire _w20561_ ;
	wire _w20562_ ;
	wire _w20563_ ;
	wire _w20564_ ;
	wire _w20565_ ;
	wire _w20566_ ;
	wire _w20567_ ;
	wire _w20568_ ;
	wire _w20569_ ;
	wire _w20570_ ;
	wire _w20571_ ;
	wire _w20572_ ;
	wire _w20573_ ;
	wire _w20574_ ;
	wire _w20575_ ;
	wire _w20576_ ;
	wire _w20577_ ;
	wire _w20578_ ;
	wire _w20579_ ;
	wire _w20580_ ;
	wire _w20581_ ;
	wire _w20582_ ;
	wire _w20583_ ;
	wire _w20584_ ;
	wire _w20585_ ;
	wire _w20586_ ;
	wire _w20587_ ;
	wire _w20588_ ;
	wire _w20589_ ;
	wire _w20590_ ;
	wire _w20591_ ;
	wire _w20592_ ;
	wire _w20593_ ;
	wire _w20594_ ;
	wire _w20595_ ;
	wire _w20596_ ;
	wire _w20597_ ;
	wire _w20598_ ;
	wire _w20599_ ;
	wire _w20600_ ;
	wire _w20601_ ;
	wire _w20602_ ;
	wire _w20603_ ;
	wire _w20604_ ;
	wire _w20605_ ;
	wire _w20606_ ;
	wire _w20607_ ;
	wire _w20608_ ;
	wire _w20609_ ;
	wire _w20610_ ;
	wire _w20611_ ;
	wire _w20612_ ;
	wire _w20613_ ;
	wire _w20614_ ;
	wire _w20615_ ;
	wire _w20616_ ;
	wire _w20617_ ;
	wire _w20618_ ;
	wire _w20619_ ;
	wire _w20620_ ;
	wire _w20621_ ;
	wire _w20622_ ;
	wire _w20623_ ;
	wire _w20624_ ;
	wire _w20625_ ;
	wire _w20626_ ;
	wire _w20627_ ;
	wire _w20628_ ;
	wire _w20629_ ;
	wire _w20630_ ;
	wire _w20631_ ;
	wire _w20632_ ;
	wire _w20633_ ;
	wire _w20634_ ;
	wire _w20635_ ;
	wire _w20636_ ;
	wire _w20637_ ;
	wire _w20638_ ;
	wire _w20639_ ;
	wire _w20640_ ;
	wire _w20641_ ;
	wire _w20642_ ;
	wire _w20643_ ;
	wire _w20644_ ;
	wire _w20645_ ;
	wire _w20646_ ;
	wire _w20647_ ;
	wire _w20648_ ;
	wire _w20649_ ;
	wire _w20650_ ;
	wire _w20651_ ;
	wire _w20652_ ;
	wire _w20653_ ;
	wire _w20654_ ;
	wire _w20655_ ;
	wire _w20656_ ;
	wire _w20657_ ;
	wire _w20658_ ;
	wire _w20659_ ;
	wire _w20660_ ;
	wire _w20661_ ;
	wire _w20662_ ;
	wire _w20663_ ;
	wire _w20664_ ;
	wire _w20665_ ;
	wire _w20666_ ;
	wire _w20667_ ;
	wire _w20668_ ;
	wire _w20669_ ;
	wire _w20670_ ;
	wire _w20671_ ;
	wire _w20672_ ;
	wire _w20673_ ;
	wire _w20674_ ;
	wire _w20675_ ;
	wire _w20676_ ;
	wire _w20677_ ;
	wire _w20678_ ;
	wire _w20679_ ;
	wire _w20680_ ;
	wire _w20681_ ;
	wire _w20682_ ;
	wire _w20683_ ;
	wire _w20684_ ;
	wire _w20685_ ;
	wire _w20686_ ;
	wire _w20687_ ;
	wire _w20688_ ;
	wire _w20689_ ;
	wire _w20690_ ;
	wire _w20691_ ;
	wire _w20692_ ;
	wire _w20693_ ;
	wire _w20694_ ;
	wire _w20695_ ;
	wire _w20696_ ;
	wire _w20697_ ;
	wire _w20698_ ;
	wire _w20699_ ;
	wire _w20700_ ;
	wire _w20701_ ;
	wire _w20702_ ;
	wire _w20703_ ;
	wire _w20704_ ;
	wire _w20705_ ;
	wire _w20706_ ;
	wire _w20707_ ;
	wire _w20708_ ;
	wire _w20709_ ;
	wire _w20710_ ;
	wire _w20711_ ;
	wire _w20712_ ;
	wire _w20713_ ;
	wire _w20714_ ;
	wire _w20715_ ;
	wire _w20716_ ;
	wire _w20717_ ;
	wire _w20718_ ;
	wire _w20719_ ;
	wire _w20720_ ;
	wire _w20721_ ;
	wire _w20722_ ;
	wire _w20723_ ;
	wire _w20724_ ;
	wire _w20725_ ;
	wire _w20726_ ;
	wire _w20727_ ;
	wire _w20728_ ;
	wire _w20729_ ;
	wire _w20730_ ;
	wire _w20731_ ;
	wire _w20732_ ;
	wire _w20733_ ;
	wire _w20734_ ;
	wire _w20735_ ;
	wire _w20736_ ;
	wire _w20737_ ;
	wire _w20738_ ;
	wire _w20739_ ;
	wire _w20740_ ;
	wire _w20741_ ;
	wire _w20742_ ;
	wire _w20743_ ;
	wire _w20744_ ;
	wire _w20745_ ;
	wire _w20746_ ;
	wire _w20747_ ;
	wire _w20748_ ;
	wire _w20749_ ;
	wire _w20750_ ;
	wire _w20751_ ;
	wire _w20752_ ;
	wire _w20753_ ;
	wire _w20754_ ;
	wire _w20755_ ;
	wire _w20756_ ;
	wire _w20757_ ;
	wire _w20758_ ;
	wire _w20759_ ;
	wire _w20760_ ;
	wire _w20761_ ;
	wire _w20762_ ;
	wire _w20763_ ;
	wire _w20764_ ;
	wire _w20765_ ;
	wire _w20766_ ;
	wire _w20767_ ;
	wire _w20768_ ;
	wire _w20769_ ;
	wire _w20770_ ;
	wire _w20771_ ;
	wire _w20772_ ;
	wire _w20773_ ;
	wire _w20774_ ;
	wire _w20775_ ;
	wire _w20776_ ;
	wire _w20777_ ;
	wire _w20778_ ;
	wire _w20779_ ;
	wire _w20780_ ;
	wire _w20781_ ;
	wire _w20782_ ;
	wire _w20783_ ;
	wire _w20784_ ;
	wire _w20785_ ;
	wire _w20786_ ;
	wire _w20787_ ;
	wire _w20788_ ;
	wire _w20789_ ;
	wire _w20790_ ;
	wire _w20791_ ;
	wire _w20792_ ;
	wire _w20793_ ;
	wire _w20794_ ;
	wire _w20795_ ;
	wire _w20796_ ;
	wire _w20797_ ;
	wire _w20798_ ;
	wire _w20799_ ;
	wire _w20800_ ;
	wire _w20801_ ;
	wire _w20802_ ;
	wire _w20803_ ;
	wire _w20804_ ;
	wire _w20805_ ;
	wire _w20806_ ;
	wire _w20807_ ;
	wire _w20808_ ;
	wire _w20809_ ;
	wire _w20810_ ;
	wire _w20811_ ;
	wire _w20812_ ;
	wire _w20813_ ;
	wire _w20814_ ;
	wire _w20815_ ;
	wire _w20816_ ;
	wire _w20817_ ;
	wire _w20818_ ;
	wire _w20819_ ;
	wire _w20820_ ;
	wire _w20821_ ;
	wire _w20822_ ;
	wire _w20823_ ;
	wire _w20824_ ;
	wire _w20825_ ;
	wire _w20826_ ;
	wire _w20827_ ;
	wire _w20828_ ;
	wire _w20829_ ;
	wire _w20830_ ;
	wire _w20831_ ;
	wire _w20832_ ;
	wire _w20833_ ;
	wire _w20834_ ;
	wire _w20835_ ;
	wire _w20836_ ;
	wire _w20837_ ;
	wire _w20838_ ;
	wire _w20839_ ;
	wire _w20840_ ;
	wire _w20841_ ;
	wire _w20842_ ;
	wire _w20843_ ;
	wire _w20844_ ;
	wire _w20845_ ;
	wire _w20846_ ;
	wire _w20847_ ;
	wire _w20848_ ;
	wire _w20849_ ;
	wire _w20850_ ;
	wire _w20851_ ;
	wire _w20852_ ;
	wire _w20853_ ;
	wire _w20854_ ;
	wire _w20855_ ;
	wire _w20856_ ;
	wire _w20857_ ;
	wire _w20858_ ;
	wire _w20859_ ;
	wire _w20860_ ;
	wire _w20861_ ;
	wire _w20862_ ;
	wire _w20863_ ;
	wire _w20864_ ;
	wire _w20865_ ;
	wire _w20866_ ;
	wire _w20867_ ;
	wire _w20868_ ;
	wire _w20869_ ;
	wire _w20870_ ;
	wire _w20871_ ;
	wire _w20872_ ;
	wire _w20873_ ;
	wire _w20874_ ;
	wire _w20875_ ;
	wire _w20876_ ;
	wire _w20877_ ;
	wire _w20878_ ;
	wire _w20879_ ;
	wire _w20880_ ;
	wire _w20881_ ;
	wire _w20882_ ;
	wire _w20883_ ;
	wire _w20884_ ;
	wire _w20885_ ;
	wire _w20886_ ;
	wire _w20887_ ;
	wire _w20888_ ;
	wire _w20889_ ;
	wire _w20890_ ;
	wire _w20891_ ;
	wire _w20892_ ;
	wire _w20893_ ;
	wire _w20894_ ;
	wire _w20895_ ;
	wire _w20896_ ;
	wire _w20897_ ;
	wire _w20898_ ;
	wire _w20899_ ;
	wire _w20900_ ;
	wire _w20901_ ;
	wire _w20902_ ;
	wire _w20903_ ;
	wire _w20904_ ;
	wire _w20905_ ;
	wire _w20906_ ;
	wire _w20907_ ;
	wire _w20908_ ;
	wire _w20909_ ;
	wire _w20910_ ;
	wire _w20911_ ;
	wire _w20912_ ;
	wire _w20913_ ;
	wire _w20914_ ;
	wire _w20915_ ;
	wire _w20916_ ;
	wire _w20917_ ;
	wire _w20918_ ;
	wire _w20919_ ;
	wire _w20920_ ;
	wire _w20921_ ;
	wire _w20922_ ;
	wire _w20923_ ;
	wire _w20924_ ;
	wire _w20925_ ;
	wire _w20926_ ;
	wire _w20927_ ;
	wire _w20928_ ;
	wire _w20929_ ;
	wire _w20930_ ;
	wire _w20931_ ;
	wire _w20932_ ;
	wire _w20933_ ;
	wire _w20934_ ;
	wire _w20935_ ;
	wire _w20936_ ;
	wire _w20937_ ;
	wire _w20938_ ;
	wire _w20939_ ;
	wire _w20940_ ;
	wire _w20941_ ;
	wire _w20942_ ;
	wire _w20943_ ;
	wire _w20944_ ;
	wire _w20945_ ;
	wire _w20946_ ;
	wire _w20947_ ;
	wire _w20948_ ;
	wire _w20949_ ;
	wire _w20950_ ;
	wire _w20951_ ;
	wire _w20952_ ;
	wire _w20953_ ;
	wire _w20954_ ;
	wire _w20955_ ;
	wire _w20956_ ;
	wire _w20957_ ;
	wire _w20958_ ;
	wire _w20959_ ;
	wire _w20960_ ;
	wire _w20961_ ;
	wire _w20962_ ;
	wire _w20963_ ;
	wire _w20964_ ;
	wire _w20965_ ;
	wire _w20966_ ;
	wire _w20967_ ;
	wire _w20968_ ;
	wire _w20969_ ;
	wire _w20970_ ;
	wire _w20971_ ;
	wire _w20972_ ;
	wire _w20973_ ;
	wire _w20974_ ;
	wire _w20975_ ;
	wire _w20976_ ;
	wire _w20977_ ;
	wire _w20978_ ;
	wire _w20979_ ;
	wire _w20980_ ;
	wire _w20981_ ;
	wire _w20982_ ;
	wire _w20983_ ;
	wire _w20984_ ;
	wire _w20985_ ;
	wire _w20986_ ;
	wire _w20987_ ;
	wire _w20988_ ;
	wire _w20989_ ;
	wire _w20990_ ;
	wire _w20991_ ;
	wire _w20992_ ;
	wire _w20993_ ;
	wire _w20994_ ;
	wire _w20995_ ;
	wire _w20996_ ;
	wire _w20997_ ;
	wire _w20998_ ;
	wire _w20999_ ;
	wire _w21000_ ;
	wire _w21001_ ;
	wire _w21002_ ;
	wire _w21003_ ;
	wire _w21004_ ;
	wire _w21005_ ;
	wire _w21006_ ;
	wire _w21007_ ;
	wire _w21008_ ;
	wire _w21009_ ;
	wire _w21010_ ;
	wire _w21011_ ;
	wire _w21012_ ;
	wire _w21013_ ;
	wire _w21014_ ;
	wire _w21015_ ;
	wire _w21016_ ;
	wire _w21017_ ;
	wire _w21018_ ;
	wire _w21019_ ;
	wire _w21020_ ;
	wire _w21021_ ;
	wire _w21022_ ;
	wire _w21023_ ;
	wire _w21024_ ;
	wire _w21025_ ;
	wire _w21026_ ;
	wire _w21027_ ;
	wire _w21028_ ;
	wire _w21029_ ;
	wire _w21030_ ;
	wire _w21031_ ;
	wire _w21032_ ;
	wire _w21033_ ;
	wire _w21034_ ;
	wire _w21035_ ;
	wire _w21036_ ;
	wire _w21037_ ;
	wire _w21038_ ;
	wire _w21039_ ;
	wire _w21040_ ;
	wire _w21041_ ;
	wire _w21042_ ;
	wire _w21043_ ;
	wire _w21044_ ;
	wire _w21045_ ;
	wire _w21046_ ;
	wire _w21047_ ;
	wire _w21048_ ;
	wire _w21049_ ;
	wire _w21050_ ;
	wire _w21051_ ;
	wire _w21052_ ;
	wire _w21053_ ;
	wire _w21054_ ;
	wire _w21055_ ;
	wire _w21056_ ;
	wire _w21057_ ;
	wire _w21058_ ;
	wire _w21059_ ;
	wire _w21060_ ;
	wire _w21061_ ;
	wire _w21062_ ;
	wire _w21063_ ;
	wire _w21064_ ;
	wire _w21065_ ;
	wire _w21066_ ;
	wire _w21067_ ;
	wire _w21068_ ;
	wire _w21069_ ;
	wire _w21070_ ;
	wire _w21071_ ;
	wire _w21072_ ;
	wire _w21073_ ;
	wire _w21074_ ;
	wire _w21075_ ;
	wire _w21076_ ;
	wire _w21077_ ;
	wire _w21078_ ;
	wire _w21079_ ;
	wire _w21080_ ;
	wire _w21081_ ;
	wire _w21082_ ;
	wire _w21083_ ;
	wire _w21084_ ;
	wire _w21085_ ;
	wire _w21086_ ;
	wire _w21087_ ;
	wire _w21088_ ;
	wire _w21089_ ;
	wire _w21090_ ;
	wire _w21091_ ;
	wire _w21092_ ;
	wire _w21093_ ;
	wire _w21094_ ;
	wire _w21095_ ;
	wire _w21096_ ;
	wire _w21097_ ;
	wire _w21098_ ;
	wire _w21099_ ;
	wire _w21100_ ;
	wire _w21101_ ;
	wire _w21102_ ;
	wire _w21103_ ;
	wire _w21104_ ;
	wire _w21105_ ;
	wire _w21106_ ;
	wire _w21107_ ;
	wire _w21108_ ;
	wire _w21109_ ;
	wire _w21110_ ;
	wire _w21111_ ;
	wire _w21112_ ;
	wire _w21113_ ;
	wire _w21114_ ;
	wire _w21115_ ;
	wire _w21116_ ;
	wire _w21117_ ;
	wire _w21118_ ;
	wire _w21119_ ;
	wire _w21120_ ;
	wire _w21121_ ;
	wire _w21122_ ;
	wire _w21123_ ;
	wire _w21124_ ;
	wire _w21125_ ;
	wire _w21126_ ;
	wire _w21127_ ;
	wire _w21128_ ;
	wire _w21129_ ;
	wire _w21130_ ;
	wire _w21131_ ;
	wire _w21132_ ;
	wire _w21133_ ;
	wire _w21134_ ;
	wire _w21135_ ;
	wire _w21136_ ;
	wire _w21137_ ;
	wire _w21138_ ;
	wire _w21139_ ;
	wire _w21140_ ;
	wire _w21141_ ;
	wire _w21142_ ;
	wire _w21143_ ;
	wire _w21144_ ;
	wire _w21145_ ;
	wire _w21146_ ;
	wire _w21147_ ;
	wire _w21148_ ;
	wire _w21149_ ;
	wire _w21150_ ;
	wire _w21151_ ;
	wire _w21152_ ;
	wire _w21153_ ;
	wire _w21154_ ;
	wire _w21155_ ;
	wire _w21156_ ;
	wire _w21157_ ;
	wire _w21158_ ;
	wire _w21159_ ;
	wire _w21160_ ;
	wire _w21161_ ;
	wire _w21162_ ;
	wire _w21163_ ;
	wire _w21164_ ;
	wire _w21165_ ;
	wire _w21166_ ;
	wire _w21167_ ;
	wire _w21168_ ;
	wire _w21169_ ;
	wire _w21170_ ;
	wire _w21171_ ;
	wire _w21172_ ;
	wire _w21173_ ;
	wire _w21174_ ;
	wire _w21175_ ;
	wire _w21176_ ;
	wire _w21177_ ;
	wire _w21178_ ;
	wire _w21179_ ;
	wire _w21180_ ;
	wire _w21181_ ;
	wire _w21182_ ;
	wire _w21183_ ;
	wire _w21184_ ;
	wire _w21185_ ;
	wire _w21186_ ;
	wire _w21187_ ;
	wire _w21188_ ;
	wire _w21189_ ;
	wire _w21190_ ;
	wire _w21191_ ;
	wire _w21192_ ;
	wire _w21193_ ;
	wire _w21194_ ;
	wire _w21195_ ;
	wire _w21196_ ;
	wire _w21197_ ;
	wire _w21198_ ;
	wire _w21199_ ;
	wire _w21200_ ;
	wire _w21201_ ;
	wire _w21202_ ;
	wire _w21203_ ;
	wire _w21204_ ;
	wire _w21205_ ;
	wire _w21206_ ;
	wire _w21207_ ;
	wire _w21208_ ;
	wire _w21209_ ;
	wire _w21210_ ;
	wire _w21211_ ;
	wire _w21212_ ;
	wire _w21213_ ;
	wire _w21214_ ;
	wire _w21215_ ;
	wire _w21216_ ;
	wire _w21217_ ;
	wire _w21218_ ;
	wire _w21219_ ;
	wire _w21220_ ;
	wire _w21221_ ;
	wire _w21222_ ;
	wire _w21223_ ;
	wire _w21224_ ;
	wire _w21225_ ;
	wire _w21226_ ;
	wire _w21227_ ;
	wire _w21228_ ;
	wire _w21229_ ;
	wire _w21230_ ;
	wire _w21231_ ;
	wire _w21232_ ;
	wire _w21233_ ;
	wire _w21234_ ;
	wire _w21235_ ;
	wire _w21236_ ;
	wire _w21237_ ;
	wire _w21238_ ;
	wire _w21239_ ;
	wire _w21240_ ;
	wire _w21241_ ;
	wire _w21242_ ;
	wire _w21243_ ;
	wire _w21244_ ;
	wire _w21245_ ;
	wire _w21246_ ;
	wire _w21247_ ;
	wire _w21248_ ;
	wire _w21249_ ;
	wire _w21250_ ;
	wire _w21251_ ;
	wire _w21252_ ;
	wire _w21253_ ;
	wire _w21254_ ;
	wire _w21255_ ;
	wire _w21256_ ;
	wire _w21257_ ;
	wire _w21258_ ;
	wire _w21259_ ;
	wire _w21260_ ;
	wire _w21261_ ;
	wire _w21262_ ;
	wire _w21263_ ;
	wire _w21264_ ;
	wire _w21265_ ;
	wire _w21266_ ;
	wire _w21267_ ;
	wire _w21268_ ;
	wire _w21269_ ;
	wire _w21270_ ;
	wire _w21271_ ;
	wire _w21272_ ;
	wire _w21273_ ;
	wire _w21274_ ;
	wire _w21275_ ;
	wire _w21276_ ;
	wire _w21277_ ;
	wire _w21278_ ;
	wire _w21279_ ;
	wire _w21280_ ;
	wire _w21281_ ;
	wire _w21282_ ;
	wire _w21283_ ;
	wire _w21284_ ;
	wire _w21285_ ;
	wire _w21286_ ;
	wire _w21287_ ;
	wire _w21288_ ;
	wire _w21289_ ;
	wire _w21290_ ;
	wire _w21291_ ;
	wire _w21292_ ;
	wire _w21293_ ;
	wire _w21294_ ;
	wire _w21295_ ;
	wire _w21296_ ;
	wire _w21297_ ;
	wire _w21298_ ;
	wire _w21299_ ;
	wire _w21300_ ;
	wire _w21301_ ;
	wire _w21302_ ;
	wire _w21303_ ;
	wire _w21304_ ;
	wire _w21305_ ;
	wire _w21306_ ;
	wire _w21307_ ;
	wire _w21308_ ;
	wire _w21309_ ;
	wire _w21310_ ;
	wire _w21311_ ;
	wire _w21312_ ;
	wire _w21313_ ;
	wire _w21314_ ;
	wire _w21315_ ;
	wire _w21316_ ;
	wire _w21317_ ;
	wire _w21318_ ;
	wire _w21319_ ;
	wire _w21320_ ;
	wire _w21321_ ;
	wire _w21322_ ;
	wire _w21323_ ;
	wire _w21324_ ;
	wire _w21325_ ;
	wire _w21326_ ;
	wire _w21327_ ;
	wire _w21328_ ;
	wire _w21329_ ;
	wire _w21330_ ;
	wire _w21331_ ;
	wire _w21332_ ;
	wire _w21333_ ;
	wire _w21334_ ;
	wire _w21335_ ;
	wire _w21336_ ;
	wire _w21337_ ;
	wire _w21338_ ;
	wire _w21339_ ;
	wire _w21340_ ;
	wire _w21341_ ;
	wire _w21342_ ;
	wire _w21343_ ;
	wire _w21344_ ;
	wire _w21345_ ;
	wire _w21346_ ;
	wire _w21347_ ;
	wire _w21348_ ;
	wire _w21349_ ;
	wire _w21350_ ;
	wire _w21351_ ;
	wire _w21352_ ;
	wire _w21353_ ;
	wire _w21354_ ;
	wire _w21355_ ;
	wire _w21356_ ;
	wire _w21357_ ;
	wire _w21358_ ;
	wire _w21359_ ;
	wire _w21360_ ;
	wire _w21361_ ;
	wire _w21362_ ;
	wire _w21363_ ;
	wire _w21364_ ;
	wire _w21365_ ;
	wire _w21366_ ;
	wire _w21367_ ;
	wire _w21368_ ;
	wire _w21369_ ;
	wire _w21370_ ;
	wire _w21371_ ;
	wire _w21372_ ;
	wire _w21373_ ;
	wire _w21374_ ;
	wire _w21375_ ;
	wire _w21376_ ;
	wire _w21377_ ;
	wire _w21378_ ;
	wire _w21379_ ;
	wire _w21380_ ;
	wire _w21381_ ;
	wire _w21382_ ;
	wire _w21383_ ;
	wire _w21384_ ;
	wire _w21385_ ;
	wire _w21386_ ;
	wire _w21387_ ;
	wire _w21388_ ;
	wire _w21389_ ;
	wire _w21390_ ;
	wire _w21391_ ;
	wire _w21392_ ;
	wire _w21393_ ;
	wire _w21394_ ;
	wire _w21395_ ;
	wire _w21396_ ;
	wire _w21397_ ;
	wire _w21398_ ;
	wire _w21399_ ;
	wire _w21400_ ;
	wire _w21401_ ;
	wire _w21402_ ;
	wire _w21403_ ;
	wire _w21404_ ;
	wire _w21405_ ;
	wire _w21406_ ;
	wire _w21407_ ;
	wire _w21408_ ;
	wire _w21409_ ;
	wire _w21410_ ;
	wire _w21411_ ;
	wire _w21412_ ;
	wire _w21413_ ;
	wire _w21414_ ;
	wire _w21415_ ;
	wire _w21416_ ;
	wire _w21417_ ;
	wire _w21418_ ;
	wire _w21419_ ;
	wire _w21420_ ;
	wire _w21421_ ;
	wire _w21422_ ;
	wire _w21423_ ;
	wire _w21424_ ;
	wire _w21425_ ;
	wire _w21426_ ;
	wire _w21427_ ;
	wire _w21428_ ;
	wire _w21429_ ;
	wire _w21430_ ;
	wire _w21431_ ;
	wire _w21432_ ;
	wire _w21433_ ;
	wire _w21434_ ;
	wire _w21435_ ;
	wire _w21436_ ;
	wire _w21437_ ;
	wire _w21438_ ;
	wire _w21439_ ;
	wire _w21440_ ;
	wire _w21441_ ;
	wire _w21442_ ;
	wire _w21443_ ;
	wire _w21444_ ;
	wire _w21445_ ;
	wire _w21446_ ;
	wire _w21447_ ;
	wire _w21448_ ;
	wire _w21449_ ;
	wire _w21450_ ;
	wire _w21451_ ;
	wire _w21452_ ;
	wire _w21453_ ;
	wire _w21454_ ;
	wire _w21455_ ;
	wire _w21456_ ;
	wire _w21457_ ;
	wire _w21458_ ;
	wire _w21459_ ;
	wire _w21460_ ;
	wire _w21461_ ;
	wire _w21462_ ;
	wire _w21463_ ;
	wire _w21464_ ;
	wire _w21465_ ;
	wire _w21466_ ;
	wire _w21467_ ;
	wire _w21468_ ;
	wire _w21469_ ;
	wire _w21470_ ;
	wire _w21471_ ;
	wire _w21472_ ;
	wire _w21473_ ;
	wire _w21474_ ;
	wire _w21475_ ;
	wire _w21476_ ;
	wire _w21477_ ;
	wire _w21478_ ;
	wire _w21479_ ;
	wire _w21480_ ;
	wire _w21481_ ;
	wire _w21482_ ;
	wire _w21483_ ;
	wire _w21484_ ;
	wire _w21485_ ;
	wire _w21486_ ;
	wire _w21487_ ;
	wire _w21488_ ;
	wire _w21489_ ;
	wire _w21490_ ;
	wire _w21491_ ;
	wire _w21492_ ;
	wire _w21493_ ;
	wire _w21494_ ;
	wire _w21495_ ;
	wire _w21496_ ;
	wire _w21497_ ;
	wire _w21498_ ;
	wire _w21499_ ;
	wire _w21500_ ;
	wire _w21501_ ;
	wire _w21502_ ;
	wire _w21503_ ;
	wire _w21504_ ;
	wire _w21505_ ;
	wire _w21506_ ;
	wire _w21507_ ;
	wire _w21508_ ;
	wire _w21509_ ;
	wire _w21510_ ;
	wire _w21511_ ;
	wire _w21512_ ;
	wire _w21513_ ;
	wire _w21514_ ;
	wire _w21515_ ;
	wire _w21516_ ;
	wire _w21517_ ;
	wire _w21518_ ;
	wire _w21519_ ;
	wire _w21520_ ;
	wire _w21521_ ;
	wire _w21522_ ;
	wire _w21523_ ;
	wire _w21524_ ;
	wire _w21525_ ;
	wire _w21526_ ;
	wire _w21527_ ;
	wire _w21528_ ;
	wire _w21529_ ;
	wire _w21530_ ;
	wire _w21531_ ;
	wire _w21532_ ;
	wire _w21533_ ;
	wire _w21534_ ;
	wire _w21535_ ;
	wire _w21536_ ;
	wire _w21537_ ;
	wire _w21538_ ;
	wire _w21539_ ;
	wire _w21540_ ;
	wire _w21541_ ;
	wire _w21542_ ;
	wire _w21543_ ;
	wire _w21544_ ;
	wire _w21545_ ;
	wire _w21546_ ;
	wire _w21547_ ;
	wire _w21548_ ;
	wire _w21549_ ;
	wire _w21550_ ;
	wire _w21551_ ;
	wire _w21552_ ;
	wire _w21553_ ;
	wire _w21554_ ;
	wire _w21555_ ;
	wire _w21556_ ;
	wire _w21557_ ;
	wire _w21558_ ;
	wire _w21559_ ;
	wire _w21560_ ;
	wire _w21561_ ;
	wire _w21562_ ;
	wire _w21563_ ;
	wire _w21564_ ;
	wire _w21565_ ;
	wire _w21566_ ;
	wire _w21567_ ;
	wire _w21568_ ;
	wire _w21569_ ;
	wire _w21570_ ;
	wire _w21571_ ;
	wire _w21572_ ;
	wire _w21573_ ;
	wire _w21574_ ;
	wire _w21575_ ;
	wire _w21576_ ;
	wire _w21577_ ;
	wire _w21578_ ;
	wire _w21579_ ;
	wire _w21580_ ;
	wire _w21581_ ;
	wire _w21582_ ;
	wire _w21583_ ;
	wire _w21584_ ;
	wire _w21585_ ;
	wire _w21586_ ;
	wire _w21587_ ;
	wire _w21588_ ;
	wire _w21589_ ;
	wire _w21590_ ;
	wire _w21591_ ;
	wire _w21592_ ;
	wire _w21593_ ;
	wire _w21594_ ;
	wire _w21595_ ;
	wire _w21596_ ;
	wire _w21597_ ;
	wire _w21598_ ;
	wire _w21599_ ;
	wire _w21600_ ;
	wire _w21601_ ;
	wire _w21602_ ;
	wire _w21603_ ;
	wire _w21604_ ;
	wire _w21605_ ;
	wire _w21606_ ;
	wire _w21607_ ;
	wire _w21608_ ;
	wire _w21609_ ;
	wire _w21610_ ;
	wire _w21611_ ;
	wire _w21612_ ;
	wire _w21613_ ;
	wire _w21614_ ;
	wire _w21615_ ;
	wire _w21616_ ;
	wire _w21617_ ;
	wire _w21618_ ;
	wire _w21619_ ;
	wire _w21620_ ;
	wire _w21621_ ;
	wire _w21622_ ;
	wire _w21623_ ;
	wire _w21624_ ;
	wire _w21625_ ;
	wire _w21626_ ;
	wire _w21627_ ;
	wire _w21628_ ;
	wire _w21629_ ;
	wire _w21630_ ;
	wire _w21631_ ;
	wire _w21632_ ;
	wire _w21633_ ;
	wire _w21634_ ;
	wire _w21635_ ;
	wire _w21636_ ;
	wire _w21637_ ;
	wire _w21638_ ;
	wire _w21639_ ;
	wire _w21640_ ;
	wire _w21641_ ;
	wire _w21642_ ;
	wire _w21643_ ;
	wire _w21644_ ;
	wire _w21645_ ;
	wire _w21646_ ;
	wire _w21647_ ;
	wire _w21648_ ;
	wire _w21649_ ;
	wire _w21650_ ;
	wire _w21651_ ;
	wire _w21652_ ;
	wire _w21653_ ;
	wire _w21654_ ;
	wire _w21655_ ;
	wire _w21656_ ;
	wire _w21657_ ;
	wire _w21658_ ;
	wire _w21659_ ;
	wire _w21660_ ;
	wire _w21661_ ;
	wire _w21662_ ;
	wire _w21663_ ;
	wire _w21664_ ;
	wire _w21665_ ;
	wire _w21666_ ;
	wire _w21667_ ;
	wire _w21668_ ;
	wire _w21669_ ;
	wire _w21670_ ;
	wire _w21671_ ;
	wire _w21672_ ;
	wire _w21673_ ;
	wire _w21674_ ;
	wire _w21675_ ;
	wire _w21676_ ;
	wire _w21677_ ;
	wire _w21678_ ;
	wire _w21679_ ;
	wire _w21680_ ;
	wire _w21681_ ;
	wire _w21682_ ;
	wire _w21683_ ;
	wire _w21684_ ;
	wire _w21685_ ;
	wire _w21686_ ;
	wire _w21687_ ;
	wire _w21688_ ;
	wire _w21689_ ;
	wire _w21690_ ;
	wire _w21691_ ;
	wire _w21692_ ;
	wire _w21693_ ;
	wire _w21694_ ;
	wire _w21695_ ;
	wire _w21696_ ;
	wire _w21697_ ;
	wire _w21698_ ;
	wire _w21699_ ;
	wire _w21700_ ;
	wire _w21701_ ;
	wire _w21702_ ;
	wire _w21703_ ;
	wire _w21704_ ;
	wire _w21705_ ;
	wire _w21706_ ;
	wire _w21707_ ;
	wire _w21708_ ;
	wire _w21709_ ;
	wire _w21710_ ;
	wire _w21711_ ;
	wire _w21712_ ;
	wire _w21713_ ;
	wire _w21714_ ;
	wire _w21715_ ;
	wire _w21716_ ;
	wire _w21717_ ;
	wire _w21718_ ;
	wire _w21719_ ;
	wire _w21720_ ;
	wire _w21721_ ;
	wire _w21722_ ;
	wire _w21723_ ;
	wire _w21724_ ;
	wire _w21725_ ;
	wire _w21726_ ;
	wire _w21727_ ;
	wire _w21728_ ;
	wire _w21729_ ;
	wire _w21730_ ;
	wire _w21731_ ;
	wire _w21732_ ;
	wire _w21733_ ;
	wire _w21734_ ;
	wire _w21735_ ;
	wire _w21736_ ;
	wire _w21737_ ;
	wire _w21738_ ;
	wire _w21739_ ;
	wire _w21740_ ;
	wire _w21741_ ;
	wire _w21742_ ;
	wire _w21743_ ;
	wire _w21744_ ;
	wire _w21745_ ;
	wire _w21746_ ;
	wire _w21747_ ;
	wire _w21748_ ;
	wire _w21749_ ;
	wire _w21750_ ;
	wire _w21751_ ;
	wire _w21752_ ;
	wire _w21753_ ;
	wire _w21754_ ;
	wire _w21755_ ;
	wire _w21756_ ;
	wire _w21757_ ;
	wire _w21758_ ;
	wire _w21759_ ;
	wire _w21760_ ;
	wire _w21761_ ;
	wire _w21762_ ;
	wire _w21763_ ;
	wire _w21764_ ;
	wire _w21765_ ;
	wire _w21766_ ;
	wire _w21767_ ;
	wire _w21768_ ;
	wire _w21769_ ;
	wire _w21770_ ;
	wire _w21771_ ;
	wire _w21772_ ;
	wire _w21773_ ;
	wire _w21774_ ;
	wire _w21775_ ;
	wire _w21776_ ;
	wire _w21777_ ;
	wire _w21778_ ;
	wire _w21779_ ;
	wire _w21780_ ;
	wire _w21781_ ;
	wire _w21782_ ;
	wire _w21783_ ;
	wire _w21784_ ;
	wire _w21785_ ;
	wire _w21786_ ;
	wire _w21787_ ;
	wire _w21788_ ;
	wire _w21789_ ;
	wire _w21790_ ;
	wire _w21791_ ;
	wire _w21792_ ;
	wire _w21793_ ;
	wire _w21794_ ;
	wire _w21795_ ;
	wire _w21796_ ;
	wire _w21797_ ;
	wire _w21798_ ;
	wire _w21799_ ;
	wire _w21800_ ;
	wire _w21801_ ;
	wire _w21802_ ;
	wire _w21803_ ;
	wire _w21804_ ;
	wire _w21805_ ;
	wire _w21806_ ;
	wire _w21807_ ;
	wire _w21808_ ;
	wire _w21809_ ;
	wire _w21810_ ;
	wire _w21811_ ;
	wire _w21812_ ;
	wire _w21813_ ;
	wire _w21814_ ;
	wire _w21815_ ;
	wire _w21816_ ;
	wire _w21817_ ;
	wire _w21818_ ;
	wire _w21819_ ;
	wire _w21820_ ;
	wire _w21821_ ;
	wire _w21822_ ;
	wire _w21823_ ;
	wire _w21824_ ;
	wire _w21825_ ;
	wire _w21826_ ;
	wire _w21827_ ;
	wire _w21828_ ;
	wire _w21829_ ;
	wire _w21830_ ;
	wire _w21831_ ;
	wire _w21832_ ;
	wire _w21833_ ;
	wire _w21834_ ;
	wire _w21835_ ;
	wire _w21836_ ;
	wire _w21837_ ;
	wire _w21838_ ;
	wire _w21839_ ;
	wire _w21840_ ;
	wire _w21841_ ;
	wire _w21842_ ;
	wire _w21843_ ;
	wire _w21844_ ;
	wire _w21845_ ;
	wire _w21846_ ;
	wire _w21847_ ;
	wire _w21848_ ;
	wire _w21849_ ;
	wire _w21850_ ;
	wire _w21851_ ;
	wire _w21852_ ;
	wire _w21853_ ;
	wire _w21854_ ;
	wire _w21855_ ;
	wire _w21856_ ;
	wire _w21857_ ;
	wire _w21858_ ;
	wire _w21859_ ;
	wire _w21860_ ;
	wire _w21861_ ;
	wire _w21862_ ;
	wire _w21863_ ;
	wire _w21864_ ;
	wire _w21865_ ;
	wire _w21866_ ;
	wire _w21867_ ;
	wire _w21868_ ;
	wire _w21869_ ;
	wire _w21870_ ;
	wire _w21871_ ;
	wire _w21872_ ;
	wire _w21873_ ;
	wire _w21874_ ;
	wire _w21875_ ;
	wire _w21876_ ;
	wire _w21877_ ;
	wire _w21878_ ;
	wire _w21879_ ;
	wire _w21880_ ;
	wire _w21881_ ;
	wire _w21882_ ;
	wire _w21883_ ;
	wire _w21884_ ;
	wire _w21885_ ;
	wire _w21886_ ;
	wire _w21887_ ;
	wire _w21888_ ;
	wire _w21889_ ;
	wire _w21890_ ;
	wire _w21891_ ;
	wire _w21892_ ;
	wire _w21893_ ;
	wire _w21894_ ;
	wire _w21895_ ;
	wire _w21896_ ;
	wire _w21897_ ;
	wire _w21898_ ;
	wire _w21899_ ;
	wire _w21900_ ;
	wire _w21901_ ;
	wire _w21902_ ;
	wire _w21903_ ;
	wire _w21904_ ;
	wire _w21905_ ;
	wire _w21906_ ;
	wire _w21907_ ;
	wire _w21908_ ;
	wire _w21909_ ;
	wire _w21910_ ;
	wire _w21911_ ;
	wire _w21912_ ;
	wire _w21913_ ;
	wire _w21914_ ;
	wire _w21915_ ;
	wire _w21916_ ;
	wire _w21917_ ;
	wire _w21918_ ;
	wire _w21919_ ;
	wire _w21920_ ;
	wire _w21921_ ;
	wire _w21922_ ;
	wire _w21923_ ;
	wire _w21924_ ;
	wire _w21925_ ;
	wire _w21926_ ;
	wire _w21927_ ;
	wire _w21928_ ;
	wire _w21929_ ;
	wire _w21930_ ;
	wire _w21931_ ;
	wire _w21932_ ;
	wire _w21933_ ;
	wire _w21934_ ;
	wire _w21935_ ;
	wire _w21936_ ;
	wire _w21937_ ;
	wire _w21938_ ;
	wire _w21939_ ;
	wire _w21940_ ;
	wire _w21941_ ;
	wire _w21942_ ;
	wire _w21943_ ;
	wire _w21944_ ;
	wire _w21945_ ;
	wire _w21946_ ;
	wire _w21947_ ;
	wire _w21948_ ;
	wire _w21949_ ;
	wire _w21950_ ;
	wire _w21951_ ;
	wire _w21952_ ;
	wire _w21953_ ;
	wire _w21954_ ;
	wire _w21955_ ;
	wire _w21956_ ;
	wire _w21957_ ;
	wire _w21958_ ;
	wire _w21959_ ;
	wire _w21960_ ;
	wire _w21961_ ;
	wire _w21962_ ;
	wire _w21963_ ;
	wire _w21964_ ;
	wire _w21965_ ;
	wire _w21966_ ;
	wire _w21967_ ;
	wire _w21968_ ;
	wire _w21969_ ;
	wire _w21970_ ;
	wire _w21971_ ;
	wire _w21972_ ;
	wire _w21973_ ;
	wire _w21974_ ;
	wire _w21975_ ;
	wire _w21976_ ;
	wire _w21977_ ;
	wire _w21978_ ;
	wire _w21979_ ;
	wire _w21980_ ;
	wire _w21981_ ;
	wire _w21982_ ;
	wire _w21983_ ;
	wire _w21984_ ;
	wire _w21985_ ;
	wire _w21986_ ;
	wire _w21987_ ;
	wire _w21988_ ;
	wire _w21989_ ;
	wire _w21990_ ;
	wire _w21991_ ;
	wire _w21992_ ;
	wire _w21993_ ;
	wire _w21994_ ;
	wire _w21995_ ;
	wire _w21996_ ;
	wire _w21997_ ;
	wire _w21998_ ;
	wire _w21999_ ;
	wire _w22000_ ;
	wire _w22001_ ;
	wire _w22002_ ;
	wire _w22003_ ;
	wire _w22004_ ;
	wire _w22005_ ;
	wire _w22006_ ;
	wire _w22007_ ;
	wire _w22008_ ;
	wire _w22009_ ;
	wire _w22010_ ;
	wire _w22011_ ;
	wire _w22012_ ;
	wire _w22013_ ;
	wire _w22014_ ;
	wire _w22015_ ;
	wire _w22016_ ;
	wire _w22017_ ;
	wire _w22018_ ;
	wire _w22019_ ;
	wire _w22020_ ;
	wire _w22021_ ;
	wire _w22022_ ;
	wire _w22023_ ;
	wire _w22024_ ;
	wire _w22025_ ;
	wire _w22026_ ;
	wire _w22027_ ;
	wire _w22028_ ;
	wire _w22029_ ;
	wire _w22030_ ;
	wire _w22031_ ;
	wire _w22032_ ;
	wire _w22033_ ;
	wire _w22034_ ;
	wire _w22035_ ;
	wire _w22036_ ;
	wire _w22037_ ;
	wire _w22038_ ;
	wire _w22039_ ;
	wire _w22040_ ;
	wire _w22041_ ;
	wire _w22042_ ;
	wire _w22043_ ;
	wire _w22044_ ;
	wire _w22045_ ;
	wire _w22046_ ;
	wire _w22047_ ;
	wire _w22048_ ;
	wire _w22049_ ;
	wire _w22050_ ;
	wire _w22051_ ;
	wire _w22052_ ;
	wire _w22053_ ;
	wire _w22054_ ;
	wire _w22055_ ;
	wire _w22056_ ;
	wire _w22057_ ;
	wire _w22058_ ;
	wire _w22059_ ;
	wire _w22060_ ;
	wire _w22061_ ;
	wire _w22062_ ;
	wire _w22063_ ;
	wire _w22064_ ;
	wire _w22065_ ;
	wire _w22066_ ;
	wire _w22067_ ;
	wire _w22068_ ;
	wire _w22069_ ;
	wire _w22070_ ;
	wire _w22071_ ;
	wire _w22072_ ;
	wire _w22073_ ;
	wire _w22074_ ;
	wire _w22075_ ;
	wire _w22076_ ;
	wire _w22077_ ;
	wire _w22078_ ;
	wire _w22079_ ;
	wire _w22080_ ;
	wire _w22081_ ;
	wire _w22082_ ;
	wire _w22083_ ;
	wire _w22084_ ;
	wire _w22085_ ;
	wire _w22086_ ;
	wire _w22087_ ;
	wire _w22088_ ;
	wire _w22089_ ;
	wire _w22090_ ;
	wire _w22091_ ;
	wire _w22092_ ;
	wire _w22093_ ;
	wire _w22094_ ;
	wire _w22095_ ;
	wire _w22096_ ;
	wire _w22097_ ;
	wire _w22098_ ;
	wire _w22099_ ;
	wire _w22100_ ;
	wire _w22101_ ;
	wire _w22102_ ;
	wire _w22103_ ;
	wire _w22104_ ;
	wire _w22105_ ;
	wire _w22106_ ;
	wire _w22107_ ;
	wire _w22108_ ;
	wire _w22109_ ;
	wire _w22110_ ;
	wire _w22111_ ;
	wire _w22112_ ;
	wire _w22113_ ;
	wire _w22114_ ;
	wire _w22115_ ;
	wire _w22116_ ;
	wire _w22117_ ;
	wire _w22118_ ;
	wire _w22119_ ;
	wire _w22120_ ;
	wire _w22121_ ;
	wire _w22122_ ;
	wire _w22123_ ;
	wire _w22124_ ;
	wire _w22125_ ;
	wire _w22126_ ;
	wire _w22127_ ;
	wire _w22128_ ;
	wire _w22129_ ;
	wire _w22130_ ;
	wire _w22131_ ;
	wire _w22132_ ;
	wire _w22133_ ;
	wire _w22134_ ;
	wire _w22135_ ;
	wire _w22136_ ;
	wire _w22137_ ;
	wire _w22138_ ;
	wire _w22139_ ;
	wire _w22140_ ;
	wire _w22141_ ;
	wire _w22142_ ;
	wire _w22143_ ;
	wire _w22144_ ;
	wire _w22145_ ;
	wire _w22146_ ;
	wire _w22147_ ;
	wire _w22148_ ;
	wire _w22149_ ;
	wire _w22150_ ;
	wire _w22151_ ;
	wire _w22152_ ;
	wire _w22153_ ;
	wire _w22154_ ;
	wire _w22155_ ;
	wire _w22156_ ;
	wire _w22157_ ;
	wire _w22158_ ;
	wire _w22159_ ;
	wire _w22160_ ;
	wire _w22161_ ;
	wire _w22162_ ;
	wire _w22163_ ;
	wire _w22164_ ;
	wire _w22165_ ;
	wire _w22166_ ;
	wire _w22167_ ;
	wire _w22168_ ;
	wire _w22169_ ;
	wire _w22170_ ;
	wire _w22171_ ;
	wire _w22172_ ;
	wire _w22173_ ;
	wire _w22174_ ;
	wire _w22175_ ;
	wire _w22176_ ;
	wire _w22177_ ;
	wire _w22178_ ;
	wire _w22179_ ;
	wire _w22180_ ;
	wire _w22181_ ;
	wire _w22182_ ;
	wire _w22183_ ;
	wire _w22184_ ;
	wire _w22185_ ;
	wire _w22186_ ;
	wire _w22187_ ;
	wire _w22188_ ;
	wire _w22189_ ;
	wire _w22190_ ;
	wire _w22191_ ;
	wire _w22192_ ;
	wire _w22193_ ;
	wire _w22194_ ;
	wire _w22195_ ;
	wire _w22196_ ;
	wire _w22197_ ;
	wire _w22198_ ;
	wire _w22199_ ;
	wire _w22200_ ;
	wire _w22201_ ;
	wire _w22202_ ;
	wire _w22203_ ;
	wire _w22204_ ;
	wire _w22205_ ;
	wire _w22206_ ;
	wire _w22207_ ;
	wire _w22208_ ;
	wire _w22209_ ;
	wire _w22210_ ;
	wire _w22211_ ;
	wire _w22212_ ;
	wire _w22213_ ;
	wire _w22214_ ;
	wire _w22215_ ;
	wire _w22216_ ;
	wire _w22217_ ;
	wire _w22218_ ;
	wire _w22219_ ;
	wire _w22220_ ;
	wire _w22221_ ;
	wire _w22222_ ;
	wire _w22223_ ;
	wire _w22224_ ;
	wire _w22225_ ;
	wire _w22226_ ;
	wire _w22227_ ;
	wire _w22228_ ;
	wire _w22229_ ;
	wire _w22230_ ;
	wire _w22231_ ;
	wire _w22232_ ;
	wire _w22233_ ;
	wire _w22234_ ;
	wire _w22235_ ;
	wire _w22236_ ;
	wire _w22237_ ;
	wire _w22238_ ;
	wire _w22239_ ;
	wire _w22240_ ;
	wire _w22241_ ;
	wire _w22242_ ;
	wire _w22243_ ;
	wire _w22244_ ;
	wire _w22245_ ;
	wire _w22246_ ;
	wire _w22247_ ;
	wire _w22248_ ;
	wire _w22249_ ;
	wire _w22250_ ;
	wire _w22251_ ;
	wire _w22252_ ;
	wire _w22253_ ;
	wire _w22254_ ;
	wire _w22255_ ;
	wire _w22256_ ;
	wire _w22257_ ;
	wire _w22258_ ;
	wire _w22259_ ;
	wire _w22260_ ;
	wire _w22261_ ;
	wire _w22262_ ;
	wire _w22263_ ;
	wire _w22264_ ;
	wire _w22265_ ;
	wire _w22266_ ;
	wire _w22267_ ;
	wire _w22268_ ;
	wire _w22269_ ;
	wire _w22270_ ;
	wire _w22271_ ;
	wire _w22272_ ;
	wire _w22273_ ;
	wire _w22274_ ;
	wire _w22275_ ;
	wire _w22276_ ;
	wire _w22277_ ;
	wire _w22278_ ;
	wire _w22279_ ;
	wire _w22280_ ;
	wire _w22281_ ;
	wire _w22282_ ;
	wire _w22283_ ;
	wire _w22284_ ;
	wire _w22285_ ;
	wire _w22286_ ;
	wire _w22287_ ;
	wire _w22288_ ;
	wire _w22289_ ;
	wire _w22290_ ;
	wire _w22291_ ;
	wire _w22292_ ;
	wire _w22293_ ;
	wire _w22294_ ;
	wire _w22295_ ;
	wire _w22296_ ;
	wire _w22297_ ;
	wire _w22298_ ;
	wire _w22299_ ;
	wire _w22300_ ;
	wire _w22301_ ;
	wire _w22302_ ;
	wire _w22303_ ;
	wire _w22304_ ;
	wire _w22305_ ;
	wire _w22306_ ;
	wire _w22307_ ;
	wire _w22308_ ;
	wire _w22309_ ;
	wire _w22310_ ;
	wire _w22311_ ;
	wire _w22312_ ;
	wire _w22313_ ;
	wire _w22314_ ;
	wire _w22315_ ;
	wire _w22316_ ;
	wire _w22317_ ;
	wire _w22318_ ;
	wire _w22319_ ;
	wire _w22320_ ;
	wire _w22321_ ;
	wire _w22322_ ;
	wire _w22323_ ;
	wire _w22324_ ;
	wire _w22325_ ;
	wire _w22326_ ;
	wire _w22327_ ;
	wire _w22328_ ;
	wire _w22329_ ;
	wire _w22330_ ;
	wire _w22331_ ;
	wire _w22332_ ;
	wire _w22333_ ;
	wire _w22334_ ;
	wire _w22335_ ;
	wire _w22336_ ;
	wire _w22337_ ;
	wire _w22338_ ;
	wire _w22339_ ;
	wire _w22340_ ;
	wire _w22341_ ;
	wire _w22342_ ;
	wire _w22343_ ;
	wire _w22344_ ;
	wire _w22345_ ;
	wire _w22346_ ;
	wire _w22347_ ;
	wire _w22348_ ;
	wire _w22349_ ;
	wire _w22350_ ;
	wire _w22351_ ;
	wire _w22352_ ;
	wire _w22353_ ;
	wire _w22354_ ;
	wire _w22355_ ;
	wire _w22356_ ;
	wire _w22357_ ;
	wire _w22358_ ;
	wire _w22359_ ;
	wire _w22360_ ;
	wire _w22361_ ;
	wire _w22362_ ;
	wire _w22363_ ;
	wire _w22364_ ;
	wire _w22365_ ;
	wire _w22366_ ;
	wire _w22367_ ;
	wire _w22368_ ;
	wire _w22369_ ;
	wire _w22370_ ;
	wire _w22371_ ;
	wire _w22372_ ;
	wire _w22373_ ;
	wire _w22374_ ;
	wire _w22375_ ;
	wire _w22376_ ;
	wire _w22377_ ;
	wire _w22378_ ;
	wire _w22379_ ;
	wire _w22380_ ;
	wire _w22381_ ;
	wire _w22382_ ;
	wire _w22383_ ;
	wire _w22384_ ;
	wire _w22385_ ;
	wire _w22386_ ;
	wire _w22387_ ;
	wire _w22388_ ;
	wire _w22389_ ;
	wire _w22390_ ;
	wire _w22391_ ;
	wire _w22392_ ;
	wire _w22393_ ;
	wire _w22394_ ;
	wire _w22395_ ;
	wire _w22396_ ;
	wire _w22397_ ;
	wire _w22398_ ;
	wire _w22399_ ;
	wire _w22400_ ;
	wire _w22401_ ;
	wire _w22402_ ;
	wire _w22403_ ;
	wire _w22404_ ;
	wire _w22405_ ;
	wire _w22406_ ;
	wire _w22407_ ;
	wire _w22408_ ;
	wire _w22409_ ;
	wire _w22410_ ;
	wire _w22411_ ;
	wire _w22412_ ;
	wire _w22413_ ;
	wire _w22414_ ;
	wire _w22415_ ;
	wire _w22416_ ;
	wire _w22417_ ;
	wire _w22418_ ;
	wire _w22419_ ;
	wire _w22420_ ;
	wire _w22421_ ;
	wire _w22422_ ;
	wire _w22423_ ;
	wire _w22424_ ;
	wire _w22425_ ;
	wire _w22426_ ;
	wire _w22427_ ;
	wire _w22428_ ;
	wire _w22429_ ;
	wire _w22430_ ;
	wire _w22431_ ;
	wire _w22432_ ;
	wire _w22433_ ;
	wire _w22434_ ;
	wire _w22435_ ;
	wire _w22436_ ;
	wire _w22437_ ;
	wire _w22438_ ;
	wire _w22439_ ;
	wire _w22440_ ;
	wire _w22441_ ;
	wire _w22442_ ;
	wire _w22443_ ;
	wire _w22444_ ;
	wire _w22445_ ;
	wire _w22446_ ;
	wire _w22447_ ;
	wire _w22448_ ;
	wire _w22449_ ;
	wire _w22450_ ;
	wire _w22451_ ;
	wire _w22452_ ;
	wire _w22453_ ;
	wire _w22454_ ;
	wire _w22455_ ;
	wire _w22456_ ;
	wire _w22457_ ;
	wire _w22458_ ;
	wire _w22459_ ;
	wire _w22460_ ;
	wire _w22461_ ;
	wire _w22462_ ;
	wire _w22463_ ;
	wire _w22464_ ;
	wire _w22465_ ;
	wire _w22466_ ;
	wire _w22467_ ;
	wire _w22468_ ;
	wire _w22469_ ;
	wire _w22470_ ;
	wire _w22471_ ;
	wire _w22472_ ;
	wire _w22473_ ;
	wire _w22474_ ;
	wire _w22475_ ;
	wire _w22476_ ;
	wire _w22477_ ;
	wire _w22478_ ;
	wire _w22479_ ;
	wire _w22480_ ;
	wire _w22481_ ;
	wire _w22482_ ;
	wire _w22483_ ;
	wire _w22484_ ;
	wire _w22485_ ;
	wire _w22486_ ;
	wire _w22487_ ;
	wire _w22488_ ;
	wire _w22489_ ;
	wire _w22490_ ;
	wire _w22491_ ;
	wire _w22492_ ;
	wire _w22493_ ;
	wire _w22494_ ;
	wire _w22495_ ;
	wire _w22496_ ;
	wire _w22497_ ;
	wire _w22498_ ;
	wire _w22499_ ;
	wire _w22500_ ;
	wire _w22501_ ;
	wire _w22502_ ;
	wire _w22503_ ;
	wire _w22504_ ;
	wire _w22505_ ;
	wire _w22506_ ;
	wire _w22507_ ;
	wire _w22508_ ;
	wire _w22509_ ;
	wire _w22510_ ;
	wire _w22511_ ;
	wire _w22512_ ;
	wire _w22513_ ;
	wire _w22514_ ;
	wire _w22515_ ;
	wire _w22516_ ;
	wire _w22517_ ;
	wire _w22518_ ;
	wire _w22519_ ;
	wire _w22520_ ;
	wire _w22521_ ;
	wire _w22522_ ;
	wire _w22523_ ;
	wire _w22524_ ;
	wire _w22525_ ;
	wire _w22526_ ;
	wire _w22527_ ;
	wire _w22528_ ;
	wire _w22529_ ;
	wire _w22530_ ;
	wire _w22531_ ;
	wire _w22532_ ;
	wire _w22533_ ;
	wire _w22534_ ;
	wire _w22535_ ;
	wire _w22536_ ;
	wire _w22537_ ;
	wire _w22538_ ;
	wire _w22539_ ;
	wire _w22540_ ;
	wire _w22541_ ;
	wire _w22542_ ;
	wire _w22543_ ;
	wire _w22544_ ;
	wire _w22545_ ;
	wire _w22546_ ;
	wire _w22547_ ;
	wire _w22548_ ;
	wire _w22549_ ;
	wire _w22550_ ;
	wire _w22551_ ;
	wire _w22552_ ;
	wire _w22553_ ;
	wire _w22554_ ;
	wire _w22555_ ;
	wire _w22556_ ;
	wire _w22557_ ;
	wire _w22558_ ;
	wire _w22559_ ;
	wire _w22560_ ;
	wire _w22561_ ;
	wire _w22562_ ;
	wire _w22563_ ;
	wire _w22564_ ;
	wire _w22565_ ;
	wire _w22566_ ;
	wire _w22567_ ;
	wire _w22568_ ;
	wire _w22569_ ;
	wire _w22570_ ;
	wire _w22571_ ;
	wire _w22572_ ;
	wire _w22573_ ;
	wire _w22574_ ;
	wire _w22575_ ;
	wire _w22576_ ;
	wire _w22577_ ;
	wire _w22578_ ;
	wire _w22579_ ;
	wire _w22580_ ;
	wire _w22581_ ;
	wire _w22582_ ;
	wire _w22583_ ;
	wire _w22584_ ;
	wire _w22585_ ;
	wire _w22586_ ;
	wire _w22587_ ;
	wire _w22588_ ;
	wire _w22589_ ;
	wire _w22590_ ;
	wire _w22591_ ;
	wire _w22592_ ;
	wire _w22593_ ;
	wire _w22594_ ;
	wire _w22595_ ;
	wire _w22596_ ;
	wire _w22597_ ;
	wire _w22598_ ;
	wire _w22599_ ;
	wire _w22600_ ;
	wire _w22601_ ;
	wire _w22602_ ;
	wire _w22603_ ;
	wire _w22604_ ;
	wire _w22605_ ;
	wire _w22606_ ;
	wire _w22607_ ;
	wire _w22608_ ;
	wire _w22609_ ;
	wire _w22610_ ;
	wire _w22611_ ;
	wire _w22612_ ;
	wire _w22613_ ;
	wire _w22614_ ;
	wire _w22615_ ;
	wire _w22616_ ;
	wire _w22617_ ;
	wire _w22618_ ;
	wire _w22619_ ;
	wire _w22620_ ;
	wire _w22621_ ;
	wire _w22622_ ;
	wire _w22623_ ;
	wire _w22624_ ;
	wire _w22625_ ;
	wire _w22626_ ;
	wire _w22627_ ;
	wire _w22628_ ;
	wire _w22629_ ;
	wire _w22630_ ;
	wire _w22631_ ;
	wire _w22632_ ;
	wire _w22633_ ;
	wire _w22634_ ;
	wire _w22635_ ;
	wire _w22636_ ;
	wire _w22637_ ;
	wire _w22638_ ;
	wire _w22639_ ;
	wire _w22640_ ;
	wire _w22641_ ;
	wire _w22642_ ;
	wire _w22643_ ;
	wire _w22644_ ;
	wire _w22645_ ;
	wire _w22646_ ;
	wire _w22647_ ;
	wire _w22648_ ;
	wire _w22649_ ;
	wire _w22650_ ;
	wire _w22651_ ;
	wire _w22652_ ;
	wire _w22653_ ;
	wire _w22654_ ;
	wire _w22655_ ;
	wire _w22656_ ;
	wire _w22657_ ;
	wire _w22658_ ;
	wire _w22659_ ;
	wire _w22660_ ;
	wire _w22661_ ;
	wire _w22662_ ;
	wire _w22663_ ;
	wire _w22664_ ;
	wire _w22665_ ;
	wire _w22666_ ;
	wire _w22667_ ;
	wire _w22668_ ;
	wire _w22669_ ;
	wire _w22670_ ;
	wire _w22671_ ;
	wire _w22672_ ;
	wire _w22673_ ;
	wire _w22674_ ;
	wire _w22675_ ;
	wire _w22676_ ;
	wire _w22677_ ;
	wire _w22678_ ;
	wire _w22679_ ;
	wire _w22680_ ;
	wire _w22681_ ;
	wire _w22682_ ;
	wire _w22683_ ;
	wire _w22684_ ;
	wire _w22685_ ;
	wire _w22686_ ;
	wire _w22687_ ;
	wire _w22688_ ;
	wire _w22689_ ;
	wire _w22690_ ;
	wire _w22691_ ;
	wire _w22692_ ;
	wire _w22693_ ;
	wire _w22694_ ;
	wire _w22695_ ;
	wire _w22696_ ;
	wire _w22697_ ;
	wire _w22698_ ;
	wire _w22699_ ;
	wire _w22700_ ;
	wire _w22701_ ;
	wire _w22702_ ;
	wire _w22703_ ;
	wire _w22704_ ;
	wire _w22705_ ;
	wire _w22706_ ;
	wire _w22707_ ;
	wire _w22708_ ;
	wire _w22709_ ;
	wire _w22710_ ;
	wire _w22711_ ;
	wire _w22712_ ;
	wire _w22713_ ;
	wire _w22714_ ;
	wire _w22715_ ;
	wire _w22716_ ;
	wire _w22717_ ;
	wire _w22718_ ;
	wire _w22719_ ;
	wire _w22720_ ;
	wire _w22721_ ;
	wire _w22722_ ;
	wire _w22723_ ;
	wire _w22724_ ;
	wire _w22725_ ;
	wire _w22726_ ;
	wire _w22727_ ;
	wire _w22728_ ;
	wire _w22729_ ;
	wire _w22730_ ;
	wire _w22731_ ;
	wire _w22732_ ;
	wire _w22733_ ;
	wire _w22734_ ;
	wire _w22735_ ;
	wire _w22736_ ;
	wire _w22737_ ;
	wire _w22738_ ;
	wire _w22739_ ;
	wire _w22740_ ;
	wire _w22741_ ;
	wire _w22742_ ;
	wire _w22743_ ;
	wire _w22744_ ;
	wire _w22745_ ;
	wire _w22746_ ;
	wire _w22747_ ;
	wire _w22748_ ;
	wire _w22749_ ;
	wire _w22750_ ;
	wire _w22751_ ;
	wire _w22752_ ;
	wire _w22753_ ;
	wire _w22754_ ;
	wire _w22755_ ;
	wire _w22756_ ;
	wire _w22757_ ;
	wire _w22758_ ;
	wire _w22759_ ;
	wire _w22760_ ;
	wire _w22761_ ;
	wire _w22762_ ;
	wire _w22763_ ;
	wire _w22764_ ;
	wire _w22765_ ;
	wire _w22766_ ;
	wire _w22767_ ;
	wire _w22768_ ;
	wire _w22769_ ;
	wire _w22770_ ;
	wire _w22771_ ;
	wire _w22772_ ;
	wire _w22773_ ;
	wire _w22774_ ;
	wire _w22775_ ;
	wire _w22776_ ;
	wire _w22777_ ;
	wire _w22778_ ;
	wire _w22779_ ;
	wire _w22780_ ;
	wire _w22781_ ;
	wire _w22782_ ;
	wire _w22783_ ;
	wire _w22784_ ;
	wire _w22785_ ;
	wire _w22786_ ;
	wire _w22787_ ;
	wire _w22788_ ;
	wire _w22789_ ;
	wire _w22790_ ;
	wire _w22791_ ;
	wire _w22792_ ;
	wire _w22793_ ;
	wire _w22794_ ;
	wire _w22795_ ;
	wire _w22796_ ;
	wire _w22797_ ;
	wire _w22798_ ;
	wire _w22799_ ;
	wire _w22800_ ;
	wire _w22801_ ;
	wire _w22802_ ;
	wire _w22803_ ;
	wire _w22804_ ;
	wire _w22805_ ;
	wire _w22806_ ;
	wire _w22807_ ;
	wire _w22808_ ;
	wire _w22809_ ;
	wire _w22810_ ;
	wire _w22811_ ;
	wire _w22812_ ;
	wire _w22813_ ;
	wire _w22814_ ;
	wire _w22815_ ;
	wire _w22816_ ;
	wire _w22817_ ;
	wire _w22818_ ;
	wire _w22819_ ;
	wire _w22820_ ;
	wire _w22821_ ;
	wire _w22822_ ;
	wire _w22823_ ;
	wire _w22824_ ;
	wire _w22825_ ;
	wire _w22826_ ;
	wire _w22827_ ;
	wire _w22828_ ;
	wire _w22829_ ;
	wire _w22830_ ;
	wire _w22831_ ;
	wire _w22832_ ;
	wire _w22833_ ;
	wire _w22834_ ;
	wire _w22835_ ;
	wire _w22836_ ;
	wire _w22837_ ;
	wire _w22838_ ;
	wire _w22839_ ;
	wire _w22840_ ;
	wire _w22841_ ;
	wire _w22842_ ;
	wire _w22843_ ;
	wire _w22844_ ;
	wire _w22845_ ;
	wire _w22846_ ;
	wire _w22847_ ;
	wire _w22848_ ;
	wire _w22849_ ;
	wire _w22850_ ;
	wire _w22851_ ;
	wire _w22852_ ;
	wire _w22853_ ;
	wire _w22854_ ;
	wire _w22855_ ;
	wire _w22856_ ;
	wire _w22857_ ;
	wire _w22858_ ;
	wire _w22859_ ;
	wire _w22860_ ;
	wire _w22861_ ;
	wire _w22862_ ;
	wire _w22863_ ;
	wire _w22864_ ;
	wire _w22865_ ;
	wire _w22866_ ;
	wire _w22867_ ;
	wire _w22868_ ;
	wire _w22869_ ;
	wire _w22870_ ;
	wire _w22871_ ;
	wire _w22872_ ;
	wire _w22873_ ;
	wire _w22874_ ;
	wire _w22875_ ;
	wire _w22876_ ;
	wire _w22877_ ;
	wire _w22878_ ;
	wire _w22879_ ;
	wire _w22880_ ;
	wire _w22881_ ;
	wire _w22882_ ;
	wire _w22883_ ;
	wire _w22884_ ;
	wire _w22885_ ;
	wire _w22886_ ;
	wire _w22887_ ;
	wire _w22888_ ;
	wire _w22889_ ;
	wire _w22890_ ;
	wire _w22891_ ;
	wire _w22892_ ;
	wire _w22893_ ;
	wire _w22894_ ;
	wire _w22895_ ;
	wire _w22896_ ;
	wire _w22897_ ;
	wire _w22898_ ;
	wire _w22899_ ;
	wire _w22900_ ;
	wire _w22901_ ;
	wire _w22902_ ;
	wire _w22903_ ;
	wire _w22904_ ;
	wire _w22905_ ;
	wire _w22906_ ;
	wire _w22907_ ;
	wire _w22908_ ;
	wire _w22909_ ;
	wire _w22910_ ;
	wire _w22911_ ;
	wire _w22912_ ;
	wire _w22913_ ;
	wire _w22914_ ;
	wire _w22915_ ;
	wire _w22916_ ;
	wire _w22917_ ;
	wire _w22918_ ;
	wire _w22919_ ;
	wire _w22920_ ;
	wire _w22921_ ;
	wire _w22922_ ;
	wire _w22923_ ;
	wire _w22924_ ;
	wire _w22925_ ;
	wire _w22926_ ;
	wire _w22927_ ;
	wire _w22928_ ;
	wire _w22929_ ;
	wire _w22930_ ;
	wire _w22931_ ;
	wire _w22932_ ;
	wire _w22933_ ;
	wire _w22934_ ;
	wire _w22935_ ;
	wire _w22936_ ;
	wire _w22937_ ;
	wire _w22938_ ;
	wire _w22939_ ;
	wire _w22940_ ;
	wire _w22941_ ;
	wire _w22942_ ;
	wire _w22943_ ;
	wire _w22944_ ;
	wire _w22945_ ;
	wire _w22946_ ;
	wire _w22947_ ;
	wire _w22948_ ;
	wire _w22949_ ;
	wire _w22950_ ;
	wire _w22951_ ;
	wire _w22952_ ;
	wire _w22953_ ;
	wire _w22954_ ;
	wire _w22955_ ;
	wire _w22956_ ;
	wire _w22957_ ;
	wire _w22958_ ;
	wire _w22959_ ;
	wire _w22960_ ;
	wire _w22961_ ;
	wire _w22962_ ;
	wire _w22963_ ;
	wire _w22964_ ;
	wire _w22965_ ;
	wire _w22966_ ;
	wire _w22967_ ;
	wire _w22968_ ;
	wire _w22969_ ;
	wire _w22970_ ;
	wire _w22971_ ;
	wire _w22972_ ;
	wire _w22973_ ;
	wire _w22974_ ;
	wire _w22975_ ;
	wire _w22976_ ;
	wire _w22977_ ;
	wire _w22978_ ;
	wire _w22979_ ;
	wire _w22980_ ;
	wire _w22981_ ;
	wire _w22982_ ;
	wire _w22983_ ;
	wire _w22984_ ;
	wire _w22985_ ;
	wire _w22986_ ;
	wire _w22987_ ;
	wire _w22988_ ;
	wire _w22989_ ;
	wire _w22990_ ;
	wire _w22991_ ;
	wire _w22992_ ;
	wire _w22993_ ;
	wire _w22994_ ;
	wire _w22995_ ;
	wire _w22996_ ;
	wire _w22997_ ;
	wire _w22998_ ;
	wire _w22999_ ;
	wire _w23000_ ;
	wire _w23001_ ;
	wire _w23002_ ;
	wire _w23003_ ;
	wire _w23004_ ;
	wire _w23005_ ;
	wire _w23006_ ;
	wire _w23007_ ;
	wire _w23008_ ;
	wire _w23009_ ;
	wire _w23010_ ;
	wire _w23011_ ;
	wire _w23012_ ;
	wire _w23013_ ;
	wire _w23014_ ;
	wire _w23015_ ;
	wire _w23016_ ;
	wire _w23017_ ;
	wire _w23018_ ;
	wire _w23019_ ;
	wire _w23020_ ;
	wire _w23021_ ;
	wire _w23022_ ;
	wire _w23023_ ;
	wire _w23024_ ;
	wire _w23025_ ;
	wire _w23026_ ;
	wire _w23027_ ;
	wire _w23028_ ;
	wire _w23029_ ;
	wire _w23030_ ;
	wire _w23031_ ;
	wire _w23032_ ;
	wire _w23033_ ;
	wire _w23034_ ;
	wire _w23035_ ;
	wire _w23036_ ;
	wire _w23037_ ;
	wire _w23038_ ;
	wire _w23039_ ;
	wire _w23040_ ;
	wire _w23041_ ;
	wire _w23042_ ;
	wire _w23043_ ;
	wire _w23044_ ;
	wire _w23045_ ;
	wire _w23046_ ;
	wire _w23047_ ;
	wire _w23048_ ;
	wire _w23049_ ;
	wire _w23050_ ;
	wire _w23051_ ;
	wire _w23052_ ;
	wire _w23053_ ;
	wire _w23054_ ;
	wire _w23055_ ;
	wire _w23056_ ;
	wire _w23057_ ;
	wire _w23058_ ;
	wire _w23059_ ;
	wire _w23060_ ;
	wire _w23061_ ;
	wire _w23062_ ;
	wire _w23063_ ;
	wire _w23064_ ;
	wire _w23065_ ;
	wire _w23066_ ;
	wire _w23067_ ;
	wire _w23068_ ;
	wire _w23069_ ;
	wire _w23070_ ;
	wire _w23071_ ;
	wire _w23072_ ;
	wire _w23073_ ;
	wire _w23074_ ;
	wire _w23075_ ;
	wire _w23076_ ;
	wire _w23077_ ;
	wire _w23078_ ;
	wire _w23079_ ;
	wire _w23080_ ;
	wire _w23081_ ;
	wire _w23082_ ;
	wire _w23083_ ;
	wire _w23084_ ;
	wire _w23085_ ;
	wire _w23086_ ;
	wire _w23087_ ;
	wire _w23088_ ;
	wire _w23089_ ;
	wire _w23090_ ;
	wire _w23091_ ;
	wire _w23092_ ;
	wire _w23093_ ;
	wire _w23094_ ;
	wire _w23095_ ;
	wire _w23096_ ;
	wire _w23097_ ;
	wire _w23098_ ;
	wire _w23099_ ;
	wire _w23100_ ;
	wire _w23101_ ;
	wire _w23102_ ;
	wire _w23103_ ;
	wire _w23104_ ;
	wire _w23105_ ;
	wire _w23106_ ;
	wire _w23107_ ;
	wire _w23108_ ;
	wire _w23109_ ;
	wire _w23110_ ;
	wire _w23111_ ;
	wire _w23112_ ;
	wire _w23113_ ;
	wire _w23114_ ;
	wire _w23115_ ;
	wire _w23116_ ;
	wire _w23117_ ;
	wire _w23118_ ;
	wire _w23119_ ;
	wire _w23120_ ;
	wire _w23121_ ;
	wire _w23122_ ;
	wire _w23123_ ;
	wire _w23124_ ;
	wire _w23125_ ;
	wire _w23126_ ;
	wire _w23127_ ;
	wire _w23128_ ;
	wire _w23129_ ;
	wire _w23130_ ;
	wire _w23131_ ;
	wire _w23132_ ;
	wire _w23133_ ;
	wire _w23134_ ;
	wire _w23135_ ;
	wire _w23136_ ;
	wire _w23137_ ;
	wire _w23138_ ;
	wire _w23139_ ;
	wire _w23140_ ;
	wire _w23141_ ;
	wire _w23142_ ;
	wire _w23143_ ;
	wire _w23144_ ;
	wire _w23145_ ;
	wire _w23146_ ;
	wire _w23147_ ;
	wire _w23148_ ;
	wire _w23149_ ;
	wire _w23150_ ;
	wire _w23151_ ;
	wire _w23152_ ;
	wire _w23153_ ;
	wire _w23154_ ;
	wire _w23155_ ;
	wire _w23156_ ;
	wire _w23157_ ;
	wire _w23158_ ;
	wire _w23159_ ;
	wire _w23160_ ;
	wire _w23161_ ;
	wire _w23162_ ;
	wire _w23163_ ;
	wire _w23164_ ;
	wire _w23165_ ;
	wire _w23166_ ;
	wire _w23167_ ;
	wire _w23168_ ;
	wire _w23169_ ;
	wire _w23170_ ;
	wire _w23171_ ;
	wire _w23172_ ;
	wire _w23173_ ;
	wire _w23174_ ;
	wire _w23175_ ;
	wire _w23176_ ;
	wire _w23177_ ;
	wire _w23178_ ;
	wire _w23179_ ;
	wire _w23180_ ;
	wire _w23181_ ;
	wire _w23182_ ;
	wire _w23183_ ;
	wire _w23184_ ;
	wire _w23185_ ;
	wire _w23186_ ;
	wire _w23187_ ;
	wire _w23188_ ;
	wire _w23189_ ;
	wire _w23190_ ;
	wire _w23191_ ;
	wire _w23192_ ;
	wire _w23193_ ;
	wire _w23194_ ;
	wire _w23195_ ;
	wire _w23196_ ;
	wire _w23197_ ;
	wire _w23198_ ;
	wire _w23199_ ;
	wire _w23200_ ;
	wire _w23201_ ;
	wire _w23202_ ;
	wire _w23203_ ;
	wire _w23204_ ;
	wire _w23205_ ;
	wire _w23206_ ;
	wire _w23207_ ;
	wire _w23208_ ;
	wire _w23209_ ;
	wire _w23210_ ;
	wire _w23211_ ;
	wire _w23212_ ;
	wire _w23213_ ;
	wire _w23214_ ;
	wire _w23215_ ;
	wire _w23216_ ;
	wire _w23217_ ;
	wire _w23218_ ;
	wire _w23219_ ;
	wire _w23220_ ;
	wire _w23221_ ;
	wire _w23222_ ;
	wire _w23223_ ;
	wire _w23224_ ;
	wire _w23225_ ;
	wire _w23226_ ;
	wire _w23227_ ;
	wire _w23228_ ;
	wire _w23229_ ;
	wire _w23230_ ;
	wire _w23231_ ;
	wire _w23232_ ;
	wire _w23233_ ;
	wire _w23234_ ;
	wire _w23235_ ;
	wire _w23236_ ;
	wire _w23237_ ;
	wire _w23238_ ;
	wire _w23239_ ;
	wire _w23240_ ;
	wire _w23241_ ;
	wire _w23242_ ;
	wire _w23243_ ;
	wire _w23244_ ;
	wire _w23245_ ;
	wire _w23246_ ;
	wire _w23247_ ;
	wire _w23248_ ;
	wire _w23249_ ;
	wire _w23250_ ;
	wire _w23251_ ;
	wire _w23252_ ;
	wire _w23253_ ;
	wire _w23254_ ;
	wire _w23255_ ;
	wire _w23256_ ;
	wire _w23257_ ;
	wire _w23258_ ;
	wire _w23259_ ;
	wire _w23260_ ;
	wire _w23261_ ;
	wire _w23262_ ;
	wire _w23263_ ;
	wire _w23264_ ;
	wire _w23265_ ;
	wire _w23266_ ;
	wire _w23267_ ;
	wire _w23268_ ;
	wire _w23269_ ;
	wire _w23270_ ;
	wire _w23271_ ;
	wire _w23272_ ;
	wire _w23273_ ;
	wire _w23274_ ;
	wire _w23275_ ;
	wire _w23276_ ;
	wire _w23277_ ;
	wire _w23278_ ;
	wire _w23279_ ;
	wire _w23280_ ;
	wire _w23281_ ;
	wire _w23282_ ;
	wire _w23283_ ;
	wire _w23284_ ;
	wire _w23285_ ;
	wire _w23286_ ;
	wire _w23287_ ;
	wire _w23288_ ;
	wire _w23289_ ;
	wire _w23290_ ;
	wire _w23291_ ;
	wire _w23292_ ;
	wire _w23293_ ;
	wire _w23294_ ;
	wire _w23295_ ;
	wire _w23296_ ;
	wire _w23297_ ;
	wire _w23298_ ;
	wire _w23299_ ;
	wire _w23300_ ;
	wire _w23301_ ;
	wire _w23302_ ;
	wire _w23303_ ;
	wire _w23304_ ;
	wire _w23305_ ;
	wire _w23306_ ;
	wire _w23307_ ;
	wire _w23308_ ;
	wire _w23309_ ;
	wire _w23310_ ;
	wire _w23311_ ;
	wire _w23312_ ;
	wire _w23313_ ;
	wire _w23314_ ;
	wire _w23315_ ;
	wire _w23316_ ;
	wire _w23317_ ;
	wire _w23318_ ;
	wire _w23319_ ;
	wire _w23320_ ;
	wire _w23321_ ;
	wire _w23322_ ;
	wire _w23323_ ;
	wire _w23324_ ;
	wire _w23325_ ;
	wire _w23326_ ;
	wire _w23327_ ;
	wire _w23328_ ;
	wire _w23329_ ;
	wire _w23330_ ;
	wire _w23331_ ;
	wire _w23332_ ;
	wire _w23333_ ;
	wire _w23334_ ;
	wire _w23335_ ;
	wire _w23336_ ;
	wire _w23337_ ;
	wire _w23338_ ;
	wire _w23339_ ;
	wire _w23340_ ;
	wire _w23341_ ;
	wire _w23342_ ;
	wire _w23343_ ;
	wire _w23344_ ;
	wire _w23345_ ;
	wire _w23346_ ;
	wire _w23347_ ;
	wire _w23348_ ;
	wire _w23349_ ;
	wire _w23350_ ;
	wire _w23351_ ;
	wire _w23352_ ;
	wire _w23353_ ;
	wire _w23354_ ;
	wire _w23355_ ;
	wire _w23356_ ;
	wire _w23357_ ;
	wire _w23358_ ;
	wire _w23359_ ;
	wire _w23360_ ;
	wire _w23361_ ;
	wire _w23362_ ;
	wire _w23363_ ;
	wire _w23364_ ;
	wire _w23365_ ;
	wire _w23366_ ;
	wire _w23367_ ;
	wire _w23368_ ;
	wire _w23369_ ;
	wire _w23370_ ;
	wire _w23371_ ;
	wire _w23372_ ;
	wire _w23373_ ;
	wire _w23374_ ;
	wire _w23375_ ;
	wire _w23376_ ;
	wire _w23377_ ;
	wire _w23378_ ;
	wire _w23379_ ;
	wire _w23380_ ;
	wire _w23381_ ;
	wire _w23382_ ;
	wire _w23383_ ;
	wire _w23384_ ;
	wire _w23385_ ;
	wire _w23386_ ;
	wire _w23387_ ;
	wire _w23388_ ;
	wire _w23389_ ;
	wire _w23390_ ;
	wire _w23391_ ;
	wire _w23392_ ;
	wire _w23393_ ;
	wire _w23394_ ;
	wire _w23395_ ;
	wire _w23396_ ;
	wire _w23397_ ;
	wire _w23398_ ;
	wire _w23399_ ;
	wire _w23400_ ;
	wire _w23401_ ;
	wire _w23402_ ;
	wire _w23403_ ;
	wire _w23404_ ;
	wire _w23405_ ;
	wire _w23406_ ;
	wire _w23407_ ;
	wire _w23408_ ;
	wire _w23409_ ;
	wire _w23410_ ;
	wire _w23411_ ;
	wire _w23412_ ;
	wire _w23413_ ;
	wire _w23414_ ;
	wire _w23415_ ;
	wire _w23416_ ;
	wire _w23417_ ;
	wire _w23418_ ;
	wire _w23419_ ;
	wire _w23420_ ;
	wire _w23421_ ;
	wire _w23422_ ;
	wire _w23423_ ;
	wire _w23424_ ;
	wire _w23425_ ;
	wire _w23426_ ;
	wire _w23427_ ;
	wire _w23428_ ;
	wire _w23429_ ;
	wire _w23430_ ;
	wire _w23431_ ;
	wire _w23432_ ;
	wire _w23433_ ;
	wire _w23434_ ;
	wire _w23435_ ;
	wire _w23436_ ;
	wire _w23437_ ;
	wire _w23438_ ;
	wire _w23439_ ;
	wire _w23440_ ;
	wire _w23441_ ;
	wire _w23442_ ;
	wire _w23443_ ;
	wire _w23444_ ;
	wire _w23445_ ;
	wire _w23446_ ;
	wire _w23447_ ;
	wire _w23448_ ;
	wire _w23449_ ;
	wire _w23450_ ;
	wire _w23451_ ;
	wire _w23452_ ;
	wire _w23453_ ;
	wire _w23454_ ;
	wire _w23455_ ;
	wire _w23456_ ;
	wire _w23457_ ;
	wire _w23458_ ;
	wire _w23459_ ;
	wire _w23460_ ;
	wire _w23461_ ;
	wire _w23462_ ;
	wire _w23463_ ;
	wire _w23464_ ;
	wire _w23465_ ;
	wire _w23466_ ;
	wire _w23467_ ;
	wire _w23468_ ;
	wire _w23469_ ;
	wire _w23470_ ;
	wire _w23471_ ;
	wire _w23472_ ;
	wire _w23473_ ;
	wire _w23474_ ;
	wire _w23475_ ;
	wire _w23476_ ;
	wire _w23477_ ;
	wire _w23478_ ;
	wire _w23479_ ;
	wire _w23480_ ;
	wire _w23481_ ;
	wire _w23482_ ;
	wire _w23483_ ;
	wire _w23484_ ;
	wire _w23485_ ;
	wire _w23486_ ;
	wire _w23487_ ;
	wire _w23488_ ;
	wire _w23489_ ;
	wire _w23490_ ;
	wire _w23491_ ;
	wire _w23492_ ;
	wire _w23493_ ;
	wire _w23494_ ;
	wire _w23495_ ;
	wire _w23496_ ;
	wire _w23497_ ;
	wire _w23498_ ;
	wire _w23499_ ;
	wire _w23500_ ;
	wire _w23501_ ;
	wire _w23502_ ;
	wire _w23503_ ;
	wire _w23504_ ;
	wire _w23505_ ;
	wire _w23506_ ;
	wire _w23507_ ;
	wire _w23508_ ;
	wire _w23509_ ;
	wire _w23510_ ;
	wire _w23511_ ;
	wire _w23512_ ;
	wire _w23513_ ;
	wire _w23514_ ;
	wire _w23515_ ;
	wire _w23516_ ;
	wire _w23517_ ;
	wire _w23518_ ;
	wire _w23519_ ;
	wire _w23520_ ;
	wire _w23521_ ;
	wire _w23522_ ;
	wire _w23523_ ;
	wire _w23524_ ;
	wire _w23525_ ;
	wire _w23526_ ;
	wire _w23527_ ;
	wire _w23528_ ;
	wire _w23529_ ;
	wire _w23530_ ;
	wire _w23531_ ;
	wire _w23532_ ;
	wire _w23533_ ;
	wire _w23534_ ;
	wire _w23535_ ;
	wire _w23536_ ;
	wire _w23537_ ;
	wire _w23538_ ;
	wire _w23539_ ;
	wire _w23540_ ;
	wire _w23541_ ;
	wire _w23542_ ;
	wire _w23543_ ;
	wire _w23544_ ;
	wire _w23545_ ;
	wire _w23546_ ;
	wire _w23547_ ;
	wire _w23548_ ;
	wire _w23549_ ;
	wire _w23550_ ;
	wire _w23551_ ;
	wire _w23552_ ;
	wire _w23553_ ;
	wire _w23554_ ;
	wire _w23555_ ;
	wire _w23556_ ;
	wire _w23557_ ;
	wire _w23558_ ;
	wire _w23559_ ;
	wire _w23560_ ;
	wire _w23561_ ;
	wire _w23562_ ;
	wire _w23563_ ;
	wire _w23564_ ;
	wire _w23565_ ;
	wire _w23566_ ;
	wire _w23567_ ;
	wire _w23568_ ;
	wire _w23569_ ;
	wire _w23570_ ;
	wire _w23571_ ;
	wire _w23572_ ;
	wire _w23573_ ;
	wire _w23574_ ;
	wire _w23575_ ;
	wire _w23576_ ;
	wire _w23577_ ;
	wire _w23578_ ;
	wire _w23579_ ;
	wire _w23580_ ;
	wire _w23581_ ;
	wire _w23582_ ;
	wire _w23583_ ;
	wire _w23584_ ;
	wire _w23585_ ;
	wire _w23586_ ;
	wire _w23587_ ;
	wire _w23588_ ;
	wire _w23589_ ;
	wire _w23590_ ;
	wire _w23591_ ;
	wire _w23592_ ;
	wire _w23593_ ;
	wire _w23594_ ;
	wire _w23595_ ;
	wire _w23596_ ;
	wire _w23597_ ;
	wire _w23598_ ;
	wire _w23599_ ;
	wire _w23600_ ;
	wire _w23601_ ;
	wire _w23602_ ;
	wire _w23603_ ;
	wire _w23604_ ;
	wire _w23605_ ;
	wire _w23606_ ;
	wire _w23607_ ;
	wire _w23608_ ;
	wire _w23609_ ;
	wire _w23610_ ;
	wire _w23611_ ;
	wire _w23612_ ;
	wire _w23613_ ;
	wire _w23614_ ;
	wire _w23615_ ;
	wire _w23616_ ;
	wire _w23617_ ;
	wire _w23618_ ;
	wire _w23619_ ;
	wire _w23620_ ;
	wire _w23621_ ;
	wire _w23622_ ;
	wire _w23623_ ;
	wire _w23624_ ;
	wire _w23625_ ;
	wire _w23626_ ;
	wire _w23627_ ;
	wire _w23628_ ;
	wire _w23629_ ;
	wire _w23630_ ;
	wire _w23631_ ;
	wire _w23632_ ;
	wire _w23633_ ;
	wire _w23634_ ;
	wire _w23635_ ;
	wire _w23636_ ;
	wire _w23637_ ;
	wire _w23638_ ;
	wire _w23639_ ;
	wire _w23640_ ;
	wire _w23641_ ;
	wire _w23642_ ;
	wire _w23643_ ;
	wire _w23644_ ;
	wire _w23645_ ;
	wire _w23646_ ;
	wire _w23647_ ;
	wire _w23648_ ;
	wire _w23649_ ;
	wire _w23650_ ;
	wire _w23651_ ;
	wire _w23652_ ;
	wire _w23653_ ;
	wire _w23654_ ;
	wire _w23655_ ;
	wire _w23656_ ;
	wire _w23657_ ;
	wire _w23658_ ;
	wire _w23659_ ;
	wire _w23660_ ;
	wire _w23661_ ;
	wire _w23662_ ;
	wire _w23663_ ;
	wire _w23664_ ;
	wire _w23665_ ;
	wire _w23666_ ;
	wire _w23667_ ;
	wire _w23668_ ;
	wire _w23669_ ;
	wire _w23670_ ;
	wire _w23671_ ;
	wire _w23672_ ;
	wire _w23673_ ;
	wire _w23674_ ;
	wire _w23675_ ;
	wire _w23676_ ;
	wire _w23677_ ;
	wire _w23678_ ;
	wire _w23679_ ;
	wire _w23680_ ;
	wire _w23681_ ;
	wire _w23682_ ;
	wire _w23683_ ;
	wire _w23684_ ;
	wire _w23685_ ;
	wire _w23686_ ;
	wire _w23687_ ;
	wire _w23688_ ;
	wire _w23689_ ;
	wire _w23690_ ;
	wire _w23691_ ;
	wire _w23692_ ;
	wire _w23693_ ;
	wire _w23694_ ;
	wire _w23695_ ;
	wire _w23696_ ;
	wire _w23697_ ;
	wire _w23698_ ;
	wire _w23699_ ;
	wire _w23700_ ;
	wire _w23701_ ;
	wire _w23702_ ;
	wire _w23703_ ;
	wire _w23704_ ;
	wire _w23705_ ;
	wire _w23706_ ;
	wire _w23707_ ;
	wire _w23708_ ;
	wire _w23709_ ;
	wire _w23710_ ;
	wire _w23711_ ;
	wire _w23712_ ;
	wire _w23713_ ;
	wire _w23714_ ;
	wire _w23715_ ;
	wire _w23716_ ;
	wire _w23717_ ;
	wire _w23718_ ;
	wire _w23719_ ;
	wire _w23720_ ;
	wire _w23721_ ;
	wire _w23722_ ;
	wire _w23723_ ;
	wire _w23724_ ;
	wire _w23725_ ;
	wire _w23726_ ;
	wire _w23727_ ;
	wire _w23728_ ;
	wire _w23729_ ;
	wire _w23730_ ;
	wire _w23731_ ;
	wire _w23732_ ;
	wire _w23733_ ;
	wire _w23734_ ;
	wire _w23735_ ;
	wire _w23736_ ;
	wire _w23737_ ;
	wire _w23738_ ;
	wire _w23739_ ;
	wire _w23740_ ;
	wire _w23741_ ;
	wire _w23742_ ;
	wire _w23743_ ;
	wire _w23744_ ;
	wire _w23745_ ;
	wire _w23746_ ;
	wire _w23747_ ;
	wire _w23748_ ;
	wire _w23749_ ;
	wire _w23750_ ;
	wire _w23751_ ;
	wire _w23752_ ;
	wire _w23753_ ;
	wire _w23754_ ;
	wire _w23755_ ;
	wire _w23756_ ;
	wire _w23757_ ;
	wire _w23758_ ;
	wire _w23759_ ;
	wire _w23760_ ;
	wire _w23761_ ;
	wire _w23762_ ;
	wire _w23763_ ;
	wire _w23764_ ;
	wire _w23765_ ;
	wire _w23766_ ;
	wire _w23767_ ;
	wire _w23768_ ;
	wire _w23769_ ;
	wire _w23770_ ;
	wire _w23771_ ;
	wire _w23772_ ;
	wire _w23773_ ;
	wire _w23774_ ;
	wire _w23775_ ;
	wire _w23776_ ;
	wire _w23777_ ;
	wire _w23778_ ;
	wire _w23779_ ;
	wire _w23780_ ;
	wire _w23781_ ;
	wire _w23782_ ;
	wire _w23783_ ;
	wire _w23784_ ;
	wire _w23785_ ;
	wire _w23786_ ;
	wire _w23787_ ;
	wire _w23788_ ;
	wire _w23789_ ;
	wire _w23790_ ;
	wire _w23791_ ;
	wire _w23792_ ;
	wire _w23793_ ;
	wire _w23794_ ;
	wire _w23795_ ;
	wire _w23796_ ;
	wire _w23797_ ;
	wire _w23798_ ;
	wire _w23799_ ;
	wire _w23800_ ;
	wire _w23801_ ;
	wire _w23802_ ;
	wire _w23803_ ;
	wire _w23804_ ;
	wire _w23805_ ;
	wire _w23806_ ;
	wire _w23807_ ;
	wire _w23808_ ;
	wire _w23809_ ;
	wire _w23810_ ;
	wire _w23811_ ;
	wire _w23812_ ;
	wire _w23813_ ;
	wire _w23814_ ;
	wire _w23815_ ;
	wire _w23816_ ;
	wire _w23817_ ;
	wire _w23818_ ;
	wire _w23819_ ;
	wire _w23820_ ;
	wire _w23821_ ;
	wire _w23822_ ;
	wire _w23823_ ;
	wire _w23824_ ;
	wire _w23825_ ;
	wire _w23826_ ;
	wire _w23827_ ;
	wire _w23828_ ;
	wire _w23829_ ;
	wire _w23830_ ;
	wire _w23831_ ;
	wire _w23832_ ;
	wire _w23833_ ;
	wire _w23834_ ;
	wire _w23835_ ;
	wire _w23836_ ;
	wire _w23837_ ;
	wire _w23838_ ;
	wire _w23839_ ;
	wire _w23840_ ;
	wire _w23841_ ;
	wire _w23842_ ;
	wire _w23843_ ;
	wire _w23844_ ;
	wire _w23845_ ;
	wire _w23846_ ;
	wire _w23847_ ;
	wire _w23848_ ;
	wire _w23849_ ;
	wire _w23850_ ;
	wire _w23851_ ;
	wire _w23852_ ;
	wire _w23853_ ;
	wire _w23854_ ;
	wire _w23855_ ;
	wire _w23856_ ;
	wire _w23857_ ;
	wire _w23858_ ;
	wire _w23859_ ;
	wire _w23860_ ;
	wire _w23861_ ;
	wire _w23862_ ;
	wire _w23863_ ;
	wire _w23864_ ;
	wire _w23865_ ;
	wire _w23866_ ;
	wire _w23867_ ;
	wire _w23868_ ;
	wire _w23869_ ;
	wire _w23870_ ;
	wire _w23871_ ;
	wire _w23872_ ;
	wire _w23873_ ;
	wire _w23874_ ;
	wire _w23875_ ;
	wire _w23876_ ;
	wire _w23877_ ;
	wire _w23878_ ;
	wire _w23879_ ;
	wire _w23880_ ;
	wire _w23881_ ;
	wire _w23882_ ;
	wire _w23883_ ;
	wire _w23884_ ;
	wire _w23885_ ;
	wire _w23886_ ;
	wire _w23887_ ;
	wire _w23888_ ;
	wire _w23889_ ;
	wire _w23890_ ;
	wire _w23891_ ;
	wire _w23892_ ;
	wire _w23893_ ;
	wire _w23894_ ;
	wire _w23895_ ;
	wire _w23896_ ;
	wire _w23897_ ;
	wire _w23898_ ;
	wire _w23899_ ;
	wire _w23900_ ;
	wire _w23901_ ;
	wire _w23902_ ;
	wire _w23903_ ;
	wire _w23904_ ;
	wire _w23905_ ;
	wire _w23906_ ;
	wire _w23907_ ;
	wire _w23908_ ;
	wire _w23909_ ;
	wire _w23910_ ;
	wire _w23911_ ;
	wire _w23912_ ;
	wire _w23913_ ;
	wire _w23914_ ;
	wire _w23915_ ;
	wire _w23916_ ;
	wire _w23917_ ;
	wire _w23918_ ;
	wire _w23919_ ;
	wire _w23920_ ;
	wire _w23921_ ;
	wire _w23922_ ;
	wire _w23923_ ;
	wire _w23924_ ;
	wire _w23925_ ;
	wire _w23926_ ;
	wire _w23927_ ;
	wire _w23928_ ;
	wire _w23929_ ;
	wire _w23930_ ;
	wire _w23931_ ;
	wire _w23932_ ;
	wire _w23933_ ;
	wire _w23934_ ;
	wire _w23935_ ;
	wire _w23936_ ;
	wire _w23937_ ;
	wire _w23938_ ;
	wire _w23939_ ;
	wire _w23940_ ;
	wire _w23941_ ;
	wire _w23942_ ;
	wire _w23943_ ;
	wire _w23944_ ;
	wire _w23945_ ;
	wire _w23946_ ;
	wire _w23947_ ;
	wire _w23948_ ;
	wire _w23949_ ;
	wire _w23950_ ;
	wire _w23951_ ;
	wire _w23952_ ;
	wire _w23953_ ;
	wire _w23954_ ;
	wire _w23955_ ;
	wire _w23956_ ;
	wire _w23957_ ;
	wire _w23958_ ;
	wire _w23959_ ;
	wire _w23960_ ;
	wire _w23961_ ;
	wire _w23962_ ;
	wire _w23963_ ;
	wire _w23964_ ;
	wire _w23965_ ;
	wire _w23966_ ;
	wire _w23967_ ;
	wire _w23968_ ;
	wire _w23969_ ;
	wire _w23970_ ;
	wire _w23971_ ;
	wire _w23972_ ;
	wire _w23973_ ;
	wire _w23974_ ;
	wire _w23975_ ;
	wire _w23976_ ;
	wire _w23977_ ;
	wire _w23978_ ;
	wire _w23979_ ;
	wire _w23980_ ;
	wire _w23981_ ;
	wire _w23982_ ;
	wire _w23983_ ;
	wire _w23984_ ;
	wire _w23985_ ;
	wire _w23986_ ;
	wire _w23987_ ;
	wire _w23988_ ;
	wire _w23989_ ;
	wire _w23990_ ;
	wire _w23991_ ;
	wire _w23992_ ;
	wire _w23993_ ;
	wire _w23994_ ;
	wire _w23995_ ;
	wire _w23996_ ;
	wire _w23997_ ;
	wire _w23998_ ;
	wire _w23999_ ;
	wire _w24000_ ;
	wire _w24001_ ;
	wire _w24002_ ;
	wire _w24003_ ;
	wire _w24004_ ;
	wire _w24005_ ;
	wire _w24006_ ;
	wire _w24007_ ;
	wire _w24008_ ;
	wire _w24009_ ;
	wire _w24010_ ;
	wire _w24011_ ;
	wire _w24012_ ;
	wire _w24013_ ;
	wire _w24014_ ;
	wire _w24015_ ;
	wire _w24016_ ;
	wire _w24017_ ;
	wire _w24018_ ;
	wire _w24019_ ;
	wire _w24020_ ;
	wire _w24021_ ;
	wire _w24022_ ;
	wire _w24023_ ;
	wire _w24024_ ;
	wire _w24025_ ;
	wire _w24026_ ;
	wire _w24027_ ;
	wire _w24028_ ;
	wire _w24029_ ;
	wire _w24030_ ;
	wire _w24031_ ;
	wire _w24032_ ;
	wire _w24033_ ;
	wire _w24034_ ;
	wire _w24035_ ;
	wire _w24036_ ;
	wire _w24037_ ;
	wire _w24038_ ;
	wire _w24039_ ;
	wire _w24040_ ;
	wire _w24041_ ;
	wire _w24042_ ;
	wire _w24043_ ;
	wire _w24044_ ;
	wire _w24045_ ;
	wire _w24046_ ;
	wire _w24047_ ;
	wire _w24048_ ;
	wire _w24049_ ;
	wire _w24050_ ;
	wire _w24051_ ;
	wire _w24052_ ;
	wire _w24053_ ;
	wire _w24054_ ;
	wire _w24055_ ;
	wire _w24056_ ;
	wire _w24057_ ;
	wire _w24058_ ;
	wire _w24059_ ;
	wire _w24060_ ;
	wire _w24061_ ;
	wire _w24062_ ;
	wire _w24063_ ;
	wire _w24064_ ;
	wire _w24065_ ;
	wire _w24066_ ;
	wire _w24067_ ;
	wire _w24068_ ;
	wire _w24069_ ;
	wire _w24070_ ;
	wire _w24071_ ;
	wire _w24072_ ;
	wire _w24073_ ;
	wire _w24074_ ;
	wire _w24075_ ;
	wire _w24076_ ;
	wire _w24077_ ;
	wire _w24078_ ;
	wire _w24079_ ;
	wire _w24080_ ;
	wire _w24081_ ;
	wire _w24082_ ;
	wire _w24083_ ;
	wire _w24084_ ;
	wire _w24085_ ;
	wire _w24086_ ;
	wire _w24087_ ;
	wire _w24088_ ;
	wire _w24089_ ;
	wire _w24090_ ;
	wire _w24091_ ;
	wire _w24092_ ;
	wire _w24093_ ;
	wire _w24094_ ;
	wire _w24095_ ;
	wire _w24096_ ;
	wire _w24097_ ;
	wire _w24098_ ;
	wire _w24099_ ;
	wire _w24100_ ;
	wire _w24101_ ;
	wire _w24102_ ;
	wire _w24103_ ;
	wire _w24104_ ;
	wire _w24105_ ;
	wire _w24106_ ;
	wire _w24107_ ;
	wire _w24108_ ;
	wire _w24109_ ;
	wire _w24110_ ;
	wire _w24111_ ;
	wire _w24112_ ;
	wire _w24113_ ;
	wire _w24114_ ;
	wire _w24115_ ;
	wire _w24116_ ;
	wire _w24117_ ;
	wire _w24118_ ;
	wire _w24119_ ;
	wire _w24120_ ;
	wire _w24121_ ;
	wire _w24122_ ;
	wire _w24123_ ;
	wire _w24124_ ;
	wire _w24125_ ;
	wire _w24126_ ;
	wire _w24127_ ;
	wire _w24128_ ;
	wire _w24129_ ;
	wire _w24130_ ;
	wire _w24131_ ;
	wire _w24132_ ;
	wire _w24133_ ;
	wire _w24134_ ;
	wire _w24135_ ;
	wire _w24136_ ;
	wire _w24137_ ;
	wire _w24138_ ;
	wire _w24139_ ;
	wire _w24140_ ;
	wire _w24141_ ;
	wire _w24142_ ;
	wire _w24143_ ;
	wire _w24144_ ;
	wire _w24145_ ;
	wire _w24146_ ;
	wire _w24147_ ;
	wire _w24148_ ;
	wire _w24149_ ;
	wire _w24150_ ;
	wire _w24151_ ;
	wire _w24152_ ;
	wire _w24153_ ;
	wire _w24154_ ;
	wire _w24155_ ;
	wire _w24156_ ;
	wire _w24157_ ;
	wire _w24158_ ;
	wire _w24159_ ;
	wire _w24160_ ;
	wire _w24161_ ;
	wire _w24162_ ;
	wire _w24163_ ;
	wire _w24164_ ;
	wire _w24165_ ;
	wire _w24166_ ;
	wire _w24167_ ;
	wire _w24168_ ;
	wire _w24169_ ;
	wire _w24170_ ;
	wire _w24171_ ;
	wire _w24172_ ;
	wire _w24173_ ;
	wire _w24174_ ;
	wire _w24175_ ;
	wire _w24176_ ;
	wire _w24177_ ;
	wire _w24178_ ;
	wire _w24179_ ;
	wire _w24180_ ;
	wire _w24181_ ;
	wire _w24182_ ;
	wire _w24183_ ;
	wire _w24184_ ;
	wire _w24185_ ;
	wire _w24186_ ;
	wire _w24187_ ;
	wire _w24188_ ;
	wire _w24189_ ;
	wire _w24190_ ;
	wire _w24191_ ;
	wire _w24192_ ;
	wire _w24193_ ;
	wire _w24194_ ;
	wire _w24195_ ;
	wire _w24196_ ;
	wire _w24197_ ;
	wire _w24198_ ;
	wire _w24199_ ;
	wire _w24200_ ;
	wire _w24201_ ;
	wire _w24202_ ;
	wire _w24203_ ;
	wire _w24204_ ;
	wire _w24205_ ;
	wire _w24206_ ;
	wire _w24207_ ;
	wire _w24208_ ;
	wire _w24209_ ;
	wire _w24210_ ;
	wire _w24211_ ;
	wire _w24212_ ;
	wire _w24213_ ;
	wire _w24214_ ;
	wire _w24215_ ;
	wire _w24216_ ;
	wire _w24217_ ;
	wire _w24218_ ;
	wire _w24219_ ;
	wire _w24220_ ;
	wire _w24221_ ;
	wire _w24222_ ;
	wire _w24223_ ;
	wire _w24224_ ;
	wire _w24225_ ;
	wire _w24226_ ;
	wire _w24227_ ;
	wire _w24228_ ;
	wire _w24229_ ;
	wire _w24230_ ;
	wire _w24231_ ;
	wire _w24232_ ;
	wire _w24233_ ;
	wire _w24234_ ;
	wire _w24235_ ;
	wire _w24236_ ;
	wire _w24237_ ;
	wire _w24238_ ;
	wire _w24239_ ;
	wire _w24240_ ;
	wire _w24241_ ;
	wire _w24242_ ;
	wire _w24243_ ;
	wire _w24244_ ;
	wire _w24245_ ;
	wire _w24246_ ;
	wire _w24247_ ;
	wire _w24248_ ;
	wire _w24249_ ;
	wire _w24250_ ;
	wire _w24251_ ;
	wire _w24252_ ;
	wire _w24253_ ;
	wire _w24254_ ;
	wire _w24255_ ;
	wire _w24256_ ;
	wire _w24257_ ;
	wire _w24258_ ;
	wire _w24259_ ;
	wire _w24260_ ;
	wire _w24261_ ;
	wire _w24262_ ;
	wire _w24263_ ;
	wire _w24264_ ;
	wire _w24265_ ;
	wire _w24266_ ;
	wire _w24267_ ;
	wire _w24268_ ;
	wire _w24269_ ;
	wire _w24270_ ;
	wire _w24271_ ;
	wire _w24272_ ;
	wire _w24273_ ;
	wire _w24274_ ;
	wire _w24275_ ;
	wire _w24276_ ;
	wire _w24277_ ;
	wire _w24278_ ;
	wire _w24279_ ;
	wire _w24280_ ;
	wire _w24281_ ;
	wire _w24282_ ;
	wire _w24283_ ;
	wire _w24284_ ;
	wire _w24285_ ;
	wire _w24286_ ;
	wire _w24287_ ;
	wire _w24288_ ;
	wire _w24289_ ;
	wire _w24290_ ;
	wire _w24291_ ;
	wire _w24292_ ;
	wire _w24293_ ;
	wire _w24294_ ;
	wire _w24295_ ;
	wire _w24296_ ;
	wire _w24297_ ;
	wire _w24298_ ;
	wire _w24299_ ;
	wire _w24300_ ;
	wire _w24301_ ;
	wire _w24302_ ;
	wire _w24303_ ;
	wire _w24304_ ;
	wire _w24305_ ;
	wire _w24306_ ;
	wire _w24307_ ;
	wire _w24308_ ;
	wire _w24309_ ;
	wire _w24310_ ;
	wire _w24311_ ;
	wire _w24312_ ;
	wire _w24313_ ;
	wire _w24314_ ;
	wire _w24315_ ;
	wire _w24316_ ;
	wire _w24317_ ;
	wire _w24318_ ;
	wire _w24319_ ;
	wire _w24320_ ;
	wire _w24321_ ;
	wire _w24322_ ;
	wire _w24323_ ;
	wire _w24324_ ;
	wire _w24325_ ;
	wire _w24326_ ;
	wire _w24327_ ;
	wire _w24328_ ;
	wire _w24329_ ;
	wire _w24330_ ;
	wire _w24331_ ;
	wire _w24332_ ;
	wire _w24333_ ;
	wire _w24334_ ;
	wire _w24335_ ;
	wire _w24336_ ;
	wire _w24337_ ;
	wire _w24338_ ;
	wire _w24339_ ;
	wire _w24340_ ;
	wire _w24341_ ;
	wire _w24342_ ;
	wire _w24343_ ;
	wire _w24344_ ;
	wire _w24345_ ;
	wire _w24346_ ;
	wire _w24347_ ;
	wire _w24348_ ;
	wire _w24349_ ;
	wire _w24350_ ;
	wire _w24351_ ;
	wire _w24352_ ;
	wire _w24353_ ;
	wire _w24354_ ;
	wire _w24355_ ;
	wire _w24356_ ;
	wire _w24357_ ;
	wire _w24358_ ;
	wire _w24359_ ;
	wire _w24360_ ;
	wire _w24361_ ;
	wire _w24362_ ;
	wire _w24363_ ;
	wire _w24364_ ;
	wire _w24365_ ;
	wire _w24366_ ;
	wire _w24367_ ;
	wire _w24368_ ;
	wire _w24369_ ;
	wire _w24370_ ;
	wire _w24371_ ;
	wire _w24372_ ;
	wire _w24373_ ;
	wire _w24374_ ;
	wire _w24375_ ;
	wire _w24376_ ;
	wire _w24377_ ;
	wire _w24378_ ;
	wire _w24379_ ;
	wire _w24380_ ;
	wire _w24381_ ;
	wire _w24382_ ;
	wire _w24383_ ;
	wire _w24384_ ;
	wire _w24385_ ;
	wire _w24386_ ;
	wire _w24387_ ;
	wire _w24388_ ;
	wire _w24389_ ;
	wire _w24390_ ;
	wire _w24391_ ;
	wire _w24392_ ;
	wire _w24393_ ;
	wire _w24394_ ;
	wire _w24395_ ;
	wire _w24396_ ;
	wire _w24397_ ;
	wire _w24398_ ;
	wire _w24399_ ;
	wire _w24400_ ;
	wire _w24401_ ;
	wire _w24402_ ;
	wire _w24403_ ;
	wire _w24404_ ;
	wire _w24405_ ;
	wire _w24406_ ;
	wire _w24407_ ;
	wire _w24408_ ;
	wire _w24409_ ;
	wire _w24410_ ;
	wire _w24411_ ;
	wire _w24412_ ;
	wire _w24413_ ;
	wire _w24414_ ;
	wire _w24415_ ;
	wire _w24416_ ;
	wire _w24417_ ;
	wire _w24418_ ;
	wire _w24419_ ;
	wire _w24420_ ;
	wire _w24421_ ;
	wire _w24422_ ;
	wire _w24423_ ;
	wire _w24424_ ;
	wire _w24425_ ;
	wire _w24426_ ;
	wire _w24427_ ;
	wire _w24428_ ;
	wire _w24429_ ;
	wire _w24430_ ;
	wire _w24431_ ;
	wire _w24432_ ;
	wire _w24433_ ;
	wire _w24434_ ;
	wire _w24435_ ;
	wire _w24436_ ;
	wire _w24437_ ;
	wire _w24438_ ;
	wire _w24439_ ;
	wire _w24440_ ;
	wire _w24441_ ;
	wire _w24442_ ;
	wire _w24443_ ;
	wire _w24444_ ;
	wire _w24445_ ;
	wire _w24446_ ;
	wire _w24447_ ;
	wire _w24448_ ;
	wire _w24449_ ;
	wire _w24450_ ;
	wire _w24451_ ;
	wire _w24452_ ;
	wire _w24453_ ;
	wire _w24454_ ;
	wire _w24455_ ;
	wire _w24456_ ;
	wire _w24457_ ;
	wire _w24458_ ;
	wire _w24459_ ;
	wire _w24460_ ;
	wire _w24461_ ;
	wire _w24462_ ;
	wire _w24463_ ;
	wire _w24464_ ;
	wire _w24465_ ;
	wire _w24466_ ;
	wire _w24467_ ;
	wire _w24468_ ;
	wire _w24469_ ;
	wire _w24470_ ;
	wire _w24471_ ;
	wire _w24472_ ;
	wire _w24473_ ;
	wire _w24474_ ;
	wire _w24475_ ;
	wire _w24476_ ;
	wire _w24477_ ;
	wire _w24478_ ;
	wire _w24479_ ;
	wire _w24480_ ;
	wire _w24481_ ;
	wire _w24482_ ;
	wire _w24483_ ;
	wire _w24484_ ;
	wire _w24485_ ;
	wire _w24486_ ;
	wire _w24487_ ;
	wire _w24488_ ;
	wire _w24489_ ;
	wire _w24490_ ;
	wire _w24491_ ;
	wire _w24492_ ;
	wire _w24493_ ;
	wire _w24494_ ;
	wire _w24495_ ;
	wire _w24496_ ;
	wire _w24497_ ;
	wire _w24498_ ;
	wire _w24499_ ;
	wire _w24500_ ;
	wire _w24501_ ;
	wire _w24502_ ;
	wire _w24503_ ;
	wire _w24504_ ;
	wire _w24505_ ;
	wire _w24506_ ;
	wire _w24507_ ;
	wire _w24508_ ;
	wire _w24509_ ;
	wire _w24510_ ;
	wire _w24511_ ;
	wire _w24512_ ;
	wire _w24513_ ;
	wire _w24514_ ;
	wire _w24515_ ;
	wire _w24516_ ;
	wire _w24517_ ;
	wire _w24518_ ;
	wire _w24519_ ;
	wire _w24520_ ;
	wire _w24521_ ;
	wire _w24522_ ;
	wire _w24523_ ;
	wire _w24524_ ;
	wire _w24525_ ;
	wire _w24526_ ;
	wire _w24527_ ;
	wire _w24528_ ;
	wire _w24529_ ;
	wire _w24530_ ;
	wire _w24531_ ;
	wire _w24532_ ;
	wire _w24533_ ;
	wire _w24534_ ;
	wire _w24535_ ;
	wire _w24536_ ;
	wire _w24537_ ;
	wire _w24538_ ;
	wire _w24539_ ;
	wire _w24540_ ;
	wire _w24541_ ;
	wire _w24542_ ;
	wire _w24543_ ;
	wire _w24544_ ;
	wire _w24545_ ;
	wire _w24546_ ;
	wire _w24547_ ;
	wire _w24548_ ;
	wire _w24549_ ;
	wire _w24550_ ;
	wire _w24551_ ;
	wire _w24552_ ;
	wire _w24553_ ;
	wire _w24554_ ;
	wire _w24555_ ;
	wire _w24556_ ;
	wire _w24557_ ;
	wire _w24558_ ;
	wire _w24559_ ;
	wire _w24560_ ;
	wire _w24561_ ;
	wire _w24562_ ;
	wire _w24563_ ;
	wire _w24564_ ;
	wire _w24565_ ;
	wire _w24566_ ;
	wire _w24567_ ;
	wire _w24568_ ;
	wire _w24569_ ;
	wire _w24570_ ;
	wire _w24571_ ;
	wire _w24572_ ;
	wire _w24573_ ;
	wire _w24574_ ;
	wire _w24575_ ;
	wire _w24576_ ;
	wire _w24577_ ;
	wire _w24578_ ;
	wire _w24579_ ;
	wire _w24580_ ;
	wire _w24581_ ;
	wire _w24582_ ;
	wire _w24583_ ;
	wire _w24584_ ;
	wire _w24585_ ;
	wire _w24586_ ;
	wire _w24587_ ;
	wire _w24588_ ;
	wire _w24589_ ;
	wire _w24590_ ;
	wire _w24591_ ;
	wire _w24592_ ;
	wire _w24593_ ;
	wire _w24594_ ;
	wire _w24595_ ;
	wire _w24596_ ;
	wire _w24597_ ;
	wire _w24598_ ;
	wire _w24599_ ;
	wire _w24600_ ;
	wire _w24601_ ;
	wire _w24602_ ;
	wire _w24603_ ;
	wire _w24604_ ;
	wire _w24605_ ;
	wire _w24606_ ;
	wire _w24607_ ;
	wire _w24608_ ;
	wire _w24609_ ;
	wire _w24610_ ;
	wire _w24611_ ;
	wire _w24612_ ;
	wire _w24613_ ;
	wire _w24614_ ;
	wire _w24615_ ;
	wire _w24616_ ;
	wire _w24617_ ;
	wire _w24618_ ;
	wire _w24619_ ;
	wire _w24620_ ;
	wire _w24621_ ;
	wire _w24622_ ;
	wire _w24623_ ;
	wire _w24624_ ;
	wire _w24625_ ;
	wire _w24626_ ;
	wire _w24627_ ;
	wire _w24628_ ;
	wire _w24629_ ;
	wire _w24630_ ;
	wire _w24631_ ;
	wire _w24632_ ;
	wire _w24633_ ;
	wire _w24634_ ;
	wire _w24635_ ;
	wire _w24636_ ;
	wire _w24637_ ;
	wire _w24638_ ;
	wire _w24639_ ;
	wire _w24640_ ;
	wire _w24641_ ;
	wire _w24642_ ;
	wire _w24643_ ;
	wire _w24644_ ;
	wire _w24645_ ;
	wire _w24646_ ;
	wire _w24647_ ;
	wire _w24648_ ;
	wire _w24649_ ;
	wire _w24650_ ;
	wire _w24651_ ;
	wire _w24652_ ;
	wire _w24653_ ;
	wire _w24654_ ;
	wire _w24655_ ;
	wire _w24656_ ;
	wire _w24657_ ;
	wire _w24658_ ;
	wire _w24659_ ;
	wire _w24660_ ;
	wire _w24661_ ;
	wire _w24662_ ;
	wire _w24663_ ;
	wire _w24664_ ;
	wire _w24665_ ;
	wire _w24666_ ;
	wire _w24667_ ;
	wire _w24668_ ;
	wire _w24669_ ;
	wire _w24670_ ;
	wire _w24671_ ;
	wire _w24672_ ;
	wire _w24673_ ;
	wire _w24674_ ;
	wire _w24675_ ;
	wire _w24676_ ;
	wire _w24677_ ;
	wire _w24678_ ;
	wire _w24679_ ;
	wire _w24680_ ;
	wire _w24681_ ;
	wire _w24682_ ;
	wire _w24683_ ;
	wire _w24684_ ;
	wire _w24685_ ;
	wire _w24686_ ;
	wire _w24687_ ;
	wire _w24688_ ;
	wire _w24689_ ;
	wire _w24690_ ;
	wire _w24691_ ;
	wire _w24692_ ;
	wire _w24693_ ;
	wire _w24694_ ;
	wire _w24695_ ;
	wire _w24696_ ;
	wire _w24697_ ;
	wire _w24698_ ;
	wire _w24699_ ;
	wire _w24700_ ;
	wire _w24701_ ;
	wire _w24702_ ;
	wire _w24703_ ;
	wire _w24704_ ;
	wire _w24705_ ;
	wire _w24706_ ;
	wire _w24707_ ;
	wire _w24708_ ;
	wire _w24709_ ;
	wire _w24710_ ;
	wire _w24711_ ;
	wire _w24712_ ;
	wire _w24713_ ;
	wire _w24714_ ;
	wire _w24715_ ;
	wire _w24716_ ;
	wire _w24717_ ;
	wire _w24718_ ;
	wire _w24719_ ;
	wire _w24720_ ;
	wire _w24721_ ;
	wire _w24722_ ;
	wire _w24723_ ;
	wire _w24724_ ;
	wire _w24725_ ;
	wire _w24726_ ;
	wire _w24727_ ;
	wire _w24728_ ;
	wire _w24729_ ;
	wire _w24730_ ;
	wire _w24731_ ;
	wire _w24732_ ;
	wire _w24733_ ;
	wire _w24734_ ;
	wire _w24735_ ;
	wire _w24736_ ;
	wire _w24737_ ;
	wire _w24738_ ;
	wire _w24739_ ;
	wire _w24740_ ;
	wire _w24741_ ;
	wire _w24742_ ;
	wire _w24743_ ;
	wire _w24744_ ;
	wire _w24745_ ;
	wire _w24746_ ;
	wire _w24747_ ;
	wire _w24748_ ;
	wire _w24749_ ;
	wire _w24750_ ;
	wire _w24751_ ;
	wire _w24752_ ;
	wire _w24753_ ;
	wire _w24754_ ;
	wire _w24755_ ;
	wire _w24756_ ;
	wire _w24757_ ;
	wire _w24758_ ;
	wire _w24759_ ;
	wire _w24760_ ;
	wire _w24761_ ;
	wire _w24762_ ;
	wire _w24763_ ;
	wire _w24764_ ;
	wire _w24765_ ;
	wire _w24766_ ;
	wire _w24767_ ;
	wire _w24768_ ;
	wire _w24769_ ;
	wire _w24770_ ;
	wire _w24771_ ;
	wire _w24772_ ;
	wire _w24773_ ;
	wire _w24774_ ;
	wire _w24775_ ;
	wire _w24776_ ;
	wire _w24777_ ;
	wire _w24778_ ;
	wire _w24779_ ;
	wire _w24780_ ;
	wire _w24781_ ;
	wire _w24782_ ;
	wire _w24783_ ;
	wire _w24784_ ;
	wire _w24785_ ;
	wire _w24786_ ;
	wire _w24787_ ;
	wire _w24788_ ;
	wire _w24789_ ;
	wire _w24790_ ;
	wire _w24791_ ;
	wire _w24792_ ;
	wire _w24793_ ;
	wire _w24794_ ;
	wire _w24795_ ;
	wire _w24796_ ;
	wire _w24797_ ;
	wire _w24798_ ;
	wire _w24799_ ;
	wire _w24800_ ;
	wire _w24801_ ;
	wire _w24802_ ;
	wire _w24803_ ;
	wire _w24804_ ;
	wire _w24805_ ;
	wire _w24806_ ;
	wire _w24807_ ;
	wire _w24808_ ;
	wire _w24809_ ;
	wire _w24810_ ;
	wire _w24811_ ;
	wire _w24812_ ;
	wire _w24813_ ;
	wire _w24814_ ;
	wire _w24815_ ;
	wire _w24816_ ;
	wire _w24817_ ;
	wire _w24818_ ;
	wire _w24819_ ;
	wire _w24820_ ;
	wire _w24821_ ;
	wire _w24822_ ;
	wire _w24823_ ;
	wire _w24824_ ;
	wire _w24825_ ;
	wire _w24826_ ;
	wire _w24827_ ;
	wire _w24828_ ;
	wire _w24829_ ;
	wire _w24830_ ;
	wire _w24831_ ;
	wire _w24832_ ;
	wire _w24833_ ;
	wire _w24834_ ;
	wire _w24835_ ;
	wire _w24836_ ;
	wire _w24837_ ;
	wire _w24838_ ;
	wire _w24839_ ;
	wire _w24840_ ;
	wire _w24841_ ;
	wire _w24842_ ;
	wire _w24843_ ;
	wire _w24844_ ;
	wire _w24845_ ;
	wire _w24846_ ;
	wire _w24847_ ;
	wire _w24848_ ;
	wire _w24849_ ;
	wire _w24850_ ;
	wire _w24851_ ;
	wire _w24852_ ;
	wire _w24853_ ;
	wire _w24854_ ;
	wire _w24855_ ;
	wire _w24856_ ;
	wire _w24857_ ;
	wire _w24858_ ;
	wire _w24859_ ;
	wire _w24860_ ;
	wire _w24861_ ;
	wire _w24862_ ;
	wire _w24863_ ;
	wire _w24864_ ;
	wire _w24865_ ;
	wire _w24866_ ;
	wire _w24867_ ;
	wire _w24868_ ;
	wire _w24869_ ;
	wire _w24870_ ;
	wire _w24871_ ;
	wire _w24872_ ;
	wire _w24873_ ;
	wire _w24874_ ;
	wire _w24875_ ;
	wire _w24876_ ;
	wire _w24877_ ;
	wire _w24878_ ;
	wire _w24879_ ;
	wire _w24880_ ;
	wire _w24881_ ;
	wire _w24882_ ;
	wire _w24883_ ;
	wire _w24884_ ;
	wire _w24885_ ;
	wire _w24886_ ;
	wire _w24887_ ;
	wire _w24888_ ;
	wire _w24889_ ;
	wire _w24890_ ;
	wire _w24891_ ;
	wire _w24892_ ;
	wire _w24893_ ;
	wire _w24894_ ;
	wire _w24895_ ;
	wire _w24896_ ;
	wire _w24897_ ;
	wire _w24898_ ;
	wire _w24899_ ;
	wire _w24900_ ;
	wire _w24901_ ;
	wire _w24902_ ;
	wire _w24903_ ;
	wire _w24904_ ;
	wire _w24905_ ;
	wire _w24906_ ;
	wire _w24907_ ;
	wire _w24908_ ;
	wire _w24909_ ;
	wire _w24910_ ;
	wire _w24911_ ;
	wire _w24912_ ;
	wire _w24913_ ;
	wire _w24914_ ;
	wire _w24915_ ;
	wire _w24916_ ;
	wire _w24917_ ;
	wire _w24918_ ;
	wire _w24919_ ;
	wire _w24920_ ;
	wire _w24921_ ;
	wire _w24922_ ;
	wire _w24923_ ;
	wire _w24924_ ;
	wire _w24925_ ;
	wire _w24926_ ;
	wire _w24927_ ;
	wire _w24928_ ;
	wire _w24929_ ;
	wire _w24930_ ;
	wire _w24931_ ;
	wire _w24932_ ;
	wire _w24933_ ;
	wire _w24934_ ;
	wire _w24935_ ;
	wire _w24936_ ;
	wire _w24937_ ;
	wire _w24938_ ;
	wire _w24939_ ;
	wire _w24940_ ;
	wire _w24941_ ;
	wire _w24942_ ;
	wire _w24943_ ;
	wire _w24944_ ;
	wire _w24945_ ;
	wire _w24946_ ;
	wire _w24947_ ;
	wire _w24948_ ;
	wire _w24949_ ;
	wire _w24950_ ;
	wire _w24951_ ;
	wire _w24952_ ;
	wire _w24953_ ;
	wire _w24954_ ;
	wire _w24955_ ;
	wire _w24956_ ;
	wire _w24957_ ;
	wire _w24958_ ;
	wire _w24959_ ;
	wire _w24960_ ;
	wire _w24961_ ;
	wire _w24962_ ;
	wire _w24963_ ;
	wire _w24964_ ;
	wire _w24965_ ;
	wire _w24966_ ;
	wire _w24967_ ;
	wire _w24968_ ;
	wire _w24969_ ;
	wire _w24970_ ;
	wire _w24971_ ;
	wire _w24972_ ;
	wire _w24973_ ;
	wire _w24974_ ;
	wire _w24975_ ;
	wire _w24976_ ;
	wire _w24977_ ;
	wire _w24978_ ;
	wire _w24979_ ;
	wire _w24980_ ;
	wire _w24981_ ;
	wire _w24982_ ;
	wire _w24983_ ;
	wire _w24984_ ;
	wire _w24985_ ;
	wire _w24986_ ;
	wire _w24987_ ;
	wire _w24988_ ;
	wire _w24989_ ;
	wire _w24990_ ;
	wire _w24991_ ;
	wire _w24992_ ;
	wire _w24993_ ;
	wire _w24994_ ;
	wire _w24995_ ;
	wire _w24996_ ;
	wire _w24997_ ;
	wire _w24998_ ;
	wire _w24999_ ;
	wire _w25000_ ;
	wire _w25001_ ;
	wire _w25002_ ;
	wire _w25003_ ;
	wire _w25004_ ;
	wire _w25005_ ;
	wire _w25006_ ;
	wire _w25007_ ;
	wire _w25008_ ;
	wire _w25009_ ;
	wire _w25010_ ;
	wire _w25011_ ;
	wire _w25012_ ;
	wire _w25013_ ;
	wire _w25014_ ;
	wire _w25015_ ;
	wire _w25016_ ;
	wire _w25017_ ;
	wire _w25018_ ;
	wire _w25019_ ;
	wire _w25020_ ;
	wire _w25021_ ;
	wire _w25022_ ;
	wire _w25023_ ;
	wire _w25024_ ;
	wire _w25025_ ;
	wire _w25026_ ;
	wire _w25027_ ;
	wire _w25028_ ;
	wire _w25029_ ;
	wire _w25030_ ;
	wire _w25031_ ;
	wire _w25032_ ;
	wire _w25033_ ;
	wire _w25034_ ;
	wire _w25035_ ;
	wire _w25036_ ;
	wire _w25037_ ;
	wire _w25038_ ;
	wire _w25039_ ;
	wire _w25040_ ;
	wire _w25041_ ;
	wire _w25042_ ;
	wire _w25043_ ;
	wire _w25044_ ;
	wire _w25045_ ;
	wire _w25046_ ;
	wire _w25047_ ;
	wire _w25048_ ;
	wire _w25049_ ;
	wire _w25050_ ;
	wire _w25051_ ;
	wire _w25052_ ;
	wire _w25053_ ;
	wire _w25054_ ;
	wire _w25055_ ;
	wire _w25056_ ;
	wire _w25057_ ;
	wire _w25058_ ;
	wire _w25059_ ;
	wire _w25060_ ;
	wire _w25061_ ;
	wire _w25062_ ;
	wire _w25063_ ;
	wire _w25064_ ;
	wire _w25065_ ;
	wire _w25066_ ;
	wire _w25067_ ;
	wire _w25068_ ;
	wire _w25069_ ;
	wire _w25070_ ;
	wire _w25071_ ;
	wire _w25072_ ;
	wire _w25073_ ;
	wire _w25074_ ;
	wire _w25075_ ;
	wire _w25076_ ;
	wire _w25077_ ;
	wire _w25078_ ;
	wire _w25079_ ;
	wire _w25080_ ;
	wire _w25081_ ;
	wire _w25082_ ;
	wire _w25083_ ;
	wire _w25084_ ;
	wire _w25085_ ;
	wire _w25086_ ;
	wire _w25087_ ;
	wire _w25088_ ;
	wire _w25089_ ;
	wire _w25090_ ;
	wire _w25091_ ;
	wire _w25092_ ;
	wire _w25093_ ;
	wire _w25094_ ;
	wire _w25095_ ;
	wire _w25096_ ;
	wire _w25097_ ;
	wire _w25098_ ;
	wire _w25099_ ;
	wire _w25100_ ;
	wire _w25101_ ;
	wire _w25102_ ;
	wire _w25103_ ;
	wire _w25104_ ;
	wire _w25105_ ;
	wire _w25106_ ;
	wire _w25107_ ;
	wire _w25108_ ;
	wire _w25109_ ;
	wire _w25110_ ;
	wire _w25111_ ;
	wire _w25112_ ;
	wire _w25113_ ;
	wire _w25114_ ;
	wire _w25115_ ;
	wire _w25116_ ;
	wire _w25117_ ;
	wire _w25118_ ;
	wire _w25119_ ;
	wire _w25120_ ;
	wire _w25121_ ;
	wire _w25122_ ;
	wire _w25123_ ;
	wire _w25124_ ;
	wire _w25125_ ;
	wire _w25126_ ;
	wire _w25127_ ;
	wire _w25128_ ;
	wire _w25129_ ;
	wire _w25130_ ;
	wire _w25131_ ;
	wire _w25132_ ;
	wire _w25133_ ;
	wire _w25134_ ;
	wire _w25135_ ;
	wire _w25136_ ;
	wire _w25137_ ;
	wire _w25138_ ;
	wire _w25139_ ;
	wire _w25140_ ;
	wire _w25141_ ;
	wire _w25142_ ;
	wire _w25143_ ;
	wire _w25144_ ;
	wire _w25145_ ;
	wire _w25146_ ;
	wire _w25147_ ;
	wire _w25148_ ;
	wire _w25149_ ;
	wire _w25150_ ;
	wire _w25151_ ;
	wire _w25152_ ;
	wire _w25153_ ;
	wire _w25154_ ;
	wire _w25155_ ;
	wire _w25156_ ;
	wire _w25157_ ;
	wire _w25158_ ;
	wire _w25159_ ;
	wire _w25160_ ;
	wire _w25161_ ;
	wire _w25162_ ;
	wire _w25163_ ;
	wire _w25164_ ;
	wire _w25165_ ;
	wire _w25166_ ;
	wire _w25167_ ;
	wire _w25168_ ;
	wire _w25169_ ;
	wire _w25170_ ;
	wire _w25171_ ;
	wire _w25172_ ;
	wire _w25173_ ;
	wire _w25174_ ;
	wire _w25175_ ;
	wire _w25176_ ;
	wire _w25177_ ;
	wire _w25178_ ;
	wire _w25179_ ;
	wire _w25180_ ;
	wire _w25181_ ;
	wire _w25182_ ;
	wire _w25183_ ;
	wire _w25184_ ;
	wire _w25185_ ;
	wire _w25186_ ;
	wire _w25187_ ;
	wire _w25188_ ;
	wire _w25189_ ;
	wire _w25190_ ;
	wire _w25191_ ;
	wire _w25192_ ;
	wire _w25193_ ;
	wire _w25194_ ;
	wire _w25195_ ;
	wire _w25196_ ;
	wire _w25197_ ;
	wire _w25198_ ;
	wire _w25199_ ;
	wire _w25200_ ;
	wire _w25201_ ;
	wire _w25202_ ;
	wire _w25203_ ;
	wire _w25204_ ;
	wire _w25205_ ;
	wire _w25206_ ;
	wire _w25207_ ;
	wire _w25208_ ;
	wire _w25209_ ;
	wire _w25210_ ;
	wire _w25211_ ;
	wire _w25212_ ;
	wire _w25213_ ;
	wire _w25214_ ;
	wire _w25215_ ;
	wire _w25216_ ;
	wire _w25217_ ;
	wire _w25218_ ;
	wire _w25219_ ;
	wire _w25220_ ;
	wire _w25221_ ;
	wire _w25222_ ;
	wire _w25223_ ;
	wire _w25224_ ;
	wire _w25225_ ;
	wire _w25226_ ;
	wire _w25227_ ;
	wire _w25228_ ;
	wire _w25229_ ;
	wire _w25230_ ;
	wire _w25231_ ;
	wire _w25232_ ;
	wire _w25233_ ;
	wire _w25234_ ;
	wire _w25235_ ;
	wire _w25236_ ;
	wire _w25237_ ;
	wire _w25238_ ;
	wire _w25239_ ;
	wire _w25240_ ;
	wire _w25241_ ;
	wire _w25242_ ;
	wire _w25243_ ;
	wire _w25244_ ;
	wire _w25245_ ;
	wire _w25246_ ;
	wire _w25247_ ;
	wire _w25248_ ;
	wire _w25249_ ;
	wire _w25250_ ;
	wire _w25251_ ;
	wire _w25252_ ;
	wire _w25253_ ;
	wire _w25254_ ;
	wire _w25255_ ;
	wire _w25256_ ;
	wire _w25257_ ;
	wire _w25258_ ;
	wire _w25259_ ;
	wire _w25260_ ;
	wire _w25261_ ;
	wire _w25262_ ;
	wire _w25263_ ;
	wire _w25264_ ;
	wire _w25265_ ;
	wire _w25266_ ;
	wire _w25267_ ;
	wire _w25268_ ;
	wire _w25269_ ;
	wire _w25270_ ;
	wire _w25271_ ;
	wire _w25272_ ;
	wire _w25273_ ;
	wire _w25274_ ;
	wire _w25275_ ;
	wire _w25276_ ;
	wire _w25277_ ;
	wire _w25278_ ;
	wire _w25279_ ;
	wire _w25280_ ;
	wire _w25281_ ;
	wire _w25282_ ;
	wire _w25283_ ;
	wire _w25284_ ;
	wire _w25285_ ;
	wire _w25286_ ;
	wire _w25287_ ;
	wire _w25288_ ;
	wire _w25289_ ;
	wire _w25290_ ;
	wire _w25291_ ;
	wire _w25292_ ;
	wire _w25293_ ;
	wire _w25294_ ;
	wire _w25295_ ;
	wire _w25296_ ;
	wire _w25297_ ;
	wire _w25298_ ;
	wire _w25299_ ;
	wire _w25300_ ;
	wire _w25301_ ;
	wire _w25302_ ;
	wire _w25303_ ;
	wire _w25304_ ;
	wire _w25305_ ;
	wire _w25306_ ;
	wire _w25307_ ;
	wire _w25308_ ;
	wire _w25309_ ;
	wire _w25310_ ;
	wire _w25311_ ;
	wire _w25312_ ;
	wire _w25313_ ;
	wire _w25314_ ;
	wire _w25315_ ;
	wire _w25316_ ;
	wire _w25317_ ;
	wire _w25318_ ;
	wire _w25319_ ;
	wire _w25320_ ;
	wire _w25321_ ;
	wire _w25322_ ;
	wire _w25323_ ;
	wire _w25324_ ;
	wire _w25325_ ;
	wire _w25326_ ;
	wire _w25327_ ;
	wire _w25328_ ;
	wire _w25329_ ;
	wire _w25330_ ;
	wire _w25331_ ;
	wire _w25332_ ;
	wire _w25333_ ;
	wire _w25334_ ;
	wire _w25335_ ;
	wire _w25336_ ;
	wire _w25337_ ;
	wire _w25338_ ;
	wire _w25339_ ;
	wire _w25340_ ;
	wire _w25341_ ;
	wire _w25342_ ;
	wire _w25343_ ;
	wire _w25344_ ;
	wire _w25345_ ;
	wire _w25346_ ;
	wire _w25347_ ;
	wire _w25348_ ;
	wire _w25349_ ;
	wire _w25350_ ;
	wire _w25351_ ;
	wire _w25352_ ;
	wire _w25353_ ;
	wire _w25354_ ;
	wire _w25355_ ;
	wire _w25356_ ;
	wire _w25357_ ;
	wire _w25358_ ;
	wire _w25359_ ;
	wire _w25360_ ;
	wire _w25361_ ;
	wire _w25362_ ;
	wire _w25363_ ;
	wire _w25364_ ;
	wire _w25365_ ;
	wire _w25366_ ;
	wire _w25367_ ;
	wire _w25368_ ;
	wire _w25369_ ;
	wire _w25370_ ;
	wire _w25371_ ;
	wire _w25372_ ;
	wire _w25373_ ;
	wire _w25374_ ;
	wire _w25375_ ;
	wire _w25376_ ;
	wire _w25377_ ;
	wire _w25378_ ;
	wire _w25379_ ;
	wire _w25380_ ;
	wire _w25381_ ;
	wire _w25382_ ;
	wire _w25383_ ;
	wire _w25384_ ;
	wire _w25385_ ;
	wire _w25386_ ;
	wire _w25387_ ;
	wire _w25388_ ;
	wire _w25389_ ;
	wire _w25390_ ;
	wire _w25391_ ;
	wire _w25392_ ;
	wire _w25393_ ;
	wire _w25394_ ;
	wire _w25395_ ;
	wire _w25396_ ;
	wire _w25397_ ;
	wire _w25398_ ;
	wire _w25399_ ;
	wire _w25400_ ;
	wire _w25401_ ;
	wire _w25402_ ;
	wire _w25403_ ;
	wire _w25404_ ;
	wire _w25405_ ;
	wire _w25406_ ;
	wire _w25407_ ;
	wire _w25408_ ;
	wire _w25409_ ;
	wire _w25410_ ;
	wire _w25411_ ;
	wire _w25412_ ;
	wire _w25413_ ;
	wire _w25414_ ;
	wire _w25415_ ;
	wire _w25416_ ;
	wire _w25417_ ;
	wire _w25418_ ;
	wire _w25419_ ;
	wire _w25420_ ;
	wire _w25421_ ;
	wire _w25422_ ;
	wire _w25423_ ;
	wire _w25424_ ;
	wire _w25425_ ;
	wire _w25426_ ;
	wire _w25427_ ;
	wire _w25428_ ;
	wire _w25429_ ;
	wire _w25430_ ;
	wire _w25431_ ;
	wire _w25432_ ;
	wire _w25433_ ;
	wire _w25434_ ;
	wire _w25435_ ;
	wire _w25436_ ;
	wire _w25437_ ;
	wire _w25438_ ;
	wire _w25439_ ;
	wire _w25440_ ;
	wire _w25441_ ;
	wire _w25442_ ;
	wire _w25443_ ;
	wire _w25444_ ;
	wire _w25445_ ;
	wire _w25446_ ;
	wire _w25447_ ;
	wire _w25448_ ;
	wire _w25449_ ;
	wire _w25450_ ;
	wire _w25451_ ;
	wire _w25452_ ;
	wire _w25453_ ;
	wire _w25454_ ;
	wire _w25455_ ;
	wire _w25456_ ;
	wire _w25457_ ;
	wire _w25458_ ;
	wire _w25459_ ;
	wire _w25460_ ;
	wire _w25461_ ;
	wire _w25462_ ;
	wire _w25463_ ;
	wire _w25464_ ;
	wire _w25465_ ;
	wire _w25466_ ;
	wire _w25467_ ;
	wire _w25468_ ;
	wire _w25469_ ;
	wire _w25470_ ;
	wire _w25471_ ;
	wire _w25472_ ;
	wire _w25473_ ;
	wire _w25474_ ;
	wire _w25475_ ;
	wire _w25476_ ;
	wire _w25477_ ;
	wire _w25478_ ;
	wire _w25479_ ;
	wire _w25480_ ;
	wire _w25481_ ;
	wire _w25482_ ;
	wire _w25483_ ;
	wire _w25484_ ;
	wire _w25485_ ;
	wire _w25486_ ;
	wire _w25487_ ;
	wire _w25488_ ;
	wire _w25489_ ;
	wire _w25490_ ;
	wire _w25491_ ;
	wire _w25492_ ;
	wire _w25493_ ;
	wire _w25494_ ;
	wire _w25495_ ;
	wire _w25496_ ;
	wire _w25497_ ;
	wire _w25498_ ;
	wire _w25499_ ;
	wire _w25500_ ;
	wire _w25501_ ;
	wire _w25502_ ;
	wire _w25503_ ;
	wire _w25504_ ;
	wire _w25505_ ;
	wire _w25506_ ;
	wire _w25507_ ;
	wire _w25508_ ;
	wire _w25509_ ;
	wire _w25510_ ;
	wire _w25511_ ;
	wire _w25512_ ;
	wire _w25513_ ;
	wire _w25514_ ;
	wire _w25515_ ;
	wire _w25516_ ;
	wire _w25517_ ;
	wire _w25518_ ;
	wire _w25519_ ;
	wire _w25520_ ;
	wire _w25521_ ;
	wire _w25522_ ;
	wire _w25523_ ;
	wire _w25524_ ;
	wire _w25525_ ;
	wire _w25526_ ;
	wire _w25527_ ;
	wire _w25528_ ;
	wire _w25529_ ;
	wire _w25530_ ;
	wire _w25531_ ;
	wire _w25532_ ;
	wire _w25533_ ;
	wire _w25534_ ;
	wire _w25535_ ;
	wire _w25536_ ;
	wire _w25537_ ;
	wire _w25538_ ;
	wire _w25539_ ;
	wire _w25540_ ;
	wire _w25541_ ;
	wire _w25542_ ;
	wire _w25543_ ;
	wire _w25544_ ;
	wire _w25545_ ;
	wire _w25546_ ;
	wire _w25547_ ;
	wire _w25548_ ;
	wire _w25549_ ;
	wire _w25550_ ;
	wire _w25551_ ;
	wire _w25552_ ;
	wire _w25553_ ;
	wire _w25554_ ;
	wire _w25555_ ;
	wire _w25556_ ;
	wire _w25557_ ;
	wire _w25558_ ;
	wire _w25559_ ;
	wire _w25560_ ;
	wire _w25561_ ;
	wire _w25562_ ;
	wire _w25563_ ;
	wire _w25564_ ;
	wire _w25565_ ;
	wire _w25566_ ;
	wire _w25567_ ;
	wire _w25568_ ;
	wire _w25569_ ;
	wire _w25570_ ;
	wire _w25571_ ;
	wire _w25572_ ;
	wire _w25573_ ;
	wire _w25574_ ;
	wire _w25575_ ;
	wire _w25576_ ;
	wire _w25577_ ;
	wire _w25578_ ;
	wire _w25579_ ;
	wire _w25580_ ;
	wire _w25581_ ;
	wire _w25582_ ;
	wire _w25583_ ;
	wire _w25584_ ;
	wire _w25585_ ;
	wire _w25586_ ;
	wire _w25587_ ;
	wire _w25588_ ;
	wire _w25589_ ;
	wire _w25590_ ;
	wire _w25591_ ;
	wire _w25592_ ;
	wire _w25593_ ;
	wire _w25594_ ;
	wire _w25595_ ;
	wire _w25596_ ;
	wire _w25597_ ;
	wire _w25598_ ;
	wire _w25599_ ;
	wire _w25600_ ;
	wire _w25601_ ;
	wire _w25602_ ;
	wire _w25603_ ;
	wire _w25604_ ;
	wire _w25605_ ;
	wire _w25606_ ;
	wire _w25607_ ;
	wire _w25608_ ;
	wire _w25609_ ;
	wire _w25610_ ;
	wire _w25611_ ;
	wire _w25612_ ;
	wire _w25613_ ;
	wire _w25614_ ;
	wire _w25615_ ;
	wire _w25616_ ;
	wire _w25617_ ;
	wire _w25618_ ;
	wire _w25619_ ;
	wire _w25620_ ;
	wire _w25621_ ;
	wire _w25622_ ;
	wire _w25623_ ;
	wire _w25624_ ;
	wire _w25625_ ;
	wire _w25626_ ;
	wire _w25627_ ;
	wire _w25628_ ;
	wire _w25629_ ;
	wire _w25630_ ;
	wire _w25631_ ;
	wire _w25632_ ;
	wire _w25633_ ;
	wire _w25634_ ;
	wire _w25635_ ;
	wire _w25636_ ;
	wire _w25637_ ;
	wire _w25638_ ;
	wire _w25639_ ;
	wire _w25640_ ;
	wire _w25641_ ;
	wire _w25642_ ;
	wire _w25643_ ;
	wire _w25644_ ;
	wire _w25645_ ;
	wire _w25646_ ;
	wire _w25647_ ;
	wire _w25648_ ;
	wire _w25649_ ;
	wire _w25650_ ;
	wire _w25651_ ;
	wire _w25652_ ;
	wire _w25653_ ;
	wire _w25654_ ;
	wire _w25655_ ;
	wire _w25656_ ;
	wire _w25657_ ;
	wire _w25658_ ;
	wire _w25659_ ;
	wire _w25660_ ;
	wire _w25661_ ;
	wire _w25662_ ;
	wire _w25663_ ;
	wire _w25664_ ;
	wire _w25665_ ;
	wire _w25666_ ;
	wire _w25667_ ;
	wire _w25668_ ;
	wire _w25669_ ;
	wire _w25670_ ;
	wire _w25671_ ;
	wire _w25672_ ;
	wire _w25673_ ;
	wire _w25674_ ;
	wire _w25675_ ;
	wire _w25676_ ;
	wire _w25677_ ;
	wire _w25678_ ;
	wire _w25679_ ;
	wire _w25680_ ;
	wire _w25681_ ;
	wire _w25682_ ;
	wire _w25683_ ;
	wire _w25684_ ;
	wire _w25685_ ;
	wire _w25686_ ;
	wire _w25687_ ;
	wire _w25688_ ;
	wire _w25689_ ;
	wire _w25690_ ;
	wire _w25691_ ;
	wire _w25692_ ;
	wire _w25693_ ;
	wire _w25694_ ;
	wire _w25695_ ;
	wire _w25696_ ;
	wire _w25697_ ;
	wire _w25698_ ;
	wire _w25699_ ;
	wire _w25700_ ;
	wire _w25701_ ;
	wire _w25702_ ;
	wire _w25703_ ;
	wire _w25704_ ;
	wire _w25705_ ;
	wire _w25706_ ;
	wire _w25707_ ;
	wire _w25708_ ;
	wire _w25709_ ;
	wire _w25710_ ;
	wire _w25711_ ;
	wire _w25712_ ;
	wire _w25713_ ;
	wire _w25714_ ;
	wire _w25715_ ;
	wire _w25716_ ;
	wire _w25717_ ;
	wire _w25718_ ;
	wire _w25719_ ;
	wire _w25720_ ;
	wire _w25721_ ;
	wire _w25722_ ;
	wire _w25723_ ;
	wire _w25724_ ;
	wire _w25725_ ;
	wire _w25726_ ;
	wire _w25727_ ;
	wire _w25728_ ;
	wire _w25729_ ;
	wire _w25730_ ;
	wire _w25731_ ;
	wire _w25732_ ;
	wire _w25733_ ;
	wire _w25734_ ;
	wire _w25735_ ;
	wire _w25736_ ;
	wire _w25737_ ;
	wire _w25738_ ;
	wire _w25739_ ;
	wire _w25740_ ;
	wire _w25741_ ;
	wire _w25742_ ;
	wire _w25743_ ;
	wire _w25744_ ;
	wire _w25745_ ;
	wire _w25746_ ;
	wire _w25747_ ;
	wire _w25748_ ;
	wire _w25749_ ;
	wire _w25750_ ;
	wire _w25751_ ;
	wire _w25752_ ;
	wire _w25753_ ;
	wire _w25754_ ;
	wire _w25755_ ;
	wire _w25756_ ;
	wire _w25757_ ;
	wire _w25758_ ;
	wire _w25759_ ;
	wire _w25760_ ;
	wire _w25761_ ;
	wire _w25762_ ;
	wire _w25763_ ;
	wire _w25764_ ;
	wire _w25765_ ;
	wire _w25766_ ;
	wire _w25767_ ;
	wire _w25768_ ;
	wire _w25769_ ;
	wire _w25770_ ;
	wire _w25771_ ;
	wire _w25772_ ;
	wire _w25773_ ;
	wire _w25774_ ;
	wire _w25775_ ;
	wire _w25776_ ;
	wire _w25777_ ;
	wire _w25778_ ;
	wire _w25779_ ;
	wire _w25780_ ;
	wire _w25781_ ;
	wire _w25782_ ;
	wire _w25783_ ;
	wire _w25784_ ;
	wire _w25785_ ;
	wire _w25786_ ;
	wire _w25787_ ;
	wire _w25788_ ;
	wire _w25789_ ;
	wire _w25790_ ;
	wire _w25791_ ;
	wire _w25792_ ;
	wire _w25793_ ;
	wire _w25794_ ;
	wire _w25795_ ;
	wire _w25796_ ;
	wire _w25797_ ;
	wire _w25798_ ;
	wire _w25799_ ;
	wire _w25800_ ;
	wire _w25801_ ;
	wire _w25802_ ;
	wire _w25803_ ;
	wire _w25804_ ;
	wire _w25805_ ;
	wire _w25806_ ;
	wire _w25807_ ;
	wire _w25808_ ;
	wire _w25809_ ;
	wire _w25810_ ;
	wire _w25811_ ;
	wire _w25812_ ;
	wire _w25813_ ;
	wire _w25814_ ;
	wire _w25815_ ;
	wire _w25816_ ;
	wire _w25817_ ;
	wire _w25818_ ;
	wire _w25819_ ;
	wire _w25820_ ;
	wire _w25821_ ;
	wire _w25822_ ;
	wire _w25823_ ;
	wire _w25824_ ;
	wire _w25825_ ;
	wire _w25826_ ;
	wire _w25827_ ;
	wire _w25828_ ;
	wire _w25829_ ;
	wire _w25830_ ;
	wire _w25831_ ;
	wire _w25832_ ;
	wire _w25833_ ;
	wire _w25834_ ;
	wire _w25835_ ;
	wire _w25836_ ;
	wire _w25837_ ;
	wire _w25838_ ;
	wire _w25839_ ;
	wire _w25840_ ;
	wire _w25841_ ;
	wire _w25842_ ;
	wire _w25843_ ;
	wire _w25844_ ;
	wire _w25845_ ;
	wire _w25846_ ;
	wire _w25847_ ;
	wire _w25848_ ;
	wire _w25849_ ;
	wire _w25850_ ;
	wire _w25851_ ;
	wire _w25852_ ;
	wire _w25853_ ;
	wire _w25854_ ;
	wire _w25855_ ;
	wire _w25856_ ;
	wire _w25857_ ;
	wire _w25858_ ;
	wire _w25859_ ;
	wire _w25860_ ;
	wire _w25861_ ;
	wire _w25862_ ;
	wire _w25863_ ;
	wire _w25864_ ;
	wire _w25865_ ;
	wire _w25866_ ;
	wire _w25867_ ;
	wire _w25868_ ;
	wire _w25869_ ;
	wire _w25870_ ;
	wire _w25871_ ;
	wire _w25872_ ;
	wire _w25873_ ;
	wire _w25874_ ;
	wire _w25875_ ;
	wire _w25876_ ;
	wire _w25877_ ;
	wire _w25878_ ;
	wire _w25879_ ;
	wire _w25880_ ;
	wire _w25881_ ;
	wire _w25882_ ;
	wire _w25883_ ;
	wire _w25884_ ;
	wire _w25885_ ;
	wire _w25886_ ;
	wire _w25887_ ;
	wire _w25888_ ;
	wire _w25889_ ;
	wire _w25890_ ;
	wire _w25891_ ;
	wire _w25892_ ;
	wire _w25893_ ;
	wire _w25894_ ;
	wire _w25895_ ;
	wire _w25896_ ;
	wire _w25897_ ;
	wire _w25898_ ;
	wire _w25899_ ;
	wire _w25900_ ;
	wire _w25901_ ;
	wire _w25902_ ;
	wire _w25903_ ;
	wire _w25904_ ;
	wire _w25905_ ;
	wire _w25906_ ;
	wire _w25907_ ;
	wire _w25908_ ;
	wire _w25909_ ;
	wire _w25910_ ;
	wire _w25911_ ;
	wire _w25912_ ;
	wire _w25913_ ;
	wire _w25914_ ;
	wire _w25915_ ;
	wire _w25916_ ;
	wire _w25917_ ;
	wire _w25918_ ;
	wire _w25919_ ;
	wire _w25920_ ;
	wire _w25921_ ;
	wire _w25922_ ;
	wire _w25923_ ;
	wire _w25924_ ;
	wire _w25925_ ;
	wire _w25926_ ;
	wire _w25927_ ;
	wire _w25928_ ;
	wire _w25929_ ;
	wire _w25930_ ;
	wire _w25931_ ;
	wire _w25932_ ;
	wire _w25933_ ;
	wire _w25934_ ;
	wire _w25935_ ;
	wire _w25936_ ;
	wire _w25937_ ;
	wire _w25938_ ;
	wire _w25939_ ;
	wire _w25940_ ;
	wire _w25941_ ;
	wire _w25942_ ;
	wire _w25943_ ;
	wire _w25944_ ;
	wire _w25945_ ;
	wire _w25946_ ;
	wire _w25947_ ;
	wire _w25948_ ;
	wire _w25949_ ;
	wire _w25950_ ;
	wire _w25951_ ;
	wire _w25952_ ;
	wire _w25953_ ;
	wire _w25954_ ;
	wire _w25955_ ;
	wire _w25956_ ;
	wire _w25957_ ;
	wire _w25958_ ;
	wire _w25959_ ;
	wire _w25960_ ;
	wire _w25961_ ;
	wire _w25962_ ;
	wire _w25963_ ;
	wire _w25964_ ;
	wire _w25965_ ;
	wire _w25966_ ;
	wire _w25967_ ;
	wire _w25968_ ;
	wire _w25969_ ;
	wire _w25970_ ;
	wire _w25971_ ;
	wire _w25972_ ;
	wire _w25973_ ;
	wire _w25974_ ;
	wire _w25975_ ;
	wire _w25976_ ;
	wire _w25977_ ;
	wire _w25978_ ;
	wire _w25979_ ;
	wire _w25980_ ;
	wire _w25981_ ;
	wire _w25982_ ;
	wire _w25983_ ;
	wire _w25984_ ;
	wire _w25985_ ;
	wire _w25986_ ;
	wire _w25987_ ;
	wire _w25988_ ;
	wire _w25989_ ;
	wire _w25990_ ;
	wire _w25991_ ;
	wire _w25992_ ;
	wire _w25993_ ;
	wire _w25994_ ;
	wire _w25995_ ;
	wire _w25996_ ;
	wire _w25997_ ;
	wire _w25998_ ;
	wire _w25999_ ;
	wire _w26000_ ;
	wire _w26001_ ;
	wire _w26002_ ;
	wire _w26003_ ;
	wire _w26004_ ;
	wire _w26005_ ;
	wire _w26006_ ;
	wire _w26007_ ;
	wire _w26008_ ;
	wire _w26009_ ;
	wire _w26010_ ;
	wire _w26011_ ;
	wire _w26012_ ;
	wire _w26013_ ;
	wire _w26014_ ;
	wire _w26015_ ;
	wire _w26016_ ;
	wire _w26017_ ;
	wire _w26018_ ;
	wire _w26019_ ;
	wire _w26020_ ;
	wire _w26021_ ;
	wire _w26022_ ;
	wire _w26023_ ;
	wire _w26024_ ;
	wire _w26025_ ;
	wire _w26026_ ;
	wire _w26027_ ;
	wire _w26028_ ;
	wire _w26029_ ;
	wire _w26030_ ;
	wire _w26031_ ;
	wire _w26032_ ;
	wire _w26033_ ;
	wire _w26034_ ;
	wire _w26035_ ;
	wire _w26036_ ;
	wire _w26037_ ;
	wire _w26038_ ;
	wire _w26039_ ;
	wire _w26040_ ;
	wire _w26041_ ;
	wire _w26042_ ;
	wire _w26043_ ;
	wire _w26044_ ;
	wire _w26045_ ;
	wire _w26046_ ;
	wire _w26047_ ;
	wire _w26048_ ;
	wire _w26049_ ;
	wire _w26050_ ;
	wire _w26051_ ;
	wire _w26052_ ;
	wire _w26053_ ;
	wire _w26054_ ;
	wire _w26055_ ;
	wire _w26056_ ;
	wire _w26057_ ;
	wire _w26058_ ;
	wire _w26059_ ;
	wire _w26060_ ;
	wire _w26061_ ;
	wire _w26062_ ;
	wire _w26063_ ;
	wire _w26064_ ;
	wire _w26065_ ;
	wire _w26066_ ;
	wire _w26067_ ;
	wire _w26068_ ;
	wire _w26069_ ;
	wire _w26070_ ;
	wire _w26071_ ;
	wire _w26072_ ;
	wire _w26073_ ;
	wire _w26074_ ;
	wire _w26075_ ;
	wire _w26076_ ;
	wire _w26077_ ;
	wire _w26078_ ;
	wire _w26079_ ;
	wire _w26080_ ;
	wire _w26081_ ;
	wire _w26082_ ;
	wire _w26083_ ;
	wire _w26084_ ;
	wire _w26085_ ;
	wire _w26086_ ;
	wire _w26087_ ;
	wire _w26088_ ;
	wire _w26089_ ;
	wire _w26090_ ;
	wire _w26091_ ;
	wire _w26092_ ;
	wire _w26093_ ;
	wire _w26094_ ;
	wire _w26095_ ;
	wire _w26096_ ;
	wire _w26097_ ;
	wire _w26098_ ;
	wire _w26099_ ;
	wire _w26100_ ;
	wire _w26101_ ;
	wire _w26102_ ;
	wire _w26103_ ;
	wire _w26104_ ;
	wire _w26105_ ;
	wire _w26106_ ;
	wire _w26107_ ;
	wire _w26108_ ;
	wire _w26109_ ;
	wire _w26110_ ;
	wire _w26111_ ;
	wire _w26112_ ;
	wire _w26113_ ;
	wire _w26114_ ;
	wire _w26115_ ;
	wire _w26116_ ;
	wire _w26117_ ;
	wire _w26118_ ;
	wire _w26119_ ;
	wire _w26120_ ;
	wire _w26121_ ;
	wire _w26122_ ;
	wire _w26123_ ;
	wire _w26124_ ;
	wire _w26125_ ;
	wire _w26126_ ;
	wire _w26127_ ;
	wire _w26128_ ;
	wire _w26129_ ;
	wire _w26130_ ;
	wire _w26131_ ;
	wire _w26132_ ;
	wire _w26133_ ;
	wire _w26134_ ;
	wire _w26135_ ;
	wire _w26136_ ;
	wire _w26137_ ;
	wire _w26138_ ;
	wire _w26139_ ;
	wire _w26140_ ;
	wire _w26141_ ;
	wire _w26142_ ;
	wire _w26143_ ;
	wire _w26144_ ;
	wire _w26145_ ;
	wire _w26146_ ;
	wire _w26147_ ;
	wire _w26148_ ;
	wire _w26149_ ;
	wire _w26150_ ;
	wire _w26151_ ;
	wire _w26152_ ;
	wire _w26153_ ;
	wire _w26154_ ;
	wire _w26155_ ;
	wire _w26156_ ;
	wire _w26157_ ;
	wire _w26158_ ;
	wire _w26159_ ;
	wire _w26160_ ;
	wire _w26161_ ;
	wire _w26162_ ;
	wire _w26163_ ;
	wire _w26164_ ;
	wire _w26165_ ;
	wire _w26166_ ;
	wire _w26167_ ;
	wire _w26168_ ;
	wire _w26169_ ;
	wire _w26170_ ;
	wire _w26171_ ;
	wire _w26172_ ;
	wire _w26173_ ;
	wire _w26174_ ;
	wire _w26175_ ;
	wire _w26176_ ;
	wire _w26177_ ;
	wire _w26178_ ;
	wire _w26179_ ;
	wire _w26180_ ;
	wire _w26181_ ;
	wire _w26182_ ;
	wire _w26183_ ;
	wire _w26184_ ;
	wire _w26185_ ;
	wire _w26186_ ;
	wire _w26187_ ;
	wire _w26188_ ;
	wire _w26189_ ;
	wire _w26190_ ;
	wire _w26191_ ;
	wire _w26192_ ;
	wire _w26193_ ;
	wire _w26194_ ;
	wire _w26195_ ;
	wire _w26196_ ;
	wire _w26197_ ;
	wire _w26198_ ;
	wire _w26199_ ;
	wire _w26200_ ;
	wire _w26201_ ;
	wire _w26202_ ;
	wire _w26203_ ;
	wire _w26204_ ;
	wire _w26205_ ;
	wire _w26206_ ;
	wire _w26207_ ;
	wire _w26208_ ;
	wire _w26209_ ;
	wire _w26210_ ;
	wire _w26211_ ;
	wire _w26212_ ;
	wire _w26213_ ;
	wire _w26214_ ;
	wire _w26215_ ;
	wire _w26216_ ;
	wire _w26217_ ;
	wire _w26218_ ;
	wire _w26219_ ;
	wire _w26220_ ;
	wire _w26221_ ;
	wire _w26222_ ;
	wire _w26223_ ;
	wire _w26224_ ;
	wire _w26225_ ;
	wire _w26226_ ;
	wire _w26227_ ;
	wire _w26228_ ;
	wire _w26229_ ;
	wire _w26230_ ;
	wire _w26231_ ;
	wire _w26232_ ;
	wire _w26233_ ;
	wire _w26234_ ;
	wire _w26235_ ;
	wire _w26236_ ;
	wire _w26237_ ;
	wire _w26238_ ;
	wire _w26239_ ;
	wire _w26240_ ;
	wire _w26241_ ;
	wire _w26242_ ;
	wire _w26243_ ;
	wire _w26244_ ;
	wire _w26245_ ;
	wire _w26246_ ;
	wire _w26247_ ;
	wire _w26248_ ;
	wire _w26249_ ;
	wire _w26250_ ;
	wire _w26251_ ;
	wire _w26252_ ;
	wire _w26253_ ;
	wire _w26254_ ;
	wire _w26255_ ;
	wire _w26256_ ;
	wire _w26257_ ;
	wire _w26258_ ;
	wire _w26259_ ;
	wire _w26260_ ;
	wire _w26261_ ;
	wire _w26262_ ;
	wire _w26263_ ;
	wire _w26264_ ;
	wire _w26265_ ;
	wire _w26266_ ;
	wire _w26267_ ;
	wire _w26268_ ;
	wire _w26269_ ;
	wire _w26270_ ;
	wire _w26271_ ;
	wire _w26272_ ;
	wire _w26273_ ;
	wire _w26274_ ;
	wire _w26275_ ;
	wire _w26276_ ;
	wire _w26277_ ;
	wire _w26278_ ;
	wire _w26279_ ;
	wire _w26280_ ;
	wire _w26281_ ;
	wire _w26282_ ;
	wire _w26283_ ;
	wire _w26284_ ;
	wire _w26285_ ;
	wire _w26286_ ;
	wire _w26287_ ;
	wire _w26288_ ;
	wire _w26289_ ;
	wire _w26290_ ;
	wire _w26291_ ;
	wire _w26292_ ;
	wire _w26293_ ;
	wire _w26294_ ;
	wire _w26295_ ;
	wire _w26296_ ;
	wire _w26297_ ;
	wire _w26298_ ;
	wire _w26299_ ;
	wire _w26300_ ;
	wire _w26301_ ;
	wire _w26302_ ;
	wire _w26303_ ;
	wire _w26304_ ;
	wire _w26305_ ;
	wire _w26306_ ;
	wire _w26307_ ;
	wire _w26308_ ;
	wire _w26309_ ;
	wire _w26310_ ;
	wire _w26311_ ;
	wire _w26312_ ;
	wire _w26313_ ;
	wire _w26314_ ;
	wire _w26315_ ;
	wire _w26316_ ;
	wire _w26317_ ;
	wire _w26318_ ;
	wire _w26319_ ;
	wire _w26320_ ;
	wire _w26321_ ;
	wire _w26322_ ;
	wire _w26323_ ;
	wire _w26324_ ;
	wire _w26325_ ;
	wire _w26326_ ;
	wire _w26327_ ;
	wire _w26328_ ;
	wire _w26329_ ;
	wire _w26330_ ;
	wire _w26331_ ;
	wire _w26332_ ;
	wire _w26333_ ;
	wire _w26334_ ;
	wire _w26335_ ;
	wire _w26336_ ;
	wire _w26337_ ;
	wire _w26338_ ;
	wire _w26339_ ;
	wire _w26340_ ;
	wire _w26341_ ;
	wire _w26342_ ;
	wire _w26343_ ;
	wire _w26344_ ;
	wire _w26345_ ;
	wire _w26346_ ;
	wire _w26347_ ;
	wire _w26348_ ;
	wire _w26349_ ;
	wire _w26350_ ;
	wire _w26351_ ;
	wire _w26352_ ;
	wire _w26353_ ;
	wire _w26354_ ;
	wire _w26355_ ;
	wire _w26356_ ;
	wire _w26357_ ;
	wire _w26358_ ;
	wire _w26359_ ;
	wire _w26360_ ;
	wire _w26361_ ;
	wire _w26362_ ;
	wire _w26363_ ;
	wire _w26364_ ;
	wire _w26365_ ;
	wire _w26366_ ;
	wire _w26367_ ;
	wire _w26368_ ;
	wire _w26369_ ;
	wire _w26370_ ;
	wire _w26371_ ;
	wire _w26372_ ;
	wire _w26373_ ;
	wire _w26374_ ;
	wire _w26375_ ;
	wire _w26376_ ;
	wire _w26377_ ;
	wire _w26378_ ;
	wire _w26379_ ;
	wire _w26380_ ;
	wire _w26381_ ;
	wire _w26382_ ;
	wire _w26383_ ;
	wire _w26384_ ;
	wire _w26385_ ;
	wire _w26386_ ;
	wire _w26387_ ;
	wire _w26388_ ;
	wire _w26389_ ;
	wire _w26390_ ;
	wire _w26391_ ;
	wire _w26392_ ;
	wire _w26393_ ;
	wire _w26394_ ;
	wire _w26395_ ;
	wire _w26396_ ;
	wire _w26397_ ;
	wire _w26398_ ;
	wire _w26399_ ;
	wire _w26400_ ;
	wire _w26401_ ;
	wire _w26402_ ;
	wire _w26403_ ;
	wire _w26404_ ;
	wire _w26405_ ;
	wire _w26406_ ;
	wire _w26407_ ;
	wire _w26408_ ;
	wire _w26409_ ;
	wire _w26410_ ;
	wire _w26411_ ;
	wire _w26412_ ;
	wire _w26413_ ;
	wire _w26414_ ;
	wire _w26415_ ;
	wire _w26416_ ;
	wire _w26417_ ;
	wire _w26418_ ;
	wire _w26419_ ;
	wire _w26420_ ;
	wire _w26421_ ;
	wire _w26422_ ;
	wire _w26423_ ;
	wire _w26424_ ;
	wire _w26425_ ;
	wire _w26426_ ;
	wire _w26427_ ;
	wire _w26428_ ;
	wire _w26429_ ;
	wire _w26430_ ;
	wire _w26431_ ;
	wire _w26432_ ;
	wire _w26433_ ;
	wire _w26434_ ;
	wire _w26435_ ;
	wire _w26436_ ;
	wire _w26437_ ;
	wire _w26438_ ;
	wire _w26439_ ;
	wire _w26440_ ;
	wire _w26441_ ;
	wire _w26442_ ;
	wire _w26443_ ;
	wire _w26444_ ;
	wire _w26445_ ;
	wire _w26446_ ;
	wire _w26447_ ;
	wire _w26448_ ;
	wire _w26449_ ;
	wire _w26450_ ;
	wire _w26451_ ;
	wire _w26452_ ;
	wire _w26453_ ;
	wire _w26454_ ;
	wire _w26455_ ;
	wire _w26456_ ;
	wire _w26457_ ;
	wire _w26458_ ;
	wire _w26459_ ;
	wire _w26460_ ;
	wire _w26461_ ;
	wire _w26462_ ;
	wire _w26463_ ;
	wire _w26464_ ;
	wire _w26465_ ;
	wire _w26466_ ;
	wire _w26467_ ;
	wire _w26468_ ;
	wire _w26469_ ;
	wire _w26470_ ;
	wire _w26471_ ;
	wire _w26472_ ;
	wire _w26473_ ;
	wire _w26474_ ;
	wire _w26475_ ;
	wire _w26476_ ;
	wire _w26477_ ;
	wire _w26478_ ;
	wire _w26479_ ;
	wire _w26480_ ;
	wire _w26481_ ;
	wire _w26482_ ;
	wire _w26483_ ;
	wire _w26484_ ;
	wire _w26485_ ;
	wire _w26486_ ;
	wire _w26487_ ;
	wire _w26488_ ;
	wire _w26489_ ;
	wire _w26490_ ;
	wire _w26491_ ;
	wire _w26492_ ;
	wire _w26493_ ;
	wire _w26494_ ;
	wire _w26495_ ;
	wire _w26496_ ;
	wire _w26497_ ;
	wire _w26498_ ;
	wire _w26499_ ;
	wire _w26500_ ;
	wire _w26501_ ;
	wire _w26502_ ;
	wire _w26503_ ;
	wire _w26504_ ;
	wire _w26505_ ;
	wire _w26506_ ;
	wire _w26507_ ;
	wire _w26508_ ;
	wire _w26509_ ;
	wire _w26510_ ;
	wire _w26511_ ;
	wire _w26512_ ;
	wire _w26513_ ;
	wire _w26514_ ;
	wire _w26515_ ;
	wire _w26516_ ;
	wire _w26517_ ;
	wire _w26518_ ;
	wire _w26519_ ;
	wire _w26520_ ;
	wire _w26521_ ;
	wire _w26522_ ;
	wire _w26523_ ;
	wire _w26524_ ;
	wire _w26525_ ;
	wire _w26526_ ;
	wire _w26527_ ;
	wire _w26528_ ;
	wire _w26529_ ;
	wire _w26530_ ;
	wire _w26531_ ;
	wire _w26532_ ;
	wire _w26533_ ;
	wire _w26534_ ;
	wire _w26535_ ;
	wire _w26536_ ;
	wire _w26537_ ;
	wire _w26538_ ;
	wire _w26539_ ;
	wire _w26540_ ;
	wire _w26541_ ;
	wire _w26542_ ;
	wire _w26543_ ;
	wire _w26544_ ;
	wire _w26545_ ;
	wire _w26546_ ;
	wire _w26547_ ;
	wire _w26548_ ;
	wire _w26549_ ;
	wire _w26550_ ;
	wire _w26551_ ;
	wire _w26552_ ;
	wire _w26553_ ;
	wire _w26554_ ;
	wire _w26555_ ;
	wire _w26556_ ;
	wire _w26557_ ;
	wire _w26558_ ;
	wire _w26559_ ;
	wire _w26560_ ;
	wire _w26561_ ;
	wire _w26562_ ;
	wire _w26563_ ;
	wire _w26564_ ;
	wire _w26565_ ;
	wire _w26566_ ;
	wire _w26567_ ;
	wire _w26568_ ;
	wire _w26569_ ;
	wire _w26570_ ;
	wire _w26571_ ;
	wire _w26572_ ;
	wire _w26573_ ;
	wire _w26574_ ;
	wire _w26575_ ;
	wire _w26576_ ;
	wire _w26577_ ;
	wire _w26578_ ;
	wire _w26579_ ;
	LUT4 #(
		.INIT('hc963)
	) name0 (
		decrypt_pad,
		\u1_R3_reg[1]/NET0131 ,
		\u1_uk_K_r3_reg[12]/NET0131 ,
		\u1_uk_K_r3_reg[3]/NET0131 ,
		_w5827_
	);
	LUT4 #(
		.INIT('hc693)
	) name1 (
		decrypt_pad,
		\u1_R3_reg[32]/NET0131 ,
		\u1_uk_K_r3_reg[39]/NET0131 ,
		\u1_uk_K_r3_reg[48]/NET0131 ,
		_w5828_
	);
	LUT4 #(
		.INIT('hc963)
	) name2 (
		decrypt_pad,
		\u1_R3_reg[5]/NET0131 ,
		\u1_uk_K_r3_reg[10]/NET0131 ,
		\u1_uk_K_r3_reg[33]/NET0131 ,
		_w5829_
	);
	LUT3 #(
		.INIT('h80)
	) name3 (
		_w5828_,
		_w5827_,
		_w5829_,
		_w5830_
	);
	LUT3 #(
		.INIT('h7d)
	) name4 (
		_w5828_,
		_w5827_,
		_w5829_,
		_w5831_
	);
	LUT4 #(
		.INIT('hc693)
	) name5 (
		decrypt_pad,
		\u1_R3_reg[2]/NET0131 ,
		\u1_uk_K_r3_reg[18]/NET0131 ,
		\u1_uk_K_r3_reg[27]/NET0131 ,
		_w5832_
	);
	LUT4 #(
		.INIT('h0440)
	) name6 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w5833_
	);
	LUT4 #(
		.INIT('hc693)
	) name7 (
		decrypt_pad,
		\u1_R3_reg[3]/NET0131 ,
		\u1_uk_K_r3_reg[27]/NET0131 ,
		\u1_uk_K_r3_reg[4]/NET0131 ,
		_w5834_
	);
	LUT3 #(
		.INIT('h40)
	) name8 (
		_w5833_,
		_w5831_,
		_w5834_,
		_w5835_
	);
	LUT3 #(
		.INIT('h21)
	) name9 (
		_w5828_,
		_w5827_,
		_w5829_,
		_w5836_
	);
	LUT4 #(
		.INIT('h00fe)
	) name10 (
		_w5828_,
		_w5832_,
		_w5829_,
		_w5834_,
		_w5837_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w5836_,
		_w5837_,
		_w5838_
	);
	LUT4 #(
		.INIT('h0080)
	) name12 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w5839_
	);
	LUT4 #(
		.INIT('hc963)
	) name13 (
		decrypt_pad,
		\u1_R3_reg[4]/NET0131 ,
		\u1_uk_K_r3_reg[39]/NET0131 ,
		\u1_uk_K_r3_reg[5]/NET0131 ,
		_w5840_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w5828_,
		_w5827_,
		_w5841_
	);
	LUT4 #(
		.INIT('h1000)
	) name15 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w5842_
	);
	LUT3 #(
		.INIT('h01)
	) name16 (
		_w5839_,
		_w5840_,
		_w5842_,
		_w5843_
	);
	LUT3 #(
		.INIT('he0)
	) name17 (
		_w5835_,
		_w5838_,
		_w5843_,
		_w5844_
	);
	LUT4 #(
		.INIT('h005e)
	) name18 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5834_,
		_w5845_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w5828_,
		_w5829_,
		_w5846_
	);
	LUT4 #(
		.INIT('h0200)
	) name20 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w5847_
	);
	LUT4 #(
		.INIT('hab00)
	) name21 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5834_,
		_w5848_
	);
	LUT3 #(
		.INIT('h45)
	) name22 (
		_w5845_,
		_w5847_,
		_w5848_,
		_w5849_
	);
	LUT4 #(
		.INIT('h0008)
	) name23 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w5850_
	);
	LUT3 #(
		.INIT('h80)
	) name24 (
		_w5827_,
		_w5832_,
		_w5829_,
		_w5851_
	);
	LUT4 #(
		.INIT('h7f00)
	) name25 (
		_w5827_,
		_w5832_,
		_w5829_,
		_w5840_,
		_w5852_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w5850_,
		_w5852_,
		_w5853_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w5849_,
		_w5853_,
		_w5854_
	);
	LUT3 #(
		.INIT('ha9)
	) name28 (
		\u1_L3_reg[17]/NET0131 ,
		_w5844_,
		_w5854_,
		_w5855_
	);
	LUT4 #(
		.INIT('hc963)
	) name29 (
		decrypt_pad,
		\u2_R13_reg[27]/P0001 ,
		\u2_uk_K_r13_reg[45]/NET0131 ,
		\u2_uk_K_r13_reg[7]/NET0131 ,
		_w5856_
	);
	LUT4 #(
		.INIT('hc963)
	) name30 (
		decrypt_pad,
		\u2_R13_reg[24]/NET0131 ,
		\u2_uk_K_r13_reg[43]/NET0131 ,
		\u2_uk_K_r13_reg[9]/NET0131 ,
		_w5857_
	);
	LUT4 #(
		.INIT('hc693)
	) name31 (
		decrypt_pad,
		\u2_R13_reg[26]/NET0131 ,
		\u2_uk_K_r13_reg[29]/NET0131 ,
		\u2_uk_K_r13_reg[8]/NET0131 ,
		_w5858_
	);
	LUT4 #(
		.INIT('hc963)
	) name32 (
		decrypt_pad,
		\u2_R13_reg[25]/NET0131 ,
		\u2_uk_K_r13_reg[23]/NET0131 ,
		\u2_uk_K_r13_reg[44]/NET0131 ,
		_w5859_
	);
	LUT4 #(
		.INIT('hc693)
	) name33 (
		decrypt_pad,
		\u2_R13_reg[29]/NET0131 ,
		\u2_uk_K_r13_reg[45]/NET0131 ,
		\u2_uk_K_r13_reg[51]/NET0131 ,
		_w5860_
	);
	LUT4 #(
		.INIT('hb7f7)
	) name34 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w5861_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		_w5856_,
		_w5861_,
		_w5862_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		_w5860_,
		_w5856_,
		_w5863_
	);
	LUT3 #(
		.INIT('h34)
	) name37 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5864_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w5863_,
		_w5864_,
		_w5865_
	);
	LUT4 #(
		.INIT('h0200)
	) name39 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w5866_
	);
	LUT4 #(
		.INIT('h0001)
	) name40 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w5867_
	);
	LUT4 #(
		.INIT('hc963)
	) name41 (
		decrypt_pad,
		\u2_R13_reg[28]/NET0131 ,
		\u2_uk_K_r13_reg[28]/NET0131 ,
		\u2_uk_K_r13_reg[49]/NET0131 ,
		_w5868_
	);
	LUT3 #(
		.INIT('h10)
	) name42 (
		_w5867_,
		_w5866_,
		_w5868_,
		_w5869_
	);
	LUT3 #(
		.INIT('h10)
	) name43 (
		_w5865_,
		_w5862_,
		_w5869_,
		_w5870_
	);
	LUT3 #(
		.INIT('hab)
	) name44 (
		_w5857_,
		_w5859_,
		_w5860_,
		_w5871_
	);
	LUT4 #(
		.INIT('h000d)
	) name45 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w5872_
	);
	LUT3 #(
		.INIT('h0b)
	) name46 (
		_w5858_,
		_w5860_,
		_w5856_,
		_w5873_
	);
	LUT3 #(
		.INIT('h40)
	) name47 (
		_w5872_,
		_w5871_,
		_w5873_,
		_w5874_
	);
	LUT4 #(
		.INIT('hddad)
	) name48 (
		_w5857_,
		_w5859_,
		_w5860_,
		_w5856_,
		_w5875_
	);
	LUT4 #(
		.INIT('h9000)
	) name49 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w5876_
	);
	LUT4 #(
		.INIT('h0302)
	) name50 (
		_w5858_,
		_w5868_,
		_w5876_,
		_w5875_,
		_w5877_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w5874_,
		_w5877_,
		_w5878_
	);
	LUT4 #(
		.INIT('h0020)
	) name52 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w5879_
	);
	LUT4 #(
		.INIT('h0004)
	) name53 (
		_w5866_,
		_w5856_,
		_w5872_,
		_w5879_,
		_w5880_
	);
	LUT4 #(
		.INIT('hff90)
	) name54 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5856_,
		_w5881_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w5880_,
		_w5881_,
		_w5882_
	);
	LUT4 #(
		.INIT('h55a9)
	) name56 (
		\u2_L13_reg[22]/NET0131 ,
		_w5870_,
		_w5878_,
		_w5882_,
		_w5883_
	);
	LUT4 #(
		.INIT('hc693)
	) name57 (
		decrypt_pad,
		\u2_R13_reg[4]/NET0131 ,
		\u2_uk_K_r13_reg[20]/NET0131 ,
		\u2_uk_K_r13_reg[24]/NET0131 ,
		_w5884_
	);
	LUT4 #(
		.INIT('hc693)
	) name58 (
		decrypt_pad,
		\u2_R13_reg[3]/NET0131 ,
		\u2_uk_K_r13_reg[10]/NET0131 ,
		\u2_uk_K_r13_reg[46]/NET0131 ,
		_w5885_
	);
	LUT4 #(
		.INIT('hc693)
	) name59 (
		decrypt_pad,
		\u2_R13_reg[1]/NET0131 ,
		\u2_uk_K_r13_reg[18]/NET0131 ,
		\u2_uk_K_r13_reg[54]/NET0131 ,
		_w5886_
	);
	LUT4 #(
		.INIT('hc963)
	) name60 (
		decrypt_pad,
		\u2_R13_reg[5]/NET0131 ,
		\u2_uk_K_r13_reg[27]/NET0131 ,
		\u2_uk_K_r13_reg[48]/NET0131 ,
		_w5887_
	);
	LUT4 #(
		.INIT('hc963)
	) name61 (
		decrypt_pad,
		\u2_R13_reg[32]/NET0131 ,
		\u2_uk_K_r13_reg[33]/NET0131 ,
		\u2_uk_K_r13_reg[54]/NET0131 ,
		_w5888_
	);
	LUT4 #(
		.INIT('hc963)
	) name62 (
		decrypt_pad,
		\u2_R13_reg[2]/NET0131 ,
		\u2_uk_K_r13_reg[12]/NET0131 ,
		\u2_uk_K_r13_reg[33]/NET0131 ,
		_w5889_
	);
	LUT4 #(
		.INIT('hb8bb)
	) name63 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w5890_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		_w5885_,
		_w5890_,
		_w5891_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		_w5887_,
		_w5888_,
		_w5892_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		_w5885_,
		_w5889_,
		_w5893_
	);
	LUT3 #(
		.INIT('hc4)
	) name67 (
		_w5885_,
		_w5886_,
		_w5889_,
		_w5894_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w5886_,
		_w5889_,
		_w5895_
	);
	LUT4 #(
		.INIT('h4340)
	) name69 (
		_w5885_,
		_w5886_,
		_w5888_,
		_w5889_,
		_w5896_
	);
	LUT4 #(
		.INIT('h0010)
	) name70 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w5897_
	);
	LUT4 #(
		.INIT('h0301)
	) name71 (
		_w5892_,
		_w5896_,
		_w5897_,
		_w5894_,
		_w5898_
	);
	LUT3 #(
		.INIT('h8a)
	) name72 (
		_w5884_,
		_w5891_,
		_w5898_,
		_w5899_
	);
	LUT3 #(
		.INIT('h10)
	) name73 (
		_w5886_,
		_w5887_,
		_w5889_,
		_w5900_
	);
	LUT4 #(
		.INIT('heff4)
	) name74 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w5901_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w5885_,
		_w5901_,
		_w5902_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w5885_,
		_w5886_,
		_w5903_
	);
	LUT2 #(
		.INIT('h6)
	) name77 (
		_w5887_,
		_w5888_,
		_w5904_
	);
	LUT3 #(
		.INIT('h60)
	) name78 (
		_w5887_,
		_w5888_,
		_w5889_,
		_w5905_
	);
	LUT3 #(
		.INIT('h43)
	) name79 (
		_w5885_,
		_w5886_,
		_w5887_,
		_w5906_
	);
	LUT3 #(
		.INIT('h09)
	) name80 (
		_w5887_,
		_w5888_,
		_w5889_,
		_w5907_
	);
	LUT4 #(
		.INIT('h7077)
	) name81 (
		_w5903_,
		_w5905_,
		_w5906_,
		_w5907_,
		_w5908_
	);
	LUT3 #(
		.INIT('h45)
	) name82 (
		_w5884_,
		_w5902_,
		_w5908_,
		_w5909_
	);
	LUT4 #(
		.INIT('h7bdd)
	) name83 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w5910_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w5885_,
		_w5910_,
		_w5911_
	);
	LUT3 #(
		.INIT('h02)
	) name85 (
		_w5885_,
		_w5887_,
		_w5888_,
		_w5912_
	);
	LUT4 #(
		.INIT('h0020)
	) name86 (
		_w5885_,
		_w5886_,
		_w5888_,
		_w5889_,
		_w5913_
	);
	LUT3 #(
		.INIT('h07)
	) name87 (
		_w5895_,
		_w5912_,
		_w5913_,
		_w5914_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w5911_,
		_w5914_,
		_w5915_
	);
	LUT4 #(
		.INIT('h5655)
	) name89 (
		\u2_L13_reg[31]/NET0131 ,
		_w5909_,
		_w5899_,
		_w5915_,
		_w5916_
	);
	LUT4 #(
		.INIT('hc693)
	) name90 (
		decrypt_pad,
		\u2_R13_reg[23]/NET0131 ,
		\u2_uk_K_r13_reg[16]/NET0131 ,
		\u2_uk_K_r13_reg[50]/NET0131 ,
		_w5917_
	);
	LUT4 #(
		.INIT('hc693)
	) name91 (
		decrypt_pad,
		\u2_R13_reg[22]/NET0131 ,
		\u2_uk_K_r13_reg[31]/NET0131 ,
		\u2_uk_K_r13_reg[37]/NET0131 ,
		_w5918_
	);
	LUT4 #(
		.INIT('hc963)
	) name92 (
		decrypt_pad,
		\u2_R13_reg[20]/NET0131 ,
		\u2_uk_K_r13_reg[0]/NET0131 ,
		\u2_uk_K_r13_reg[21]/NET0131 ,
		_w5919_
	);
	LUT4 #(
		.INIT('hc963)
	) name93 (
		decrypt_pad,
		\u2_R13_reg[25]/NET0131 ,
		\u2_uk_K_r13_reg[16]/NET0131 ,
		\u2_uk_K_r13_reg[37]/NET0131 ,
		_w5920_
	);
	LUT4 #(
		.INIT('hc963)
	) name94 (
		decrypt_pad,
		\u2_R13_reg[21]/NET0131 ,
		\u2_uk_K_r13_reg[15]/NET0131 ,
		\u2_uk_K_r13_reg[36]/NET0131 ,
		_w5921_
	);
	LUT3 #(
		.INIT('h20)
	) name95 (
		_w5919_,
		_w5921_,
		_w5920_,
		_w5922_
	);
	LUT4 #(
		.INIT('h168a)
	) name96 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w5923_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w5917_,
		_w5923_,
		_w5924_
	);
	LUT4 #(
		.INIT('hc963)
	) name98 (
		decrypt_pad,
		\u2_R13_reg[24]/NET0131 ,
		\u2_uk_K_r13_reg[21]/NET0131 ,
		\u2_uk_K_r13_reg[42]/NET0131 ,
		_w5925_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name99 (
		_w5917_,
		_w5918_,
		_w5919_,
		_w5921_,
		_w5926_
	);
	LUT4 #(
		.INIT('h0004)
	) name100 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w5927_
	);
	LUT4 #(
		.INIT('h3ffb)
	) name101 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w5928_
	);
	LUT3 #(
		.INIT('h2a)
	) name102 (
		_w5925_,
		_w5926_,
		_w5928_,
		_w5929_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w5924_,
		_w5929_,
		_w5930_
	);
	LUT4 #(
		.INIT('h0040)
	) name104 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w5931_
	);
	LUT4 #(
		.INIT('h0800)
	) name105 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w5932_
	);
	LUT4 #(
		.INIT('h0200)
	) name106 (
		_w5917_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w5933_
	);
	LUT3 #(
		.INIT('h01)
	) name107 (
		_w5932_,
		_w5933_,
		_w5931_,
		_w5934_
	);
	LUT4 #(
		.INIT('h1400)
	) name108 (
		_w5917_,
		_w5918_,
		_w5919_,
		_w5921_,
		_w5935_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w5917_,
		_w5918_,
		_w5936_
	);
	LUT4 #(
		.INIT('h0080)
	) name110 (
		_w5917_,
		_w5918_,
		_w5919_,
		_w5921_,
		_w5937_
	);
	LUT4 #(
		.INIT('h0010)
	) name111 (
		_w5917_,
		_w5918_,
		_w5919_,
		_w5920_,
		_w5938_
	);
	LUT4 #(
		.INIT('hfded)
	) name112 (
		_w5917_,
		_w5918_,
		_w5919_,
		_w5920_,
		_w5939_
	);
	LUT3 #(
		.INIT('h10)
	) name113 (
		_w5935_,
		_w5937_,
		_w5939_,
		_w5940_
	);
	LUT3 #(
		.INIT('h15)
	) name114 (
		_w5925_,
		_w5934_,
		_w5940_,
		_w5941_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name115 (
		_w5917_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w5942_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w5918_,
		_w5942_,
		_w5943_
	);
	LUT4 #(
		.INIT('h0010)
	) name117 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w5944_
	);
	LUT4 #(
		.INIT('h77ef)
	) name118 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w5945_
	);
	LUT3 #(
		.INIT('h01)
	) name119 (
		_w5919_,
		_w5921_,
		_w5920_,
		_w5946_
	);
	LUT4 #(
		.INIT('he4f5)
	) name120 (
		_w5917_,
		_w5918_,
		_w5945_,
		_w5946_,
		_w5947_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		_w5943_,
		_w5947_,
		_w5948_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name122 (
		\u2_L13_reg[11]/NET0131 ,
		_w5941_,
		_w5930_,
		_w5948_,
		_w5949_
	);
	LUT4 #(
		.INIT('hc963)
	) name123 (
		decrypt_pad,
		\u2_R13_reg[31]/P0001 ,
		\u2_uk_K_r13_reg[42]/NET0131 ,
		\u2_uk_K_r13_reg[8]/NET0131 ,
		_w5950_
	);
	LUT4 #(
		.INIT('hc963)
	) name124 (
		decrypt_pad,
		\u2_R13_reg[30]/NET0131 ,
		\u2_uk_K_r13_reg[30]/NET0131 ,
		\u2_uk_K_r13_reg[51]/NET0131 ,
		_w5951_
	);
	LUT4 #(
		.INIT('hc963)
	) name125 (
		decrypt_pad,
		\u2_R13_reg[29]/NET0131 ,
		\u2_uk_K_r13_reg[29]/NET0131 ,
		\u2_uk_K_r13_reg[50]/NET0131 ,
		_w5952_
	);
	LUT4 #(
		.INIT('hc693)
	) name126 (
		decrypt_pad,
		\u2_R13_reg[28]/NET0131 ,
		\u2_uk_K_r13_reg[23]/NET0131 ,
		\u2_uk_K_r13_reg[2]/NET0131 ,
		_w5953_
	);
	LUT3 #(
		.INIT('h01)
	) name127 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5954_
	);
	LUT4 #(
		.INIT('h5554)
	) name128 (
		_w5950_,
		_w5951_,
		_w5952_,
		_w5953_,
		_w5955_
	);
	LUT4 #(
		.INIT('hc963)
	) name129 (
		decrypt_pad,
		\u2_R13_reg[1]/NET0131 ,
		\u2_uk_K_r13_reg[14]/NET0131 ,
		\u2_uk_K_r13_reg[35]/NET0131 ,
		_w5956_
	);
	LUT4 #(
		.INIT('h0040)
	) name130 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w5957_
	);
	LUT4 #(
		.INIT('h509c)
	) name131 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w5958_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w5952_,
		_w5956_,
		_w5959_
	);
	LUT4 #(
		.INIT('h0800)
	) name133 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w5960_
	);
	LUT4 #(
		.INIT('h001b)
	) name134 (
		_w5950_,
		_w5954_,
		_w5958_,
		_w5960_,
		_w5961_
	);
	LUT4 #(
		.INIT('hc693)
	) name135 (
		decrypt_pad,
		\u2_R13_reg[32]/NET0131 ,
		\u2_uk_K_r13_reg[14]/NET0131 ,
		\u2_uk_K_r13_reg[52]/NET0131 ,
		_w5962_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w5961_,
		_w5962_,
		_w5963_
	);
	LUT4 #(
		.INIT('h0001)
	) name137 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w5964_
	);
	LUT4 #(
		.INIT('h0200)
	) name138 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w5965_
	);
	LUT4 #(
		.INIT('hedf7)
	) name139 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w5966_
	);
	LUT3 #(
		.INIT('h20)
	) name140 (
		_w5950_,
		_w5964_,
		_w5966_,
		_w5967_
	);
	LUT4 #(
		.INIT('h2000)
	) name141 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5962_,
		_w5968_
	);
	LUT3 #(
		.INIT('h01)
	) name142 (
		_w5950_,
		_w5957_,
		_w5968_,
		_w5969_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w5967_,
		_w5969_,
		_w5970_
	);
	LUT4 #(
		.INIT('h0020)
	) name144 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w5971_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name145 (
		_w5950_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w5972_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		_w5951_,
		_w5953_,
		_w5973_
	);
	LUT3 #(
		.INIT('h02)
	) name147 (
		_w5951_,
		_w5953_,
		_w5956_,
		_w5974_
	);
	LUT3 #(
		.INIT('h15)
	) name148 (
		_w5950_,
		_w5952_,
		_w5956_,
		_w5975_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name149 (
		_w5971_,
		_w5972_,
		_w5974_,
		_w5975_,
		_w5976_
	);
	LUT3 #(
		.INIT('h10)
	) name150 (
		_w5950_,
		_w5951_,
		_w5953_,
		_w5977_
	);
	LUT4 #(
		.INIT('h8000)
	) name151 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w5978_
	);
	LUT3 #(
		.INIT('h01)
	) name152 (
		_w5957_,
		_w5977_,
		_w5978_,
		_w5979_
	);
	LUT3 #(
		.INIT('h45)
	) name153 (
		_w5962_,
		_w5976_,
		_w5979_,
		_w5980_
	);
	LUT4 #(
		.INIT('haaa9)
	) name154 (
		\u2_L13_reg[5]/NET0131 ,
		_w5963_,
		_w5970_,
		_w5980_,
		_w5981_
	);
	LUT4 #(
		.INIT('hc963)
	) name155 (
		decrypt_pad,
		\u2_R13_reg[16]/NET0131 ,
		\u2_uk_K_r13_reg[26]/NET0131 ,
		\u2_uk_K_r13_reg[47]/NET0131 ,
		_w5982_
	);
	LUT4 #(
		.INIT('hc963)
	) name156 (
		decrypt_pad,
		\u2_R13_reg[14]/NET0131 ,
		\u2_uk_K_r13_reg[10]/NET0131 ,
		\u2_uk_K_r13_reg[6]/NET0131 ,
		_w5983_
	);
	LUT4 #(
		.INIT('hc963)
	) name157 (
		decrypt_pad,
		\u2_R13_reg[15]/NET0131 ,
		\u2_uk_K_r13_reg[18]/NET0131 ,
		\u2_uk_K_r13_reg[39]/NET0131 ,
		_w5984_
	);
	LUT4 #(
		.INIT('hc693)
	) name158 (
		decrypt_pad,
		\u2_R13_reg[12]/NET0131 ,
		\u2_uk_K_r13_reg[11]/NET0131 ,
		\u2_uk_K_r13_reg[47]/NET0131 ,
		_w5985_
	);
	LUT4 #(
		.INIT('hc693)
	) name159 (
		decrypt_pad,
		\u2_R13_reg[17]/NET0131 ,
		\u2_uk_K_r13_reg[27]/NET0131 ,
		\u2_uk_K_r13_reg[6]/NET0131 ,
		_w5986_
	);
	LUT4 #(
		.INIT('hc963)
	) name160 (
		decrypt_pad,
		\u2_R13_reg[13]/NET0131 ,
		\u2_uk_K_r13_reg[41]/NET0131 ,
		\u2_uk_K_r13_reg[5]/NET0131 ,
		_w5987_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		_w5987_,
		_w5984_,
		_w5988_
	);
	LUT3 #(
		.INIT('h8a)
	) name162 (
		_w5985_,
		_w5987_,
		_w5984_,
		_w5989_
	);
	LUT4 #(
		.INIT('h2757)
	) name163 (
		_w5985_,
		_w5987_,
		_w5986_,
		_w5984_,
		_w5990_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w5983_,
		_w5990_,
		_w5991_
	);
	LUT3 #(
		.INIT('h8a)
	) name165 (
		_w5985_,
		_w5983_,
		_w5986_,
		_w5992_
	);
	LUT4 #(
		.INIT('h0001)
	) name166 (
		_w5985_,
		_w5987_,
		_w5986_,
		_w5984_,
		_w5993_
	);
	LUT4 #(
		.INIT('h0040)
	) name167 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w5994_
	);
	LUT4 #(
		.INIT('hffbe)
	) name168 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w5995_
	);
	LUT4 #(
		.INIT('h1300)
	) name169 (
		_w5992_,
		_w5993_,
		_w5988_,
		_w5995_,
		_w5996_
	);
	LUT3 #(
		.INIT('h45)
	) name170 (
		_w5982_,
		_w5991_,
		_w5996_,
		_w5997_
	);
	LUT4 #(
		.INIT('h9000)
	) name171 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w5998_
	);
	LUT4 #(
		.INIT('h0400)
	) name172 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w5999_
	);
	LUT4 #(
		.INIT('h6b5d)
	) name173 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w6000_
	);
	LUT3 #(
		.INIT('h0b)
	) name174 (
		_w5998_,
		_w5984_,
		_w6000_,
		_w6001_
	);
	LUT4 #(
		.INIT('h2e00)
	) name175 (
		_w5985_,
		_w5987_,
		_w5986_,
		_w5984_,
		_w6002_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		_w5992_,
		_w6002_,
		_w6003_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name177 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w6004_
	);
	LUT2 #(
		.INIT('h9)
	) name178 (
		_w5985_,
		_w5983_,
		_w6005_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w5987_,
		_w5984_,
		_w6006_
	);
	LUT4 #(
		.INIT('h8a00)
	) name180 (
		_w5987_,
		_w5983_,
		_w5986_,
		_w5984_,
		_w6007_
	);
	LUT4 #(
		.INIT('he0ee)
	) name181 (
		_w5984_,
		_w6004_,
		_w6005_,
		_w6007_,
		_w6008_
	);
	LUT4 #(
		.INIT('h5700)
	) name182 (
		_w5982_,
		_w6001_,
		_w6003_,
		_w6008_,
		_w6009_
	);
	LUT3 #(
		.INIT('h65)
	) name183 (
		\u2_L13_reg[10]/NET0131 ,
		_w5997_,
		_w6009_,
		_w6010_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name184 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6011_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		_w5856_,
		_w6011_,
		_w6012_
	);
	LUT4 #(
		.INIT('h1428)
	) name186 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6013_
	);
	LUT4 #(
		.INIT('h00d0)
	) name187 (
		_w5866_,
		_w5856_,
		_w5868_,
		_w6013_,
		_w6014_
	);
	LUT4 #(
		.INIT('hef00)
	) name188 (
		_w5857_,
		_w5859_,
		_w5860_,
		_w5856_,
		_w6015_
	);
	LUT2 #(
		.INIT('h6)
	) name189 (
		_w5859_,
		_w5860_,
		_w6016_
	);
	LUT3 #(
		.INIT('h07)
	) name190 (
		_w5858_,
		_w5857_,
		_w5856_,
		_w6017_
	);
	LUT3 #(
		.INIT('h15)
	) name191 (
		_w6015_,
		_w6016_,
		_w6017_,
		_w6018_
	);
	LUT4 #(
		.INIT('h2014)
	) name192 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6019_
	);
	LUT4 #(
		.INIT('h0800)
	) name193 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6020_
	);
	LUT4 #(
		.INIT('h0002)
	) name194 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6021_
	);
	LUT4 #(
		.INIT('h0001)
	) name195 (
		_w5868_,
		_w6019_,
		_w6020_,
		_w6021_,
		_w6022_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name196 (
		_w6012_,
		_w6014_,
		_w6018_,
		_w6022_,
		_w6023_
	);
	LUT2 #(
		.INIT('h6)
	) name197 (
		\u2_L13_reg[12]/NET0131 ,
		_w6023_,
		_w6024_
	);
	LUT4 #(
		.INIT('hc693)
	) name198 (
		decrypt_pad,
		\u2_R13_reg[20]/NET0131 ,
		\u2_uk_K_r13_reg[30]/NET0131 ,
		\u2_uk_K_r13_reg[9]/NET0131 ,
		_w6025_
	);
	LUT4 #(
		.INIT('hc693)
	) name199 (
		decrypt_pad,
		\u2_R13_reg[19]/NET0131 ,
		\u2_uk_K_r13_reg[15]/NET0131 ,
		\u2_uk_K_r13_reg[49]/NET0131 ,
		_w6026_
	);
	LUT4 #(
		.INIT('hc693)
	) name200 (
		decrypt_pad,
		\u2_R13_reg[18]/NET0131 ,
		\u2_uk_K_r13_reg[28]/NET0131 ,
		\u2_uk_K_r13_reg[7]/NET0131 ,
		_w6027_
	);
	LUT4 #(
		.INIT('hc693)
	) name201 (
		decrypt_pad,
		\u2_R13_reg[17]/NET0131 ,
		\u2_uk_K_r13_reg[38]/NET0131 ,
		\u2_uk_K_r13_reg[44]/NET0131 ,
		_w6028_
	);
	LUT4 #(
		.INIT('hc963)
	) name202 (
		decrypt_pad,
		\u2_R13_reg[16]/NET0131 ,
		\u2_uk_K_r13_reg[22]/NET0131 ,
		\u2_uk_K_r13_reg[43]/NET0131 ,
		_w6029_
	);
	LUT4 #(
		.INIT('hc693)
	) name203 (
		decrypt_pad,
		\u2_R13_reg[21]/NET0131 ,
		\u2_uk_K_r13_reg[0]/NET0131 ,
		\u2_uk_K_r13_reg[38]/NET0131 ,
		_w6030_
	);
	LUT3 #(
		.INIT('h80)
	) name204 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6031_
	);
	LUT4 #(
		.INIT('h0080)
	) name205 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6032_
	);
	LUT4 #(
		.INIT('h0004)
	) name206 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6033_
	);
	LUT3 #(
		.INIT('h20)
	) name207 (
		_w6028_,
		_w6030_,
		_w6027_,
		_w6034_
	);
	LUT4 #(
		.INIT('he56b)
	) name208 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6035_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		_w6026_,
		_w6035_,
		_w6036_
	);
	LUT4 #(
		.INIT('h4000)
	) name210 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6037_
	);
	LUT4 #(
		.INIT('h30d0)
	) name211 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6038_
	);
	LUT4 #(
		.INIT('h0002)
	) name212 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6039_
	);
	LUT3 #(
		.INIT('hd0)
	) name213 (
		_w6029_,
		_w6030_,
		_w6026_,
		_w6040_
	);
	LUT4 #(
		.INIT('h4544)
	) name214 (
		_w6038_,
		_w6039_,
		_w6034_,
		_w6040_,
		_w6041_
	);
	LUT4 #(
		.INIT('h5554)
	) name215 (
		_w6025_,
		_w6037_,
		_w6041_,
		_w6036_,
		_w6042_
	);
	LUT4 #(
		.INIT('hc727)
	) name216 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6043_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w6043_,
		_w6026_,
		_w6044_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w6027_,
		_w6026_,
		_w6045_
	);
	LUT3 #(
		.INIT('hde)
	) name219 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6046_
	);
	LUT2 #(
		.INIT('h2)
	) name220 (
		_w6045_,
		_w6046_,
		_w6047_
	);
	LUT4 #(
		.INIT('h0048)
	) name221 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6048_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		_w6027_,
		_w6026_,
		_w6049_
	);
	LUT4 #(
		.INIT('h0400)
	) name223 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6050_
	);
	LUT4 #(
		.INIT('h0015)
	) name224 (
		_w6048_,
		_w6031_,
		_w6049_,
		_w6050_,
		_w6051_
	);
	LUT4 #(
		.INIT('hef00)
	) name225 (
		_w6044_,
		_w6047_,
		_w6051_,
		_w6025_,
		_w6052_
	);
	LUT4 #(
		.INIT('h0008)
	) name226 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6053_
	);
	LUT4 #(
		.INIT('hfef7)
	) name227 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6054_
	);
	LUT4 #(
		.INIT('h1000)
	) name228 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6055_
	);
	LUT4 #(
		.INIT('hedff)
	) name229 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6056_
	);
	LUT3 #(
		.INIT('hd8)
	) name230 (
		_w6026_,
		_w6054_,
		_w6056_,
		_w6057_
	);
	LUT4 #(
		.INIT('h5655)
	) name231 (
		\u2_L13_reg[14]/NET0131 ,
		_w6052_,
		_w6042_,
		_w6057_,
		_w6058_
	);
	LUT3 #(
		.INIT('ha8)
	) name232 (
		_w5886_,
		_w5888_,
		_w5889_,
		_w6059_
	);
	LUT3 #(
		.INIT('h41)
	) name233 (
		_w5885_,
		_w5887_,
		_w5888_,
		_w6060_
	);
	LUT4 #(
		.INIT('h8200)
	) name234 (
		_w5885_,
		_w5886_,
		_w5887_,
		_w5888_,
		_w6061_
	);
	LUT4 #(
		.INIT('h2400)
	) name235 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6062_
	);
	LUT4 #(
		.INIT('h1011)
	) name236 (
		_w6061_,
		_w6062_,
		_w6059_,
		_w6060_,
		_w6063_
	);
	LUT3 #(
		.INIT('hed)
	) name237 (
		_w5887_,
		_w5888_,
		_w5889_,
		_w6064_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		_w5903_,
		_w6064_,
		_w6065_
	);
	LUT4 #(
		.INIT('h0040)
	) name239 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6066_
	);
	LUT4 #(
		.INIT('hf0b5)
	) name240 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6067_
	);
	LUT4 #(
		.INIT('h5001)
	) name241 (
		_w5885_,
		_w5886_,
		_w5888_,
		_w5889_,
		_w6068_
	);
	LUT4 #(
		.INIT('h0020)
	) name242 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6069_
	);
	LUT4 #(
		.INIT('h77df)
	) name243 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6070_
	);
	LUT4 #(
		.INIT('h0d00)
	) name244 (
		_w5885_,
		_w6067_,
		_w6068_,
		_w6070_,
		_w6071_
	);
	LUT4 #(
		.INIT('h0e04)
	) name245 (
		_w5884_,
		_w6063_,
		_w6065_,
		_w6071_,
		_w6072_
	);
	LUT2 #(
		.INIT('h9)
	) name246 (
		\u2_L13_reg[17]/NET0131 ,
		_w6072_,
		_w6073_
	);
	LUT3 #(
		.INIT('h04)
	) name247 (
		_w5998_,
		_w5984_,
		_w5994_,
		_w6074_
	);
	LUT3 #(
		.INIT('h71)
	) name248 (
		_w5985_,
		_w5983_,
		_w5986_,
		_w6075_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		_w5982_,
		_w5987_,
		_w6076_
	);
	LUT4 #(
		.INIT('h0090)
	) name250 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w6077_
	);
	LUT4 #(
		.INIT('h0015)
	) name251 (
		_w5984_,
		_w6075_,
		_w6076_,
		_w6077_,
		_w6078_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w6074_,
		_w6078_,
		_w6079_
	);
	LUT4 #(
		.INIT('h8000)
	) name253 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w6080_
	);
	LUT3 #(
		.INIT('h01)
	) name254 (
		_w5982_,
		_w5999_,
		_w6080_,
		_w6081_
	);
	LUT4 #(
		.INIT('h0700)
	) name255 (
		_w5985_,
		_w5987_,
		_w5986_,
		_w5984_,
		_w6082_
	);
	LUT3 #(
		.INIT('h53)
	) name256 (
		_w5987_,
		_w5983_,
		_w5986_,
		_w6083_
	);
	LUT4 #(
		.INIT('h135f)
	) name257 (
		_w6005_,
		_w5989_,
		_w6082_,
		_w6083_,
		_w6084_
	);
	LUT3 #(
		.INIT('h0d)
	) name258 (
		_w5985_,
		_w5983_,
		_w5986_,
		_w6085_
	);
	LUT2 #(
		.INIT('h2)
	) name259 (
		_w5988_,
		_w6085_,
		_w6086_
	);
	LUT4 #(
		.INIT('h0080)
	) name260 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w6087_
	);
	LUT3 #(
		.INIT('h10)
	) name261 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w6088_
	);
	LUT3 #(
		.INIT('h02)
	) name262 (
		_w5982_,
		_w6087_,
		_w6088_,
		_w6089_
	);
	LUT4 #(
		.INIT('h7077)
	) name263 (
		_w6081_,
		_w6084_,
		_w6086_,
		_w6089_,
		_w6090_
	);
	LUT3 #(
		.INIT('h56)
	) name264 (
		\u2_L13_reg[1]/NET0131 ,
		_w6079_,
		_w6090_,
		_w6091_
	);
	LUT2 #(
		.INIT('h2)
	) name265 (
		_w5951_,
		_w5952_,
		_w6092_
	);
	LUT4 #(
		.INIT('h9d80)
	) name266 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6093_
	);
	LUT4 #(
		.INIT('h2000)
	) name267 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6094_
	);
	LUT3 #(
		.INIT('h04)
	) name268 (
		_w5951_,
		_w5953_,
		_w5956_,
		_w6095_
	);
	LUT4 #(
		.INIT('hddd8)
	) name269 (
		_w5950_,
		_w6093_,
		_w6094_,
		_w6095_,
		_w6096_
	);
	LUT4 #(
		.INIT('h0082)
	) name270 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6097_
	);
	LUT4 #(
		.INIT('h0100)
	) name271 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6098_
	);
	LUT3 #(
		.INIT('h02)
	) name272 (
		_w5962_,
		_w6097_,
		_w6098_,
		_w6099_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w6096_,
		_w6099_,
		_w6100_
	);
	LUT4 #(
		.INIT('h0004)
	) name274 (
		_w5950_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6101_
	);
	LUT3 #(
		.INIT('h01)
	) name275 (
		_w5962_,
		_w5964_,
		_w6101_,
		_w6102_
	);
	LUT3 #(
		.INIT('h23)
	) name276 (
		_w5950_,
		_w5952_,
		_w5956_,
		_w6103_
	);
	LUT3 #(
		.INIT('h51)
	) name277 (
		_w5971_,
		_w5973_,
		_w6103_,
		_w6104_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name278 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6105_
	);
	LUT4 #(
		.INIT('hceff)
	) name279 (
		_w5950_,
		_w5951_,
		_w5952_,
		_w5953_,
		_w6106_
	);
	LUT4 #(
		.INIT('hf531)
	) name280 (
		_w5950_,
		_w5956_,
		_w6105_,
		_w6106_,
		_w6107_
	);
	LUT3 #(
		.INIT('h80)
	) name281 (
		_w6102_,
		_w6104_,
		_w6107_,
		_w6108_
	);
	LUT4 #(
		.INIT('h0002)
	) name282 (
		_w5950_,
		_w5951_,
		_w5952_,
		_w5953_,
		_w6109_
	);
	LUT3 #(
		.INIT('h07)
	) name283 (
		_w5959_,
		_w5977_,
		_w6109_,
		_w6110_
	);
	LUT4 #(
		.INIT('ha955)
	) name284 (
		\u2_L13_reg[21]/NET0131 ,
		_w6100_,
		_w6108_,
		_w6110_,
		_w6111_
	);
	LUT4 #(
		.INIT('h085d)
	) name285 (
		_w5987_,
		_w5983_,
		_w5986_,
		_w5984_,
		_w6112_
	);
	LUT3 #(
		.INIT('h45)
	) name286 (
		_w5985_,
		_w5983_,
		_w5986_,
		_w6113_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		_w6112_,
		_w6113_,
		_w6114_
	);
	LUT4 #(
		.INIT('h54ff)
	) name288 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w6115_
	);
	LUT3 #(
		.INIT('h0d)
	) name289 (
		_w5985_,
		_w5983_,
		_w5984_,
		_w6116_
	);
	LUT4 #(
		.INIT('h2022)
	) name290 (
		_w5982_,
		_w6087_,
		_w6115_,
		_w6116_,
		_w6117_
	);
	LUT2 #(
		.INIT('h2)
	) name291 (
		_w6006_,
		_w6075_,
		_w6118_
	);
	LUT3 #(
		.INIT('h02)
	) name292 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w6119_
	);
	LUT3 #(
		.INIT('h01)
	) name293 (
		_w5982_,
		_w5999_,
		_w6119_,
		_w6120_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name294 (
		_w6114_,
		_w6117_,
		_w6118_,
		_w6120_,
		_w6121_
	);
	LUT4 #(
		.INIT('hefcc)
	) name295 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w6122_
	);
	LUT3 #(
		.INIT('h08)
	) name296 (
		_w5985_,
		_w5987_,
		_w5986_,
		_w6123_
	);
	LUT4 #(
		.INIT('h0806)
	) name297 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w6124_
	);
	LUT4 #(
		.INIT('h0302)
	) name298 (
		_w5982_,
		_w5984_,
		_w6124_,
		_w6122_,
		_w6125_
	);
	LUT4 #(
		.INIT('h0200)
	) name299 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w6126_
	);
	LUT3 #(
		.INIT('h02)
	) name300 (
		_w5984_,
		_w5999_,
		_w6126_,
		_w6127_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w6125_,
		_w6127_,
		_w6128_
	);
	LUT3 #(
		.INIT('h56)
	) name302 (
		\u2_L13_reg[26]/NET0131 ,
		_w6121_,
		_w6128_,
		_w6129_
	);
	LUT4 #(
		.INIT('h6c6a)
	) name303 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6130_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name304 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6131_
	);
	LUT4 #(
		.INIT('hf75f)
	) name305 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6132_
	);
	LUT4 #(
		.INIT('hd800)
	) name306 (
		_w6026_,
		_w6130_,
		_w6131_,
		_w6132_,
		_w6133_
	);
	LUT2 #(
		.INIT('h2)
	) name307 (
		_w6025_,
		_w6133_,
		_w6134_
	);
	LUT4 #(
		.INIT('h51f3)
	) name308 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6135_
	);
	LUT3 #(
		.INIT('h07)
	) name309 (
		_w6028_,
		_w6029_,
		_w6026_,
		_w6136_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w6135_,
		_w6136_,
		_w6137_
	);
	LUT4 #(
		.INIT('h0200)
	) name311 (
		_w6028_,
		_w6030_,
		_w6027_,
		_w6026_,
		_w6138_
	);
	LUT4 #(
		.INIT('h0001)
	) name312 (
		_w6028_,
		_w6029_,
		_w6027_,
		_w6026_,
		_w6139_
	);
	LUT4 #(
		.INIT('h2000)
	) name313 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6140_
	);
	LUT3 #(
		.INIT('h01)
	) name314 (
		_w6139_,
		_w6140_,
		_w6138_,
		_w6141_
	);
	LUT4 #(
		.INIT('hf6ef)
	) name315 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6142_
	);
	LUT4 #(
		.INIT('h0040)
	) name316 (
		_w6028_,
		_w6029_,
		_w6027_,
		_w6026_,
		_w6143_
	);
	LUT4 #(
		.INIT('h0031)
	) name317 (
		_w6026_,
		_w6032_,
		_w6142_,
		_w6143_,
		_w6144_
	);
	LUT4 #(
		.INIT('hba00)
	) name318 (
		_w6025_,
		_w6137_,
		_w6141_,
		_w6144_,
		_w6145_
	);
	LUT3 #(
		.INIT('h65)
	) name319 (
		\u2_L13_reg[25]/NET0131 ,
		_w6134_,
		_w6145_,
		_w6146_
	);
	LUT4 #(
		.INIT('h3fd2)
	) name320 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6147_
	);
	LUT4 #(
		.INIT('hab6f)
	) name321 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6148_
	);
	LUT4 #(
		.INIT('h0200)
	) name322 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6149_
	);
	LUT4 #(
		.INIT('h00e4)
	) name323 (
		_w5917_,
		_w6148_,
		_w6147_,
		_w6149_,
		_w6150_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w5925_,
		_w6150_,
		_w6151_
	);
	LUT4 #(
		.INIT('hcf6f)
	) name325 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6152_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		_w5917_,
		_w6152_,
		_w6153_
	);
	LUT4 #(
		.INIT('h0102)
	) name327 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6154_
	);
	LUT4 #(
		.INIT('h77dc)
	) name328 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6155_
	);
	LUT4 #(
		.INIT('h0302)
	) name329 (
		_w5917_,
		_w5938_,
		_w5932_,
		_w6155_,
		_w6156_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name330 (
		_w5925_,
		_w6153_,
		_w6154_,
		_w6156_,
		_w6157_
	);
	LUT4 #(
		.INIT('h2000)
	) name331 (
		_w5917_,
		_w5918_,
		_w5921_,
		_w5920_,
		_w6158_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w5927_,
		_w6158_,
		_w6159_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name333 (
		\u2_L13_reg[29]/NET0131 ,
		_w6157_,
		_w6151_,
		_w6159_,
		_w6160_
	);
	LUT4 #(
		.INIT('hc693)
	) name334 (
		decrypt_pad,
		\u2_R13_reg[5]/NET0131 ,
		\u2_uk_K_r13_reg[13]/NET0131 ,
		\u2_uk_K_r13_reg[17]/NET0131 ,
		_w6161_
	);
	LUT4 #(
		.INIT('hc963)
	) name335 (
		decrypt_pad,
		\u2_R13_reg[4]/NET0131 ,
		\u2_uk_K_r13_reg[13]/NET0131 ,
		\u2_uk_K_r13_reg[34]/NET0131 ,
		_w6162_
	);
	LUT4 #(
		.INIT('hc693)
	) name336 (
		decrypt_pad,
		\u2_R13_reg[9]/NET0131 ,
		\u2_uk_K_r13_reg[26]/NET0131 ,
		\u2_uk_K_r13_reg[5]/NET0131 ,
		_w6163_
	);
	LUT4 #(
		.INIT('hc963)
	) name337 (
		decrypt_pad,
		\u2_R13_reg[6]/NET0131 ,
		\u2_uk_K_r13_reg[40]/NET0131 ,
		\u2_uk_K_r13_reg[4]/NET0131 ,
		_w6164_
	);
	LUT4 #(
		.INIT('hc038)
	) name338 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6165_
	);
	LUT4 #(
		.INIT('hc963)
	) name339 (
		decrypt_pad,
		\u2_R13_reg[7]/NET0131 ,
		\u2_uk_K_r13_reg[34]/NET0131 ,
		\u2_uk_K_r13_reg[55]/NET0131 ,
		_w6166_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		_w6165_,
		_w6166_,
		_w6167_
	);
	LUT4 #(
		.INIT('h0c05)
	) name341 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6168_
	);
	LUT4 #(
		.INIT('h0080)
	) name342 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6169_
	);
	LUT4 #(
		.INIT('h00fd)
	) name343 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6166_,
		_w6170_
	);
	LUT3 #(
		.INIT('h10)
	) name344 (
		_w6168_,
		_w6169_,
		_w6170_,
		_w6171_
	);
	LUT3 #(
		.INIT('h40)
	) name345 (
		_w6161_,
		_w6162_,
		_w6163_,
		_w6172_
	);
	LUT4 #(
		.INIT('h00bf)
	) name346 (
		_w6161_,
		_w6162_,
		_w6163_,
		_w6166_,
		_w6173_
	);
	LUT2 #(
		.INIT('h4)
	) name347 (
		_w6164_,
		_w6162_,
		_w6174_
	);
	LUT4 #(
		.INIT('h0200)
	) name348 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6175_
	);
	LUT4 #(
		.INIT('hc963)
	) name349 (
		decrypt_pad,
		\u2_R13_reg[8]/NET0131 ,
		\u2_uk_K_r13_reg[25]/P0001 ,
		\u2_uk_K_r13_reg[46]/NET0131 ,
		_w6176_
	);
	LUT4 #(
		.INIT('h4500)
	) name350 (
		_w6175_,
		_w6173_,
		_w6174_,
		_w6176_,
		_w6177_
	);
	LUT3 #(
		.INIT('he0)
	) name351 (
		_w6167_,
		_w6171_,
		_w6177_,
		_w6178_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		_w6166_,
		_w6168_,
		_w6179_
	);
	LUT4 #(
		.INIT('h3c2f)
	) name353 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6180_
	);
	LUT3 #(
		.INIT('h40)
	) name354 (
		_w6169_,
		_w6170_,
		_w6180_,
		_w6181_
	);
	LUT4 #(
		.INIT('h2002)
	) name355 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6182_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w6169_,
		_w6176_,
		_w6183_
	);
	LUT3 #(
		.INIT('h01)
	) name357 (
		_w6169_,
		_w6176_,
		_w6182_,
		_w6184_
	);
	LUT3 #(
		.INIT('he0)
	) name358 (
		_w6179_,
		_w6181_,
		_w6184_,
		_w6185_
	);
	LUT3 #(
		.INIT('ha9)
	) name359 (
		\u2_L13_reg[28]/NET0131 ,
		_w6178_,
		_w6185_,
		_w6186_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name360 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6187_
	);
	LUT4 #(
		.INIT('h7f7c)
	) name361 (
		_w6164_,
		_w6166_,
		_w6172_,
		_w6187_,
		_w6188_
	);
	LUT4 #(
		.INIT('h0144)
	) name362 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6189_
	);
	LUT4 #(
		.INIT('h0800)
	) name363 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6190_
	);
	LUT4 #(
		.INIT('h0010)
	) name364 (
		_w6164_,
		_w6161_,
		_w6163_,
		_w6166_,
		_w6191_
	);
	LUT3 #(
		.INIT('h01)
	) name365 (
		_w6189_,
		_w6190_,
		_w6191_,
		_w6192_
	);
	LUT3 #(
		.INIT('h15)
	) name366 (
		_w6176_,
		_w6188_,
		_w6192_,
		_w6193_
	);
	LUT3 #(
		.INIT('h01)
	) name367 (
		_w6164_,
		_w6161_,
		_w6163_,
		_w6194_
	);
	LUT4 #(
		.INIT('h0010)
	) name368 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6195_
	);
	LUT4 #(
		.INIT('h9fe4)
	) name369 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6196_
	);
	LUT4 #(
		.INIT('h0900)
	) name370 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6197_
	);
	LUT4 #(
		.INIT('h0501)
	) name371 (
		_w6166_,
		_w6176_,
		_w6197_,
		_w6196_,
		_w6198_
	);
	LUT3 #(
		.INIT('h2a)
	) name372 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6199_
	);
	LUT4 #(
		.INIT('hae00)
	) name373 (
		_w6161_,
		_w6162_,
		_w6163_,
		_w6176_,
		_w6200_
	);
	LUT4 #(
		.INIT('h0002)
	) name374 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6201_
	);
	LUT4 #(
		.INIT('hbf00)
	) name375 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6166_,
		_w6202_
	);
	LUT4 #(
		.INIT('h4500)
	) name376 (
		_w6201_,
		_w6199_,
		_w6200_,
		_w6202_,
		_w6203_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w6198_,
		_w6203_,
		_w6204_
	);
	LUT3 #(
		.INIT('h56)
	) name378 (
		\u2_L13_reg[2]/NET0131 ,
		_w6193_,
		_w6204_,
		_w6205_
	);
	LUT4 #(
		.INIT('he63f)
	) name379 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6206_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		_w5917_,
		_w6206_,
		_w6207_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name381 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6208_
	);
	LUT4 #(
		.INIT('h1000)
	) name382 (
		_w5917_,
		_w5918_,
		_w5919_,
		_w5920_,
		_w6209_
	);
	LUT4 #(
		.INIT('h0032)
	) name383 (
		_w5917_,
		_w5927_,
		_w6208_,
		_w6209_,
		_w6210_
	);
	LUT3 #(
		.INIT('h45)
	) name384 (
		_w5925_,
		_w6207_,
		_w6210_,
		_w6211_
	);
	LUT4 #(
		.INIT('heeae)
	) name385 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6212_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		_w5917_,
		_w6212_,
		_w6213_
	);
	LUT3 #(
		.INIT('h80)
	) name387 (
		_w5918_,
		_w5921_,
		_w5920_,
		_w6214_
	);
	LUT4 #(
		.INIT('h2000)
	) name388 (
		_w5917_,
		_w5918_,
		_w5919_,
		_w5920_,
		_w6215_
	);
	LUT3 #(
		.INIT('h01)
	) name389 (
		_w5944_,
		_w6214_,
		_w6215_,
		_w6216_
	);
	LUT3 #(
		.INIT('hb6)
	) name390 (
		_w5919_,
		_w5921_,
		_w5920_,
		_w6217_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name391 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6218_
	);
	LUT4 #(
		.INIT('h4445)
	) name392 (
		_w5917_,
		_w5918_,
		_w5919_,
		_w5920_,
		_w6219_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name393 (
		_w5936_,
		_w6217_,
		_w6218_,
		_w6219_,
		_w6220_
	);
	LUT4 #(
		.INIT('h7500)
	) name394 (
		_w5925_,
		_w6213_,
		_w6216_,
		_w6220_,
		_w6221_
	);
	LUT3 #(
		.INIT('h65)
	) name395 (
		\u2_L13_reg[4]/NET0131 ,
		_w6211_,
		_w6221_,
		_w6222_
	);
	LUT3 #(
		.INIT('h02)
	) name396 (
		_w6164_,
		_w6161_,
		_w6163_,
		_w6223_
	);
	LUT4 #(
		.INIT('hdf00)
	) name397 (
		_w6164_,
		_w6162_,
		_w6163_,
		_w6166_,
		_w6224_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name398 (
		_w6173_,
		_w6194_,
		_w6223_,
		_w6224_,
		_w6225_
	);
	LUT4 #(
		.INIT('h0004)
	) name399 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6226_
	);
	LUT4 #(
		.INIT('h0002)
	) name400 (
		_w6176_,
		_w6190_,
		_w6191_,
		_w6226_,
		_w6227_
	);
	LUT4 #(
		.INIT('h0600)
	) name401 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6228_
	);
	LUT3 #(
		.INIT('h02)
	) name402 (
		_w6161_,
		_w6162_,
		_w6163_,
		_w6229_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w6166_,
		_w6176_,
		_w6230_
	);
	LUT4 #(
		.INIT('h0100)
	) name404 (
		_w6195_,
		_w6229_,
		_w6228_,
		_w6230_,
		_w6231_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name405 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6232_
	);
	LUT4 #(
		.INIT('hf400)
	) name406 (
		_w6225_,
		_w6227_,
		_w6231_,
		_w6232_,
		_w6233_
	);
	LUT4 #(
		.INIT('h1141)
	) name407 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6234_
	);
	LUT4 #(
		.INIT('ha022)
	) name408 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6235_
	);
	LUT4 #(
		.INIT('h0400)
	) name409 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6236_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		_w6166_,
		_w6176_,
		_w6237_
	);
	LUT4 #(
		.INIT('h0100)
	) name411 (
		_w6235_,
		_w6236_,
		_w6234_,
		_w6237_,
		_w6238_
	);
	LUT3 #(
		.INIT('h56)
	) name412 (
		\u2_L13_reg[13]/NET0131 ,
		_w6233_,
		_w6238_,
		_w6239_
	);
	LUT4 #(
		.INIT('h7343)
	) name413 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6240_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		_w5917_,
		_w6240_,
		_w6241_
	);
	LUT4 #(
		.INIT('h1001)
	) name415 (
		_w5917_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6242_
	);
	LUT4 #(
		.INIT('h8000)
	) name416 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6243_
	);
	LUT3 #(
		.INIT('h01)
	) name417 (
		_w5925_,
		_w6243_,
		_w6242_,
		_w6244_
	);
	LUT4 #(
		.INIT('h2000)
	) name418 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6245_
	);
	LUT3 #(
		.INIT('h04)
	) name419 (
		_w5917_,
		_w5919_,
		_w5921_,
		_w6246_
	);
	LUT4 #(
		.INIT('haa8a)
	) name420 (
		_w5925_,
		_w5918_,
		_w5921_,
		_w5920_,
		_w6247_
	);
	LUT3 #(
		.INIT('h10)
	) name421 (
		_w6245_,
		_w6246_,
		_w6247_,
		_w6248_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name422 (
		_w5918_,
		_w5919_,
		_w5921_,
		_w5920_,
		_w6249_
	);
	LUT3 #(
		.INIT('h31)
	) name423 (
		_w5917_,
		_w6154_,
		_w6249_,
		_w6250_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name424 (
		_w6241_,
		_w6244_,
		_w6248_,
		_w6250_,
		_w6251_
	);
	LUT4 #(
		.INIT('hefcc)
	) name425 (
		_w5917_,
		_w5918_,
		_w5922_,
		_w5942_,
		_w6252_
	);
	LUT3 #(
		.INIT('h65)
	) name426 (
		\u2_L13_reg[19]/P0001 ,
		_w6251_,
		_w6252_,
		_w6253_
	);
	LUT4 #(
		.INIT('h5040)
	) name427 (
		_w5885_,
		_w5886_,
		_w5888_,
		_w5889_,
		_w6254_
	);
	LUT4 #(
		.INIT('hfcf4)
	) name428 (
		_w5885_,
		_w5886_,
		_w5887_,
		_w5888_,
		_w6255_
	);
	LUT3 #(
		.INIT('h45)
	) name429 (
		_w5900_,
		_w6254_,
		_w6255_,
		_w6256_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		_w5885_,
		_w5886_,
		_w6257_
	);
	LUT4 #(
		.INIT('h8c00)
	) name431 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6258_
	);
	LUT2 #(
		.INIT('h4)
	) name432 (
		_w6257_,
		_w6258_,
		_w6259_
	);
	LUT3 #(
		.INIT('h54)
	) name433 (
		_w5884_,
		_w6256_,
		_w6259_,
		_w6260_
	);
	LUT4 #(
		.INIT('h8808)
	) name434 (
		_w5885_,
		_w5886_,
		_w5888_,
		_w5889_,
		_w6261_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		_w5904_,
		_w6261_,
		_w6262_
	);
	LUT3 #(
		.INIT('h07)
	) name436 (
		_w5895_,
		_w5912_,
		_w6066_,
		_w6263_
	);
	LUT3 #(
		.INIT('h8a)
	) name437 (
		_w5884_,
		_w6262_,
		_w6263_,
		_w6264_
	);
	LUT4 #(
		.INIT('he9f9)
	) name438 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6265_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		_w5884_,
		_w5885_,
		_w6266_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w6265_,
		_w6266_,
		_w6267_
	);
	LUT4 #(
		.INIT('h7fdb)
	) name441 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6268_
	);
	LUT3 #(
		.INIT('had)
	) name442 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w6269_
	);
	LUT4 #(
		.INIT('hfad8)
	) name443 (
		_w5885_,
		_w5889_,
		_w6268_,
		_w6269_,
		_w6270_
	);
	LUT2 #(
		.INIT('h4)
	) name444 (
		_w6267_,
		_w6270_,
		_w6271_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name445 (
		\u2_L13_reg[23]/P0001 ,
		_w6260_,
		_w6264_,
		_w6271_,
		_w6272_
	);
	LUT4 #(
		.INIT('h0004)
	) name446 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6273_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name447 (
		_w5950_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6274_
	);
	LUT3 #(
		.INIT('hd7)
	) name448 (
		_w5952_,
		_w5953_,
		_w5956_,
		_w6275_
	);
	LUT4 #(
		.INIT('h45cf)
	) name449 (
		_w5955_,
		_w6273_,
		_w6274_,
		_w6275_,
		_w6276_
	);
	LUT4 #(
		.INIT('he6df)
	) name450 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6277_
	);
	LUT3 #(
		.INIT('h8a)
	) name451 (
		_w5962_,
		_w6276_,
		_w6277_,
		_w6278_
	);
	LUT4 #(
		.INIT('h004c)
	) name452 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6279_
	);
	LUT4 #(
		.INIT('h20aa)
	) name453 (
		_w5950_,
		_w5951_,
		_w5952_,
		_w5956_,
		_w6280_
	);
	LUT4 #(
		.INIT('hcd00)
	) name454 (
		_w5962_,
		_w6092_,
		_w6279_,
		_w6280_,
		_w6281_
	);
	LUT4 #(
		.INIT('hefb7)
	) name455 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w6282_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		_w5950_,
		_w6282_,
		_w6283_
	);
	LUT4 #(
		.INIT('h4000)
	) name457 (
		_w5950_,
		_w5951_,
		_w5953_,
		_w5956_,
		_w6284_
	);
	LUT4 #(
		.INIT('h5554)
	) name458 (
		_w5962_,
		_w5965_,
		_w6101_,
		_w6284_,
		_w6285_
	);
	LUT3 #(
		.INIT('h01)
	) name459 (
		_w6283_,
		_w6285_,
		_w6281_,
		_w6286_
	);
	LUT3 #(
		.INIT('h65)
	) name460 (
		\u2_L13_reg[27]/NET0131 ,
		_w6278_,
		_w6286_,
		_w6287_
	);
	LUT4 #(
		.INIT('h0080)
	) name461 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6288_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w5856_,
		_w6020_,
		_w6289_
	);
	LUT3 #(
		.INIT('h48)
	) name463 (
		_w5857_,
		_w5859_,
		_w5860_,
		_w6290_
	);
	LUT4 #(
		.INIT('h0134)
	) name464 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6291_
	);
	LUT3 #(
		.INIT('h01)
	) name465 (
		_w5856_,
		_w6020_,
		_w6291_,
		_w6292_
	);
	LUT3 #(
		.INIT('hc4)
	) name466 (
		_w5858_,
		_w5857_,
		_w5860_,
		_w6293_
	);
	LUT4 #(
		.INIT('h008b)
	) name467 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6294_
	);
	LUT4 #(
		.INIT('hbf00)
	) name468 (
		_w5858_,
		_w5859_,
		_w5860_,
		_w5856_,
		_w6295_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		_w6294_,
		_w6295_,
		_w6296_
	);
	LUT4 #(
		.INIT('h888a)
	) name470 (
		_w5868_,
		_w6288_,
		_w6292_,
		_w6296_,
		_w6297_
	);
	LUT3 #(
		.INIT('h04)
	) name471 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w6298_
	);
	LUT3 #(
		.INIT('h09)
	) name472 (
		_w5859_,
		_w5860_,
		_w5856_,
		_w6299_
	);
	LUT2 #(
		.INIT('h4)
	) name473 (
		_w6298_,
		_w6299_,
		_w6300_
	);
	LUT4 #(
		.INIT('hbf8c)
	) name474 (
		_w5858_,
		_w5859_,
		_w5860_,
		_w5856_,
		_w6301_
	);
	LUT3 #(
		.INIT('h15)
	) name475 (
		_w5879_,
		_w6293_,
		_w6301_,
		_w6302_
	);
	LUT4 #(
		.INIT('h9fdf)
	) name476 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6303_
	);
	LUT4 #(
		.INIT('h7544)
	) name477 (
		_w5866_,
		_w5856_,
		_w5868_,
		_w6303_,
		_w6304_
	);
	LUT4 #(
		.INIT('hba00)
	) name478 (
		_w5868_,
		_w6300_,
		_w6302_,
		_w6304_,
		_w6305_
	);
	LUT3 #(
		.INIT('h65)
	) name479 (
		\u2_L13_reg[32]/NET0131 ,
		_w6297_,
		_w6305_,
		_w6306_
	);
	LUT4 #(
		.INIT('hc693)
	) name480 (
		decrypt_pad,
		\u2_R13_reg[12]/NET0131 ,
		\u2_uk_K_r13_reg[24]/NET0131 ,
		\u2_uk_K_r13_reg[3]/NET0131 ,
		_w6307_
	);
	LUT4 #(
		.INIT('hc963)
	) name481 (
		decrypt_pad,
		\u2_R13_reg[11]/NET0131 ,
		\u2_uk_K_r13_reg[20]/NET0131 ,
		\u2_uk_K_r13_reg[41]/NET0131 ,
		_w6308_
	);
	LUT4 #(
		.INIT('hc963)
	) name482 (
		decrypt_pad,
		\u2_R13_reg[9]/NET0131 ,
		\u2_uk_K_r13_reg[11]/NET0131 ,
		\u2_uk_K_r13_reg[32]/NET0131 ,
		_w6309_
	);
	LUT4 #(
		.INIT('hc963)
	) name483 (
		decrypt_pad,
		\u2_R13_reg[10]/NET0131 ,
		\u2_uk_K_r13_reg[19]/NET0131 ,
		\u2_uk_K_r13_reg[40]/NET0131 ,
		_w6310_
	);
	LUT4 #(
		.INIT('hc963)
	) name484 (
		decrypt_pad,
		\u2_R13_reg[8]/NET0131 ,
		\u2_uk_K_r13_reg[39]/NET0131 ,
		\u2_uk_K_r13_reg[3]/NET0131 ,
		_w6311_
	);
	LUT4 #(
		.INIT('hc693)
	) name485 (
		decrypt_pad,
		\u2_R13_reg[13]/NET0131 ,
		\u2_uk_K_r13_reg[12]/NET0131 ,
		\u2_uk_K_r13_reg[48]/NET0131 ,
		_w6312_
	);
	LUT4 #(
		.INIT('h4000)
	) name486 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6313_
	);
	LUT2 #(
		.INIT('h4)
	) name487 (
		_w6308_,
		_w6313_,
		_w6314_
	);
	LUT2 #(
		.INIT('h6)
	) name488 (
		_w6311_,
		_w6312_,
		_w6315_
	);
	LUT4 #(
		.INIT('h9990)
	) name489 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6316_
	);
	LUT4 #(
		.INIT('h0990)
	) name490 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6317_
	);
	LUT2 #(
		.INIT('h4)
	) name491 (
		_w6311_,
		_w6308_,
		_w6318_
	);
	LUT4 #(
		.INIT('h000b)
	) name492 (
		_w6311_,
		_w6308_,
		_w6309_,
		_w6310_,
		_w6319_
	);
	LUT2 #(
		.INIT('h2)
	) name493 (
		_w6308_,
		_w6310_,
		_w6320_
	);
	LUT4 #(
		.INIT('h0040)
	) name494 (
		_w6311_,
		_w6308_,
		_w6309_,
		_w6310_,
		_w6321_
	);
	LUT4 #(
		.INIT('h2000)
	) name495 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6322_
	);
	LUT4 #(
		.INIT('h0007)
	) name496 (
		_w6315_,
		_w6319_,
		_w6321_,
		_w6322_,
		_w6323_
	);
	LUT4 #(
		.INIT('h5455)
	) name497 (
		_w6307_,
		_w6317_,
		_w6314_,
		_w6323_,
		_w6324_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w6307_,
		_w6310_,
		_w6325_
	);
	LUT3 #(
		.INIT('h10)
	) name499 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6326_
	);
	LUT4 #(
		.INIT('h93d3)
	) name500 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6327_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		_w6307_,
		_w6308_,
		_w6328_
	);
	LUT4 #(
		.INIT('h7077)
	) name502 (
		_w6325_,
		_w6326_,
		_w6327_,
		_w6328_,
		_w6329_
	);
	LUT4 #(
		.INIT('h0001)
	) name503 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6330_
	);
	LUT4 #(
		.INIT('hf3fe)
	) name504 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6331_
	);
	LUT2 #(
		.INIT('h2)
	) name505 (
		_w6307_,
		_w6308_,
		_w6332_
	);
	LUT3 #(
		.INIT('h80)
	) name506 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6333_
	);
	LUT3 #(
		.INIT('h08)
	) name507 (
		_w6312_,
		_w6309_,
		_w6310_,
		_w6334_
	);
	LUT2 #(
		.INIT('h2)
	) name508 (
		_w6311_,
		_w6309_,
		_w6335_
	);
	LUT3 #(
		.INIT('h02)
	) name509 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6336_
	);
	LUT4 #(
		.INIT('h7d3d)
	) name510 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6337_
	);
	LUT4 #(
		.INIT('hf3d1)
	) name511 (
		_w6307_,
		_w6308_,
		_w6331_,
		_w6337_,
		_w6338_
	);
	LUT2 #(
		.INIT('h8)
	) name512 (
		_w6329_,
		_w6338_,
		_w6339_
	);
	LUT3 #(
		.INIT('h65)
	) name513 (
		\u2_L13_reg[6]/NET0131 ,
		_w6324_,
		_w6339_,
		_w6340_
	);
	LUT2 #(
		.INIT('h2)
	) name514 (
		_w5856_,
		_w5868_,
		_w6341_
	);
	LUT4 #(
		.INIT('h2080)
	) name515 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6342_
	);
	LUT4 #(
		.INIT('h936e)
	) name516 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6343_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		_w6341_,
		_w6343_,
		_w6344_
	);
	LUT4 #(
		.INIT('h4410)
	) name518 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6345_
	);
	LUT2 #(
		.INIT('h9)
	) name519 (
		_w5856_,
		_w5868_,
		_w6346_
	);
	LUT4 #(
		.INIT('h0100)
	) name520 (
		_w6020_,
		_w6342_,
		_w6345_,
		_w6346_,
		_w6347_
	);
	LUT3 #(
		.INIT('h54)
	) name521 (
		_w6021_,
		_w6344_,
		_w6347_,
		_w6348_
	);
	LUT4 #(
		.INIT('h20a8)
	) name522 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5860_,
		_w6349_
	);
	LUT4 #(
		.INIT('hfe00)
	) name523 (
		_w5858_,
		_w5857_,
		_w5859_,
		_w5868_,
		_w6350_
	);
	LUT3 #(
		.INIT('h10)
	) name524 (
		_w6290_,
		_w6349_,
		_w6350_,
		_w6351_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w6289_,
		_w6351_,
		_w6352_
	);
	LUT3 #(
		.INIT('ha9)
	) name526 (
		\u2_L13_reg[7]/NET0131 ,
		_w6348_,
		_w6352_,
		_w6353_
	);
	LUT4 #(
		.INIT('h9f8f)
	) name527 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6354_
	);
	LUT4 #(
		.INIT('h7f7b)
	) name528 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6355_
	);
	LUT4 #(
		.INIT('hf6dd)
	) name529 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6356_
	);
	LUT4 #(
		.INIT('hd800)
	) name530 (
		_w6026_,
		_w6355_,
		_w6354_,
		_w6356_,
		_w6357_
	);
	LUT4 #(
		.INIT('h0001)
	) name531 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6358_
	);
	LUT4 #(
		.INIT('hbfbe)
	) name532 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6359_
	);
	LUT3 #(
		.INIT('h02)
	) name533 (
		_w6029_,
		_w6027_,
		_w6026_,
		_w6360_
	);
	LUT4 #(
		.INIT('h00c4)
	) name534 (
		_w6026_,
		_w6056_,
		_w6359_,
		_w6360_,
		_w6361_
	);
	LUT4 #(
		.INIT('he5df)
	) name535 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6362_
	);
	LUT4 #(
		.INIT('haf23)
	) name536 (
		_w6030_,
		_w6026_,
		_w6143_,
		_w6362_,
		_w6363_
	);
	LUT4 #(
		.INIT('hd800)
	) name537 (
		_w6025_,
		_w6361_,
		_w6357_,
		_w6363_,
		_w6364_
	);
	LUT2 #(
		.INIT('h9)
	) name538 (
		\u2_L13_reg[8]/NET0131 ,
		_w6364_,
		_w6365_
	);
	LUT3 #(
		.INIT('h84)
	) name539 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6366_
	);
	LUT4 #(
		.INIT('h5ba5)
	) name540 (
		_w6311_,
		_w6308_,
		_w6312_,
		_w6309_,
		_w6367_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w6310_,
		_w6367_,
		_w6368_
	);
	LUT4 #(
		.INIT('h0102)
	) name542 (
		_w6311_,
		_w6308_,
		_w6312_,
		_w6310_,
		_w6369_
	);
	LUT3 #(
		.INIT('h02)
	) name543 (
		_w6307_,
		_w6313_,
		_w6369_,
		_w6370_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name544 (
		_w6311_,
		_w6308_,
		_w6312_,
		_w6309_,
		_w6371_
	);
	LUT3 #(
		.INIT('h70)
	) name545 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6372_
	);
	LUT4 #(
		.INIT('h844c)
	) name546 (
		_w6311_,
		_w6308_,
		_w6312_,
		_w6309_,
		_w6373_
	);
	LUT4 #(
		.INIT('h3332)
	) name547 (
		_w6311_,
		_w6308_,
		_w6312_,
		_w6310_,
		_w6374_
	);
	LUT3 #(
		.INIT('h23)
	) name548 (
		_w6366_,
		_w6373_,
		_w6374_,
		_w6375_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		_w6307_,
		_w6330_,
		_w6376_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name550 (
		_w6368_,
		_w6370_,
		_w6375_,
		_w6376_,
		_w6377_
	);
	LUT4 #(
		.INIT('hdeff)
	) name551 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6378_
	);
	LUT4 #(
		.INIT('h0200)
	) name552 (
		_w6311_,
		_w6308_,
		_w6309_,
		_w6310_,
		_w6379_
	);
	LUT3 #(
		.INIT('h0d)
	) name553 (
		_w6308_,
		_w6378_,
		_w6379_,
		_w6380_
	);
	LUT3 #(
		.INIT('h65)
	) name554 (
		\u2_L13_reg[16]/NET0131 ,
		_w6377_,
		_w6380_,
		_w6381_
	);
	LUT4 #(
		.INIT('h0009)
	) name555 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6382_
	);
	LUT4 #(
		.INIT('h9bd6)
	) name556 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6383_
	);
	LUT3 #(
		.INIT('h54)
	) name557 (
		_w6307_,
		_w6308_,
		_w6383_,
		_w6384_
	);
	LUT2 #(
		.INIT('h4)
	) name558 (
		_w6308_,
		_w6316_,
		_w6385_
	);
	LUT3 #(
		.INIT('h2a)
	) name559 (
		_w6307_,
		_w6315_,
		_w6319_,
		_w6386_
	);
	LUT3 #(
		.INIT('h0b)
	) name560 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6387_
	);
	LUT4 #(
		.INIT('hc800)
	) name561 (
		_w6311_,
		_w6308_,
		_w6312_,
		_w6310_,
		_w6388_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name562 (
		_w6320_,
		_w6335_,
		_w6387_,
		_w6388_,
		_w6389_
	);
	LUT4 #(
		.INIT('h4555)
	) name563 (
		_w6384_,
		_w6385_,
		_w6386_,
		_w6389_,
		_w6390_
	);
	LUT4 #(
		.INIT('he4ab)
	) name564 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6391_
	);
	LUT4 #(
		.INIT('h0200)
	) name565 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6392_
	);
	LUT4 #(
		.INIT('h5504)
	) name566 (
		_w6307_,
		_w6308_,
		_w6391_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w6318_,
		_w6334_,
		_w6394_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name568 (
		_w6308_,
		_w6310_,
		_w6336_,
		_w6333_,
		_w6395_
	);
	LUT3 #(
		.INIT('h10)
	) name569 (
		_w6393_,
		_w6394_,
		_w6395_,
		_w6396_
	);
	LUT3 #(
		.INIT('h65)
	) name570 (
		\u2_L13_reg[24]/NET0131 ,
		_w6390_,
		_w6396_,
		_w6397_
	);
	LUT4 #(
		.INIT('h75cf)
	) name571 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6398_
	);
	LUT2 #(
		.INIT('h2)
	) name572 (
		_w6308_,
		_w6398_,
		_w6399_
	);
	LUT4 #(
		.INIT('h0400)
	) name573 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6400_
	);
	LUT3 #(
		.INIT('hb1)
	) name574 (
		_w6311_,
		_w6309_,
		_w6310_,
		_w6401_
	);
	LUT3 #(
		.INIT('h45)
	) name575 (
		_w6308_,
		_w6312_,
		_w6309_,
		_w6402_
	);
	LUT4 #(
		.INIT('h0045)
	) name576 (
		_w6382_,
		_w6401_,
		_w6402_,
		_w6400_,
		_w6403_
	);
	LUT3 #(
		.INIT('h45)
	) name577 (
		_w6307_,
		_w6399_,
		_w6403_,
		_w6404_
	);
	LUT4 #(
		.INIT('h0440)
	) name578 (
		_w6311_,
		_w6308_,
		_w6312_,
		_w6310_,
		_w6405_
	);
	LUT4 #(
		.INIT('haa80)
	) name579 (
		_w6307_,
		_w6320_,
		_w6336_,
		_w6405_,
		_w6406_
	);
	LUT4 #(
		.INIT('hba00)
	) name580 (
		_w6308_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6407_
	);
	LUT2 #(
		.INIT('h4)
	) name581 (
		_w6371_,
		_w6407_,
		_w6408_
	);
	LUT4 #(
		.INIT('h45ef)
	) name582 (
		_w6311_,
		_w6312_,
		_w6309_,
		_w6310_,
		_w6409_
	);
	LUT4 #(
		.INIT('h5f13)
	) name583 (
		_w6325_,
		_w6332_,
		_w6372_,
		_w6409_,
		_w6410_
	);
	LUT3 #(
		.INIT('h10)
	) name584 (
		_w6406_,
		_w6408_,
		_w6410_,
		_w6411_
	);
	LUT3 #(
		.INIT('h9a)
	) name585 (
		\u2_L13_reg[30]/NET0131 ,
		_w6404_,
		_w6411_,
		_w6412_
	);
	LUT3 #(
		.INIT('hb0)
	) name586 (
		_w6028_,
		_w6027_,
		_w6026_,
		_w6413_
	);
	LUT4 #(
		.INIT('h0cbc)
	) name587 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6414_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w6413_,
		_w6414_,
		_w6415_
	);
	LUT4 #(
		.INIT('hf7c7)
	) name589 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6027_,
		_w6416_
	);
	LUT3 #(
		.INIT('h31)
	) name590 (
		_w6026_,
		_w6025_,
		_w6416_,
		_w6417_
	);
	LUT3 #(
		.INIT('ha2)
	) name591 (
		_w6029_,
		_w6030_,
		_w6027_,
		_w6418_
	);
	LUT4 #(
		.INIT('hce00)
	) name592 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6026_,
		_w6419_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		_w6418_,
		_w6419_,
		_w6420_
	);
	LUT4 #(
		.INIT('h0020)
	) name594 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w6026_,
		_w6421_
	);
	LUT4 #(
		.INIT('h0004)
	) name595 (
		_w6050_,
		_w6025_,
		_w6032_,
		_w6421_,
		_w6422_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name596 (
		_w6415_,
		_w6417_,
		_w6420_,
		_w6422_,
		_w6423_
	);
	LUT4 #(
		.INIT('h0001)
	) name597 (
		_w6026_,
		_w6053_,
		_w6037_,
		_w6358_,
		_w6424_
	);
	LUT3 #(
		.INIT('h02)
	) name598 (
		_w6026_,
		_w6055_,
		_w6033_,
		_w6425_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		_w6424_,
		_w6425_,
		_w6426_
	);
	LUT3 #(
		.INIT('h56)
	) name600 (
		\u2_L13_reg[3]/NET0131 ,
		_w6423_,
		_w6426_,
		_w6427_
	);
	LUT4 #(
		.INIT('h9600)
	) name601 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6428_
	);
	LUT3 #(
		.INIT('h19)
	) name602 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w6429_
	);
	LUT4 #(
		.INIT('h0013)
	) name603 (
		_w5893_,
		_w6069_,
		_w6429_,
		_w6428_,
		_w6430_
	);
	LUT4 #(
		.INIT('h0141)
	) name604 (
		_w5885_,
		_w5886_,
		_w5887_,
		_w5888_,
		_w6431_
	);
	LUT3 #(
		.INIT('h08)
	) name605 (
		_w5886_,
		_w5888_,
		_w5889_,
		_w6432_
	);
	LUT3 #(
		.INIT('h28)
	) name606 (
		_w5885_,
		_w5886_,
		_w5887_,
		_w6433_
	);
	LUT4 #(
		.INIT('hbe7f)
	) name607 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6434_
	);
	LUT4 #(
		.INIT('h0b00)
	) name608 (
		_w6432_,
		_w6433_,
		_w6431_,
		_w6434_,
		_w6435_
	);
	LUT4 #(
		.INIT('hf77f)
	) name609 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w6436_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		_w5885_,
		_w6436_,
		_w6437_
	);
	LUT4 #(
		.INIT('h0e04)
	) name611 (
		_w5884_,
		_w6435_,
		_w6437_,
		_w6430_,
		_w6438_
	);
	LUT2 #(
		.INIT('h9)
	) name612 (
		\u2_L13_reg[9]/NET0131 ,
		_w6438_,
		_w6439_
	);
	LUT4 #(
		.INIT('h1a00)
	) name613 (
		_w6161_,
		_w6162_,
		_w6163_,
		_w6166_,
		_w6440_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		_w6164_,
		_w6163_,
		_w6441_
	);
	LUT4 #(
		.INIT('h00c4)
	) name615 (
		_w6161_,
		_w6162_,
		_w6163_,
		_w6166_,
		_w6442_
	);
	LUT4 #(
		.INIT('h2022)
	) name616 (
		_w6176_,
		_w6201_,
		_w6441_,
		_w6442_,
		_w6443_
	);
	LUT2 #(
		.INIT('h2)
	) name617 (
		_w6161_,
		_w6166_,
		_w6444_
	);
	LUT4 #(
		.INIT('he000)
	) name618 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6445_
	);
	LUT4 #(
		.INIT('h0109)
	) name619 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6166_,
		_w6446_
	);
	LUT4 #(
		.INIT('h0405)
	) name620 (
		_w6194_,
		_w6444_,
		_w6446_,
		_w6445_,
		_w6447_
	);
	LUT4 #(
		.INIT('h45cf)
	) name621 (
		_w6183_,
		_w6440_,
		_w6443_,
		_w6447_,
		_w6448_
	);
	LUT4 #(
		.INIT('h0020)
	) name622 (
		_w6161_,
		_w6162_,
		_w6163_,
		_w6166_,
		_w6449_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name623 (
		_w6164_,
		_w6161_,
		_w6162_,
		_w6163_,
		_w6450_
	);
	LUT3 #(
		.INIT('h31)
	) name624 (
		_w6166_,
		_w6449_,
		_w6450_,
		_w6451_
	);
	LUT3 #(
		.INIT('h65)
	) name625 (
		\u2_L13_reg[18]/P0001 ,
		_w6448_,
		_w6451_,
		_w6452_
	);
	LUT4 #(
		.INIT('hc963)
	) name626 (
		decrypt_pad,
		\u2_R12_reg[4]/NET0131 ,
		\u2_uk_K_r12_reg[10]/P0001 ,
		\u2_uk_K_r12_reg[34]/NET0131 ,
		_w6453_
	);
	LUT4 #(
		.INIT('hc693)
	) name627 (
		decrypt_pad,
		\u2_R12_reg[1]/NET0131 ,
		\u2_uk_K_r12_reg[32]/NET0131 ,
		\u2_uk_K_r12_reg[40]/NET0131 ,
		_w6454_
	);
	LUT4 #(
		.INIT('hc693)
	) name628 (
		decrypt_pad,
		\u2_R12_reg[3]/NET0131 ,
		\u2_uk_K_r12_reg[24]/NET0131 ,
		\u2_uk_K_r12_reg[32]/NET0131 ,
		_w6455_
	);
	LUT4 #(
		.INIT('hc693)
	) name629 (
		decrypt_pad,
		\u2_R12_reg[2]/NET0131 ,
		\u2_uk_K_r12_reg[47]/NET0131 ,
		\u2_uk_K_r12_reg[55]/NET0131 ,
		_w6456_
	);
	LUT4 #(
		.INIT('hc963)
	) name630 (
		decrypt_pad,
		\u2_R12_reg[5]/NET0131 ,
		\u2_uk_K_r12_reg[13]/NET0131 ,
		\u2_uk_K_r12_reg[5]/NET0131 ,
		_w6457_
	);
	LUT4 #(
		.INIT('hc693)
	) name631 (
		decrypt_pad,
		\u2_R12_reg[32]/NET0131 ,
		\u2_uk_K_r12_reg[11]/NET0131 ,
		\u2_uk_K_r12_reg[19]/NET0131 ,
		_w6458_
	);
	LUT4 #(
		.INIT('hff7c)
	) name632 (
		_w6455_,
		_w6456_,
		_w6457_,
		_w6458_,
		_w6459_
	);
	LUT2 #(
		.INIT('h2)
	) name633 (
		_w6454_,
		_w6459_,
		_w6460_
	);
	LUT4 #(
		.INIT('h2000)
	) name634 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6461_
	);
	LUT4 #(
		.INIT('h9bff)
	) name635 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6462_
	);
	LUT4 #(
		.INIT('h0400)
	) name636 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6463_
	);
	LUT3 #(
		.INIT('h0d)
	) name637 (
		_w6455_,
		_w6462_,
		_w6463_,
		_w6464_
	);
	LUT3 #(
		.INIT('h45)
	) name638 (
		_w6453_,
		_w6460_,
		_w6464_,
		_w6465_
	);
	LUT3 #(
		.INIT('h02)
	) name639 (
		_w6456_,
		_w6457_,
		_w6458_,
		_w6466_
	);
	LUT4 #(
		.INIT('hf3d1)
	) name640 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6467_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		_w6455_,
		_w6467_,
		_w6468_
	);
	LUT2 #(
		.INIT('h4)
	) name642 (
		_w6455_,
		_w6454_,
		_w6469_
	);
	LUT4 #(
		.INIT('haafc)
	) name643 (
		_w6455_,
		_w6456_,
		_w6457_,
		_w6454_,
		_w6470_
	);
	LUT2 #(
		.INIT('h2)
	) name644 (
		_w6455_,
		_w6456_,
		_w6471_
	);
	LUT3 #(
		.INIT('hd0)
	) name645 (
		_w6455_,
		_w6456_,
		_w6454_,
		_w6472_
	);
	LUT3 #(
		.INIT('h0e)
	) name646 (
		_w6456_,
		_w6457_,
		_w6458_,
		_w6473_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name647 (
		_w6458_,
		_w6470_,
		_w6472_,
		_w6473_,
		_w6474_
	);
	LUT3 #(
		.INIT('h8a)
	) name648 (
		_w6453_,
		_w6468_,
		_w6474_,
		_w6475_
	);
	LUT4 #(
		.INIT('hfdae)
	) name649 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6476_
	);
	LUT4 #(
		.INIT('h0008)
	) name650 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6477_
	);
	LUT4 #(
		.INIT('h6fe7)
	) name651 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6478_
	);
	LUT4 #(
		.INIT('h0155)
	) name652 (
		_w6455_,
		_w6476_,
		_w6453_,
		_w6478_,
		_w6479_
	);
	LUT2 #(
		.INIT('h2)
	) name653 (
		_w6455_,
		_w6454_,
		_w6480_
	);
	LUT4 #(
		.INIT('h0200)
	) name654 (
		_w6455_,
		_w6456_,
		_w6454_,
		_w6458_,
		_w6481_
	);
	LUT3 #(
		.INIT('h07)
	) name655 (
		_w6466_,
		_w6480_,
		_w6481_,
		_w6482_
	);
	LUT2 #(
		.INIT('h4)
	) name656 (
		_w6479_,
		_w6482_,
		_w6483_
	);
	LUT4 #(
		.INIT('h5655)
	) name657 (
		\u2_L12_reg[31]/NET0131 ,
		_w6475_,
		_w6465_,
		_w6483_,
		_w6484_
	);
	LUT4 #(
		.INIT('hc693)
	) name658 (
		decrypt_pad,
		\u2_R12_reg[23]/NET0131 ,
		\u2_uk_K_r12_reg[30]/NET0131 ,
		\u2_uk_K_r12_reg[36]/NET0131 ,
		_w6485_
	);
	LUT4 #(
		.INIT('hc963)
	) name659 (
		decrypt_pad,
		\u2_R12_reg[22]/NET0131 ,
		\u2_uk_K_r12_reg[23]/NET0131 ,
		\u2_uk_K_r12_reg[45]/NET0131 ,
		_w6486_
	);
	LUT4 #(
		.INIT('hc693)
	) name660 (
		decrypt_pad,
		\u2_R12_reg[20]/NET0131 ,
		\u2_uk_K_r12_reg[35]/NET0131 ,
		\u2_uk_K_r12_reg[45]/NET0131 ,
		_w6487_
	);
	LUT4 #(
		.INIT('hc963)
	) name661 (
		decrypt_pad,
		\u2_R12_reg[25]/NET0131 ,
		\u2_uk_K_r12_reg[2]/NET0131 ,
		\u2_uk_K_r12_reg[51]/NET0131 ,
		_w6488_
	);
	LUT4 #(
		.INIT('hc963)
	) name662 (
		decrypt_pad,
		\u2_R12_reg[21]/NET0131 ,
		\u2_uk_K_r12_reg[1]/NET0131 ,
		\u2_uk_K_r12_reg[50]/NET0131 ,
		_w6489_
	);
	LUT3 #(
		.INIT('h20)
	) name663 (
		_w6487_,
		_w6489_,
		_w6488_,
		_w6490_
	);
	LUT4 #(
		.INIT('h168a)
	) name664 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6491_
	);
	LUT2 #(
		.INIT('h1)
	) name665 (
		_w6485_,
		_w6491_,
		_w6492_
	);
	LUT4 #(
		.INIT('hc693)
	) name666 (
		decrypt_pad,
		\u2_R12_reg[24]/NET0131 ,
		\u2_uk_K_r12_reg[1]/NET0131 ,
		\u2_uk_K_r12_reg[7]/P0001 ,
		_w6493_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name667 (
		_w6485_,
		_w6486_,
		_w6487_,
		_w6489_,
		_w6494_
	);
	LUT4 #(
		.INIT('h0004)
	) name668 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6495_
	);
	LUT4 #(
		.INIT('h3ffb)
	) name669 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6496_
	);
	LUT3 #(
		.INIT('h2a)
	) name670 (
		_w6493_,
		_w6494_,
		_w6496_,
		_w6497_
	);
	LUT2 #(
		.INIT('h4)
	) name671 (
		_w6492_,
		_w6497_,
		_w6498_
	);
	LUT4 #(
		.INIT('h0040)
	) name672 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6499_
	);
	LUT4 #(
		.INIT('h0800)
	) name673 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6500_
	);
	LUT4 #(
		.INIT('h0200)
	) name674 (
		_w6485_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6501_
	);
	LUT3 #(
		.INIT('h01)
	) name675 (
		_w6500_,
		_w6501_,
		_w6499_,
		_w6502_
	);
	LUT4 #(
		.INIT('h1400)
	) name676 (
		_w6485_,
		_w6486_,
		_w6487_,
		_w6489_,
		_w6503_
	);
	LUT2 #(
		.INIT('h8)
	) name677 (
		_w6485_,
		_w6486_,
		_w6504_
	);
	LUT4 #(
		.INIT('h0080)
	) name678 (
		_w6485_,
		_w6486_,
		_w6487_,
		_w6489_,
		_w6505_
	);
	LUT4 #(
		.INIT('h0010)
	) name679 (
		_w6485_,
		_w6486_,
		_w6487_,
		_w6488_,
		_w6506_
	);
	LUT4 #(
		.INIT('hfded)
	) name680 (
		_w6485_,
		_w6486_,
		_w6487_,
		_w6488_,
		_w6507_
	);
	LUT3 #(
		.INIT('h10)
	) name681 (
		_w6503_,
		_w6505_,
		_w6507_,
		_w6508_
	);
	LUT3 #(
		.INIT('h15)
	) name682 (
		_w6493_,
		_w6502_,
		_w6508_,
		_w6509_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name683 (
		_w6485_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6510_
	);
	LUT2 #(
		.INIT('h1)
	) name684 (
		_w6486_,
		_w6510_,
		_w6511_
	);
	LUT4 #(
		.INIT('h0010)
	) name685 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6512_
	);
	LUT4 #(
		.INIT('h77ef)
	) name686 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6513_
	);
	LUT3 #(
		.INIT('h01)
	) name687 (
		_w6487_,
		_w6489_,
		_w6488_,
		_w6514_
	);
	LUT4 #(
		.INIT('he4f5)
	) name688 (
		_w6485_,
		_w6486_,
		_w6513_,
		_w6514_,
		_w6515_
	);
	LUT2 #(
		.INIT('h4)
	) name689 (
		_w6511_,
		_w6515_,
		_w6516_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name690 (
		\u2_L12_reg[11]/NET0131 ,
		_w6509_,
		_w6498_,
		_w6516_,
		_w6517_
	);
	LUT4 #(
		.INIT('hc963)
	) name691 (
		decrypt_pad,
		\u2_R12_reg[28]/NET0131 ,
		\u2_uk_K_r12_reg[14]/NET0131 ,
		\u2_uk_K_r12_reg[8]/NET0131 ,
		_w6518_
	);
	LUT4 #(
		.INIT('hc693)
	) name692 (
		decrypt_pad,
		\u2_R12_reg[27]/NET0131 ,
		\u2_uk_K_r12_reg[21]/NET0131 ,
		\u2_uk_K_r12_reg[31]/NET0131 ,
		_w6519_
	);
	LUT4 #(
		.INIT('hc693)
	) name693 (
		decrypt_pad,
		\u2_R12_reg[26]/NET0131 ,
		\u2_uk_K_r12_reg[43]/NET0131 ,
		\u2_uk_K_r12_reg[49]/NET0131 ,
		_w6520_
	);
	LUT4 #(
		.INIT('hc693)
	) name694 (
		decrypt_pad,
		\u2_R12_reg[24]/NET0131 ,
		\u2_uk_K_r12_reg[23]/NET0131 ,
		\u2_uk_K_r12_reg[29]/NET0131 ,
		_w6521_
	);
	LUT4 #(
		.INIT('hc693)
	) name695 (
		decrypt_pad,
		\u2_R12_reg[29]/NET0131 ,
		\u2_uk_K_r12_reg[0]/NET0131 ,
		\u2_uk_K_r12_reg[37]/NET0131 ,
		_w6522_
	);
	LUT4 #(
		.INIT('hc693)
	) name696 (
		decrypt_pad,
		\u2_R12_reg[25]/NET0131 ,
		\u2_uk_K_r12_reg[31]/NET0131 ,
		\u2_uk_K_r12_reg[9]/NET0131 ,
		_w6523_
	);
	LUT4 #(
		.INIT('h0004)
	) name697 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6524_
	);
	LUT4 #(
		.INIT('h27fb)
	) name698 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6525_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w6519_,
		_w6525_,
		_w6526_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w6519_,
		_w6522_,
		_w6527_
	);
	LUT3 #(
		.INIT('h10)
	) name701 (
		_w6520_,
		_w6523_,
		_w6521_,
		_w6528_
	);
	LUT2 #(
		.INIT('h4)
	) name702 (
		_w6527_,
		_w6528_,
		_w6529_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		_w6520_,
		_w6521_,
		_w6530_
	);
	LUT3 #(
		.INIT('h3b)
	) name704 (
		_w6519_,
		_w6522_,
		_w6523_,
		_w6531_
	);
	LUT4 #(
		.INIT('h8000)
	) name705 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6532_
	);
	LUT3 #(
		.INIT('h0d)
	) name706 (
		_w6530_,
		_w6531_,
		_w6532_,
		_w6533_
	);
	LUT4 #(
		.INIT('h5455)
	) name707 (
		_w6518_,
		_w6526_,
		_w6529_,
		_w6533_,
		_w6534_
	);
	LUT3 #(
		.INIT('hd3)
	) name708 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6535_
	);
	LUT2 #(
		.INIT('h8)
	) name709 (
		_w6519_,
		_w6521_,
		_w6536_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		_w6535_,
		_w6536_,
		_w6537_
	);
	LUT3 #(
		.INIT('he3)
	) name711 (
		_w6520_,
		_w6523_,
		_w6521_,
		_w6538_
	);
	LUT4 #(
		.INIT('h0008)
	) name712 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6539_
	);
	LUT4 #(
		.INIT('hfff6)
	) name713 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6540_
	);
	LUT3 #(
		.INIT('hd0)
	) name714 (
		_w6527_,
		_w6538_,
		_w6540_,
		_w6541_
	);
	LUT2 #(
		.INIT('h6)
	) name715 (
		_w6520_,
		_w6521_,
		_w6542_
	);
	LUT4 #(
		.INIT('h4010)
	) name716 (
		_w6519_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6543_
	);
	LUT2 #(
		.INIT('h4)
	) name717 (
		_w6522_,
		_w6520_,
		_w6544_
	);
	LUT4 #(
		.INIT('h0040)
	) name718 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6545_
	);
	LUT4 #(
		.INIT('hfab6)
	) name719 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6546_
	);
	LUT3 #(
		.INIT('h31)
	) name720 (
		_w6519_,
		_w6543_,
		_w6546_,
		_w6547_
	);
	LUT4 #(
		.INIT('h7500)
	) name721 (
		_w6518_,
		_w6537_,
		_w6541_,
		_w6547_,
		_w6548_
	);
	LUT3 #(
		.INIT('h65)
	) name722 (
		\u2_L12_reg[22]/NET0131 ,
		_w6534_,
		_w6548_,
		_w6549_
	);
	LUT4 #(
		.INIT('hc693)
	) name723 (
		decrypt_pad,
		\u2_R12_reg[14]/NET0131 ,
		\u2_uk_K_r12_reg[20]/NET0131 ,
		\u2_uk_K_r12_reg[53]/NET0131 ,
		_w6550_
	);
	LUT4 #(
		.INIT('hc693)
	) name724 (
		decrypt_pad,
		\u2_R12_reg[13]/NET0131 ,
		\u2_uk_K_r12_reg[19]/NET0131 ,
		\u2_uk_K_r12_reg[27]/NET0131 ,
		_w6551_
	);
	LUT4 #(
		.INIT('hc693)
	) name725 (
		decrypt_pad,
		\u2_R12_reg[12]/NET0131 ,
		\u2_uk_K_r12_reg[25]/NET0131 ,
		\u2_uk_K_r12_reg[33]/NET0131 ,
		_w6552_
	);
	LUT4 #(
		.INIT('hc963)
	) name726 (
		decrypt_pad,
		\u2_R12_reg[17]/NET0131 ,
		\u2_uk_K_r12_reg[17]/NET0131 ,
		\u2_uk_K_r12_reg[41]/NET0131 ,
		_w6553_
	);
	LUT3 #(
		.INIT('h80)
	) name727 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6554_
	);
	LUT4 #(
		.INIT('hc963)
	) name728 (
		decrypt_pad,
		\u2_R12_reg[15]/NET0131 ,
		\u2_uk_K_r12_reg[4]/NET0131 ,
		\u2_uk_K_r12_reg[53]/NET0131 ,
		_w6555_
	);
	LUT4 #(
		.INIT('h0001)
	) name729 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6553_,
		_w6556_
	);
	LUT4 #(
		.INIT('h5ffe)
	) name730 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6553_,
		_w6557_
	);
	LUT2 #(
		.INIT('h2)
	) name731 (
		_w6550_,
		_w6557_,
		_w6558_
	);
	LUT4 #(
		.INIT('h0080)
	) name732 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6553_,
		_w6559_
	);
	LUT2 #(
		.INIT('h4)
	) name733 (
		_w6552_,
		_w6553_,
		_w6560_
	);
	LUT3 #(
		.INIT('h20)
	) name734 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6561_
	);
	LUT4 #(
		.INIT('h0020)
	) name735 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6562_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w6559_,
		_w6562_,
		_w6563_
	);
	LUT4 #(
		.INIT('h0400)
	) name737 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6553_,
		_w6564_
	);
	LUT2 #(
		.INIT('h9)
	) name738 (
		_w6551_,
		_w6552_,
		_w6565_
	);
	LUT4 #(
		.INIT('h0012)
	) name739 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6550_,
		_w6566_
	);
	LUT4 #(
		.INIT('hc963)
	) name740 (
		decrypt_pad,
		\u2_R12_reg[16]/NET0131 ,
		\u2_uk_K_r12_reg[12]/NET0131 ,
		\u2_uk_K_r12_reg[4]/NET0131 ,
		_w6567_
	);
	LUT3 #(
		.INIT('h04)
	) name741 (
		_w6566_,
		_w6567_,
		_w6564_,
		_w6568_
	);
	LUT3 #(
		.INIT('h40)
	) name742 (
		_w6558_,
		_w6563_,
		_w6568_,
		_w6569_
	);
	LUT4 #(
		.INIT('h0040)
	) name743 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6570_
	);
	LUT4 #(
		.INIT('h0004)
	) name744 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6553_,
		_w6571_
	);
	LUT3 #(
		.INIT('h80)
	) name745 (
		_w6551_,
		_w6555_,
		_w6550_,
		_w6572_
	);
	LUT4 #(
		.INIT('h0800)
	) name746 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6550_,
		_w6573_
	);
	LUT3 #(
		.INIT('h01)
	) name747 (
		_w6571_,
		_w6573_,
		_w6570_,
		_w6574_
	);
	LUT4 #(
		.INIT('h0200)
	) name748 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6575_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name749 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6576_
	);
	LUT4 #(
		.INIT('ha3af)
	) name750 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6577_
	);
	LUT4 #(
		.INIT('h1302)
	) name751 (
		_w6555_,
		_w6567_,
		_w6554_,
		_w6577_,
		_w6578_
	);
	LUT3 #(
		.INIT('h80)
	) name752 (
		_w6576_,
		_w6574_,
		_w6578_,
		_w6579_
	);
	LUT4 #(
		.INIT('h0400)
	) name753 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6580_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name754 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6581_
	);
	LUT2 #(
		.INIT('h2)
	) name755 (
		_w6555_,
		_w6581_,
		_w6582_
	);
	LUT4 #(
		.INIT('hf2f3)
	) name756 (
		_w6555_,
		_w6559_,
		_w6550_,
		_w6561_,
		_w6583_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		_w6582_,
		_w6583_,
		_w6584_
	);
	LUT4 #(
		.INIT('ha955)
	) name758 (
		\u2_L12_reg[20]/NET0131 ,
		_w6569_,
		_w6579_,
		_w6584_,
		_w6585_
	);
	LUT4 #(
		.INIT('h1000)
	) name759 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6586_
	);
	LUT2 #(
		.INIT('h2)
	) name760 (
		_w6453_,
		_w6586_,
		_w6587_
	);
	LUT4 #(
		.INIT('hfb05)
	) name761 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6588_
	);
	LUT3 #(
		.INIT('h80)
	) name762 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6589_
	);
	LUT4 #(
		.INIT('h4401)
	) name763 (
		_w6455_,
		_w6456_,
		_w6454_,
		_w6458_,
		_w6590_
	);
	LUT4 #(
		.INIT('h000d)
	) name764 (
		_w6455_,
		_w6588_,
		_w6589_,
		_w6590_,
		_w6591_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		_w6587_,
		_w6591_,
		_w6592_
	);
	LUT4 #(
		.INIT('h3c9f)
	) name766 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6593_
	);
	LUT2 #(
		.INIT('h2)
	) name767 (
		_w6455_,
		_w6593_,
		_w6594_
	);
	LUT4 #(
		.INIT('hf3ec)
	) name768 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6595_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		_w6455_,
		_w6595_,
		_w6596_
	);
	LUT3 #(
		.INIT('h01)
	) name770 (
		_w6477_,
		_w6453_,
		_w6461_,
		_w6597_
	);
	LUT3 #(
		.INIT('h10)
	) name771 (
		_w6596_,
		_w6594_,
		_w6597_,
		_w6598_
	);
	LUT3 #(
		.INIT('ha9)
	) name772 (
		\u2_L12_reg[17]/NET0131 ,
		_w6592_,
		_w6598_,
		_w6599_
	);
	LUT4 #(
		.INIT('h3fd2)
	) name773 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6600_
	);
	LUT4 #(
		.INIT('hab6f)
	) name774 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6601_
	);
	LUT4 #(
		.INIT('h0200)
	) name775 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6602_
	);
	LUT4 #(
		.INIT('h00e4)
	) name776 (
		_w6485_,
		_w6601_,
		_w6600_,
		_w6602_,
		_w6603_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w6493_,
		_w6603_,
		_w6604_
	);
	LUT4 #(
		.INIT('hcf6f)
	) name778 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6605_
	);
	LUT2 #(
		.INIT('h2)
	) name779 (
		_w6485_,
		_w6605_,
		_w6606_
	);
	LUT4 #(
		.INIT('h0102)
	) name780 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6607_
	);
	LUT4 #(
		.INIT('h77dc)
	) name781 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6608_
	);
	LUT4 #(
		.INIT('h0302)
	) name782 (
		_w6485_,
		_w6506_,
		_w6500_,
		_w6608_,
		_w6609_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name783 (
		_w6493_,
		_w6606_,
		_w6607_,
		_w6609_,
		_w6610_
	);
	LUT4 #(
		.INIT('h2000)
	) name784 (
		_w6485_,
		_w6486_,
		_w6489_,
		_w6488_,
		_w6611_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w6495_,
		_w6611_,
		_w6612_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name786 (
		\u2_L12_reg[29]/NET0131 ,
		_w6610_,
		_w6604_,
		_w6612_,
		_w6613_
	);
	LUT4 #(
		.INIT('hc693)
	) name787 (
		decrypt_pad,
		\u2_R12_reg[6]/NET0131 ,
		\u2_uk_K_r12_reg[18]/NET0131 ,
		\u2_uk_K_r12_reg[26]/NET0131 ,
		_w6614_
	);
	LUT4 #(
		.INIT('hc693)
	) name788 (
		decrypt_pad,
		\u2_R12_reg[9]/NET0131 ,
		\u2_uk_K_r12_reg[40]/NET0131 ,
		\u2_uk_K_r12_reg[48]/NET0131 ,
		_w6615_
	);
	LUT4 #(
		.INIT('hc693)
	) name789 (
		decrypt_pad,
		\u2_R12_reg[5]/NET0131 ,
		\u2_uk_K_r12_reg[27]/NET0131 ,
		\u2_uk_K_r12_reg[3]/NET0131 ,
		_w6616_
	);
	LUT2 #(
		.INIT('h4)
	) name790 (
		_w6615_,
		_w6616_,
		_w6617_
	);
	LUT4 #(
		.INIT('hc963)
	) name791 (
		decrypt_pad,
		\u2_R12_reg[4]/NET0131 ,
		\u2_uk_K_r12_reg[24]/NET0131 ,
		\u2_uk_K_r12_reg[48]/NET0131 ,
		_w6618_
	);
	LUT2 #(
		.INIT('h2)
	) name792 (
		_w6615_,
		_w6616_,
		_w6619_
	);
	LUT4 #(
		.INIT('h0406)
	) name793 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6620_
	);
	LUT4 #(
		.INIT('hc693)
	) name794 (
		decrypt_pad,
		\u2_R12_reg[7]/NET0131 ,
		\u2_uk_K_r12_reg[12]/NET0131 ,
		\u2_uk_K_r12_reg[20]/NET0131 ,
		_w6621_
	);
	LUT3 #(
		.INIT('h80)
	) name795 (
		_w6621_,
		_w6614_,
		_w6618_,
		_w6622_
	);
	LUT4 #(
		.INIT('hc963)
	) name796 (
		decrypt_pad,
		\u2_R12_reg[8]/NET0131 ,
		\u2_uk_K_r12_reg[11]/NET0131 ,
		\u2_uk_K_r12_reg[3]/NET0131 ,
		_w6623_
	);
	LUT4 #(
		.INIT('h0013)
	) name797 (
		_w6619_,
		_w6620_,
		_w6622_,
		_w6623_,
		_w6624_
	);
	LUT2 #(
		.INIT('h2)
	) name798 (
		_w6615_,
		_w6618_,
		_w6625_
	);
	LUT4 #(
		.INIT('hf070)
	) name799 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6626_
	);
	LUT3 #(
		.INIT('h0e)
	) name800 (
		_w6621_,
		_w6616_,
		_w6614_,
		_w6627_
	);
	LUT4 #(
		.INIT('hff04)
	) name801 (
		_w6621_,
		_w6615_,
		_w6616_,
		_w6614_,
		_w6628_
	);
	LUT4 #(
		.INIT('h2fdd)
	) name802 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6629_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name803 (
		_w6621_,
		_w6626_,
		_w6628_,
		_w6629_,
		_w6630_
	);
	LUT2 #(
		.INIT('h8)
	) name804 (
		_w6624_,
		_w6630_,
		_w6631_
	);
	LUT4 #(
		.INIT('h51f5)
	) name805 (
		_w6621_,
		_w6615_,
		_w6614_,
		_w6618_,
		_w6632_
	);
	LUT2 #(
		.INIT('h2)
	) name806 (
		_w6616_,
		_w6632_,
		_w6633_
	);
	LUT3 #(
		.INIT('h8a)
	) name807 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6634_
	);
	LUT3 #(
		.INIT('hae)
	) name808 (
		_w6621_,
		_w6616_,
		_w6614_,
		_w6635_
	);
	LUT2 #(
		.INIT('h9)
	) name809 (
		_w6615_,
		_w6618_,
		_w6636_
	);
	LUT3 #(
		.INIT('h10)
	) name810 (
		_w6635_,
		_w6634_,
		_w6636_,
		_w6637_
	);
	LUT3 #(
		.INIT('h01)
	) name811 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6638_
	);
	LUT4 #(
		.INIT('h0100)
	) name812 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6639_
	);
	LUT2 #(
		.INIT('h2)
	) name813 (
		_w6623_,
		_w6639_,
		_w6640_
	);
	LUT3 #(
		.INIT('h10)
	) name814 (
		_w6637_,
		_w6633_,
		_w6640_,
		_w6641_
	);
	LUT3 #(
		.INIT('h04)
	) name815 (
		_w6616_,
		_w6614_,
		_w6618_,
		_w6642_
	);
	LUT4 #(
		.INIT('h0010)
	) name816 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6643_
	);
	LUT4 #(
		.INIT('hf3ef)
	) name817 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6644_
	);
	LUT3 #(
		.INIT('h0b)
	) name818 (
		_w6616_,
		_w6614_,
		_w6618_,
		_w6645_
	);
	LUT4 #(
		.INIT('h4404)
	) name819 (
		_w6621_,
		_w6615_,
		_w6616_,
		_w6614_,
		_w6646_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name820 (
		_w6621_,
		_w6644_,
		_w6645_,
		_w6646_,
		_w6647_
	);
	LUT4 #(
		.INIT('ha955)
	) name821 (
		\u2_L12_reg[2]/NET0131 ,
		_w6631_,
		_w6641_,
		_w6647_,
		_w6648_
	);
	LUT4 #(
		.INIT('hc693)
	) name822 (
		decrypt_pad,
		\u2_R12_reg[32]/NET0131 ,
		\u2_uk_K_r12_reg[28]/NET0131 ,
		\u2_uk_K_r12_reg[38]/NET0131 ,
		_w6649_
	);
	LUT4 #(
		.INIT('hc693)
	) name823 (
		decrypt_pad,
		\u2_R12_reg[31]/P0001 ,
		\u2_uk_K_r12_reg[22]/NET0131 ,
		\u2_uk_K_r12_reg[28]/NET0131 ,
		_w6650_
	);
	LUT4 #(
		.INIT('hc963)
	) name824 (
		decrypt_pad,
		\u2_R12_reg[30]/NET0131 ,
		\u2_uk_K_r12_reg[16]/NET0131 ,
		\u2_uk_K_r12_reg[38]/NET0131 ,
		_w6651_
	);
	LUT4 #(
		.INIT('hc963)
	) name825 (
		decrypt_pad,
		\u2_R12_reg[29]/NET0131 ,
		\u2_uk_K_r12_reg[15]/NET0131 ,
		\u2_uk_K_r12_reg[9]/NET0131 ,
		_w6652_
	);
	LUT4 #(
		.INIT('hc693)
	) name826 (
		decrypt_pad,
		\u2_R12_reg[28]/NET0131 ,
		\u2_uk_K_r12_reg[37]/NET0131 ,
		\u2_uk_K_r12_reg[43]/NET0131 ,
		_w6653_
	);
	LUT4 #(
		.INIT('hc963)
	) name827 (
		decrypt_pad,
		\u2_R12_reg[1]/NET0131 ,
		\u2_uk_K_r12_reg[0]/NET0131 ,
		\u2_uk_K_r12_reg[49]/NET0131 ,
		_w6654_
	);
	LUT4 #(
		.INIT('ha6f3)
	) name828 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6655_
	);
	LUT3 #(
		.INIT('h01)
	) name829 (
		_w6651_,
		_w6652_,
		_w6653_,
		_w6656_
	);
	LUT4 #(
		.INIT('h0080)
	) name830 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6657_
	);
	LUT4 #(
		.INIT('h008d)
	) name831 (
		_w6650_,
		_w6655_,
		_w6656_,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		_w6649_,
		_w6658_,
		_w6659_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name833 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6660_
	);
	LUT2 #(
		.INIT('h2)
	) name834 (
		_w6650_,
		_w6660_,
		_w6661_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name835 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6650_,
		_w6662_
	);
	LUT2 #(
		.INIT('h4)
	) name836 (
		_w6662_,
		_w6653_,
		_w6663_
	);
	LUT3 #(
		.INIT('h23)
	) name837 (
		_w6654_,
		_w6650_,
		_w6653_,
		_w6664_
	);
	LUT3 #(
		.INIT('hca)
	) name838 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6665_
	);
	LUT3 #(
		.INIT('h20)
	) name839 (
		_w6652_,
		_w6654_,
		_w6653_,
		_w6666_
	);
	LUT4 #(
		.INIT('h0400)
	) name840 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6667_
	);
	LUT3 #(
		.INIT('h07)
	) name841 (
		_w6664_,
		_w6665_,
		_w6667_,
		_w6668_
	);
	LUT4 #(
		.INIT('h00ef)
	) name842 (
		_w6663_,
		_w6661_,
		_w6668_,
		_w6649_,
		_w6669_
	);
	LUT4 #(
		.INIT('heff7)
	) name843 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6670_
	);
	LUT4 #(
		.INIT('h0020)
	) name844 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6671_
	);
	LUT4 #(
		.INIT('h0001)
	) name845 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6672_
	);
	LUT4 #(
		.INIT('hefd6)
	) name846 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6673_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		_w6650_,
		_w6673_,
		_w6674_
	);
	LUT3 #(
		.INIT('h40)
	) name848 (
		_w6652_,
		_w6653_,
		_w6649_,
		_w6675_
	);
	LUT4 #(
		.INIT('hcdef)
	) name849 (
		_w6651_,
		_w6650_,
		_w6666_,
		_w6675_,
		_w6676_
	);
	LUT2 #(
		.INIT('h4)
	) name850 (
		_w6674_,
		_w6676_,
		_w6677_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name851 (
		\u2_L12_reg[5]/NET0131 ,
		_w6669_,
		_w6659_,
		_w6677_,
		_w6678_
	);
	LUT4 #(
		.INIT('he63f)
	) name852 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6679_
	);
	LUT2 #(
		.INIT('h2)
	) name853 (
		_w6485_,
		_w6679_,
		_w6680_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name854 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6681_
	);
	LUT4 #(
		.INIT('h1000)
	) name855 (
		_w6485_,
		_w6486_,
		_w6487_,
		_w6488_,
		_w6682_
	);
	LUT4 #(
		.INIT('h0032)
	) name856 (
		_w6485_,
		_w6495_,
		_w6681_,
		_w6682_,
		_w6683_
	);
	LUT3 #(
		.INIT('h45)
	) name857 (
		_w6493_,
		_w6680_,
		_w6683_,
		_w6684_
	);
	LUT4 #(
		.INIT('heeae)
	) name858 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6685_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w6485_,
		_w6685_,
		_w6686_
	);
	LUT3 #(
		.INIT('h80)
	) name860 (
		_w6486_,
		_w6489_,
		_w6488_,
		_w6687_
	);
	LUT4 #(
		.INIT('h2000)
	) name861 (
		_w6485_,
		_w6486_,
		_w6487_,
		_w6488_,
		_w6688_
	);
	LUT3 #(
		.INIT('h01)
	) name862 (
		_w6512_,
		_w6687_,
		_w6688_,
		_w6689_
	);
	LUT3 #(
		.INIT('hb6)
	) name863 (
		_w6487_,
		_w6489_,
		_w6488_,
		_w6690_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name864 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6691_
	);
	LUT4 #(
		.INIT('h4445)
	) name865 (
		_w6485_,
		_w6486_,
		_w6487_,
		_w6488_,
		_w6692_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name866 (
		_w6504_,
		_w6690_,
		_w6691_,
		_w6692_,
		_w6693_
	);
	LUT4 #(
		.INIT('h7500)
	) name867 (
		_w6493_,
		_w6686_,
		_w6689_,
		_w6693_,
		_w6694_
	);
	LUT3 #(
		.INIT('h65)
	) name868 (
		\u2_L12_reg[4]/NET0131 ,
		_w6684_,
		_w6694_,
		_w6695_
	);
	LUT4 #(
		.INIT('hf3db)
	) name869 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6696_
	);
	LUT4 #(
		.INIT('h8000)
	) name870 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6697_
	);
	LUT4 #(
		.INIT('h6fff)
	) name871 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6698_
	);
	LUT4 #(
		.INIT('hfdbd)
	) name872 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6699_
	);
	LUT4 #(
		.INIT('hc480)
	) name873 (
		_w6555_,
		_w6698_,
		_w6699_,
		_w6696_,
		_w6700_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		_w6567_,
		_w6700_,
		_w6701_
	);
	LUT3 #(
		.INIT('h08)
	) name875 (
		_w6551_,
		_w6552_,
		_w6550_,
		_w6702_
	);
	LUT4 #(
		.INIT('h0040)
	) name876 (
		_w6555_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6703_
	);
	LUT3 #(
		.INIT('h01)
	) name877 (
		_w6556_,
		_w6702_,
		_w6703_,
		_w6704_
	);
	LUT2 #(
		.INIT('h2)
	) name878 (
		_w6553_,
		_w6550_,
		_w6705_
	);
	LUT3 #(
		.INIT('h40)
	) name879 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6706_
	);
	LUT4 #(
		.INIT('h0020)
	) name880 (
		_w6555_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6707_
	);
	LUT3 #(
		.INIT('h0b)
	) name881 (
		_w6705_,
		_w6706_,
		_w6707_,
		_w6708_
	);
	LUT4 #(
		.INIT('h1555)
	) name882 (
		_w6567_,
		_w6576_,
		_w6704_,
		_w6708_,
		_w6709_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name883 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6710_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w6555_,
		_w6710_,
		_w6711_
	);
	LUT3 #(
		.INIT('h0d)
	) name885 (
		_w6559_,
		_w6550_,
		_w6573_,
		_w6712_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w6711_,
		_w6712_,
		_w6713_
	);
	LUT4 #(
		.INIT('h5655)
	) name887 (
		\u2_L12_reg[10]/NET0131 ,
		_w6709_,
		_w6701_,
		_w6713_,
		_w6714_
	);
	LUT3 #(
		.INIT('h0b)
	) name888 (
		_w6520_,
		_w6523_,
		_w6521_,
		_w6715_
	);
	LUT3 #(
		.INIT('hc8)
	) name889 (
		_w6519_,
		_w6522_,
		_w6523_,
		_w6716_
	);
	LUT4 #(
		.INIT('h0804)
	) name890 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6717_
	);
	LUT4 #(
		.INIT('h0111)
	) name891 (
		_w6518_,
		_w6717_,
		_w6715_,
		_w6716_,
		_w6718_
	);
	LUT2 #(
		.INIT('h6)
	) name892 (
		_w6522_,
		_w6523_,
		_w6719_
	);
	LUT4 #(
		.INIT('h125a)
	) name893 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6720_
	);
	LUT4 #(
		.INIT('h0110)
	) name894 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6721_
	);
	LUT3 #(
		.INIT('h0e)
	) name895 (
		_w6519_,
		_w6720_,
		_w6721_,
		_w6722_
	);
	LUT2 #(
		.INIT('h8)
	) name896 (
		_w6718_,
		_w6722_,
		_w6723_
	);
	LUT4 #(
		.INIT('h0ffe)
	) name897 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6724_
	);
	LUT2 #(
		.INIT('h2)
	) name898 (
		_w6519_,
		_w6724_,
		_w6725_
	);
	LUT4 #(
		.INIT('h0440)
	) name899 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6726_
	);
	LUT3 #(
		.INIT('hc8)
	) name900 (
		_w6519_,
		_w6520_,
		_w6523_,
		_w6727_
	);
	LUT4 #(
		.INIT('h00a8)
	) name901 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6728_
	);
	LUT4 #(
		.INIT('h0200)
	) name902 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6729_
	);
	LUT4 #(
		.INIT('h2022)
	) name903 (
		_w6518_,
		_w6729_,
		_w6727_,
		_w6728_,
		_w6730_
	);
	LUT3 #(
		.INIT('h10)
	) name904 (
		_w6726_,
		_w6725_,
		_w6730_,
		_w6731_
	);
	LUT3 #(
		.INIT('ha9)
	) name905 (
		\u2_L12_reg[12]/NET0131 ,
		_w6723_,
		_w6731_,
		_w6732_
	);
	LUT4 #(
		.INIT('hfe9b)
	) name906 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6733_
	);
	LUT4 #(
		.INIT('h4000)
	) name907 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6734_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name908 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6735_
	);
	LUT4 #(
		.INIT('h0155)
	) name909 (
		_w6621_,
		_w6623_,
		_w6733_,
		_w6735_,
		_w6736_
	);
	LUT4 #(
		.INIT('hd9ee)
	) name910 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6737_
	);
	LUT2 #(
		.INIT('h2)
	) name911 (
		_w6621_,
		_w6737_,
		_w6738_
	);
	LUT2 #(
		.INIT('h8)
	) name912 (
		_w6627_,
		_w6625_,
		_w6739_
	);
	LUT3 #(
		.INIT('h0b)
	) name913 (
		_w6617_,
		_w6622_,
		_w6623_,
		_w6740_
	);
	LUT3 #(
		.INIT('h10)
	) name914 (
		_w6738_,
		_w6739_,
		_w6740_,
		_w6741_
	);
	LUT4 #(
		.INIT('h3210)
	) name915 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6742_
	);
	LUT3 #(
		.INIT('h08)
	) name916 (
		_w6615_,
		_w6614_,
		_w6618_,
		_w6743_
	);
	LUT4 #(
		.INIT('hfad8)
	) name917 (
		_w6621_,
		_w6638_,
		_w6742_,
		_w6743_,
		_w6744_
	);
	LUT4 #(
		.INIT('h0004)
	) name918 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6745_
	);
	LUT4 #(
		.INIT('h00b0)
	) name919 (
		_w6626_,
		_w6628_,
		_w6623_,
		_w6745_,
		_w6746_
	);
	LUT3 #(
		.INIT('h20)
	) name920 (
		_w6735_,
		_w6744_,
		_w6746_,
		_w6747_
	);
	LUT4 #(
		.INIT('h999a)
	) name921 (
		\u2_L12_reg[13]/NET0131 ,
		_w6736_,
		_w6741_,
		_w6747_,
		_w6748_
	);
	LUT4 #(
		.INIT('hcc04)
	) name922 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6749_
	);
	LUT4 #(
		.INIT('h33cb)
	) name923 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6750_
	);
	LUT4 #(
		.INIT('h0100)
	) name924 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6751_
	);
	LUT4 #(
		.INIT('h3302)
	) name925 (
		_w6650_,
		_w6649_,
		_w6750_,
		_w6751_,
		_w6752_
	);
	LUT4 #(
		.INIT('h0020)
	) name926 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6650_,
		_w6753_
	);
	LUT4 #(
		.INIT('hbbf7)
	) name927 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6754_
	);
	LUT4 #(
		.INIT('h0010)
	) name928 (
		_w6652_,
		_w6654_,
		_w6650_,
		_w6653_,
		_w6755_
	);
	LUT4 #(
		.INIT('h2000)
	) name929 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6756_
	);
	LUT4 #(
		.INIT('h0100)
	) name930 (
		_w6755_,
		_w6756_,
		_w6753_,
		_w6754_,
		_w6757_
	);
	LUT2 #(
		.INIT('h4)
	) name931 (
		_w6651_,
		_w6649_,
		_w6758_
	);
	LUT4 #(
		.INIT('hccf7)
	) name932 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6759_
	);
	LUT4 #(
		.INIT('h4445)
	) name933 (
		_w6650_,
		_w6672_,
		_w6758_,
		_w6759_,
		_w6760_
	);
	LUT3 #(
		.INIT('h0b)
	) name934 (
		_w6651_,
		_w6652_,
		_w6650_,
		_w6761_
	);
	LUT3 #(
		.INIT('h40)
	) name935 (
		_w6651_,
		_w6652_,
		_w6650_,
		_w6762_
	);
	LUT4 #(
		.INIT('h00d0)
	) name936 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6763_
	);
	LUT3 #(
		.INIT('h10)
	) name937 (
		_w6762_,
		_w6761_,
		_w6763_,
		_w6764_
	);
	LUT4 #(
		.INIT('h0301)
	) name938 (
		_w6649_,
		_w6760_,
		_w6764_,
		_w6757_,
		_w6765_
	);
	LUT3 #(
		.INIT('h65)
	) name939 (
		\u2_L12_reg[15]/NET0131 ,
		_w6752_,
		_w6765_,
		_w6766_
	);
	LUT4 #(
		.INIT('hc693)
	) name940 (
		decrypt_pad,
		\u2_R12_reg[20]/NET0131 ,
		\u2_uk_K_r12_reg[44]/P0001 ,
		\u2_uk_K_r12_reg[50]/NET0131 ,
		_w6767_
	);
	LUT4 #(
		.INIT('hc693)
	) name941 (
		decrypt_pad,
		\u2_R12_reg[19]/NET0131 ,
		\u2_uk_K_r12_reg[29]/NET0131 ,
		\u2_uk_K_r12_reg[35]/NET0131 ,
		_w6768_
	);
	LUT4 #(
		.INIT('hc963)
	) name942 (
		decrypt_pad,
		\u2_R12_reg[17]/NET0131 ,
		\u2_uk_K_r12_reg[30]/NET0131 ,
		\u2_uk_K_r12_reg[52]/NET0131 ,
		_w6769_
	);
	LUT4 #(
		.INIT('hc693)
	) name943 (
		decrypt_pad,
		\u2_R12_reg[16]/NET0131 ,
		\u2_uk_K_r12_reg[2]/NET0131 ,
		\u2_uk_K_r12_reg[8]/NET0131 ,
		_w6770_
	);
	LUT4 #(
		.INIT('hc693)
	) name944 (
		decrypt_pad,
		\u2_R12_reg[21]/NET0131 ,
		\u2_uk_K_r12_reg[14]/NET0131 ,
		\u2_uk_K_r12_reg[51]/NET0131 ,
		_w6771_
	);
	LUT4 #(
		.INIT('hc693)
	) name945 (
		decrypt_pad,
		\u2_R12_reg[18]/NET0131 ,
		\u2_uk_K_r12_reg[42]/NET0131 ,
		\u2_uk_K_r12_reg[52]/NET0131 ,
		_w6772_
	);
	LUT3 #(
		.INIT('h20)
	) name946 (
		_w6772_,
		_w6770_,
		_w6771_,
		_w6773_
	);
	LUT4 #(
		.INIT('hc25f)
	) name947 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6774_
	);
	LUT2 #(
		.INIT('h2)
	) name948 (
		_w6768_,
		_w6774_,
		_w6775_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w6772_,
		_w6768_,
		_w6776_
	);
	LUT3 #(
		.INIT('h20)
	) name950 (
		_w6769_,
		_w6770_,
		_w6771_,
		_w6777_
	);
	LUT3 #(
		.INIT('hde)
	) name951 (
		_w6769_,
		_w6770_,
		_w6771_,
		_w6778_
	);
	LUT2 #(
		.INIT('h2)
	) name952 (
		_w6776_,
		_w6778_,
		_w6779_
	);
	LUT3 #(
		.INIT('hc4)
	) name953 (
		_w6769_,
		_w6772_,
		_w6768_,
		_w6780_
	);
	LUT4 #(
		.INIT('hd000)
	) name954 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6781_
	);
	LUT4 #(
		.INIT('h0020)
	) name955 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6782_
	);
	LUT2 #(
		.INIT('h2)
	) name956 (
		_w6770_,
		_w6771_,
		_w6783_
	);
	LUT4 #(
		.INIT('h0040)
	) name957 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6784_
	);
	LUT4 #(
		.INIT('hff9f)
	) name958 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6785_
	);
	LUT3 #(
		.INIT('hb0)
	) name959 (
		_w6780_,
		_w6781_,
		_w6785_,
		_w6786_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name960 (
		_w6767_,
		_w6779_,
		_w6775_,
		_w6786_,
		_w6787_
	);
	LUT3 #(
		.INIT('h80)
	) name961 (
		_w6769_,
		_w6770_,
		_w6771_,
		_w6788_
	);
	LUT4 #(
		.INIT('h2000)
	) name962 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6789_
	);
	LUT4 #(
		.INIT('h0010)
	) name963 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6790_
	);
	LUT4 #(
		.INIT('hda67)
	) name964 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6791_
	);
	LUT3 #(
		.INIT('h02)
	) name965 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6792_
	);
	LUT4 #(
		.INIT('h3df8)
	) name966 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6793_
	);
	LUT4 #(
		.INIT('h4000)
	) name967 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6794_
	);
	LUT4 #(
		.INIT('hbffd)
	) name968 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6795_
	);
	LUT4 #(
		.INIT('he400)
	) name969 (
		_w6768_,
		_w6791_,
		_w6793_,
		_w6795_,
		_w6796_
	);
	LUT4 #(
		.INIT('h0408)
	) name970 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6797_
	);
	LUT4 #(
		.INIT('hffdb)
	) name971 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6798_
	);
	LUT3 #(
		.INIT('hb1)
	) name972 (
		_w6768_,
		_w6797_,
		_w6798_,
		_w6799_
	);
	LUT3 #(
		.INIT('he0)
	) name973 (
		_w6767_,
		_w6796_,
		_w6799_,
		_w6800_
	);
	LUT3 #(
		.INIT('h65)
	) name974 (
		\u2_L12_reg[14]/NET0131 ,
		_w6787_,
		_w6800_,
		_w6801_
	);
	LUT4 #(
		.INIT('h7343)
	) name975 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6802_
	);
	LUT2 #(
		.INIT('h2)
	) name976 (
		_w6485_,
		_w6802_,
		_w6803_
	);
	LUT4 #(
		.INIT('h1001)
	) name977 (
		_w6485_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6804_
	);
	LUT4 #(
		.INIT('h8000)
	) name978 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6805_
	);
	LUT3 #(
		.INIT('h01)
	) name979 (
		_w6493_,
		_w6805_,
		_w6804_,
		_w6806_
	);
	LUT4 #(
		.INIT('h2000)
	) name980 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6807_
	);
	LUT3 #(
		.INIT('h04)
	) name981 (
		_w6485_,
		_w6487_,
		_w6489_,
		_w6808_
	);
	LUT4 #(
		.INIT('haa8a)
	) name982 (
		_w6493_,
		_w6486_,
		_w6489_,
		_w6488_,
		_w6809_
	);
	LUT3 #(
		.INIT('h10)
	) name983 (
		_w6807_,
		_w6808_,
		_w6809_,
		_w6810_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name984 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6488_,
		_w6811_
	);
	LUT3 #(
		.INIT('h31)
	) name985 (
		_w6485_,
		_w6607_,
		_w6811_,
		_w6812_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name986 (
		_w6803_,
		_w6806_,
		_w6810_,
		_w6812_,
		_w6813_
	);
	LUT4 #(
		.INIT('hefcc)
	) name987 (
		_w6485_,
		_w6486_,
		_w6490_,
		_w6510_,
		_w6814_
	);
	LUT3 #(
		.INIT('h65)
	) name988 (
		\u2_L12_reg[19]/NET0131 ,
		_w6813_,
		_w6814_,
		_w6815_
	);
	LUT4 #(
		.INIT('hafab)
	) name989 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6816_
	);
	LUT2 #(
		.INIT('h2)
	) name990 (
		_w6567_,
		_w6816_,
		_w6817_
	);
	LUT3 #(
		.INIT('h20)
	) name991 (
		_w6555_,
		_w6575_,
		_w6698_,
		_w6818_
	);
	LUT4 #(
		.INIT('h0100)
	) name992 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6819_
	);
	LUT4 #(
		.INIT('h0800)
	) name993 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6820_
	);
	LUT3 #(
		.INIT('h01)
	) name994 (
		_w6555_,
		_w6820_,
		_w6819_,
		_w6821_
	);
	LUT3 #(
		.INIT('h0b)
	) name995 (
		_w6817_,
		_w6818_,
		_w6821_,
		_w6822_
	);
	LUT3 #(
		.INIT('h02)
	) name996 (
		_w6552_,
		_w6553_,
		_w6550_,
		_w6823_
	);
	LUT4 #(
		.INIT('h2333)
	) name997 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6553_,
		_w6824_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		_w6823_,
		_w6824_,
		_w6825_
	);
	LUT3 #(
		.INIT('h01)
	) name999 (
		_w6552_,
		_w6553_,
		_w6550_,
		_w6826_
	);
	LUT3 #(
		.INIT('h02)
	) name1000 (
		_w6555_,
		_w6580_,
		_w6826_,
		_w6827_
	);
	LUT4 #(
		.INIT('h0028)
	) name1001 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6828_
	);
	LUT3 #(
		.INIT('h01)
	) name1002 (
		_w6567_,
		_w6697_,
		_w6828_,
		_w6829_
	);
	LUT4 #(
		.INIT('hdf5d)
	) name1003 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6830_
	);
	LUT4 #(
		.INIT('hef00)
	) name1004 (
		_w6551_,
		_w6552_,
		_w6550_,
		_w6567_,
		_w6831_
	);
	LUT4 #(
		.INIT('h3200)
	) name1005 (
		_w6555_,
		_w6820_,
		_w6830_,
		_w6831_,
		_w6832_
	);
	LUT4 #(
		.INIT('h001f)
	) name1006 (
		_w6825_,
		_w6827_,
		_w6829_,
		_w6832_,
		_w6833_
	);
	LUT3 #(
		.INIT('h56)
	) name1007 (
		\u2_L12_reg[1]/NET0131 ,
		_w6822_,
		_w6833_,
		_w6834_
	);
	LUT4 #(
		.INIT('hf1f0)
	) name1008 (
		_w6651_,
		_w6654_,
		_w6650_,
		_w6653_,
		_w6835_
	);
	LUT4 #(
		.INIT('hef00)
	) name1009 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6650_,
		_w6836_
	);
	LUT4 #(
		.INIT('h773f)
	) name1010 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6837_
	);
	LUT4 #(
		.INIT('h0eee)
	) name1011 (
		_w6756_,
		_w6835_,
		_w6836_,
		_w6837_,
		_w6838_
	);
	LUT4 #(
		.INIT('h0802)
	) name1012 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6839_
	);
	LUT4 #(
		.INIT('h0010)
	) name1013 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6840_
	);
	LUT3 #(
		.INIT('h02)
	) name1014 (
		_w6649_,
		_w6839_,
		_w6840_,
		_w6841_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name1015 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6842_
	);
	LUT4 #(
		.INIT('h4000)
	) name1016 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6843_
	);
	LUT4 #(
		.INIT('h0002)
	) name1017 (
		_w6652_,
		_w6654_,
		_w6650_,
		_w6653_,
		_w6844_
	);
	LUT3 #(
		.INIT('h10)
	) name1018 (
		_w6843_,
		_w6844_,
		_w6842_,
		_w6845_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name1019 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6846_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1020 (
		_w6651_,
		_w6652_,
		_w6653_,
		_w6649_,
		_w6847_
	);
	LUT4 #(
		.INIT('h0400)
	) name1021 (
		_w6651_,
		_w6654_,
		_w6650_,
		_w6653_,
		_w6848_
	);
	LUT4 #(
		.INIT('hfbf7)
	) name1022 (
		_w6651_,
		_w6654_,
		_w6650_,
		_w6653_,
		_w6849_
	);
	LUT4 #(
		.INIT('hd000)
	) name1023 (
		_w6650_,
		_w6846_,
		_w6847_,
		_w6849_,
		_w6850_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name1024 (
		_w6838_,
		_w6841_,
		_w6845_,
		_w6850_,
		_w6851_
	);
	LUT4 #(
		.INIT('h0010)
	) name1025 (
		_w6651_,
		_w6652_,
		_w6650_,
		_w6653_,
		_w6852_
	);
	LUT3 #(
		.INIT('h13)
	) name1026 (
		_w6652_,
		_w6852_,
		_w6848_,
		_w6853_
	);
	LUT3 #(
		.INIT('h65)
	) name1027 (
		\u2_L12_reg[21]/NET0131 ,
		_w6851_,
		_w6853_,
		_w6854_
	);
	LUT4 #(
		.INIT('hfdc3)
	) name1028 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6855_
	);
	LUT4 #(
		.INIT('heffb)
	) name1029 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6856_
	);
	LUT4 #(
		.INIT('h0455)
	) name1030 (
		_w6455_,
		_w6453_,
		_w6855_,
		_w6856_,
		_w6857_
	);
	LUT4 #(
		.INIT('hdf3f)
	) name1031 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6858_
	);
	LUT2 #(
		.INIT('h2)
	) name1032 (
		_w6455_,
		_w6858_,
		_w6859_
	);
	LUT3 #(
		.INIT('h07)
	) name1033 (
		_w6466_,
		_w6480_,
		_w6463_,
		_w6860_
	);
	LUT3 #(
		.INIT('h8a)
	) name1034 (
		_w6453_,
		_w6859_,
		_w6860_,
		_w6861_
	);
	LUT4 #(
		.INIT('hff47)
	) name1035 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w6862_
	);
	LUT2 #(
		.INIT('h2)
	) name1036 (
		_w6455_,
		_w6862_,
		_w6863_
	);
	LUT3 #(
		.INIT('h7e)
	) name1037 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6864_
	);
	LUT3 #(
		.INIT('h40)
	) name1038 (
		_w6455_,
		_w6454_,
		_w6458_,
		_w6865_
	);
	LUT4 #(
		.INIT('h4000)
	) name1039 (
		_w6455_,
		_w6456_,
		_w6457_,
		_w6458_,
		_w6866_
	);
	LUT3 #(
		.INIT('h10)
	) name1040 (
		_w6865_,
		_w6866_,
		_w6864_,
		_w6867_
	);
	LUT4 #(
		.INIT('hbffd)
	) name1041 (
		_w6455_,
		_w6456_,
		_w6457_,
		_w6458_,
		_w6868_
	);
	LUT3 #(
		.INIT('h31)
	) name1042 (
		_w6454_,
		_w6481_,
		_w6868_,
		_w6869_
	);
	LUT4 #(
		.INIT('hba00)
	) name1043 (
		_w6453_,
		_w6863_,
		_w6867_,
		_w6869_,
		_w6870_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name1044 (
		\u2_L12_reg[23]/NET0131 ,
		_w6861_,
		_w6857_,
		_w6870_,
		_w6871_
	);
	LUT4 #(
		.INIT('h005d)
	) name1045 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6768_,
		_w6872_
	);
	LUT3 #(
		.INIT('ha8)
	) name1046 (
		_w6769_,
		_w6773_,
		_w6872_,
		_w6873_
	);
	LUT3 #(
		.INIT('hd0)
	) name1047 (
		_w6769_,
		_w6771_,
		_w6768_,
		_w6874_
	);
	LUT4 #(
		.INIT('h3301)
	) name1048 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6768_,
		_w6875_
	);
	LUT4 #(
		.INIT('h7077)
	) name1049 (
		_w6783_,
		_w6872_,
		_w6874_,
		_w6875_,
		_w6876_
	);
	LUT3 #(
		.INIT('h45)
	) name1050 (
		_w6767_,
		_w6873_,
		_w6876_,
		_w6877_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1051 (
		_w6769_,
		_w6770_,
		_w6771_,
		_w6768_,
		_w6878_
	);
	LUT4 #(
		.INIT('h001d)
	) name1052 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6879_
	);
	LUT4 #(
		.INIT('h6e00)
	) name1053 (
		_w6769_,
		_w6770_,
		_w6771_,
		_w6768_,
		_w6880_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1054 (
		_w6792_,
		_w6878_,
		_w6879_,
		_w6880_,
		_w6881_
	);
	LUT4 #(
		.INIT('hdd7f)
	) name1055 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6882_
	);
	LUT4 #(
		.INIT('hff7b)
	) name1056 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6883_
	);
	LUT4 #(
		.INIT('hfe7b)
	) name1057 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6884_
	);
	LUT4 #(
		.INIT('h0040)
	) name1058 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6768_,
		_w6885_
	);
	LUT4 #(
		.INIT('h0301)
	) name1059 (
		_w6768_,
		_w6789_,
		_w6885_,
		_w6884_,
		_w6886_
	);
	LUT4 #(
		.INIT('h7500)
	) name1060 (
		_w6767_,
		_w6881_,
		_w6882_,
		_w6886_,
		_w6887_
	);
	LUT3 #(
		.INIT('h65)
	) name1061 (
		\u2_L12_reg[25]/NET0131 ,
		_w6877_,
		_w6887_,
		_w6888_
	);
	LUT4 #(
		.INIT('h0802)
	) name1062 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6889_
	);
	LUT3 #(
		.INIT('h02)
	) name1063 (
		_w6567_,
		_w6571_,
		_w6889_,
		_w6890_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name1064 (
		_w6551_,
		_w6555_,
		_w6552_,
		_w6553_,
		_w6891_
	);
	LUT4 #(
		.INIT('h3f2f)
	) name1065 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6892_
	);
	LUT3 #(
		.INIT('h51)
	) name1066 (
		_w6555_,
		_w6552_,
		_w6550_,
		_w6893_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1067 (
		_w6550_,
		_w6891_,
		_w6892_,
		_w6893_,
		_w6894_
	);
	LUT4 #(
		.INIT('h00fb)
	) name1068 (
		_w6551_,
		_w6552_,
		_w6550_,
		_w6567_,
		_w6895_
	);
	LUT3 #(
		.INIT('hb0)
	) name1069 (
		_w6560_,
		_w6572_,
		_w6895_,
		_w6896_
	);
	LUT4 #(
		.INIT('h153f)
	) name1070 (
		_w6563_,
		_w6890_,
		_w6894_,
		_w6896_,
		_w6897_
	);
	LUT4 #(
		.INIT('h0086)
	) name1071 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6898_
	);
	LUT4 #(
		.INIT('heafa)
	) name1072 (
		_w6551_,
		_w6552_,
		_w6553_,
		_w6550_,
		_w6899_
	);
	LUT4 #(
		.INIT('h5051)
	) name1073 (
		_w6555_,
		_w6567_,
		_w6898_,
		_w6899_,
		_w6900_
	);
	LUT3 #(
		.INIT('h08)
	) name1074 (
		_w6555_,
		_w6553_,
		_w6550_,
		_w6901_
	);
	LUT2 #(
		.INIT('h4)
	) name1075 (
		_w6565_,
		_w6901_,
		_w6902_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w6900_,
		_w6902_,
		_w6903_
	);
	LUT3 #(
		.INIT('h65)
	) name1077 (
		\u2_L12_reg[26]/NET0131 ,
		_w6897_,
		_w6903_,
		_w6904_
	);
	LUT3 #(
		.INIT('h90)
	) name1078 (
		_w6615_,
		_w6616_,
		_w6618_,
		_w6905_
	);
	LUT4 #(
		.INIT('h0040)
	) name1079 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6906_
	);
	LUT3 #(
		.INIT('h8a)
	) name1080 (
		_w6621_,
		_w6614_,
		_w6618_,
		_w6907_
	);
	LUT3 #(
		.INIT('h10)
	) name1081 (
		_w6906_,
		_w6905_,
		_w6907_,
		_w6908_
	);
	LUT4 #(
		.INIT('h5545)
	) name1082 (
		_w6621_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6909_
	);
	LUT4 #(
		.INIT('hff72)
	) name1083 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6910_
	);
	LUT4 #(
		.INIT('hbf72)
	) name1084 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6911_
	);
	LUT2 #(
		.INIT('h8)
	) name1085 (
		_w6909_,
		_w6911_,
		_w6912_
	);
	LUT4 #(
		.INIT('h0220)
	) name1086 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6913_
	);
	LUT2 #(
		.INIT('h2)
	) name1087 (
		_w6623_,
		_w6913_,
		_w6914_
	);
	LUT3 #(
		.INIT('he0)
	) name1088 (
		_w6908_,
		_w6912_,
		_w6914_,
		_w6915_
	);
	LUT4 #(
		.INIT('h32dd)
	) name1089 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6916_
	);
	LUT4 #(
		.INIT('h4e5f)
	) name1090 (
		_w6621_,
		_w6642_,
		_w6910_,
		_w6916_,
		_w6917_
	);
	LUT4 #(
		.INIT('h2010)
	) name1091 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w6918_
	);
	LUT3 #(
		.INIT('h01)
	) name1092 (
		_w6623_,
		_w6734_,
		_w6918_,
		_w6919_
	);
	LUT2 #(
		.INIT('h4)
	) name1093 (
		_w6917_,
		_w6919_,
		_w6920_
	);
	LUT3 #(
		.INIT('ha9)
	) name1094 (
		\u2_L12_reg[28]/NET0131 ,
		_w6915_,
		_w6920_,
		_w6921_
	);
	LUT2 #(
		.INIT('h1)
	) name1095 (
		_w6768_,
		_w6784_,
		_w6922_
	);
	LUT4 #(
		.INIT('h0200)
	) name1096 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6923_
	);
	LUT4 #(
		.INIT('h0400)
	) name1097 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6924_
	);
	LUT4 #(
		.INIT('hf700)
	) name1098 (
		_w6769_,
		_w6772_,
		_w6771_,
		_w6768_,
		_w6925_
	);
	LUT3 #(
		.INIT('h10)
	) name1099 (
		_w6923_,
		_w6924_,
		_w6925_,
		_w6926_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w6922_,
		_w6926_,
		_w6927_
	);
	LUT4 #(
		.INIT('h0001)
	) name1101 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6928_
	);
	LUT4 #(
		.INIT('haffe)
	) name1102 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6929_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1103 (
		_w6767_,
		_w6772_,
		_w6770_,
		_w6768_,
		_w6930_
	);
	LUT4 #(
		.INIT('h3100)
	) name1104 (
		_w6768_,
		_w6797_,
		_w6929_,
		_w6930_,
		_w6931_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1105 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6932_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		_w6878_,
		_w6932_,
		_w6933_
	);
	LUT3 #(
		.INIT('h02)
	) name1107 (
		_w6768_,
		_w6790_,
		_w6788_,
		_w6934_
	);
	LUT4 #(
		.INIT('h5551)
	) name1108 (
		_w6767_,
		_w6769_,
		_w6772_,
		_w6770_,
		_w6935_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		_w6883_,
		_w6935_,
		_w6936_
	);
	LUT4 #(
		.INIT('h0155)
	) name1110 (
		_w6931_,
		_w6933_,
		_w6934_,
		_w6936_,
		_w6937_
	);
	LUT3 #(
		.INIT('h56)
	) name1111 (
		\u2_L12_reg[8]/NET0131 ,
		_w6927_,
		_w6937_,
		_w6938_
	);
	LUT4 #(
		.INIT('hf32e)
	) name1112 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6939_
	);
	LUT2 #(
		.INIT('h1)
	) name1113 (
		_w6650_,
		_w6939_,
		_w6940_
	);
	LUT3 #(
		.INIT('h8c)
	) name1114 (
		_w6654_,
		_w6650_,
		_w6653_,
		_w6941_
	);
	LUT4 #(
		.INIT('hed6f)
	) name1115 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6653_,
		_w6942_
	);
	LUT3 #(
		.INIT('h70)
	) name1116 (
		_w6749_,
		_w6941_,
		_w6942_,
		_w6943_
	);
	LUT3 #(
		.INIT('h8a)
	) name1117 (
		_w6649_,
		_w6940_,
		_w6943_,
		_w6944_
	);
	LUT4 #(
		.INIT('hf070)
	) name1118 (
		_w6651_,
		_w6652_,
		_w6650_,
		_w6653_,
		_w6945_
	);
	LUT3 #(
		.INIT('h4b)
	) name1119 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6946_
	);
	LUT2 #(
		.INIT('h8)
	) name1120 (
		_w6945_,
		_w6946_,
		_w6947_
	);
	LUT4 #(
		.INIT('h0800)
	) name1121 (
		_w6651_,
		_w6654_,
		_w6650_,
		_w6653_,
		_w6948_
	);
	LUT3 #(
		.INIT('h01)
	) name1122 (
		_w6671_,
		_w6844_,
		_w6948_,
		_w6949_
	);
	LUT4 #(
		.INIT('h0200)
	) name1123 (
		_w6651_,
		_w6652_,
		_w6654_,
		_w6650_,
		_w6950_
	);
	LUT4 #(
		.INIT('h00ba)
	) name1124 (
		_w6650_,
		_w6667_,
		_w6670_,
		_w6950_,
		_w6951_
	);
	LUT4 #(
		.INIT('hba00)
	) name1125 (
		_w6649_,
		_w6947_,
		_w6949_,
		_w6951_,
		_w6952_
	);
	LUT3 #(
		.INIT('h65)
	) name1126 (
		\u2_L12_reg[27]/NET0131 ,
		_w6944_,
		_w6952_,
		_w6953_
	);
	LUT4 #(
		.INIT('h0800)
	) name1127 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6954_
	);
	LUT4 #(
		.INIT('hf6ad)
	) name1128 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6955_
	);
	LUT2 #(
		.INIT('h1)
	) name1129 (
		_w6519_,
		_w6955_,
		_w6956_
	);
	LUT3 #(
		.INIT('he0)
	) name1130 (
		_w6519_,
		_w6523_,
		_w6521_,
		_w6957_
	);
	LUT4 #(
		.INIT('hdfda)
	) name1131 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6958_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1132 (
		_w6519_,
		_w6544_,
		_w6957_,
		_w6958_,
		_w6959_
	);
	LUT3 #(
		.INIT('h8a)
	) name1133 (
		_w6518_,
		_w6956_,
		_w6959_,
		_w6960_
	);
	LUT4 #(
		.INIT('h5455)
	) name1134 (
		_w6519_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w6961_
	);
	LUT2 #(
		.INIT('h4)
	) name1135 (
		_w6719_,
		_w6961_,
		_w6962_
	);
	LUT3 #(
		.INIT('h9b)
	) name1136 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6963_
	);
	LUT3 #(
		.INIT('h15)
	) name1137 (
		_w6545_,
		_w6957_,
		_w6963_,
		_w6964_
	);
	LUT4 #(
		.INIT('h4050)
	) name1138 (
		_w6519_,
		_w6522_,
		_w6523_,
		_w6521_,
		_w6965_
	);
	LUT2 #(
		.INIT('h2)
	) name1139 (
		_w6518_,
		_w6519_,
		_w6966_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1140 (
		_w6539_,
		_w6542_,
		_w6965_,
		_w6966_,
		_w6967_
	);
	LUT4 #(
		.INIT('hba00)
	) name1141 (
		_w6518_,
		_w6962_,
		_w6964_,
		_w6967_,
		_w6968_
	);
	LUT3 #(
		.INIT('h65)
	) name1142 (
		\u2_L12_reg[32]/NET0131 ,
		_w6960_,
		_w6968_,
		_w6969_
	);
	LUT4 #(
		.INIT('hcff5)
	) name1143 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6970_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name1144 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6971_
	);
	LUT4 #(
		.INIT('hb100)
	) name1145 (
		_w6768_,
		_w6777_,
		_w6970_,
		_w6971_,
		_w6972_
	);
	LUT2 #(
		.INIT('h2)
	) name1146 (
		_w6767_,
		_w6972_,
		_w6973_
	);
	LUT4 #(
		.INIT('hb85b)
	) name1147 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6974_
	);
	LUT2 #(
		.INIT('h1)
	) name1148 (
		_w6767_,
		_w6974_,
		_w6975_
	);
	LUT3 #(
		.INIT('h02)
	) name1149 (
		_w6768_,
		_w6790_,
		_w6924_,
		_w6976_
	);
	LUT4 #(
		.INIT('h23f0)
	) name1150 (
		_w6769_,
		_w6772_,
		_w6770_,
		_w6771_,
		_w6977_
	);
	LUT3 #(
		.INIT('h0d)
	) name1151 (
		_w6767_,
		_w6794_,
		_w6977_,
		_w6978_
	);
	LUT3 #(
		.INIT('h01)
	) name1152 (
		_w6768_,
		_w6782_,
		_w6928_,
		_w6979_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1153 (
		_w6975_,
		_w6976_,
		_w6978_,
		_w6979_,
		_w6980_
	);
	LUT3 #(
		.INIT('h56)
	) name1154 (
		\u2_L12_reg[3]/NET0131 ,
		_w6973_,
		_w6980_,
		_w6981_
	);
	LUT4 #(
		.INIT('hc693)
	) name1155 (
		decrypt_pad,
		\u2_R12_reg[12]/NET0131 ,
		\u2_uk_K_r12_reg[13]/NET0131 ,
		\u2_uk_K_r12_reg[46]/NET0131 ,
		_w6982_
	);
	LUT4 #(
		.INIT('hc693)
	) name1156 (
		decrypt_pad,
		\u2_R12_reg[13]/NET0131 ,
		\u2_uk_K_r12_reg[26]/NET0131 ,
		\u2_uk_K_r12_reg[34]/NET0131 ,
		_w6983_
	);
	LUT4 #(
		.INIT('hc693)
	) name1157 (
		decrypt_pad,
		\u2_R12_reg[8]/NET0131 ,
		\u2_uk_K_r12_reg[17]/NET0131 ,
		\u2_uk_K_r12_reg[25]/NET0131 ,
		_w6984_
	);
	LUT2 #(
		.INIT('h6)
	) name1158 (
		_w6983_,
		_w6984_,
		_w6985_
	);
	LUT4 #(
		.INIT('hc693)
	) name1159 (
		decrypt_pad,
		\u2_R12_reg[9]/NET0131 ,
		\u2_uk_K_r12_reg[46]/NET0131 ,
		\u2_uk_K_r12_reg[54]/NET0131 ,
		_w6986_
	);
	LUT4 #(
		.INIT('hc693)
	) name1160 (
		decrypt_pad,
		\u2_R12_reg[10]/NET0131 ,
		\u2_uk_K_r12_reg[54]/NET0131 ,
		\u2_uk_K_r12_reg[5]/NET0131 ,
		_w6987_
	);
	LUT4 #(
		.INIT('h2100)
	) name1161 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w6988_
	);
	LUT3 #(
		.INIT('h08)
	) name1162 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6989_
	);
	LUT4 #(
		.INIT('hc693)
	) name1163 (
		decrypt_pad,
		\u2_R12_reg[11]/NET0131 ,
		\u2_uk_K_r12_reg[55]/NET0131 ,
		\u2_uk_K_r12_reg[6]/NET0131 ,
		_w6990_
	);
	LUT2 #(
		.INIT('h2)
	) name1164 (
		_w6987_,
		_w6990_,
		_w6991_
	);
	LUT3 #(
		.INIT('h40)
	) name1165 (
		_w6983_,
		_w6986_,
		_w6987_,
		_w6992_
	);
	LUT4 #(
		.INIT('h4000)
	) name1166 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w6993_
	);
	LUT4 #(
		.INIT('h0007)
	) name1167 (
		_w6989_,
		_w6991_,
		_w6993_,
		_w6988_,
		_w6994_
	);
	LUT2 #(
		.INIT('h8)
	) name1168 (
		_w6983_,
		_w6990_,
		_w6995_
	);
	LUT3 #(
		.INIT('h46)
	) name1169 (
		_w6983_,
		_w6984_,
		_w6990_,
		_w6996_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		_w6986_,
		_w6987_,
		_w6997_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		_w6997_,
		_w6996_,
		_w6998_
	);
	LUT3 #(
		.INIT('hed)
	) name1172 (
		_w6986_,
		_w6987_,
		_w6996_,
		_w6999_
	);
	LUT3 #(
		.INIT('h15)
	) name1173 (
		_w6982_,
		_w6994_,
		_w6999_,
		_w7000_
	);
	LUT4 #(
		.INIT('h959d)
	) name1174 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7001_
	);
	LUT4 #(
		.INIT('h0001)
	) name1175 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7002_
	);
	LUT4 #(
		.INIT('hddfe)
	) name1176 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7003_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1177 (
		_w7001_,
		_w6982_,
		_w7003_,
		_w6990_,
		_w7004_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		_w6987_,
		_w6982_,
		_w7005_
	);
	LUT3 #(
		.INIT('h04)
	) name1179 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w7006_
	);
	LUT2 #(
		.INIT('h2)
	) name1180 (
		_w6982_,
		_w6990_,
		_w7007_
	);
	LUT3 #(
		.INIT('h80)
	) name1181 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w7008_
	);
	LUT4 #(
		.INIT('h6f67)
	) name1182 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7009_
	);
	LUT4 #(
		.INIT('h7707)
	) name1183 (
		_w7005_,
		_w7006_,
		_w7007_,
		_w7009_,
		_w7010_
	);
	LUT2 #(
		.INIT('h4)
	) name1184 (
		_w7004_,
		_w7010_,
		_w7011_
	);
	LUT3 #(
		.INIT('h65)
	) name1185 (
		\u2_L12_reg[6]/NET0131 ,
		_w7000_,
		_w7011_,
		_w7012_
	);
	LUT4 #(
		.INIT('h152a)
	) name1186 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w7013_
	);
	LUT4 #(
		.INIT('h6290)
	) name1187 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w7014_
	);
	LUT2 #(
		.INIT('h4)
	) name1188 (
		_w6518_,
		_w6519_,
		_w7015_
	);
	LUT2 #(
		.INIT('h9)
	) name1189 (
		_w6518_,
		_w6519_,
		_w7016_
	);
	LUT3 #(
		.INIT('h10)
	) name1190 (
		_w6524_,
		_w7014_,
		_w7016_,
		_w7017_
	);
	LUT3 #(
		.INIT('h09)
	) name1191 (
		_w6520_,
		_w6523_,
		_w6521_,
		_w7018_
	);
	LUT3 #(
		.INIT('h48)
	) name1192 (
		_w6522_,
		_w6523_,
		_w6521_,
		_w7019_
	);
	LUT3 #(
		.INIT('h40)
	) name1193 (
		_w6522_,
		_w6520_,
		_w6521_,
		_w7020_
	);
	LUT4 #(
		.INIT('h0002)
	) name1194 (
		_w6966_,
		_w7020_,
		_w7019_,
		_w7018_,
		_w7021_
	);
	LUT4 #(
		.INIT('h8044)
	) name1195 (
		_w6522_,
		_w6520_,
		_w6523_,
		_w6521_,
		_w7022_
	);
	LUT3 #(
		.INIT('h04)
	) name1196 (
		_w7013_,
		_w7015_,
		_w7022_,
		_w7023_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1197 (
		_w6954_,
		_w7017_,
		_w7021_,
		_w7023_,
		_w7024_
	);
	LUT2 #(
		.INIT('h6)
	) name1198 (
		\u2_L12_reg[7]/NET0131 ,
		_w7024_,
		_w7025_
	);
	LUT3 #(
		.INIT('hb7)
	) name1199 (
		_w6456_,
		_w6457_,
		_w6458_,
		_w7026_
	);
	LUT2 #(
		.INIT('h2)
	) name1200 (
		_w6469_,
		_w7026_,
		_w7027_
	);
	LUT4 #(
		.INIT('h8228)
	) name1201 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w7028_
	);
	LUT3 #(
		.INIT('he6)
	) name1202 (
		_w6457_,
		_w6454_,
		_w6458_,
		_w7029_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1203 (
		_w6453_,
		_w6471_,
		_w6586_,
		_w7029_,
		_w7030_
	);
	LUT4 #(
		.INIT('hd3c3)
	) name1204 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w7031_
	);
	LUT2 #(
		.INIT('h2)
	) name1205 (
		_w6455_,
		_w7031_,
		_w7032_
	);
	LUT4 #(
		.INIT('h0141)
	) name1206 (
		_w6455_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w7033_
	);
	LUT4 #(
		.INIT('h0802)
	) name1207 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w7034_
	);
	LUT4 #(
		.INIT('h4000)
	) name1208 (
		_w6456_,
		_w6457_,
		_w6454_,
		_w6458_,
		_w7035_
	);
	LUT4 #(
		.INIT('h0001)
	) name1209 (
		_w6453_,
		_w7035_,
		_w7034_,
		_w7033_,
		_w7036_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1210 (
		_w7028_,
		_w7030_,
		_w7032_,
		_w7036_,
		_w7037_
	);
	LUT3 #(
		.INIT('h56)
	) name1211 (
		\u2_L12_reg[9]/NET0131 ,
		_w7027_,
		_w7037_,
		_w7038_
	);
	LUT4 #(
		.INIT('hf700)
	) name1212 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7039_
	);
	LUT4 #(
		.INIT('h0400)
	) name1213 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6990_,
		_w7040_
	);
	LUT4 #(
		.INIT('h006d)
	) name1214 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7041_
	);
	LUT3 #(
		.INIT('h45)
	) name1215 (
		_w7039_,
		_w7040_,
		_w7041_,
		_w7042_
	);
	LUT4 #(
		.INIT('h0100)
	) name1216 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7043_
	);
	LUT3 #(
		.INIT('h14)
	) name1217 (
		_w6983_,
		_w6984_,
		_w6987_,
		_w7044_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1218 (
		_w6990_,
		_w6993_,
		_w7043_,
		_w7044_,
		_w7045_
	);
	LUT3 #(
		.INIT('ha8)
	) name1219 (
		_w6982_,
		_w7042_,
		_w7045_,
		_w7046_
	);
	LUT3 #(
		.INIT('h40)
	) name1220 (
		_w6986_,
		_w6984_,
		_w6987_,
		_w7047_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1221 (
		_w6986_,
		_w6984_,
		_w6987_,
		_w6990_,
		_w7048_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1222 (
		_w6990_,
		_w6993_,
		_w7043_,
		_w7048_,
		_w7049_
	);
	LUT4 #(
		.INIT('h7d78)
	) name1223 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7050_
	);
	LUT3 #(
		.INIT('he0)
	) name1224 (
		_w6983_,
		_w6984_,
		_w6990_,
		_w7051_
	);
	LUT4 #(
		.INIT('h6800)
	) name1225 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6990_,
		_w7052_
	);
	LUT4 #(
		.INIT('h0504)
	) name1226 (
		_w7002_,
		_w6990_,
		_w7052_,
		_w7050_,
		_w7053_
	);
	LUT3 #(
		.INIT('h32)
	) name1227 (
		_w6982_,
		_w7049_,
		_w7053_,
		_w7054_
	);
	LUT3 #(
		.INIT('h65)
	) name1228 (
		\u2_L12_reg[16]/NET0131 ,
		_w7046_,
		_w7054_,
		_w7055_
	);
	LUT4 #(
		.INIT('h2028)
	) name1229 (
		_w6621_,
		_w6615_,
		_w6616_,
		_w6618_,
		_w7056_
	);
	LUT4 #(
		.INIT('he4ff)
	) name1230 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w7057_
	);
	LUT4 #(
		.INIT('h0032)
	) name1231 (
		_w6621_,
		_w6643_,
		_w7057_,
		_w7056_,
		_w7058_
	);
	LUT4 #(
		.INIT('h0043)
	) name1232 (
		_w6621_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w7059_
	);
	LUT4 #(
		.INIT('h6000)
	) name1233 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w7060_
	);
	LUT4 #(
		.INIT('h8000)
	) name1234 (
		_w6621_,
		_w6615_,
		_w6616_,
		_w6618_,
		_w7061_
	);
	LUT4 #(
		.INIT('h0001)
	) name1235 (
		_w6638_,
		_w7061_,
		_w7060_,
		_w7059_,
		_w7062_
	);
	LUT4 #(
		.INIT('h0040)
	) name1236 (
		_w6621_,
		_w6615_,
		_w6616_,
		_w6618_,
		_w7063_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name1237 (
		_w6615_,
		_w6616_,
		_w6614_,
		_w6618_,
		_w7064_
	);
	LUT3 #(
		.INIT('h31)
	) name1238 (
		_w6621_,
		_w7063_,
		_w7064_,
		_w7065_
	);
	LUT4 #(
		.INIT('hd800)
	) name1239 (
		_w6623_,
		_w7058_,
		_w7062_,
		_w7065_,
		_w7066_
	);
	LUT2 #(
		.INIT('h9)
	) name1240 (
		\u2_L12_reg[18]/P0001 ,
		_w7066_,
		_w7067_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		_w6987_,
		_w6990_,
		_w7068_
	);
	LUT3 #(
		.INIT('h31)
	) name1242 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w7069_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		_w7068_,
		_w7069_,
		_w7070_
	);
	LUT3 #(
		.INIT('h0e)
	) name1244 (
		_w6986_,
		_w6987_,
		_w6990_,
		_w7071_
	);
	LUT3 #(
		.INIT('hb0)
	) name1245 (
		_w6986_,
		_w6984_,
		_w6987_,
		_w7072_
	);
	LUT4 #(
		.INIT('h23af)
	) name1246 (
		_w6985_,
		_w7051_,
		_w7071_,
		_w7072_,
		_w7073_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1247 (
		_w6982_,
		_w6998_,
		_w7070_,
		_w7073_,
		_w7074_
	);
	LUT4 #(
		.INIT('hcaf1)
	) name1248 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7075_
	);
	LUT4 #(
		.INIT('h1000)
	) name1249 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7076_
	);
	LUT4 #(
		.INIT('h5504)
	) name1250 (
		_w6982_,
		_w6990_,
		_w7075_,
		_w7076_,
		_w7077_
	);
	LUT4 #(
		.INIT('h0021)
	) name1251 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7078_
	);
	LUT4 #(
		.INIT('hb59e)
	) name1252 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7079_
	);
	LUT2 #(
		.INIT('h1)
	) name1253 (
		_w6982_,
		_w6990_,
		_w7080_
	);
	LUT2 #(
		.INIT('h4)
	) name1254 (
		_w7079_,
		_w7080_,
		_w7081_
	);
	LUT3 #(
		.INIT('he7)
	) name1255 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w7082_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name1256 (
		_w6987_,
		_w6990_,
		_w7008_,
		_w7082_,
		_w7083_
	);
	LUT3 #(
		.INIT('h10)
	) name1257 (
		_w7077_,
		_w7081_,
		_w7083_,
		_w7084_
	);
	LUT3 #(
		.INIT('h65)
	) name1258 (
		\u2_L12_reg[24]/NET0131 ,
		_w7074_,
		_w7084_,
		_w7085_
	);
	LUT4 #(
		.INIT('hfae5)
	) name1259 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7086_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name1260 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7087_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name1261 (
		_w6982_,
		_w6992_,
		_w7086_,
		_w7087_,
		_w7088_
	);
	LUT2 #(
		.INIT('h2)
	) name1262 (
		_w6990_,
		_w7088_,
		_w7089_
	);
	LUT4 #(
		.INIT('h0200)
	) name1263 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7090_
	);
	LUT3 #(
		.INIT('h0e)
	) name1264 (
		_w6986_,
		_w6984_,
		_w6990_,
		_w7091_
	);
	LUT4 #(
		.INIT('h0015)
	) name1265 (
		_w7078_,
		_w7087_,
		_w7091_,
		_w7090_,
		_w7092_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		_w6982_,
		_w7092_,
		_w7093_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name1267 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w6987_,
		_w7094_
	);
	LUT2 #(
		.INIT('h2)
	) name1268 (
		_w7007_,
		_w7094_,
		_w7095_
	);
	LUT3 #(
		.INIT('h4c)
	) name1269 (
		_w6983_,
		_w6986_,
		_w6984_,
		_w7096_
	);
	LUT2 #(
		.INIT('h8)
	) name1270 (
		_w7005_,
		_w7096_,
		_w7097_
	);
	LUT4 #(
		.INIT('h0040)
	) name1271 (
		_w6983_,
		_w6986_,
		_w6987_,
		_w6990_,
		_w7098_
	);
	LUT3 #(
		.INIT('h07)
	) name1272 (
		_w6995_,
		_w7047_,
		_w7098_,
		_w7099_
	);
	LUT3 #(
		.INIT('h10)
	) name1273 (
		_w7095_,
		_w7097_,
		_w7099_,
		_w7100_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name1274 (
		\u2_L12_reg[30]/NET0131 ,
		_w7089_,
		_w7093_,
		_w7100_,
		_w7101_
	);
	LUT4 #(
		.INIT('hc693)
	) name1275 (
		decrypt_pad,
		\u2_R11_reg[26]/NET0131 ,
		\u2_uk_K_r11_reg[2]/NET0131 ,
		\u2_uk_K_r11_reg[35]/NET0131 ,
		_w7102_
	);
	LUT4 #(
		.INIT('hc963)
	) name1276 (
		decrypt_pad,
		\u2_R11_reg[24]/NET0131 ,
		\u2_uk_K_r11_reg[15]/NET0131 ,
		\u2_uk_K_r11_reg[37]/NET0131 ,
		_w7103_
	);
	LUT4 #(
		.INIT('hc693)
	) name1277 (
		decrypt_pad,
		\u2_R11_reg[29]/NET0131 ,
		\u2_uk_K_r11_reg[14]/NET0131 ,
		\u2_uk_K_r11_reg[23]/NET0131 ,
		_w7104_
	);
	LUT3 #(
		.INIT('h04)
	) name1278 (
		_w7103_,
		_w7102_,
		_w7104_,
		_w7105_
	);
	LUT4 #(
		.INIT('hc693)
	) name1279 (
		decrypt_pad,
		\u2_R11_reg[27]/NET0131 ,
		\u2_uk_K_r11_reg[35]/NET0131 ,
		\u2_uk_K_r11_reg[44]/NET0131 ,
		_w7106_
	);
	LUT4 #(
		.INIT('h5f1b)
	) name1280 (
		_w7103_,
		_w7102_,
		_w7106_,
		_w7104_,
		_w7107_
	);
	LUT4 #(
		.INIT('hc693)
	) name1281 (
		decrypt_pad,
		\u2_R11_reg[25]/NET0131 ,
		\u2_uk_K_r11_reg[45]/NET0131 ,
		\u2_uk_K_r11_reg[50]/NET0131 ,
		_w7108_
	);
	LUT3 #(
		.INIT('h07)
	) name1282 (
		_w7102_,
		_w7106_,
		_w7108_,
		_w7109_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		_w7107_,
		_w7109_,
		_w7110_
	);
	LUT2 #(
		.INIT('h6)
	) name1284 (
		_w7103_,
		_w7102_,
		_w7111_
	);
	LUT3 #(
		.INIT('hd0)
	) name1285 (
		_w7106_,
		_w7108_,
		_w7104_,
		_w7112_
	);
	LUT2 #(
		.INIT('h4)
	) name1286 (
		_w7111_,
		_w7112_,
		_w7113_
	);
	LUT3 #(
		.INIT('h72)
	) name1287 (
		_w7102_,
		_w7108_,
		_w7104_,
		_w7114_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		_w7103_,
		_w7106_,
		_w7115_
	);
	LUT4 #(
		.INIT('hc963)
	) name1289 (
		decrypt_pad,
		\u2_R11_reg[28]/NET0131 ,
		\u2_uk_K_r11_reg[0]/NET0131 ,
		\u2_uk_K_r11_reg[22]/NET0131 ,
		_w7116_
	);
	LUT3 #(
		.INIT('h0b)
	) name1290 (
		_w7114_,
		_w7115_,
		_w7116_,
		_w7117_
	);
	LUT3 #(
		.INIT('h10)
	) name1291 (
		_w7110_,
		_w7113_,
		_w7117_,
		_w7118_
	);
	LUT4 #(
		.INIT('h0200)
	) name1292 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7119_
	);
	LUT2 #(
		.INIT('h4)
	) name1293 (
		_w7103_,
		_w7104_,
		_w7120_
	);
	LUT3 #(
		.INIT('h40)
	) name1294 (
		_w7103_,
		_w7108_,
		_w7104_,
		_w7121_
	);
	LUT4 #(
		.INIT('hadff)
	) name1295 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7122_
	);
	LUT2 #(
		.INIT('h1)
	) name1296 (
		_w7106_,
		_w7122_,
		_w7123_
	);
	LUT2 #(
		.INIT('h6)
	) name1297 (
		_w7102_,
		_w7108_,
		_w7124_
	);
	LUT4 #(
		.INIT('ha080)
	) name1298 (
		_w7103_,
		_w7102_,
		_w7106_,
		_w7104_,
		_w7125_
	);
	LUT2 #(
		.INIT('h8)
	) name1299 (
		_w7124_,
		_w7125_,
		_w7126_
	);
	LUT4 #(
		.INIT('h0001)
	) name1300 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7127_
	);
	LUT4 #(
		.INIT('h0400)
	) name1301 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7128_
	);
	LUT3 #(
		.INIT('h04)
	) name1302 (
		_w7128_,
		_w7116_,
		_w7127_,
		_w7129_
	);
	LUT3 #(
		.INIT('h10)
	) name1303 (
		_w7123_,
		_w7126_,
		_w7129_,
		_w7130_
	);
	LUT4 #(
		.INIT('h0040)
	) name1304 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7131_
	);
	LUT4 #(
		.INIT('hfbbf)
	) name1305 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7132_
	);
	LUT4 #(
		.INIT('hfbb5)
	) name1306 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7133_
	);
	LUT4 #(
		.INIT('h0900)
	) name1307 (
		_w7103_,
		_w7102_,
		_w7106_,
		_w7108_,
		_w7134_
	);
	LUT4 #(
		.INIT('h0004)
	) name1308 (
		_w7102_,
		_w7106_,
		_w7108_,
		_w7104_,
		_w7135_
	);
	LUT4 #(
		.INIT('h0301)
	) name1309 (
		_w7106_,
		_w7134_,
		_w7135_,
		_w7133_,
		_w7136_
	);
	LUT4 #(
		.INIT('ha955)
	) name1310 (
		\u2_L11_reg[22]/NET0131 ,
		_w7118_,
		_w7130_,
		_w7136_,
		_w7137_
	);
	LUT4 #(
		.INIT('hc693)
	) name1311 (
		decrypt_pad,
		\u2_R11_reg[3]/NET0131 ,
		\u2_uk_K_r11_reg[13]/NET0131 ,
		\u2_uk_K_r11_reg[18]/NET0131 ,
		_w7138_
	);
	LUT4 #(
		.INIT('hc693)
	) name1312 (
		decrypt_pad,
		\u2_R11_reg[4]/NET0131 ,
		\u2_uk_K_r11_reg[48]/NET0131 ,
		\u2_uk_K_r11_reg[53]/P0001 ,
		_w7139_
	);
	LUT4 #(
		.INIT('hc963)
	) name1313 (
		decrypt_pad,
		\u2_R11_reg[2]/NET0131 ,
		\u2_uk_K_r11_reg[41]/NET0131 ,
		\u2_uk_K_r11_reg[4]/NET0131 ,
		_w7140_
	);
	LUT4 #(
		.INIT('hc693)
	) name1314 (
		decrypt_pad,
		\u2_R11_reg[5]/NET0131 ,
		\u2_uk_K_r11_reg[19]/NET0131 ,
		\u2_uk_K_r11_reg[24]/NET0131 ,
		_w7141_
	);
	LUT4 #(
		.INIT('hc963)
	) name1315 (
		decrypt_pad,
		\u2_R11_reg[1]/NET0131 ,
		\u2_uk_K_r11_reg[26]/NET0131 ,
		\u2_uk_K_r11_reg[46]/NET0131 ,
		_w7142_
	);
	LUT4 #(
		.INIT('hc693)
	) name1316 (
		decrypt_pad,
		\u2_R11_reg[32]/NET0131 ,
		\u2_uk_K_r11_reg[25]/NET0131 ,
		\u2_uk_K_r11_reg[5]/NET0131 ,
		_w7143_
	);
	LUT4 #(
		.INIT('heff4)
	) name1317 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7144_
	);
	LUT3 #(
		.INIT('h80)
	) name1318 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7145_
	);
	LUT4 #(
		.INIT('h7dbd)
	) name1319 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7146_
	);
	LUT4 #(
		.INIT('h0155)
	) name1320 (
		_w7138_,
		_w7139_,
		_w7144_,
		_w7146_,
		_w7147_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name1321 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7148_
	);
	LUT2 #(
		.INIT('h2)
	) name1322 (
		_w7138_,
		_w7148_,
		_w7149_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name1323 (
		_w7138_,
		_w7142_,
		_w7141_,
		_w7140_,
		_w7150_
	);
	LUT2 #(
		.INIT('h4)
	) name1324 (
		_w7150_,
		_w7143_,
		_w7151_
	);
	LUT2 #(
		.INIT('h2)
	) name1325 (
		_w7138_,
		_w7140_,
		_w7152_
	);
	LUT3 #(
		.INIT('hc4)
	) name1326 (
		_w7138_,
		_w7142_,
		_w7140_,
		_w7153_
	);
	LUT3 #(
		.INIT('h0e)
	) name1327 (
		_w7141_,
		_w7140_,
		_w7143_,
		_w7154_
	);
	LUT3 #(
		.INIT('hb0)
	) name1328 (
		_w7153_,
		_w7154_,
		_w7139_,
		_w7155_
	);
	LUT3 #(
		.INIT('h10)
	) name1329 (
		_w7151_,
		_w7149_,
		_w7155_,
		_w7156_
	);
	LUT4 #(
		.INIT('hd3ff)
	) name1330 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7157_
	);
	LUT2 #(
		.INIT('h2)
	) name1331 (
		_w7138_,
		_w7157_,
		_w7158_
	);
	LUT2 #(
		.INIT('h8)
	) name1332 (
		_w7138_,
		_w7140_,
		_w7159_
	);
	LUT4 #(
		.INIT('h0080)
	) name1333 (
		_w7138_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7160_
	);
	LUT4 #(
		.INIT('hff7c)
	) name1334 (
		_w7138_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7161_
	);
	LUT4 #(
		.INIT('h0400)
	) name1335 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7162_
	);
	LUT4 #(
		.INIT('h0031)
	) name1336 (
		_w7142_,
		_w7139_,
		_w7161_,
		_w7162_,
		_w7163_
	);
	LUT2 #(
		.INIT('h4)
	) name1337 (
		_w7158_,
		_w7163_,
		_w7164_
	);
	LUT4 #(
		.INIT('h0200)
	) name1338 (
		_w7138_,
		_w7142_,
		_w7140_,
		_w7143_,
		_w7165_
	);
	LUT3 #(
		.INIT('h01)
	) name1339 (
		_w7142_,
		_w7141_,
		_w7143_,
		_w7166_
	);
	LUT3 #(
		.INIT('h13)
	) name1340 (
		_w7159_,
		_w7165_,
		_w7166_,
		_w7167_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1341 (
		_w7156_,
		_w7164_,
		_w7147_,
		_w7167_,
		_w7168_
	);
	LUT2 #(
		.INIT('h9)
	) name1342 (
		\u2_L11_reg[31]/NET0131 ,
		_w7168_,
		_w7169_
	);
	LUT4 #(
		.INIT('hc963)
	) name1343 (
		decrypt_pad,
		\u2_R11_reg[23]/NET0131 ,
		\u2_uk_K_r11_reg[22]/NET0131 ,
		\u2_uk_K_r11_reg[44]/NET0131 ,
		_w7170_
	);
	LUT4 #(
		.INIT('hc693)
	) name1344 (
		decrypt_pad,
		\u2_R11_reg[22]/NET0131 ,
		\u2_uk_K_r11_reg[0]/NET0131 ,
		\u2_uk_K_r11_reg[9]/NET0131 ,
		_w7171_
	);
	LUT4 #(
		.INIT('hc963)
	) name1345 (
		decrypt_pad,
		\u2_R11_reg[20]/NET0131 ,
		\u2_uk_K_r11_reg[31]/NET0131 ,
		\u2_uk_K_r11_reg[49]/NET0131 ,
		_w7172_
	);
	LUT4 #(
		.INIT('hc963)
	) name1346 (
		decrypt_pad,
		\u2_R11_reg[21]/NET0131 ,
		\u2_uk_K_r11_reg[42]/NET0131 ,
		\u2_uk_K_r11_reg[9]/NET0131 ,
		_w7173_
	);
	LUT4 #(
		.INIT('hc693)
	) name1347 (
		decrypt_pad,
		\u2_R11_reg[25]/NET0131 ,
		\u2_uk_K_r11_reg[38]/NET0131 ,
		\u2_uk_K_r11_reg[43]/NET0131 ,
		_w7174_
	);
	LUT4 #(
		.INIT('h168a)
	) name1348 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7175_
	);
	LUT2 #(
		.INIT('h1)
	) name1349 (
		_w7170_,
		_w7175_,
		_w7176_
	);
	LUT4 #(
		.INIT('hc693)
	) name1350 (
		decrypt_pad,
		\u2_R11_reg[24]/NET0131 ,
		\u2_uk_K_r11_reg[15]/NET0131 ,
		\u2_uk_K_r11_reg[52]/NET0131 ,
		_w7177_
	);
	LUT4 #(
		.INIT('h0004)
	) name1351 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7178_
	);
	LUT3 #(
		.INIT('h80)
	) name1352 (
		_w7172_,
		_w7173_,
		_w7174_,
		_w7179_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1353 (
		_w7170_,
		_w7171_,
		_w7172_,
		_w7173_,
		_w7180_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1354 (
		_w7177_,
		_w7178_,
		_w7179_,
		_w7180_,
		_w7181_
	);
	LUT2 #(
		.INIT('h4)
	) name1355 (
		_w7176_,
		_w7181_,
		_w7182_
	);
	LUT4 #(
		.INIT('h0800)
	) name1356 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7183_
	);
	LUT4 #(
		.INIT('h0040)
	) name1357 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7184_
	);
	LUT4 #(
		.INIT('h0200)
	) name1358 (
		_w7170_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7185_
	);
	LUT3 #(
		.INIT('h01)
	) name1359 (
		_w7184_,
		_w7185_,
		_w7183_,
		_w7186_
	);
	LUT4 #(
		.INIT('h1400)
	) name1360 (
		_w7170_,
		_w7171_,
		_w7172_,
		_w7173_,
		_w7187_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		_w7170_,
		_w7171_,
		_w7188_
	);
	LUT4 #(
		.INIT('h0080)
	) name1362 (
		_w7170_,
		_w7171_,
		_w7172_,
		_w7173_,
		_w7189_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		_w7170_,
		_w7171_,
		_w7190_
	);
	LUT4 #(
		.INIT('hfded)
	) name1364 (
		_w7170_,
		_w7171_,
		_w7172_,
		_w7174_,
		_w7191_
	);
	LUT3 #(
		.INIT('h10)
	) name1365 (
		_w7187_,
		_w7189_,
		_w7191_,
		_w7192_
	);
	LUT3 #(
		.INIT('hf6)
	) name1366 (
		_w7172_,
		_w7173_,
		_w7174_,
		_w7193_
	);
	LUT4 #(
		.INIT('h0100)
	) name1367 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7194_
	);
	LUT4 #(
		.INIT('h76ef)
	) name1368 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7195_
	);
	LUT4 #(
		.INIT('hfe54)
	) name1369 (
		_w7170_,
		_w7171_,
		_w7193_,
		_w7195_,
		_w7196_
	);
	LUT4 #(
		.INIT('hea00)
	) name1370 (
		_w7177_,
		_w7186_,
		_w7192_,
		_w7196_,
		_w7197_
	);
	LUT3 #(
		.INIT('h9a)
	) name1371 (
		\u2_L11_reg[11]/NET0131 ,
		_w7182_,
		_w7197_,
		_w7198_
	);
	LUT4 #(
		.INIT('hc693)
	) name1372 (
		decrypt_pad,
		\u2_R11_reg[14]/NET0131 ,
		\u2_uk_K_r11_reg[34]/NET0131 ,
		\u2_uk_K_r11_reg[39]/NET0131 ,
		_w7199_
	);
	LUT4 #(
		.INIT('hc693)
	) name1373 (
		decrypt_pad,
		\u2_R11_reg[15]/NET0131 ,
		\u2_uk_K_r11_reg[10]/NET0131 ,
		\u2_uk_K_r11_reg[47]/NET0131 ,
		_w7200_
	);
	LUT2 #(
		.INIT('h8)
	) name1374 (
		_w7199_,
		_w7200_,
		_w7201_
	);
	LUT4 #(
		.INIT('hc963)
	) name1375 (
		decrypt_pad,
		\u2_R11_reg[13]/NET0131 ,
		\u2_uk_K_r11_reg[13]/NET0131 ,
		\u2_uk_K_r11_reg[33]/NET0131 ,
		_w7202_
	);
	LUT3 #(
		.INIT('h80)
	) name1376 (
		_w7199_,
		_w7200_,
		_w7202_,
		_w7203_
	);
	LUT4 #(
		.INIT('hc963)
	) name1377 (
		decrypt_pad,
		\u2_R11_reg[12]/NET0131 ,
		\u2_uk_K_r11_reg[19]/NET0131 ,
		\u2_uk_K_r11_reg[39]/NET0131 ,
		_w7204_
	);
	LUT4 #(
		.INIT('h0080)
	) name1378 (
		_w7199_,
		_w7200_,
		_w7202_,
		_w7204_,
		_w7205_
	);
	LUT4 #(
		.INIT('hc693)
	) name1379 (
		decrypt_pad,
		\u2_R11_reg[16]/NET0131 ,
		\u2_uk_K_r11_reg[18]/NET0131 ,
		\u2_uk_K_r11_reg[55]/NET0131 ,
		_w7206_
	);
	LUT4 #(
		.INIT('hc963)
	) name1380 (
		decrypt_pad,
		\u2_R11_reg[17]/NET0131 ,
		\u2_uk_K_r11_reg[3]/NET0131 ,
		\u2_uk_K_r11_reg[55]/NET0131 ,
		_w7207_
	);
	LUT4 #(
		.INIT('h0001)
	) name1381 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7208_
	);
	LUT2 #(
		.INIT('h2)
	) name1382 (
		_w7202_,
		_w7204_,
		_w7209_
	);
	LUT4 #(
		.INIT('h0008)
	) name1383 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7210_
	);
	LUT3 #(
		.INIT('h10)
	) name1384 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7211_
	);
	LUT4 #(
		.INIT('heff7)
	) name1385 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7212_
	);
	LUT4 #(
		.INIT('h0100)
	) name1386 (
		_w7205_,
		_w7206_,
		_w7208_,
		_w7212_,
		_w7213_
	);
	LUT4 #(
		.INIT('hcc5f)
	) name1387 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7214_
	);
	LUT3 #(
		.INIT('h01)
	) name1388 (
		_w7202_,
		_w7204_,
		_w7207_,
		_w7215_
	);
	LUT4 #(
		.INIT('h8002)
	) name1389 (
		_w7200_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7216_
	);
	LUT3 #(
		.INIT('h0e)
	) name1390 (
		_w7200_,
		_w7214_,
		_w7216_,
		_w7217_
	);
	LUT2 #(
		.INIT('h9)
	) name1391 (
		_w7202_,
		_w7204_,
		_w7218_
	);
	LUT4 #(
		.INIT('h0002)
	) name1392 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7219_
	);
	LUT4 #(
		.INIT('hebe9)
	) name1393 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7220_
	);
	LUT2 #(
		.INIT('h1)
	) name1394 (
		_w7200_,
		_w7220_,
		_w7221_
	);
	LUT2 #(
		.INIT('h4)
	) name1395 (
		_w7204_,
		_w7207_,
		_w7222_
	);
	LUT4 #(
		.INIT('h0400)
	) name1396 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7223_
	);
	LUT4 #(
		.INIT('h7bff)
	) name1397 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7224_
	);
	LUT4 #(
		.INIT('h0200)
	) name1398 (
		_w7200_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7225_
	);
	LUT4 #(
		.INIT('h0080)
	) name1399 (
		_w7200_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7226_
	);
	LUT4 #(
		.INIT('h0200)
	) name1400 (
		_w7206_,
		_w7226_,
		_w7225_,
		_w7224_,
		_w7227_
	);
	LUT4 #(
		.INIT('h7077)
	) name1401 (
		_w7213_,
		_w7217_,
		_w7221_,
		_w7227_,
		_w7228_
	);
	LUT2 #(
		.INIT('h4)
	) name1402 (
		_w7199_,
		_w7226_,
		_w7229_
	);
	LUT2 #(
		.INIT('h1)
	) name1403 (
		_w7199_,
		_w7200_,
		_w7230_
	);
	LUT3 #(
		.INIT('h10)
	) name1404 (
		_w7199_,
		_w7200_,
		_w7207_,
		_w7231_
	);
	LUT4 #(
		.INIT('h0020)
	) name1405 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7232_
	);
	LUT4 #(
		.INIT('hffde)
	) name1406 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7233_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1407 (
		_w7200_,
		_w7209_,
		_w7231_,
		_w7233_,
		_w7234_
	);
	LUT2 #(
		.INIT('h4)
	) name1408 (
		_w7229_,
		_w7234_,
		_w7235_
	);
	LUT3 #(
		.INIT('h65)
	) name1409 (
		\u2_L11_reg[20]/NET0131 ,
		_w7228_,
		_w7235_,
		_w7236_
	);
	LUT4 #(
		.INIT('hc693)
	) name1410 (
		decrypt_pad,
		\u2_R11_reg[32]/NET0131 ,
		\u2_uk_K_r11_reg[42]/NET0131 ,
		\u2_uk_K_r11_reg[51]/NET0131 ,
		_w7237_
	);
	LUT4 #(
		.INIT('hc963)
	) name1411 (
		decrypt_pad,
		\u2_R11_reg[31]/P0001 ,
		\u2_uk_K_r11_reg[14]/NET0131 ,
		\u2_uk_K_r11_reg[36]/NET0131 ,
		_w7238_
	);
	LUT4 #(
		.INIT('hc963)
	) name1412 (
		decrypt_pad,
		\u2_R11_reg[29]/NET0131 ,
		\u2_uk_K_r11_reg[1]/NET0131 ,
		\u2_uk_K_r11_reg[23]/NET0131 ,
		_w7239_
	);
	LUT4 #(
		.INIT('hc963)
	) name1413 (
		decrypt_pad,
		\u2_R11_reg[30]/NET0131 ,
		\u2_uk_K_r11_reg[2]/NET0131 ,
		\u2_uk_K_r11_reg[52]/NET0131 ,
		_w7240_
	);
	LUT4 #(
		.INIT('hc963)
	) name1414 (
		decrypt_pad,
		\u2_R11_reg[28]/NET0131 ,
		\u2_uk_K_r11_reg[29]/NET0131 ,
		\u2_uk_K_r11_reg[51]/NET0131 ,
		_w7241_
	);
	LUT3 #(
		.INIT('h01)
	) name1415 (
		_w7239_,
		_w7240_,
		_w7241_,
		_w7242_
	);
	LUT4 #(
		.INIT('hc963)
	) name1416 (
		decrypt_pad,
		\u2_R11_reg[1]/NET0131 ,
		\u2_uk_K_r11_reg[45]/NET0131 ,
		\u2_uk_K_r11_reg[8]/NET0131 ,
		_w7243_
	);
	LUT4 #(
		.INIT('h0400)
	) name1417 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7244_
	);
	LUT2 #(
		.INIT('h4)
	) name1418 (
		_w7243_,
		_w7239_,
		_w7245_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1419 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7246_
	);
	LUT4 #(
		.INIT('h0080)
	) name1420 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7247_
	);
	LUT4 #(
		.INIT('h001b)
	) name1421 (
		_w7238_,
		_w7242_,
		_w7246_,
		_w7247_,
		_w7248_
	);
	LUT2 #(
		.INIT('h2)
	) name1422 (
		_w7237_,
		_w7248_,
		_w7249_
	);
	LUT4 #(
		.INIT('hefdd)
	) name1423 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7250_
	);
	LUT2 #(
		.INIT('h4)
	) name1424 (
		_w7250_,
		_w7238_,
		_w7251_
	);
	LUT4 #(
		.INIT('h8000)
	) name1425 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7252_
	);
	LUT3 #(
		.INIT('h04)
	) name1426 (
		_w7240_,
		_w7241_,
		_w7238_,
		_w7253_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w7252_,
		_w7253_,
		_w7254_
	);
	LUT3 #(
		.INIT('h51)
	) name1428 (
		_w7243_,
		_w7240_,
		_w7241_,
		_w7255_
	);
	LUT3 #(
		.INIT('h0d)
	) name1429 (
		_w7243_,
		_w7239_,
		_w7238_,
		_w7256_
	);
	LUT3 #(
		.INIT('h45)
	) name1430 (
		_w7244_,
		_w7255_,
		_w7256_,
		_w7257_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1431 (
		_w7251_,
		_w7254_,
		_w7257_,
		_w7237_,
		_w7258_
	);
	LUT4 #(
		.INIT('hffbe)
	) name1432 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7259_
	);
	LUT4 #(
		.INIT('h0020)
	) name1433 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7260_
	);
	LUT4 #(
		.INIT('hfd9e)
	) name1434 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7261_
	);
	LUT2 #(
		.INIT('h2)
	) name1435 (
		_w7238_,
		_w7261_,
		_w7262_
	);
	LUT2 #(
		.INIT('h4)
	) name1436 (
		_w7239_,
		_w7241_,
		_w7263_
	);
	LUT3 #(
		.INIT('h20)
	) name1437 (
		_w7240_,
		_w7238_,
		_w7237_,
		_w7264_
	);
	LUT4 #(
		.INIT('h0777)
	) name1438 (
		_w7253_,
		_w7245_,
		_w7263_,
		_w7264_,
		_w7265_
	);
	LUT2 #(
		.INIT('h4)
	) name1439 (
		_w7262_,
		_w7265_,
		_w7266_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name1440 (
		\u2_L11_reg[5]/NET0131 ,
		_w7258_,
		_w7249_,
		_w7266_,
		_w7267_
	);
	LUT4 #(
		.INIT('hfb4f)
	) name1441 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7268_
	);
	LUT4 #(
		.INIT('h7dff)
	) name1442 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7269_
	);
	LUT4 #(
		.INIT('heff3)
	) name1443 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7270_
	);
	LUT4 #(
		.INIT('hc480)
	) name1444 (
		_w7200_,
		_w7269_,
		_w7270_,
		_w7268_,
		_w7271_
	);
	LUT2 #(
		.INIT('h2)
	) name1445 (
		_w7206_,
		_w7271_,
		_w7272_
	);
	LUT4 #(
		.INIT('ha6a3)
	) name1446 (
		_w7199_,
		_w7200_,
		_w7202_,
		_w7207_,
		_w7273_
	);
	LUT2 #(
		.INIT('h2)
	) name1447 (
		_w7204_,
		_w7273_,
		_w7274_
	);
	LUT4 #(
		.INIT('h0400)
	) name1448 (
		_w7199_,
		_w7200_,
		_w7204_,
		_w7207_,
		_w7275_
	);
	LUT4 #(
		.INIT('h0023)
	) name1449 (
		_w7201_,
		_w7210_,
		_w7215_,
		_w7275_,
		_w7276_
	);
	LUT3 #(
		.INIT('h45)
	) name1450 (
		_w7206_,
		_w7274_,
		_w7276_,
		_w7277_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name1451 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7278_
	);
	LUT2 #(
		.INIT('h1)
	) name1452 (
		_w7200_,
		_w7278_,
		_w7279_
	);
	LUT3 #(
		.INIT('h23)
	) name1453 (
		_w7199_,
		_w7205_,
		_w7226_,
		_w7280_
	);
	LUT2 #(
		.INIT('h4)
	) name1454 (
		_w7279_,
		_w7280_,
		_w7281_
	);
	LUT4 #(
		.INIT('h5655)
	) name1455 (
		\u2_L11_reg[10]/NET0131 ,
		_w7277_,
		_w7272_,
		_w7281_,
		_w7282_
	);
	LUT2 #(
		.INIT('h4)
	) name1456 (
		_w7106_,
		_w7128_,
		_w7283_
	);
	LUT3 #(
		.INIT('h04)
	) name1457 (
		_w7131_,
		_w7116_,
		_w7119_,
		_w7284_
	);
	LUT4 #(
		.INIT('h5f5e)
	) name1458 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7285_
	);
	LUT4 #(
		.INIT('h1008)
	) name1459 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7286_
	);
	LUT3 #(
		.INIT('h0d)
	) name1460 (
		_w7106_,
		_w7285_,
		_w7286_,
		_w7287_
	);
	LUT3 #(
		.INIT('h40)
	) name1461 (
		_w7283_,
		_w7284_,
		_w7287_,
		_w7288_
	);
	LUT4 #(
		.INIT('h0012)
	) name1462 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7289_
	);
	LUT4 #(
		.INIT('h0804)
	) name1463 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7290_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1464 (
		_w7103_,
		_w7102_,
		_w7106_,
		_w7116_,
		_w7291_
	);
	LUT2 #(
		.INIT('h4)
	) name1465 (
		_w7290_,
		_w7291_,
		_w7292_
	);
	LUT3 #(
		.INIT('h53)
	) name1466 (
		_w7102_,
		_w7106_,
		_w7108_,
		_w7293_
	);
	LUT3 #(
		.INIT('h41)
	) name1467 (
		_w7106_,
		_w7108_,
		_w7104_,
		_w7294_
	);
	LUT3 #(
		.INIT('h0d)
	) name1468 (
		_w7120_,
		_w7293_,
		_w7294_,
		_w7295_
	);
	LUT3 #(
		.INIT('h40)
	) name1469 (
		_w7289_,
		_w7292_,
		_w7295_,
		_w7296_
	);
	LUT3 #(
		.INIT('ha9)
	) name1470 (
		\u2_L11_reg[12]/NET0131 ,
		_w7288_,
		_w7296_,
		_w7297_
	);
	LUT4 #(
		.INIT('hc963)
	) name1471 (
		decrypt_pad,
		\u2_R11_reg[19]/NET0131 ,
		\u2_uk_K_r11_reg[21]/NET0131 ,
		\u2_uk_K_r11_reg[43]/NET0131 ,
		_w7298_
	);
	LUT4 #(
		.INIT('hc693)
	) name1472 (
		decrypt_pad,
		\u2_R11_reg[18]/NET0131 ,
		\u2_uk_K_r11_reg[1]/NET0131 ,
		\u2_uk_K_r11_reg[38]/NET0131 ,
		_w7299_
	);
	LUT4 #(
		.INIT('hc963)
	) name1473 (
		decrypt_pad,
		\u2_R11_reg[17]/NET0131 ,
		\u2_uk_K_r11_reg[16]/NET0131 ,
		\u2_uk_K_r11_reg[7]/NET0131 ,
		_w7300_
	);
	LUT4 #(
		.INIT('hc693)
	) name1474 (
		decrypt_pad,
		\u2_R11_reg[16]/NET0131 ,
		\u2_uk_K_r11_reg[16]/NET0131 ,
		\u2_uk_K_r11_reg[49]/NET0131 ,
		_w7301_
	);
	LUT4 #(
		.INIT('hc693)
	) name1475 (
		decrypt_pad,
		\u2_R11_reg[21]/NET0131 ,
		\u2_uk_K_r11_reg[28]/NET0131 ,
		\u2_uk_K_r11_reg[37]/NET0131 ,
		_w7302_
	);
	LUT3 #(
		.INIT('h04)
	) name1476 (
		_w7300_,
		_w7301_,
		_w7302_,
		_w7303_
	);
	LUT4 #(
		.INIT('h0010)
	) name1477 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7304_
	);
	LUT3 #(
		.INIT('h10)
	) name1478 (
		_w7300_,
		_w7301_,
		_w7302_,
		_w7305_
	);
	LUT4 #(
		.INIT('h4000)
	) name1479 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7306_
	);
	LUT4 #(
		.INIT('hbc67)
	) name1480 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7307_
	);
	LUT3 #(
		.INIT('h04)
	) name1481 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7308_
	);
	LUT4 #(
		.INIT('h5bf8)
	) name1482 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7309_
	);
	LUT4 #(
		.INIT('hdffb)
	) name1483 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7310_
	);
	LUT4 #(
		.INIT('he400)
	) name1484 (
		_w7298_,
		_w7307_,
		_w7309_,
		_w7310_,
		_w7311_
	);
	LUT4 #(
		.INIT('hc693)
	) name1485 (
		decrypt_pad,
		\u2_R11_reg[20]/NET0131 ,
		\u2_uk_K_r11_reg[31]/NET0131 ,
		\u2_uk_K_r11_reg[36]/NET0131 ,
		_w7312_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		_w7311_,
		_w7312_,
		_w7313_
	);
	LUT4 #(
		.INIT('ha43f)
	) name1487 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7314_
	);
	LUT2 #(
		.INIT('h2)
	) name1488 (
		_w7298_,
		_w7314_,
		_w7315_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		_w7298_,
		_w7299_,
		_w7316_
	);
	LUT3 #(
		.INIT('h20)
	) name1490 (
		_w7300_,
		_w7301_,
		_w7302_,
		_w7317_
	);
	LUT3 #(
		.INIT('hde)
	) name1491 (
		_w7300_,
		_w7301_,
		_w7302_,
		_w7318_
	);
	LUT2 #(
		.INIT('h2)
	) name1492 (
		_w7316_,
		_w7318_,
		_w7319_
	);
	LUT2 #(
		.INIT('h9)
	) name1493 (
		_w7299_,
		_w7300_,
		_w7320_
	);
	LUT4 #(
		.INIT('h0060)
	) name1494 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7321_
	);
	LUT4 #(
		.INIT('h7000)
	) name1495 (
		_w7298_,
		_w7299_,
		_w7301_,
		_w7302_,
		_w7322_
	);
	LUT3 #(
		.INIT('h13)
	) name1496 (
		_w7320_,
		_w7321_,
		_w7322_,
		_w7323_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1497 (
		_w7312_,
		_w7315_,
		_w7319_,
		_w7323_,
		_w7324_
	);
	LUT4 #(
		.INIT('h0208)
	) name1498 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7325_
	);
	LUT4 #(
		.INIT('hffbd)
	) name1499 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7326_
	);
	LUT3 #(
		.INIT('hb1)
	) name1500 (
		_w7298_,
		_w7325_,
		_w7326_,
		_w7327_
	);
	LUT4 #(
		.INIT('h5655)
	) name1501 (
		\u2_L11_reg[14]/NET0131 ,
		_w7313_,
		_w7324_,
		_w7327_,
		_w7328_
	);
	LUT4 #(
		.INIT('h33d9)
	) name1502 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7329_
	);
	LUT4 #(
		.INIT('h0100)
	) name1503 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7330_
	);
	LUT4 #(
		.INIT('h3302)
	) name1504 (
		_w7238_,
		_w7237_,
		_w7329_,
		_w7330_,
		_w7331_
	);
	LUT4 #(
		.INIT('h0020)
	) name1505 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7238_,
		_w7332_
	);
	LUT4 #(
		.INIT('hf3bf)
	) name1506 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7333_
	);
	LUT4 #(
		.INIT('h2000)
	) name1507 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7334_
	);
	LUT4 #(
		.INIT('h0100)
	) name1508 (
		_w7243_,
		_w7239_,
		_w7241_,
		_w7238_,
		_w7335_
	);
	LUT4 #(
		.INIT('h0100)
	) name1509 (
		_w7334_,
		_w7335_,
		_w7332_,
		_w7333_,
		_w7336_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1510 (
		_w7239_,
		_w7240_,
		_w7241_,
		_w7238_,
		_w7337_
	);
	LUT4 #(
		.INIT('h0008)
	) name1511 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7338_
	);
	LUT3 #(
		.INIT('h04)
	) name1512 (
		_w7239_,
		_w7241_,
		_w7237_,
		_w7339_
	);
	LUT4 #(
		.INIT('h0200)
	) name1513 (
		_w7259_,
		_w7338_,
		_w7339_,
		_w7337_,
		_w7340_
	);
	LUT4 #(
		.INIT('h0002)
	) name1514 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7341_
	);
	LUT3 #(
		.INIT('h02)
	) name1515 (
		_w7238_,
		_w7247_,
		_w7341_,
		_w7342_
	);
	LUT4 #(
		.INIT('hddd0)
	) name1516 (
		_w7237_,
		_w7336_,
		_w7340_,
		_w7342_,
		_w7343_
	);
	LUT3 #(
		.INIT('h65)
	) name1517 (
		\u2_L11_reg[15]/NET0131 ,
		_w7331_,
		_w7343_,
		_w7344_
	);
	LUT4 #(
		.INIT('hfb05)
	) name1518 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7345_
	);
	LUT4 #(
		.INIT('h5001)
	) name1519 (
		_w7138_,
		_w7142_,
		_w7140_,
		_w7143_,
		_w7346_
	);
	LUT4 #(
		.INIT('h0200)
	) name1520 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7347_
	);
	LUT4 #(
		.INIT('h7d7f)
	) name1521 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7348_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1522 (
		_w7138_,
		_w7345_,
		_w7346_,
		_w7348_,
		_w7349_
	);
	LUT3 #(
		.INIT('hf9)
	) name1523 (
		_w7141_,
		_w7140_,
		_w7143_,
		_w7350_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		_w7138_,
		_w7142_,
		_w7351_
	);
	LUT2 #(
		.INIT('h4)
	) name1525 (
		_w7350_,
		_w7351_,
		_w7352_
	);
	LUT2 #(
		.INIT('h6)
	) name1526 (
		_w7141_,
		_w7143_,
		_w7353_
	);
	LUT4 #(
		.INIT('hbbec)
	) name1527 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7354_
	);
	LUT3 #(
		.INIT('h80)
	) name1528 (
		_w7142_,
		_w7141_,
		_w7143_,
		_w7355_
	);
	LUT3 #(
		.INIT('h6f)
	) name1529 (
		_w7142_,
		_w7141_,
		_w7143_,
		_w7356_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name1530 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7357_
	);
	LUT4 #(
		.INIT('he400)
	) name1531 (
		_w7138_,
		_w7354_,
		_w7356_,
		_w7357_,
		_w7358_
	);
	LUT4 #(
		.INIT('h3210)
	) name1532 (
		_w7139_,
		_w7352_,
		_w7358_,
		_w7349_,
		_w7359_
	);
	LUT2 #(
		.INIT('h9)
	) name1533 (
		\u2_L11_reg[17]/NET0131 ,
		_w7359_,
		_w7360_
	);
	LUT4 #(
		.INIT('hccef)
	) name1534 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7361_
	);
	LUT2 #(
		.INIT('h2)
	) name1535 (
		_w7206_,
		_w7361_,
		_w7362_
	);
	LUT3 #(
		.INIT('h20)
	) name1536 (
		_w7200_,
		_w7210_,
		_w7269_,
		_w7363_
	);
	LUT4 #(
		.INIT('h0080)
	) name1537 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7364_
	);
	LUT3 #(
		.INIT('h01)
	) name1538 (
		_w7200_,
		_w7219_,
		_w7364_,
		_w7365_
	);
	LUT3 #(
		.INIT('h0b)
	) name1539 (
		_w7362_,
		_w7363_,
		_w7365_,
		_w7366_
	);
	LUT3 #(
		.INIT('h04)
	) name1540 (
		_w7199_,
		_w7204_,
		_w7207_,
		_w7367_
	);
	LUT4 #(
		.INIT('h4555)
	) name1541 (
		_w7200_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7368_
	);
	LUT2 #(
		.INIT('h4)
	) name1542 (
		_w7367_,
		_w7368_,
		_w7369_
	);
	LUT3 #(
		.INIT('h01)
	) name1543 (
		_w7199_,
		_w7204_,
		_w7207_,
		_w7370_
	);
	LUT3 #(
		.INIT('h02)
	) name1544 (
		_w7200_,
		_w7232_,
		_w7370_,
		_w7371_
	);
	LUT4 #(
		.INIT('h0040)
	) name1545 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7372_
	);
	LUT3 #(
		.INIT('h04)
	) name1546 (
		_w7206_,
		_w7224_,
		_w7372_,
		_w7373_
	);
	LUT4 #(
		.INIT('hb3fb)
	) name1547 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7374_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1548 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7206_,
		_w7375_
	);
	LUT4 #(
		.INIT('h3200)
	) name1549 (
		_w7200_,
		_w7364_,
		_w7374_,
		_w7375_,
		_w7376_
	);
	LUT4 #(
		.INIT('h001f)
	) name1550 (
		_w7369_,
		_w7371_,
		_w7373_,
		_w7376_,
		_w7377_
	);
	LUT3 #(
		.INIT('h56)
	) name1551 (
		\u2_L11_reg[1]/NET0131 ,
		_w7366_,
		_w7377_,
		_w7378_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1552 (
		_w7243_,
		_w7240_,
		_w7241_,
		_w7238_,
		_w7379_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1553 (
		_w7239_,
		_w7240_,
		_w7241_,
		_w7238_,
		_w7380_
	);
	LUT4 #(
		.INIT('hfd75)
	) name1554 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7381_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name1555 (
		_w7334_,
		_w7379_,
		_w7380_,
		_w7381_,
		_w7382_
	);
	LUT4 #(
		.INIT('h4010)
	) name1556 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7383_
	);
	LUT3 #(
		.INIT('h02)
	) name1557 (
		_w7237_,
		_w7341_,
		_w7383_,
		_w7384_
	);
	LUT2 #(
		.INIT('h4)
	) name1558 (
		_w7382_,
		_w7384_,
		_w7385_
	);
	LUT4 #(
		.INIT('h0008)
	) name1559 (
		_w7243_,
		_w7240_,
		_w7241_,
		_w7238_,
		_w7386_
	);
	LUT4 #(
		.INIT('h0004)
	) name1560 (
		_w7243_,
		_w7239_,
		_w7241_,
		_w7238_,
		_w7387_
	);
	LUT3 #(
		.INIT('h08)
	) name1561 (
		_w7239_,
		_w7240_,
		_w7241_,
		_w7388_
	);
	LUT4 #(
		.INIT('h0001)
	) name1562 (
		_w7237_,
		_w7386_,
		_w7387_,
		_w7388_,
		_w7389_
	);
	LUT4 #(
		.INIT('heffe)
	) name1563 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7390_
	);
	LUT4 #(
		.INIT('h8bff)
	) name1564 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7391_
	);
	LUT4 #(
		.INIT('hdfcf)
	) name1565 (
		_w7239_,
		_w7240_,
		_w7241_,
		_w7238_,
		_w7392_
	);
	LUT4 #(
		.INIT('hf351)
	) name1566 (
		_w7243_,
		_w7238_,
		_w7391_,
		_w7392_,
		_w7393_
	);
	LUT3 #(
		.INIT('h80)
	) name1567 (
		_w7389_,
		_w7390_,
		_w7393_,
		_w7394_
	);
	LUT4 #(
		.INIT('h0100)
	) name1568 (
		_w7239_,
		_w7240_,
		_w7241_,
		_w7238_,
		_w7395_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		_w7243_,
		_w7241_,
		_w7396_
	);
	LUT3 #(
		.INIT('h02)
	) name1570 (
		_w7239_,
		_w7240_,
		_w7238_,
		_w7397_
	);
	LUT3 #(
		.INIT('h15)
	) name1571 (
		_w7395_,
		_w7396_,
		_w7397_,
		_w7398_
	);
	LUT4 #(
		.INIT('ha955)
	) name1572 (
		\u2_L11_reg[21]/NET0131 ,
		_w7385_,
		_w7394_,
		_w7398_,
		_w7399_
	);
	LUT4 #(
		.INIT('hc693)
	) name1573 (
		decrypt_pad,
		\u2_R11_reg[5]/NET0131 ,
		\u2_uk_K_r11_reg[41]/NET0131 ,
		\u2_uk_K_r11_reg[46]/NET0131 ,
		_w7400_
	);
	LUT4 #(
		.INIT('hc963)
	) name1574 (
		decrypt_pad,
		\u2_R11_reg[4]/NET0131 ,
		\u2_uk_K_r11_reg[10]/NET0131 ,
		\u2_uk_K_r11_reg[5]/NET0131 ,
		_w7401_
	);
	LUT4 #(
		.INIT('hc963)
	) name1575 (
		decrypt_pad,
		\u2_R11_reg[9]/NET0131 ,
		\u2_uk_K_r11_reg[34]/NET0131 ,
		\u2_uk_K_r11_reg[54]/NET0131 ,
		_w7402_
	);
	LUT4 #(
		.INIT('hc963)
	) name1576 (
		decrypt_pad,
		\u2_R11_reg[6]/NET0131 ,
		\u2_uk_K_r11_reg[12]/NET0131 ,
		\u2_uk_K_r11_reg[32]/NET0131 ,
		_w7403_
	);
	LUT4 #(
		.INIT('hc038)
	) name1577 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7404_
	);
	LUT4 #(
		.INIT('hc693)
	) name1578 (
		decrypt_pad,
		\u2_R11_reg[7]/NET0131 ,
		\u2_uk_K_r11_reg[26]/NET0131 ,
		\u2_uk_K_r11_reg[6]/NET0131 ,
		_w7405_
	);
	LUT2 #(
		.INIT('h4)
	) name1579 (
		_w7404_,
		_w7405_,
		_w7406_
	);
	LUT4 #(
		.INIT('h0c05)
	) name1580 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7407_
	);
	LUT4 #(
		.INIT('h0080)
	) name1581 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7408_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1582 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7405_,
		_w7409_
	);
	LUT3 #(
		.INIT('h10)
	) name1583 (
		_w7407_,
		_w7408_,
		_w7409_,
		_w7410_
	);
	LUT3 #(
		.INIT('h40)
	) name1584 (
		_w7400_,
		_w7401_,
		_w7402_,
		_w7411_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1585 (
		_w7400_,
		_w7401_,
		_w7402_,
		_w7405_,
		_w7412_
	);
	LUT2 #(
		.INIT('h4)
	) name1586 (
		_w7403_,
		_w7401_,
		_w7413_
	);
	LUT4 #(
		.INIT('h0200)
	) name1587 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7414_
	);
	LUT4 #(
		.INIT('hc693)
	) name1588 (
		decrypt_pad,
		\u2_R11_reg[8]/NET0131 ,
		\u2_uk_K_r11_reg[17]/NET0131 ,
		\u2_uk_K_r11_reg[54]/NET0131 ,
		_w7415_
	);
	LUT4 #(
		.INIT('h4500)
	) name1589 (
		_w7414_,
		_w7412_,
		_w7413_,
		_w7415_,
		_w7416_
	);
	LUT3 #(
		.INIT('he0)
	) name1590 (
		_w7406_,
		_w7410_,
		_w7416_,
		_w7417_
	);
	LUT2 #(
		.INIT('h2)
	) name1591 (
		_w7405_,
		_w7407_,
		_w7418_
	);
	LUT4 #(
		.INIT('h3c2f)
	) name1592 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7419_
	);
	LUT3 #(
		.INIT('h40)
	) name1593 (
		_w7408_,
		_w7409_,
		_w7419_,
		_w7420_
	);
	LUT4 #(
		.INIT('h2002)
	) name1594 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7421_
	);
	LUT2 #(
		.INIT('h1)
	) name1595 (
		_w7408_,
		_w7415_,
		_w7422_
	);
	LUT3 #(
		.INIT('h01)
	) name1596 (
		_w7408_,
		_w7415_,
		_w7421_,
		_w7423_
	);
	LUT3 #(
		.INIT('he0)
	) name1597 (
		_w7418_,
		_w7420_,
		_w7423_,
		_w7424_
	);
	LUT3 #(
		.INIT('ha9)
	) name1598 (
		\u2_L11_reg[28]/NET0131 ,
		_w7417_,
		_w7424_,
		_w7425_
	);
	LUT4 #(
		.INIT('h3fd2)
	) name1599 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7426_
	);
	LUT4 #(
		.INIT('h0200)
	) name1600 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7427_
	);
	LUT4 #(
		.INIT('h5504)
	) name1601 (
		_w7177_,
		_w7170_,
		_w7426_,
		_w7427_,
		_w7428_
	);
	LUT4 #(
		.INIT('hcf6f)
	) name1602 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7429_
	);
	LUT2 #(
		.INIT('h2)
	) name1603 (
		_w7170_,
		_w7429_,
		_w7430_
	);
	LUT3 #(
		.INIT('h28)
	) name1604 (
		_w7171_,
		_w7172_,
		_w7174_,
		_w7431_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name1605 (
		_w7170_,
		_w7171_,
		_w7173_,
		_w7174_,
		_w7432_
	);
	LUT4 #(
		.INIT('h5410)
	) name1606 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7433_
	);
	LUT3 #(
		.INIT('h01)
	) name1607 (
		_w7432_,
		_w7433_,
		_w7431_,
		_w7434_
	);
	LUT4 #(
		.INIT('hab6f)
	) name1608 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7435_
	);
	LUT2 #(
		.INIT('h1)
	) name1609 (
		_w7177_,
		_w7170_,
		_w7436_
	);
	LUT4 #(
		.INIT('h2000)
	) name1610 (
		_w7170_,
		_w7171_,
		_w7173_,
		_w7174_,
		_w7437_
	);
	LUT4 #(
		.INIT('h1011)
	) name1611 (
		_w7178_,
		_w7437_,
		_w7435_,
		_w7436_,
		_w7438_
	);
	LUT4 #(
		.INIT('h5700)
	) name1612 (
		_w7177_,
		_w7430_,
		_w7434_,
		_w7438_,
		_w7439_
	);
	LUT3 #(
		.INIT('h9a)
	) name1613 (
		\u2_L11_reg[29]/NET0131 ,
		_w7428_,
		_w7439_,
		_w7440_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name1614 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7441_
	);
	LUT4 #(
		.INIT('h7f7c)
	) name1615 (
		_w7403_,
		_w7405_,
		_w7411_,
		_w7441_,
		_w7442_
	);
	LUT4 #(
		.INIT('h0144)
	) name1616 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7443_
	);
	LUT4 #(
		.INIT('h0800)
	) name1617 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7444_
	);
	LUT4 #(
		.INIT('h0010)
	) name1618 (
		_w7403_,
		_w7400_,
		_w7402_,
		_w7405_,
		_w7445_
	);
	LUT3 #(
		.INIT('h01)
	) name1619 (
		_w7443_,
		_w7444_,
		_w7445_,
		_w7446_
	);
	LUT3 #(
		.INIT('h15)
	) name1620 (
		_w7415_,
		_w7442_,
		_w7446_,
		_w7447_
	);
	LUT3 #(
		.INIT('h01)
	) name1621 (
		_w7403_,
		_w7400_,
		_w7402_,
		_w7448_
	);
	LUT4 #(
		.INIT('h0010)
	) name1622 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7449_
	);
	LUT4 #(
		.INIT('h9fe4)
	) name1623 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7450_
	);
	LUT4 #(
		.INIT('h0900)
	) name1624 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7451_
	);
	LUT4 #(
		.INIT('h0501)
	) name1625 (
		_w7405_,
		_w7415_,
		_w7451_,
		_w7450_,
		_w7452_
	);
	LUT3 #(
		.INIT('h2a)
	) name1626 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7453_
	);
	LUT4 #(
		.INIT('hae00)
	) name1627 (
		_w7400_,
		_w7401_,
		_w7402_,
		_w7415_,
		_w7454_
	);
	LUT4 #(
		.INIT('h0002)
	) name1628 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7455_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1629 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7405_,
		_w7456_
	);
	LUT4 #(
		.INIT('h4500)
	) name1630 (
		_w7455_,
		_w7453_,
		_w7454_,
		_w7456_,
		_w7457_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w7452_,
		_w7457_,
		_w7458_
	);
	LUT3 #(
		.INIT('h56)
	) name1632 (
		\u2_L11_reg[2]/NET0131 ,
		_w7447_,
		_w7458_,
		_w7459_
	);
	LUT4 #(
		.INIT('hf13f)
	) name1633 (
		_w7200_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7460_
	);
	LUT2 #(
		.INIT('h2)
	) name1634 (
		_w7199_,
		_w7460_,
		_w7461_
	);
	LUT4 #(
		.INIT('h5eff)
	) name1635 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7462_
	);
	LUT4 #(
		.INIT('h0004)
	) name1636 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7463_
	);
	LUT4 #(
		.INIT('h0702)
	) name1637 (
		_w7200_,
		_w7215_,
		_w7463_,
		_w7462_,
		_w7464_
	);
	LUT3 #(
		.INIT('h8a)
	) name1638 (
		_w7206_,
		_w7461_,
		_w7464_,
		_w7465_
	);
	LUT2 #(
		.INIT('h1)
	) name1639 (
		_w7211_,
		_w7226_,
		_w7466_
	);
	LUT3 #(
		.INIT('h0d)
	) name1640 (
		_w7203_,
		_w7222_,
		_w7223_,
		_w7467_
	);
	LUT3 #(
		.INIT('h15)
	) name1641 (
		_w7206_,
		_w7466_,
		_w7467_,
		_w7468_
	);
	LUT3 #(
		.INIT('h79)
	) name1642 (
		_w7202_,
		_w7204_,
		_w7207_,
		_w7469_
	);
	LUT2 #(
		.INIT('h2)
	) name1643 (
		_w7230_,
		_w7469_,
		_w7470_
	);
	LUT3 #(
		.INIT('h40)
	) name1644 (
		_w7199_,
		_w7200_,
		_w7207_,
		_w7471_
	);
	LUT4 #(
		.INIT('hfdcc)
	) name1645 (
		_w7199_,
		_w7202_,
		_w7204_,
		_w7207_,
		_w7472_
	);
	LUT2 #(
		.INIT('h1)
	) name1646 (
		_w7200_,
		_w7206_,
		_w7473_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1647 (
		_w7218_,
		_w7471_,
		_w7472_,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h4)
	) name1648 (
		_w7470_,
		_w7474_,
		_w7475_
	);
	LUT4 #(
		.INIT('h5655)
	) name1649 (
		\u2_L11_reg[26]/NET0131 ,
		_w7465_,
		_w7468_,
		_w7475_,
		_w7476_
	);
	LUT4 #(
		.INIT('h3ce4)
	) name1650 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7477_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name1651 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7478_
	);
	LUT4 #(
		.INIT('hbb7f)
	) name1652 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7479_
	);
	LUT4 #(
		.INIT('he400)
	) name1653 (
		_w7298_,
		_w7478_,
		_w7477_,
		_w7479_,
		_w7480_
	);
	LUT2 #(
		.INIT('h2)
	) name1654 (
		_w7312_,
		_w7480_,
		_w7481_
	);
	LUT3 #(
		.INIT('ha2)
	) name1655 (
		_w7298_,
		_w7300_,
		_w7302_,
		_w7482_
	);
	LUT4 #(
		.INIT('h2223)
	) name1656 (
		_w7298_,
		_w7299_,
		_w7300_,
		_w7301_,
		_w7483_
	);
	LUT2 #(
		.INIT('h4)
	) name1657 (
		_w7482_,
		_w7483_,
		_w7484_
	);
	LUT4 #(
		.INIT('h0010)
	) name1658 (
		_w7298_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7485_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		_w7298_,
		_w7302_,
		_w7486_
	);
	LUT3 #(
		.INIT('h08)
	) name1660 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7487_
	);
	LUT3 #(
		.INIT('h45)
	) name1661 (
		_w7485_,
		_w7486_,
		_w7487_,
		_w7488_
	);
	LUT4 #(
		.INIT('hff7d)
	) name1662 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7489_
	);
	LUT4 #(
		.INIT('hfe7d)
	) name1663 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7490_
	);
	LUT4 #(
		.INIT('h0400)
	) name1664 (
		_w7298_,
		_w7299_,
		_w7300_,
		_w7301_,
		_w7491_
	);
	LUT4 #(
		.INIT('h0031)
	) name1665 (
		_w7298_,
		_w7306_,
		_w7490_,
		_w7491_,
		_w7492_
	);
	LUT4 #(
		.INIT('hba00)
	) name1666 (
		_w7312_,
		_w7484_,
		_w7488_,
		_w7492_,
		_w7493_
	);
	LUT3 #(
		.INIT('h65)
	) name1667 (
		\u2_L11_reg[25]/NET0131 ,
		_w7481_,
		_w7493_,
		_w7494_
	);
	LUT4 #(
		.INIT('he63f)
	) name1668 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7495_
	);
	LUT2 #(
		.INIT('h2)
	) name1669 (
		_w7170_,
		_w7495_,
		_w7496_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name1670 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7497_
	);
	LUT4 #(
		.INIT('h1000)
	) name1671 (
		_w7170_,
		_w7171_,
		_w7172_,
		_w7174_,
		_w7498_
	);
	LUT4 #(
		.INIT('h0032)
	) name1672 (
		_w7170_,
		_w7178_,
		_w7497_,
		_w7498_,
		_w7499_
	);
	LUT3 #(
		.INIT('h45)
	) name1673 (
		_w7177_,
		_w7496_,
		_w7499_,
		_w7500_
	);
	LUT4 #(
		.INIT('h77cf)
	) name1674 (
		_w7170_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7501_
	);
	LUT2 #(
		.INIT('h1)
	) name1675 (
		_w7171_,
		_w7501_,
		_w7502_
	);
	LUT4 #(
		.INIT('heeae)
	) name1676 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7503_
	);
	LUT3 #(
		.INIT('h80)
	) name1677 (
		_w7171_,
		_w7173_,
		_w7174_,
		_w7504_
	);
	LUT3 #(
		.INIT('h0e)
	) name1678 (
		_w7170_,
		_w7503_,
		_w7504_,
		_w7505_
	);
	LUT3 #(
		.INIT('hb6)
	) name1679 (
		_w7172_,
		_w7173_,
		_w7174_,
		_w7506_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name1680 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7507_
	);
	LUT4 #(
		.INIT('h4445)
	) name1681 (
		_w7170_,
		_w7171_,
		_w7172_,
		_w7174_,
		_w7508_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1682 (
		_w7188_,
		_w7506_,
		_w7507_,
		_w7508_,
		_w7509_
	);
	LUT4 #(
		.INIT('h7500)
	) name1683 (
		_w7177_,
		_w7502_,
		_w7505_,
		_w7509_,
		_w7510_
	);
	LUT3 #(
		.INIT('h65)
	) name1684 (
		\u2_L11_reg[4]/NET0131 ,
		_w7500_,
		_w7510_,
		_w7511_
	);
	LUT3 #(
		.INIT('h02)
	) name1685 (
		_w7403_,
		_w7400_,
		_w7402_,
		_w7512_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1686 (
		_w7403_,
		_w7401_,
		_w7402_,
		_w7405_,
		_w7513_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name1687 (
		_w7412_,
		_w7448_,
		_w7512_,
		_w7513_,
		_w7514_
	);
	LUT4 #(
		.INIT('h0004)
	) name1688 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7515_
	);
	LUT4 #(
		.INIT('h0002)
	) name1689 (
		_w7415_,
		_w7444_,
		_w7445_,
		_w7515_,
		_w7516_
	);
	LUT4 #(
		.INIT('h0600)
	) name1690 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7517_
	);
	LUT3 #(
		.INIT('h02)
	) name1691 (
		_w7400_,
		_w7401_,
		_w7402_,
		_w7518_
	);
	LUT2 #(
		.INIT('h1)
	) name1692 (
		_w7405_,
		_w7415_,
		_w7519_
	);
	LUT4 #(
		.INIT('h0100)
	) name1693 (
		_w7449_,
		_w7518_,
		_w7517_,
		_w7519_,
		_w7520_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name1694 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7521_
	);
	LUT4 #(
		.INIT('hf400)
	) name1695 (
		_w7514_,
		_w7516_,
		_w7520_,
		_w7521_,
		_w7522_
	);
	LUT4 #(
		.INIT('h1141)
	) name1696 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7523_
	);
	LUT4 #(
		.INIT('ha022)
	) name1697 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7524_
	);
	LUT4 #(
		.INIT('h0400)
	) name1698 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7525_
	);
	LUT2 #(
		.INIT('h2)
	) name1699 (
		_w7405_,
		_w7415_,
		_w7526_
	);
	LUT4 #(
		.INIT('h0100)
	) name1700 (
		_w7524_,
		_w7525_,
		_w7523_,
		_w7526_,
		_w7527_
	);
	LUT3 #(
		.INIT('h56)
	) name1701 (
		\u2_L11_reg[13]/NET0131 ,
		_w7522_,
		_w7527_,
		_w7528_
	);
	LUT3 #(
		.INIT('hd7)
	) name1702 (
		_w7172_,
		_w7173_,
		_w7174_,
		_w7529_
	);
	LUT2 #(
		.INIT('h2)
	) name1703 (
		_w7190_,
		_w7529_,
		_w7530_
	);
	LUT3 #(
		.INIT('h04)
	) name1704 (
		_w7170_,
		_w7172_,
		_w7173_,
		_w7531_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1705 (
		_w7177_,
		_w7171_,
		_w7173_,
		_w7174_,
		_w7532_
	);
	LUT3 #(
		.INIT('h10)
	) name1706 (
		_w7194_,
		_w7531_,
		_w7532_,
		_w7533_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name1707 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7534_
	);
	LUT4 #(
		.INIT('h2002)
	) name1708 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7535_
	);
	LUT3 #(
		.INIT('h0d)
	) name1709 (
		_w7170_,
		_w7534_,
		_w7535_,
		_w7536_
	);
	LUT4 #(
		.INIT('h4554)
	) name1710 (
		_w7170_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7537_
	);
	LUT3 #(
		.INIT('h8c)
	) name1711 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7538_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1712 (
		_w7170_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7539_
	);
	LUT4 #(
		.INIT('h3233)
	) name1713 (
		_w7194_,
		_w7537_,
		_w7538_,
		_w7539_,
		_w7540_
	);
	LUT4 #(
		.INIT('h8000)
	) name1714 (
		_w7171_,
		_w7172_,
		_w7173_,
		_w7174_,
		_w7541_
	);
	LUT2 #(
		.INIT('h1)
	) name1715 (
		_w7177_,
		_w7541_,
		_w7542_
	);
	LUT4 #(
		.INIT('h7077)
	) name1716 (
		_w7533_,
		_w7536_,
		_w7540_,
		_w7542_,
		_w7543_
	);
	LUT3 #(
		.INIT('h56)
	) name1717 (
		\u2_L11_reg[19]/NET0131 ,
		_w7530_,
		_w7543_,
		_w7544_
	);
	LUT4 #(
		.INIT('h8088)
	) name1718 (
		_w7138_,
		_w7142_,
		_w7140_,
		_w7143_,
		_w7545_
	);
	LUT2 #(
		.INIT('h8)
	) name1719 (
		_w7353_,
		_w7545_,
		_w7546_
	);
	LUT4 #(
		.INIT('h020a)
	) name1720 (
		_w7139_,
		_w7159_,
		_w7162_,
		_w7166_,
		_w7547_
	);
	LUT4 #(
		.INIT('habbb)
	) name1721 (
		_w7138_,
		_w7142_,
		_w7141_,
		_w7140_,
		_w7548_
	);
	LUT2 #(
		.INIT('h2)
	) name1722 (
		_w7143_,
		_w7548_,
		_w7549_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1723 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7139_,
		_w7550_
	);
	LUT4 #(
		.INIT('h0008)
	) name1724 (
		_w7138_,
		_w7142_,
		_w7141_,
		_w7143_,
		_w7551_
	);
	LUT4 #(
		.INIT('h0100)
	) name1725 (
		_w7160_,
		_w7145_,
		_w7551_,
		_w7550_,
		_w7552_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1726 (
		_w7546_,
		_w7547_,
		_w7549_,
		_w7552_,
		_w7553_
	);
	LUT4 #(
		.INIT('hef99)
	) name1727 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7554_
	);
	LUT4 #(
		.INIT('hfdfb)
	) name1728 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7555_
	);
	LUT4 #(
		.INIT('h0455)
	) name1729 (
		_w7138_,
		_w7139_,
		_w7554_,
		_w7555_,
		_w7556_
	);
	LUT3 #(
		.INIT('had)
	) name1730 (
		_w7142_,
		_w7141_,
		_w7143_,
		_w7557_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name1731 (
		_w7138_,
		_w7140_,
		_w7355_,
		_w7557_,
		_w7558_
	);
	LUT2 #(
		.INIT('h4)
	) name1732 (
		_w7556_,
		_w7558_,
		_w7559_
	);
	LUT3 #(
		.INIT('h9a)
	) name1733 (
		\u2_L11_reg[23]/NET0131 ,
		_w7553_,
		_w7559_,
		_w7560_
	);
	LUT4 #(
		.INIT('h8804)
	) name1734 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7561_
	);
	LUT3 #(
		.INIT('hb7)
	) name1735 (
		_w7243_,
		_w7239_,
		_w7241_,
		_w7562_
	);
	LUT4 #(
		.INIT('he4f5)
	) name1736 (
		_w7238_,
		_w7242_,
		_w7561_,
		_w7562_,
		_w7563_
	);
	LUT4 #(
		.INIT('hed7d)
	) name1737 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7564_
	);
	LUT3 #(
		.INIT('h8a)
	) name1738 (
		_w7237_,
		_w7563_,
		_w7564_,
		_w7565_
	);
	LUT4 #(
		.INIT('hfb00)
	) name1739 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7238_,
		_w7566_
	);
	LUT4 #(
		.INIT('h5d1d)
	) name1740 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7567_
	);
	LUT2 #(
		.INIT('h8)
	) name1741 (
		_w7566_,
		_w7567_,
		_w7568_
	);
	LUT4 #(
		.INIT('h0080)
	) name1742 (
		_w7243_,
		_w7240_,
		_w7241_,
		_w7238_,
		_w7569_
	);
	LUT3 #(
		.INIT('h01)
	) name1743 (
		_w7260_,
		_w7387_,
		_w7569_,
		_w7570_
	);
	LUT3 #(
		.INIT('h45)
	) name1744 (
		_w7237_,
		_w7568_,
		_w7570_,
		_w7571_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name1745 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7241_,
		_w7572_
	);
	LUT2 #(
		.INIT('h1)
	) name1746 (
		_w7238_,
		_w7572_,
		_w7573_
	);
	LUT4 #(
		.INIT('h1000)
	) name1747 (
		_w7243_,
		_w7239_,
		_w7240_,
		_w7238_,
		_w7574_
	);
	LUT3 #(
		.INIT('h07)
	) name1748 (
		_w7253_,
		_w7245_,
		_w7574_,
		_w7575_
	);
	LUT2 #(
		.INIT('h4)
	) name1749 (
		_w7573_,
		_w7575_,
		_w7576_
	);
	LUT4 #(
		.INIT('h5655)
	) name1750 (
		\u2_L11_reg[27]/NET0131 ,
		_w7571_,
		_w7565_,
		_w7576_,
		_w7577_
	);
	LUT4 #(
		.INIT('hf070)
	) name1751 (
		_w7103_,
		_w7102_,
		_w7106_,
		_w7104_,
		_w7578_
	);
	LUT4 #(
		.INIT('hcffa)
	) name1752 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7579_
	);
	LUT2 #(
		.INIT('h8)
	) name1753 (
		_w7578_,
		_w7579_,
		_w7580_
	);
	LUT4 #(
		.INIT('h0102)
	) name1754 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7581_
	);
	LUT4 #(
		.INIT('h0800)
	) name1755 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7582_
	);
	LUT4 #(
		.INIT('h3323)
	) name1756 (
		_w7103_,
		_w7106_,
		_w7108_,
		_w7104_,
		_w7583_
	);
	LUT3 #(
		.INIT('h10)
	) name1757 (
		_w7581_,
		_w7582_,
		_w7583_,
		_w7584_
	);
	LUT4 #(
		.INIT('h0080)
	) name1758 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7585_
	);
	LUT2 #(
		.INIT('h2)
	) name1759 (
		_w7116_,
		_w7585_,
		_w7586_
	);
	LUT3 #(
		.INIT('he0)
	) name1760 (
		_w7580_,
		_w7584_,
		_w7586_,
		_w7587_
	);
	LUT3 #(
		.INIT('h2a)
	) name1761 (
		_w7103_,
		_w7108_,
		_w7104_,
		_w7588_
	);
	LUT3 #(
		.INIT('hc4)
	) name1762 (
		_w7102_,
		_w7106_,
		_w7104_,
		_w7589_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		_w7588_,
		_w7589_,
		_w7590_
	);
	LUT4 #(
		.INIT('h8000)
	) name1764 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7591_
	);
	LUT4 #(
		.INIT('h0020)
	) name1765 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7592_
	);
	LUT3 #(
		.INIT('h01)
	) name1766 (
		_w7116_,
		_w7592_,
		_w7591_,
		_w7593_
	);
	LUT3 #(
		.INIT('h02)
	) name1767 (
		_w7103_,
		_w7102_,
		_w7104_,
		_w7594_
	);
	LUT3 #(
		.INIT('ha2)
	) name1768 (
		_w7132_,
		_w7294_,
		_w7594_,
		_w7595_
	);
	LUT3 #(
		.INIT('h40)
	) name1769 (
		_w7590_,
		_w7593_,
		_w7595_,
		_w7596_
	);
	LUT4 #(
		.INIT('h3020)
	) name1770 (
		_w7102_,
		_w7106_,
		_w7108_,
		_w7104_,
		_w7597_
	);
	LUT4 #(
		.INIT('h153f)
	) name1771 (
		_w7111_,
		_w7106_,
		_w7128_,
		_w7597_,
		_w7598_
	);
	LUT4 #(
		.INIT('ha955)
	) name1772 (
		\u2_L11_reg[32]/NET0131 ,
		_w7587_,
		_w7596_,
		_w7598_,
		_w7599_
	);
	LUT4 #(
		.INIT('hc693)
	) name1773 (
		decrypt_pad,
		\u2_R11_reg[12]/NET0131 ,
		\u2_uk_K_r11_reg[27]/NET0131 ,
		\u2_uk_K_r11_reg[32]/NET0131 ,
		_w7600_
	);
	LUT4 #(
		.INIT('hc963)
	) name1774 (
		decrypt_pad,
		\u2_R11_reg[13]/NET0131 ,
		\u2_uk_K_r11_reg[20]/NET0131 ,
		\u2_uk_K_r11_reg[40]/NET0131 ,
		_w7601_
	);
	LUT4 #(
		.INIT('hc963)
	) name1775 (
		decrypt_pad,
		\u2_R11_reg[8]/NET0131 ,
		\u2_uk_K_r11_reg[11]/NET0131 ,
		\u2_uk_K_r11_reg[6]/NET0131 ,
		_w7602_
	);
	LUT2 #(
		.INIT('h6)
	) name1776 (
		_w7601_,
		_w7602_,
		_w7603_
	);
	LUT4 #(
		.INIT('hc693)
	) name1777 (
		decrypt_pad,
		\u2_R11_reg[9]/NET0131 ,
		\u2_uk_K_r11_reg[3]/NET0131 ,
		\u2_uk_K_r11_reg[40]/NET0131 ,
		_w7604_
	);
	LUT4 #(
		.INIT('hc693)
	) name1778 (
		decrypt_pad,
		\u2_R11_reg[10]/NET0131 ,
		\u2_uk_K_r11_reg[11]/NET0131 ,
		\u2_uk_K_r11_reg[48]/NET0131 ,
		_w7605_
	);
	LUT4 #(
		.INIT('h2100)
	) name1779 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7606_
	);
	LUT3 #(
		.INIT('h08)
	) name1780 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7607_
	);
	LUT4 #(
		.INIT('hc693)
	) name1781 (
		decrypt_pad,
		\u2_R11_reg[11]/NET0131 ,
		\u2_uk_K_r11_reg[12]/NET0131 ,
		\u2_uk_K_r11_reg[17]/NET0131 ,
		_w7608_
	);
	LUT2 #(
		.INIT('h2)
	) name1782 (
		_w7605_,
		_w7608_,
		_w7609_
	);
	LUT3 #(
		.INIT('h40)
	) name1783 (
		_w7601_,
		_w7604_,
		_w7605_,
		_w7610_
	);
	LUT4 #(
		.INIT('h4000)
	) name1784 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7611_
	);
	LUT4 #(
		.INIT('h0007)
	) name1785 (
		_w7607_,
		_w7609_,
		_w7611_,
		_w7606_,
		_w7612_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		_w7601_,
		_w7608_,
		_w7613_
	);
	LUT3 #(
		.INIT('h46)
	) name1787 (
		_w7601_,
		_w7602_,
		_w7608_,
		_w7614_
	);
	LUT2 #(
		.INIT('h1)
	) name1788 (
		_w7604_,
		_w7605_,
		_w7615_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		_w7615_,
		_w7614_,
		_w7616_
	);
	LUT3 #(
		.INIT('hed)
	) name1790 (
		_w7604_,
		_w7605_,
		_w7614_,
		_w7617_
	);
	LUT3 #(
		.INIT('h15)
	) name1791 (
		_w7600_,
		_w7612_,
		_w7617_,
		_w7618_
	);
	LUT4 #(
		.INIT('h959d)
	) name1792 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7619_
	);
	LUT4 #(
		.INIT('h0001)
	) name1793 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7620_
	);
	LUT4 #(
		.INIT('hddfe)
	) name1794 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7621_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1795 (
		_w7619_,
		_w7600_,
		_w7621_,
		_w7608_,
		_w7622_
	);
	LUT2 #(
		.INIT('h8)
	) name1796 (
		_w7605_,
		_w7600_,
		_w7623_
	);
	LUT3 #(
		.INIT('h04)
	) name1797 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7624_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		_w7600_,
		_w7608_,
		_w7625_
	);
	LUT3 #(
		.INIT('h80)
	) name1799 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7626_
	);
	LUT4 #(
		.INIT('h6f67)
	) name1800 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7627_
	);
	LUT4 #(
		.INIT('h7707)
	) name1801 (
		_w7623_,
		_w7624_,
		_w7625_,
		_w7627_,
		_w7628_
	);
	LUT2 #(
		.INIT('h4)
	) name1802 (
		_w7622_,
		_w7628_,
		_w7629_
	);
	LUT3 #(
		.INIT('h65)
	) name1803 (
		\u2_L11_reg[6]/NET0131 ,
		_w7618_,
		_w7629_,
		_w7630_
	);
	LUT4 #(
		.INIT('h152a)
	) name1804 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7631_
	);
	LUT4 #(
		.INIT('h6290)
	) name1805 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7632_
	);
	LUT2 #(
		.INIT('h4)
	) name1806 (
		_w7106_,
		_w7116_,
		_w7633_
	);
	LUT2 #(
		.INIT('h2)
	) name1807 (
		_w7106_,
		_w7116_,
		_w7634_
	);
	LUT2 #(
		.INIT('h9)
	) name1808 (
		_w7106_,
		_w7116_,
		_w7635_
	);
	LUT3 #(
		.INIT('h10)
	) name1809 (
		_w7290_,
		_w7632_,
		_w7635_,
		_w7636_
	);
	LUT4 #(
		.INIT('h08a8)
	) name1810 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7104_,
		_w7637_
	);
	LUT3 #(
		.INIT('h41)
	) name1811 (
		_w7103_,
		_w7102_,
		_w7108_,
		_w7638_
	);
	LUT4 #(
		.INIT('h0004)
	) name1812 (
		_w7121_,
		_w7633_,
		_w7638_,
		_w7637_,
		_w7639_
	);
	LUT4 #(
		.INIT('h0010)
	) name1813 (
		_w7105_,
		_w7591_,
		_w7634_,
		_w7631_,
		_w7640_
	);
	LUT4 #(
		.INIT('haaa9)
	) name1814 (
		\u2_L11_reg[7]/NET0131 ,
		_w7639_,
		_w7640_,
		_w7636_,
		_w7641_
	);
	LUT4 #(
		.INIT('hcffe)
	) name1815 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7642_
	);
	LUT3 #(
		.INIT('h10)
	) name1816 (
		_w7298_,
		_w7299_,
		_w7301_,
		_w7643_
	);
	LUT4 #(
		.INIT('h0031)
	) name1817 (
		_w7298_,
		_w7325_,
		_w7642_,
		_w7643_,
		_w7644_
	);
	LUT2 #(
		.INIT('h2)
	) name1818 (
		_w7312_,
		_w7644_,
		_w7645_
	);
	LUT4 #(
		.INIT('h8000)
	) name1819 (
		_w7298_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7646_
	);
	LUT3 #(
		.INIT('h04)
	) name1820 (
		_w7308_,
		_w7489_,
		_w7646_,
		_w7647_
	);
	LUT4 #(
		.INIT('hc2ff)
	) name1821 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7648_
	);
	LUT3 #(
		.INIT('h72)
	) name1822 (
		_w7298_,
		_w7304_,
		_w7648_,
		_w7649_
	);
	LUT4 #(
		.INIT('hf977)
	) name1823 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7650_
	);
	LUT4 #(
		.INIT('hcf45)
	) name1824 (
		_w7298_,
		_w7302_,
		_w7491_,
		_w7650_,
		_w7651_
	);
	LUT4 #(
		.INIT('hea00)
	) name1825 (
		_w7312_,
		_w7647_,
		_w7649_,
		_w7651_,
		_w7652_
	);
	LUT3 #(
		.INIT('h65)
	) name1826 (
		\u2_L11_reg[8]/NET0131 ,
		_w7645_,
		_w7652_,
		_w7653_
	);
	LUT4 #(
		.INIT('hf700)
	) name1827 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7654_
	);
	LUT4 #(
		.INIT('h0400)
	) name1828 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7608_,
		_w7655_
	);
	LUT4 #(
		.INIT('h006d)
	) name1829 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7656_
	);
	LUT3 #(
		.INIT('h45)
	) name1830 (
		_w7654_,
		_w7655_,
		_w7656_,
		_w7657_
	);
	LUT4 #(
		.INIT('h0100)
	) name1831 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7658_
	);
	LUT3 #(
		.INIT('h14)
	) name1832 (
		_w7601_,
		_w7602_,
		_w7605_,
		_w7659_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1833 (
		_w7608_,
		_w7611_,
		_w7658_,
		_w7659_,
		_w7660_
	);
	LUT3 #(
		.INIT('ha8)
	) name1834 (
		_w7600_,
		_w7657_,
		_w7660_,
		_w7661_
	);
	LUT3 #(
		.INIT('h40)
	) name1835 (
		_w7604_,
		_w7602_,
		_w7605_,
		_w7662_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1836 (
		_w7604_,
		_w7602_,
		_w7605_,
		_w7608_,
		_w7663_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1837 (
		_w7608_,
		_w7611_,
		_w7658_,
		_w7663_,
		_w7664_
	);
	LUT4 #(
		.INIT('h7d78)
	) name1838 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7665_
	);
	LUT3 #(
		.INIT('he0)
	) name1839 (
		_w7601_,
		_w7602_,
		_w7608_,
		_w7666_
	);
	LUT4 #(
		.INIT('h6800)
	) name1840 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7608_,
		_w7667_
	);
	LUT4 #(
		.INIT('h0504)
	) name1841 (
		_w7620_,
		_w7608_,
		_w7667_,
		_w7665_,
		_w7668_
	);
	LUT3 #(
		.INIT('h32)
	) name1842 (
		_w7600_,
		_w7664_,
		_w7668_,
		_w7669_
	);
	LUT3 #(
		.INIT('h65)
	) name1843 (
		\u2_L11_reg[16]/NET0131 ,
		_w7661_,
		_w7669_,
		_w7670_
	);
	LUT2 #(
		.INIT('h4)
	) name1844 (
		_w7605_,
		_w7608_,
		_w7671_
	);
	LUT3 #(
		.INIT('h31)
	) name1845 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7672_
	);
	LUT2 #(
		.INIT('h8)
	) name1846 (
		_w7671_,
		_w7672_,
		_w7673_
	);
	LUT3 #(
		.INIT('h0e)
	) name1847 (
		_w7604_,
		_w7605_,
		_w7608_,
		_w7674_
	);
	LUT3 #(
		.INIT('hb0)
	) name1848 (
		_w7604_,
		_w7602_,
		_w7605_,
		_w7675_
	);
	LUT4 #(
		.INIT('h23af)
	) name1849 (
		_w7603_,
		_w7666_,
		_w7674_,
		_w7675_,
		_w7676_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1850 (
		_w7600_,
		_w7616_,
		_w7673_,
		_w7676_,
		_w7677_
	);
	LUT4 #(
		.INIT('hcaf1)
	) name1851 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7678_
	);
	LUT4 #(
		.INIT('h1000)
	) name1852 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7679_
	);
	LUT4 #(
		.INIT('h5504)
	) name1853 (
		_w7600_,
		_w7608_,
		_w7678_,
		_w7679_,
		_w7680_
	);
	LUT4 #(
		.INIT('h0021)
	) name1854 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7681_
	);
	LUT4 #(
		.INIT('hb59e)
	) name1855 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7682_
	);
	LUT2 #(
		.INIT('h1)
	) name1856 (
		_w7600_,
		_w7608_,
		_w7683_
	);
	LUT2 #(
		.INIT('h4)
	) name1857 (
		_w7682_,
		_w7683_,
		_w7684_
	);
	LUT3 #(
		.INIT('he7)
	) name1858 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7685_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name1859 (
		_w7605_,
		_w7608_,
		_w7626_,
		_w7685_,
		_w7686_
	);
	LUT3 #(
		.INIT('h10)
	) name1860 (
		_w7680_,
		_w7684_,
		_w7686_,
		_w7687_
	);
	LUT3 #(
		.INIT('h65)
	) name1861 (
		\u2_L11_reg[24]/NET0131 ,
		_w7677_,
		_w7687_,
		_w7688_
	);
	LUT4 #(
		.INIT('hfae5)
	) name1862 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7689_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name1863 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7690_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name1864 (
		_w7600_,
		_w7610_,
		_w7689_,
		_w7690_,
		_w7691_
	);
	LUT2 #(
		.INIT('h2)
	) name1865 (
		_w7608_,
		_w7691_,
		_w7692_
	);
	LUT4 #(
		.INIT('h0200)
	) name1866 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7693_
	);
	LUT3 #(
		.INIT('h0e)
	) name1867 (
		_w7604_,
		_w7602_,
		_w7608_,
		_w7694_
	);
	LUT4 #(
		.INIT('h0015)
	) name1868 (
		_w7681_,
		_w7690_,
		_w7694_,
		_w7693_,
		_w7695_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w7600_,
		_w7695_,
		_w7696_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name1870 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7605_,
		_w7697_
	);
	LUT2 #(
		.INIT('h2)
	) name1871 (
		_w7625_,
		_w7697_,
		_w7698_
	);
	LUT3 #(
		.INIT('h4c)
	) name1872 (
		_w7601_,
		_w7604_,
		_w7602_,
		_w7699_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		_w7623_,
		_w7699_,
		_w7700_
	);
	LUT4 #(
		.INIT('h0040)
	) name1874 (
		_w7601_,
		_w7604_,
		_w7605_,
		_w7608_,
		_w7701_
	);
	LUT3 #(
		.INIT('h07)
	) name1875 (
		_w7613_,
		_w7662_,
		_w7701_,
		_w7702_
	);
	LUT3 #(
		.INIT('h10)
	) name1876 (
		_w7698_,
		_w7700_,
		_w7702_,
		_w7703_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name1877 (
		\u2_L11_reg[30]/NET0131 ,
		_w7692_,
		_w7696_,
		_w7703_,
		_w7704_
	);
	LUT4 #(
		.INIT('haff3)
	) name1878 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7705_
	);
	LUT4 #(
		.INIT('hbfdf)
	) name1879 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7706_
	);
	LUT4 #(
		.INIT('hb100)
	) name1880 (
		_w7298_,
		_w7317_,
		_w7705_,
		_w7706_,
		_w7707_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		_w7312_,
		_w7707_,
		_w7708_
	);
	LUT4 #(
		.INIT('h45f0)
	) name1882 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7709_
	);
	LUT4 #(
		.INIT('h2202)
	) name1883 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7710_
	);
	LUT4 #(
		.INIT('hfa3f)
	) name1884 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7711_
	);
	LUT4 #(
		.INIT('h3120)
	) name1885 (
		_w7298_,
		_w7710_,
		_w7711_,
		_w7709_,
		_w7712_
	);
	LUT4 #(
		.INIT('hdfbe)
	) name1886 (
		_w7299_,
		_w7300_,
		_w7301_,
		_w7302_,
		_w7713_
	);
	LUT2 #(
		.INIT('h1)
	) name1887 (
		_w7298_,
		_w7713_,
		_w7714_
	);
	LUT4 #(
		.INIT('h57df)
	) name1888 (
		_w7298_,
		_w7299_,
		_w7303_,
		_w7305_,
		_w7715_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1889 (
		_w7312_,
		_w7712_,
		_w7714_,
		_w7715_,
		_w7716_
	);
	LUT3 #(
		.INIT('h65)
	) name1890 (
		\u2_L11_reg[3]/NET0131 ,
		_w7708_,
		_w7716_,
		_w7717_
	);
	LUT4 #(
		.INIT('h9b99)
	) name1891 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7718_
	);
	LUT3 #(
		.INIT('h19)
	) name1892 (
		_w7142_,
		_w7141_,
		_w7143_,
		_w7719_
	);
	LUT4 #(
		.INIT('h4810)
	) name1893 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7720_
	);
	LUT4 #(
		.INIT('h0b01)
	) name1894 (
		_w7138_,
		_w7719_,
		_w7720_,
		_w7718_,
		_w7721_
	);
	LUT4 #(
		.INIT('hf77f)
	) name1895 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7722_
	);
	LUT2 #(
		.INIT('h1)
	) name1896 (
		_w7138_,
		_w7722_,
		_w7723_
	);
	LUT4 #(
		.INIT('h9060)
	) name1897 (
		_w7142_,
		_w7141_,
		_w7140_,
		_w7143_,
		_w7724_
	);
	LUT4 #(
		.INIT('h0013)
	) name1898 (
		_w7152_,
		_w7347_,
		_w7719_,
		_w7724_,
		_w7725_
	);
	LUT4 #(
		.INIT('h0e04)
	) name1899 (
		_w7139_,
		_w7721_,
		_w7723_,
		_w7725_,
		_w7726_
	);
	LUT2 #(
		.INIT('h9)
	) name1900 (
		\u2_L11_reg[9]/NET0131 ,
		_w7726_,
		_w7727_
	);
	LUT4 #(
		.INIT('h1a00)
	) name1901 (
		_w7400_,
		_w7401_,
		_w7402_,
		_w7405_,
		_w7728_
	);
	LUT2 #(
		.INIT('h8)
	) name1902 (
		_w7403_,
		_w7402_,
		_w7729_
	);
	LUT4 #(
		.INIT('h00c4)
	) name1903 (
		_w7400_,
		_w7401_,
		_w7402_,
		_w7405_,
		_w7730_
	);
	LUT4 #(
		.INIT('h2022)
	) name1904 (
		_w7415_,
		_w7455_,
		_w7729_,
		_w7730_,
		_w7731_
	);
	LUT2 #(
		.INIT('h2)
	) name1905 (
		_w7400_,
		_w7405_,
		_w7732_
	);
	LUT4 #(
		.INIT('he000)
	) name1906 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7733_
	);
	LUT4 #(
		.INIT('h0109)
	) name1907 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7405_,
		_w7734_
	);
	LUT4 #(
		.INIT('h0405)
	) name1908 (
		_w7448_,
		_w7732_,
		_w7734_,
		_w7733_,
		_w7735_
	);
	LUT4 #(
		.INIT('h45cf)
	) name1909 (
		_w7422_,
		_w7728_,
		_w7731_,
		_w7735_,
		_w7736_
	);
	LUT4 #(
		.INIT('h0020)
	) name1910 (
		_w7400_,
		_w7401_,
		_w7402_,
		_w7405_,
		_w7737_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name1911 (
		_w7403_,
		_w7400_,
		_w7401_,
		_w7402_,
		_w7738_
	);
	LUT3 #(
		.INIT('h31)
	) name1912 (
		_w7405_,
		_w7737_,
		_w7738_,
		_w7739_
	);
	LUT3 #(
		.INIT('h65)
	) name1913 (
		\u2_L11_reg[18]/P0001 ,
		_w7736_,
		_w7739_,
		_w7740_
	);
	LUT4 #(
		.INIT('hc963)
	) name1914 (
		decrypt_pad,
		\u2_R10_reg[4]/NET0131 ,
		\u2_uk_K_r10_reg[39]/NET0131 ,
		\u2_uk_K_r10_reg[5]/NET0131 ,
		_w7741_
	);
	LUT4 #(
		.INIT('hc963)
	) name1915 (
		decrypt_pad,
		\u2_R10_reg[1]/NET0131 ,
		\u2_uk_K_r10_reg[12]/NET0131 ,
		\u2_uk_K_r10_reg[3]/NET0131 ,
		_w7742_
	);
	LUT4 #(
		.INIT('hc693)
	) name1916 (
		decrypt_pad,
		\u2_R10_reg[3]/NET0131 ,
		\u2_uk_K_r10_reg[27]/NET0131 ,
		\u2_uk_K_r10_reg[4]/NET0131 ,
		_w7743_
	);
	LUT4 #(
		.INIT('hc693)
	) name1917 (
		decrypt_pad,
		\u2_R10_reg[2]/NET0131 ,
		\u2_uk_K_r10_reg[18]/NET0131 ,
		\u2_uk_K_r10_reg[27]/NET0131 ,
		_w7744_
	);
	LUT4 #(
		.INIT('hc963)
	) name1918 (
		decrypt_pad,
		\u2_R10_reg[5]/NET0131 ,
		\u2_uk_K_r10_reg[10]/NET0131 ,
		\u2_uk_K_r10_reg[33]/NET0131 ,
		_w7745_
	);
	LUT4 #(
		.INIT('hc693)
	) name1919 (
		decrypt_pad,
		\u2_R10_reg[32]/NET0131 ,
		\u2_uk_K_r10_reg[39]/NET0131 ,
		\u2_uk_K_r10_reg[48]/NET0131 ,
		_w7746_
	);
	LUT4 #(
		.INIT('hff7c)
	) name1920 (
		_w7743_,
		_w7744_,
		_w7745_,
		_w7746_,
		_w7747_
	);
	LUT2 #(
		.INIT('h2)
	) name1921 (
		_w7742_,
		_w7747_,
		_w7748_
	);
	LUT4 #(
		.INIT('h2000)
	) name1922 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7749_
	);
	LUT4 #(
		.INIT('h9bff)
	) name1923 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7750_
	);
	LUT4 #(
		.INIT('h0400)
	) name1924 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7751_
	);
	LUT3 #(
		.INIT('h0d)
	) name1925 (
		_w7743_,
		_w7750_,
		_w7751_,
		_w7752_
	);
	LUT3 #(
		.INIT('h45)
	) name1926 (
		_w7741_,
		_w7748_,
		_w7752_,
		_w7753_
	);
	LUT3 #(
		.INIT('h02)
	) name1927 (
		_w7744_,
		_w7745_,
		_w7746_,
		_w7754_
	);
	LUT4 #(
		.INIT('hf3d1)
	) name1928 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7755_
	);
	LUT2 #(
		.INIT('h2)
	) name1929 (
		_w7743_,
		_w7755_,
		_w7756_
	);
	LUT2 #(
		.INIT('h4)
	) name1930 (
		_w7743_,
		_w7742_,
		_w7757_
	);
	LUT4 #(
		.INIT('haafc)
	) name1931 (
		_w7743_,
		_w7744_,
		_w7745_,
		_w7742_,
		_w7758_
	);
	LUT2 #(
		.INIT('h2)
	) name1932 (
		_w7743_,
		_w7744_,
		_w7759_
	);
	LUT3 #(
		.INIT('hd0)
	) name1933 (
		_w7743_,
		_w7744_,
		_w7742_,
		_w7760_
	);
	LUT3 #(
		.INIT('h0e)
	) name1934 (
		_w7744_,
		_w7745_,
		_w7746_,
		_w7761_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1935 (
		_w7746_,
		_w7758_,
		_w7760_,
		_w7761_,
		_w7762_
	);
	LUT3 #(
		.INIT('h8a)
	) name1936 (
		_w7741_,
		_w7756_,
		_w7762_,
		_w7763_
	);
	LUT4 #(
		.INIT('hfdae)
	) name1937 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7764_
	);
	LUT4 #(
		.INIT('h0008)
	) name1938 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7765_
	);
	LUT4 #(
		.INIT('h6fe7)
	) name1939 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7766_
	);
	LUT4 #(
		.INIT('h0155)
	) name1940 (
		_w7743_,
		_w7764_,
		_w7741_,
		_w7766_,
		_w7767_
	);
	LUT2 #(
		.INIT('h2)
	) name1941 (
		_w7743_,
		_w7742_,
		_w7768_
	);
	LUT4 #(
		.INIT('h0200)
	) name1942 (
		_w7743_,
		_w7744_,
		_w7742_,
		_w7746_,
		_w7769_
	);
	LUT3 #(
		.INIT('h07)
	) name1943 (
		_w7754_,
		_w7768_,
		_w7769_,
		_w7770_
	);
	LUT2 #(
		.INIT('h4)
	) name1944 (
		_w7767_,
		_w7770_,
		_w7771_
	);
	LUT4 #(
		.INIT('h5655)
	) name1945 (
		\u2_L10_reg[31]/NET0131 ,
		_w7763_,
		_w7753_,
		_w7771_,
		_w7772_
	);
	LUT4 #(
		.INIT('hc693)
	) name1946 (
		decrypt_pad,
		\u2_R10_reg[28]/NET0131 ,
		\u2_uk_K_r10_reg[36]/NET0131 ,
		\u2_uk_K_r10_reg[45]/P0001 ,
		_w7773_
	);
	LUT4 #(
		.INIT('hc963)
	) name1947 (
		decrypt_pad,
		\u2_R10_reg[27]/NET0131 ,
		\u2_uk_K_r10_reg[30]/NET0131 ,
		\u2_uk_K_r10_reg[49]/NET0131 ,
		_w7774_
	);
	LUT4 #(
		.INIT('hc693)
	) name1948 (
		decrypt_pad,
		\u2_R10_reg[26]/NET0131 ,
		\u2_uk_K_r10_reg[16]/NET0131 ,
		\u2_uk_K_r10_reg[21]/NET0131 ,
		_w7775_
	);
	LUT4 #(
		.INIT('hc963)
	) name1949 (
		decrypt_pad,
		\u2_R10_reg[24]/NET0131 ,
		\u2_uk_K_r10_reg[1]/NET0131 ,
		\u2_uk_K_r10_reg[51]/NET0131 ,
		_w7776_
	);
	LUT4 #(
		.INIT('hc693)
	) name1950 (
		decrypt_pad,
		\u2_R10_reg[29]/NET0131 ,
		\u2_uk_K_r10_reg[28]/NET0131 ,
		\u2_uk_K_r10_reg[9]/NET0131 ,
		_w7777_
	);
	LUT4 #(
		.INIT('hc693)
	) name1951 (
		decrypt_pad,
		\u2_R10_reg[25]/NET0131 ,
		\u2_uk_K_r10_reg[0]/NET0131 ,
		\u2_uk_K_r10_reg[36]/NET0131 ,
		_w7778_
	);
	LUT4 #(
		.INIT('h0008)
	) name1952 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w7779_
	);
	LUT4 #(
		.INIT('hdfd7)
	) name1953 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w7780_
	);
	LUT2 #(
		.INIT('h1)
	) name1954 (
		_w7774_,
		_w7780_,
		_w7781_
	);
	LUT2 #(
		.INIT('h6)
	) name1955 (
		_w7778_,
		_w7775_,
		_w7782_
	);
	LUT2 #(
		.INIT('h8)
	) name1956 (
		_w7776_,
		_w7774_,
		_w7783_
	);
	LUT4 #(
		.INIT('h80c0)
	) name1957 (
		_w7777_,
		_w7776_,
		_w7774_,
		_w7778_,
		_w7784_
	);
	LUT2 #(
		.INIT('h2)
	) name1958 (
		_w7777_,
		_w7776_,
		_w7785_
	);
	LUT2 #(
		.INIT('h4)
	) name1959 (
		_w7778_,
		_w7775_,
		_w7786_
	);
	LUT4 #(
		.INIT('h0200)
	) name1960 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w7787_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name1961 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w7788_
	);
	LUT3 #(
		.INIT('h70)
	) name1962 (
		_w7782_,
		_w7784_,
		_w7788_,
		_w7789_
	);
	LUT3 #(
		.INIT('h8a)
	) name1963 (
		_w7773_,
		_w7781_,
		_w7789_,
		_w7790_
	);
	LUT4 #(
		.INIT('h0100)
	) name1964 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w7791_
	);
	LUT4 #(
		.INIT('h36bf)
	) name1965 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w7792_
	);
	LUT2 #(
		.INIT('h1)
	) name1966 (
		_w7774_,
		_w7792_,
		_w7793_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1967 (
		_w7777_,
		_w7776_,
		_w7774_,
		_w7778_,
		_w7794_
	);
	LUT4 #(
		.INIT('h0008)
	) name1968 (
		_w7776_,
		_w7774_,
		_w7778_,
		_w7775_,
		_w7795_
	);
	LUT2 #(
		.INIT('h8)
	) name1969 (
		_w7776_,
		_w7775_,
		_w7796_
	);
	LUT2 #(
		.INIT('h6)
	) name1970 (
		_w7776_,
		_w7775_,
		_w7797_
	);
	LUT4 #(
		.INIT('h8020)
	) name1971 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w7798_
	);
	LUT4 #(
		.INIT('h000e)
	) name1972 (
		_w7794_,
		_w7775_,
		_w7795_,
		_w7798_,
		_w7799_
	);
	LUT4 #(
		.INIT('h1000)
	) name1973 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w7800_
	);
	LUT4 #(
		.INIT('he9fb)
	) name1974 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w7801_
	);
	LUT4 #(
		.INIT('h2010)
	) name1975 (
		_w7776_,
		_w7774_,
		_w7778_,
		_w7775_,
		_w7802_
	);
	LUT4 #(
		.INIT('h0004)
	) name1976 (
		_w7777_,
		_w7774_,
		_w7778_,
		_w7775_,
		_w7803_
	);
	LUT4 #(
		.INIT('h0301)
	) name1977 (
		_w7774_,
		_w7802_,
		_w7803_,
		_w7801_,
		_w7804_
	);
	LUT4 #(
		.INIT('hf400)
	) name1978 (
		_w7793_,
		_w7799_,
		_w7773_,
		_w7804_,
		_w7805_
	);
	LUT3 #(
		.INIT('h65)
	) name1979 (
		\u2_L10_reg[22]/NET0131 ,
		_w7790_,
		_w7805_,
		_w7806_
	);
	LUT4 #(
		.INIT('hc693)
	) name1980 (
		decrypt_pad,
		\u2_R10_reg[24]/NET0131 ,
		\u2_uk_K_r10_reg[29]/NET0131 ,
		\u2_uk_K_r10_reg[38]/NET0131 ,
		_w7807_
	);
	LUT4 #(
		.INIT('hc693)
	) name1981 (
		decrypt_pad,
		\u2_R10_reg[23]/NET0131 ,
		\u2_uk_K_r10_reg[31]/NET0131 ,
		\u2_uk_K_r10_reg[8]/NET0131 ,
		_w7808_
	);
	LUT4 #(
		.INIT('hc963)
	) name1982 (
		decrypt_pad,
		\u2_R10_reg[20]/NET0131 ,
		\u2_uk_K_r10_reg[44]/NET0131 ,
		\u2_uk_K_r10_reg[8]/NET0131 ,
		_w7809_
	);
	LUT4 #(
		.INIT('hc963)
	) name1983 (
		decrypt_pad,
		\u2_R10_reg[25]/NET0131 ,
		\u2_uk_K_r10_reg[29]/NET0131 ,
		\u2_uk_K_r10_reg[52]/NET0131 ,
		_w7810_
	);
	LUT4 #(
		.INIT('hc693)
	) name1984 (
		decrypt_pad,
		\u2_R10_reg[22]/NET0131 ,
		\u2_uk_K_r10_reg[14]/NET0131 ,
		\u2_uk_K_r10_reg[50]/NET0131 ,
		_w7811_
	);
	LUT4 #(
		.INIT('hc693)
	) name1985 (
		decrypt_pad,
		\u2_R10_reg[21]/NET0131 ,
		\u2_uk_K_r10_reg[23]/NET0131 ,
		\u2_uk_K_r10_reg[28]/NET0131 ,
		_w7812_
	);
	LUT4 #(
		.INIT('hed75)
	) name1986 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7813_
	);
	LUT2 #(
		.INIT('h1)
	) name1987 (
		_w7808_,
		_w7813_,
		_w7814_
	);
	LUT4 #(
		.INIT('h0004)
	) name1988 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7815_
	);
	LUT4 #(
		.INIT('h1fdb)
	) name1989 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7816_
	);
	LUT4 #(
		.INIT('h1000)
	) name1990 (
		_w7808_,
		_w7811_,
		_w7809_,
		_w7810_,
		_w7817_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name1991 (
		_w7808_,
		_w7812_,
		_w7816_,
		_w7817_,
		_w7818_
	);
	LUT3 #(
		.INIT('h8a)
	) name1992 (
		_w7807_,
		_w7814_,
		_w7818_,
		_w7819_
	);
	LUT4 #(
		.INIT('h1400)
	) name1993 (
		_w7808_,
		_w7811_,
		_w7809_,
		_w7812_,
		_w7820_
	);
	LUT4 #(
		.INIT('h0010)
	) name1994 (
		_w7808_,
		_w7811_,
		_w7809_,
		_w7810_,
		_w7821_
	);
	LUT4 #(
		.INIT('h0800)
	) name1995 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7822_
	);
	LUT4 #(
		.INIT('h0200)
	) name1996 (
		_w7808_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7823_
	);
	LUT4 #(
		.INIT('h0040)
	) name1997 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7824_
	);
	LUT4 #(
		.INIT('h0001)
	) name1998 (
		_w7823_,
		_w7824_,
		_w7821_,
		_w7822_,
		_w7825_
	);
	LUT3 #(
		.INIT('h45)
	) name1999 (
		_w7807_,
		_w7820_,
		_w7825_,
		_w7826_
	);
	LUT4 #(
		.INIT('h0019)
	) name2000 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7807_,
		_w7827_
	);
	LUT4 #(
		.INIT('h77ef)
	) name2001 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7828_
	);
	LUT3 #(
		.INIT('h8a)
	) name2002 (
		_w7808_,
		_w7827_,
		_w7828_,
		_w7829_
	);
	LUT3 #(
		.INIT('h01)
	) name2003 (
		_w7809_,
		_w7812_,
		_w7810_,
		_w7830_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name2004 (
		_w7808_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7831_
	);
	LUT4 #(
		.INIT('hefcc)
	) name2005 (
		_w7808_,
		_w7811_,
		_w7830_,
		_w7831_,
		_w7832_
	);
	LUT2 #(
		.INIT('h4)
	) name2006 (
		_w7829_,
		_w7832_,
		_w7833_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2007 (
		\u2_L10_reg[11]/NET0131 ,
		_w7826_,
		_w7819_,
		_w7833_,
		_w7834_
	);
	LUT4 #(
		.INIT('hc693)
	) name2008 (
		decrypt_pad,
		\u2_R10_reg[16]/NET0131 ,
		\u2_uk_K_r10_reg[32]/NET0131 ,
		\u2_uk_K_r10_reg[41]/NET0131 ,
		_w7835_
	);
	LUT4 #(
		.INIT('hc693)
	) name2009 (
		decrypt_pad,
		\u2_R10_reg[15]/NET0131 ,
		\u2_uk_K_r10_reg[24]/NET0131 ,
		\u2_uk_K_r10_reg[33]/NET0131 ,
		_w7836_
	);
	LUT4 #(
		.INIT('hc963)
	) name2010 (
		decrypt_pad,
		\u2_R10_reg[14]/NET0131 ,
		\u2_uk_K_r10_reg[25]/NET0131 ,
		\u2_uk_K_r10_reg[48]/NET0131 ,
		_w7837_
	);
	LUT4 #(
		.INIT('hc693)
	) name2011 (
		decrypt_pad,
		\u2_R10_reg[12]/NET0131 ,
		\u2_uk_K_r10_reg[53]/NET0131 ,
		\u2_uk_K_r10_reg[5]/NET0131 ,
		_w7838_
	);
	LUT4 #(
		.INIT('hc963)
	) name2012 (
		decrypt_pad,
		\u2_R10_reg[13]/NET0131 ,
		\u2_uk_K_r10_reg[24]/NET0131 ,
		\u2_uk_K_r10_reg[47]/NET0131 ,
		_w7839_
	);
	LUT2 #(
		.INIT('h4)
	) name2013 (
		_w7838_,
		_w7839_,
		_w7840_
	);
	LUT4 #(
		.INIT('h0006)
	) name2014 (
		_w7838_,
		_w7839_,
		_w7836_,
		_w7837_,
		_w7841_
	);
	LUT4 #(
		.INIT('hc693)
	) name2015 (
		decrypt_pad,
		\u2_R10_reg[17]/NET0131 ,
		\u2_uk_K_r10_reg[12]/NET0131 ,
		\u2_uk_K_r10_reg[46]/NET0131 ,
		_w7842_
	);
	LUT2 #(
		.INIT('h4)
	) name2016 (
		_w7838_,
		_w7842_,
		_w7843_
	);
	LUT2 #(
		.INIT('h8)
	) name2017 (
		_w7839_,
		_w7836_,
		_w7844_
	);
	LUT4 #(
		.INIT('h2000)
	) name2018 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7836_,
		_w7845_
	);
	LUT4 #(
		.INIT('hdbff)
	) name2019 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7836_,
		_w7846_
	);
	LUT2 #(
		.INIT('h4)
	) name2020 (
		_w7841_,
		_w7846_,
		_w7847_
	);
	LUT4 #(
		.INIT('h0040)
	) name2021 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w7848_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name2022 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w7849_
	);
	LUT4 #(
		.INIT('h0001)
	) name2023 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7836_,
		_w7850_
	);
	LUT3 #(
		.INIT('h4c)
	) name2024 (
		_w7837_,
		_w7849_,
		_w7850_,
		_w7851_
	);
	LUT3 #(
		.INIT('h2a)
	) name2025 (
		_w7835_,
		_w7847_,
		_w7851_,
		_w7852_
	);
	LUT4 #(
		.INIT('h8000)
	) name2026 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7836_,
		_w7853_
	);
	LUT3 #(
		.INIT('h80)
	) name2027 (
		_w7839_,
		_w7836_,
		_w7837_,
		_w7854_
	);
	LUT4 #(
		.INIT('h4000)
	) name2028 (
		_w7838_,
		_w7839_,
		_w7836_,
		_w7837_,
		_w7855_
	);
	LUT4 #(
		.INIT('h0100)
	) name2029 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7836_,
		_w7856_
	);
	LUT4 #(
		.INIT('h0008)
	) name2030 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w7857_
	);
	LUT4 #(
		.INIT('h0001)
	) name2031 (
		_w7853_,
		_w7855_,
		_w7856_,
		_w7857_,
		_w7858_
	);
	LUT4 #(
		.INIT('heffe)
	) name2032 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w7859_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name2033 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w7860_
	);
	LUT3 #(
		.INIT('hc8)
	) name2034 (
		_w7836_,
		_w7859_,
		_w7860_,
		_w7861_
	);
	LUT3 #(
		.INIT('h15)
	) name2035 (
		_w7835_,
		_w7858_,
		_w7861_,
		_w7862_
	);
	LUT4 #(
		.INIT('h0200)
	) name2036 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w7863_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name2037 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w7864_
	);
	LUT2 #(
		.INIT('h2)
	) name2038 (
		_w7836_,
		_w7864_,
		_w7865_
	);
	LUT3 #(
		.INIT('h02)
	) name2039 (
		_w7842_,
		_w7836_,
		_w7837_,
		_w7866_
	);
	LUT3 #(
		.INIT('h02)
	) name2040 (
		_w7838_,
		_w7842_,
		_w7837_,
		_w7867_
	);
	LUT4 #(
		.INIT('h135f)
	) name2041 (
		_w7840_,
		_w7844_,
		_w7866_,
		_w7867_,
		_w7868_
	);
	LUT2 #(
		.INIT('h4)
	) name2042 (
		_w7865_,
		_w7868_,
		_w7869_
	);
	LUT4 #(
		.INIT('h5655)
	) name2043 (
		\u2_L10_reg[20]/NET0131 ,
		_w7862_,
		_w7852_,
		_w7869_,
		_w7870_
	);
	LUT4 #(
		.INIT('hc963)
	) name2044 (
		decrypt_pad,
		\u2_R10_reg[8]/NET0131 ,
		\u2_uk_K_r10_reg[40]/NET0131 ,
		\u2_uk_K_r10_reg[6]/NET0131 ,
		_w7871_
	);
	LUT4 #(
		.INIT('hc963)
	) name2045 (
		decrypt_pad,
		\u2_R10_reg[7]/NET0131 ,
		\u2_uk_K_r10_reg[17]/NET0131 ,
		\u2_uk_K_r10_reg[40]/NET0131 ,
		_w7872_
	);
	LUT4 #(
		.INIT('hc963)
	) name2046 (
		decrypt_pad,
		\u2_R10_reg[5]/NET0131 ,
		\u2_uk_K_r10_reg[32]/NET0131 ,
		\u2_uk_K_r10_reg[55]/NET0131 ,
		_w7873_
	);
	LUT4 #(
		.INIT('hc693)
	) name2047 (
		decrypt_pad,
		\u2_R10_reg[4]/NET0131 ,
		\u2_uk_K_r10_reg[19]/NET0131 ,
		\u2_uk_K_r10_reg[53]/NET0131 ,
		_w7874_
	);
	LUT4 #(
		.INIT('hc693)
	) name2048 (
		decrypt_pad,
		\u2_R10_reg[9]/NET0131 ,
		\u2_uk_K_r10_reg[11]/NET0131 ,
		\u2_uk_K_r10_reg[20]/NET0131 ,
		_w7875_
	);
	LUT4 #(
		.INIT('hc693)
	) name2049 (
		decrypt_pad,
		\u2_R10_reg[6]/NET0131 ,
		\u2_uk_K_r10_reg[46]/NET0131 ,
		\u2_uk_K_r10_reg[55]/NET0131 ,
		_w7876_
	);
	LUT4 #(
		.INIT('h59fb)
	) name2050 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7877_
	);
	LUT2 #(
		.INIT('h1)
	) name2051 (
		_w7872_,
		_w7877_,
		_w7878_
	);
	LUT4 #(
		.INIT('h4000)
	) name2052 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7879_
	);
	LUT4 #(
		.INIT('h0004)
	) name2053 (
		_w7872_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7880_
	);
	LUT2 #(
		.INIT('h1)
	) name2054 (
		_w7879_,
		_w7880_,
		_w7881_
	);
	LUT4 #(
		.INIT('h0800)
	) name2055 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7882_
	);
	LUT4 #(
		.INIT('h0034)
	) name2056 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7883_
	);
	LUT3 #(
		.INIT('h07)
	) name2057 (
		_w7872_,
		_w7882_,
		_w7883_,
		_w7884_
	);
	LUT4 #(
		.INIT('h4555)
	) name2058 (
		_w7871_,
		_w7878_,
		_w7881_,
		_w7884_,
		_w7885_
	);
	LUT4 #(
		.INIT('he6ee)
	) name2059 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7886_
	);
	LUT4 #(
		.INIT('h4044)
	) name2060 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7887_
	);
	LUT3 #(
		.INIT('h51)
	) name2061 (
		_w7872_,
		_w7873_,
		_w7876_,
		_w7888_
	);
	LUT4 #(
		.INIT('hf200)
	) name2062 (
		_w7871_,
		_w7886_,
		_w7887_,
		_w7888_,
		_w7889_
	);
	LUT3 #(
		.INIT('h10)
	) name2063 (
		_w7875_,
		_w7873_,
		_w7876_,
		_w7890_
	);
	LUT4 #(
		.INIT('h0100)
	) name2064 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7891_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name2065 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7892_
	);
	LUT2 #(
		.INIT('h2)
	) name2066 (
		_w7872_,
		_w7892_,
		_w7893_
	);
	LUT4 #(
		.INIT('h0002)
	) name2067 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7894_
	);
	LUT4 #(
		.INIT('h0080)
	) name2068 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w7895_
	);
	LUT4 #(
		.INIT('h80a0)
	) name2069 (
		_w7872_,
		_w7874_,
		_w7873_,
		_w7876_,
		_w7896_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2070 (
		_w7871_,
		_w7895_,
		_w7896_,
		_w7894_,
		_w7897_
	);
	LUT3 #(
		.INIT('h01)
	) name2071 (
		_w7893_,
		_w7897_,
		_w7889_,
		_w7898_
	);
	LUT3 #(
		.INIT('h65)
	) name2072 (
		\u2_L10_reg[2]/NET0131 ,
		_w7885_,
		_w7898_,
		_w7899_
	);
	LUT4 #(
		.INIT('hab6f)
	) name2073 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7900_
	);
	LUT4 #(
		.INIT('h0200)
	) name2074 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7901_
	);
	LUT4 #(
		.INIT('h3fd2)
	) name2075 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7902_
	);
	LUT4 #(
		.INIT('h3120)
	) name2076 (
		_w7808_,
		_w7901_,
		_w7902_,
		_w7900_,
		_w7903_
	);
	LUT2 #(
		.INIT('h1)
	) name2077 (
		_w7807_,
		_w7903_,
		_w7904_
	);
	LUT4 #(
		.INIT('hcf6f)
	) name2078 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7905_
	);
	LUT2 #(
		.INIT('h2)
	) name2079 (
		_w7808_,
		_w7905_,
		_w7906_
	);
	LUT4 #(
		.INIT('h77dc)
	) name2080 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7907_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w7808_,
		_w7907_,
		_w7908_
	);
	LUT4 #(
		.INIT('h0102)
	) name2082 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7909_
	);
	LUT3 #(
		.INIT('h01)
	) name2083 (
		_w7821_,
		_w7822_,
		_w7909_,
		_w7910_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2084 (
		_w7807_,
		_w7908_,
		_w7906_,
		_w7910_,
		_w7911_
	);
	LUT4 #(
		.INIT('h2000)
	) name2085 (
		_w7808_,
		_w7811_,
		_w7812_,
		_w7810_,
		_w7912_
	);
	LUT2 #(
		.INIT('h1)
	) name2086 (
		_w7815_,
		_w7912_,
		_w7913_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2087 (
		\u2_L10_reg[29]/NET0131 ,
		_w7911_,
		_w7904_,
		_w7913_,
		_w7914_
	);
	LUT4 #(
		.INIT('hc693)
	) name2088 (
		decrypt_pad,
		\u2_R10_reg[32]/NET0131 ,
		\u2_uk_K_r10_reg[1]/NET0131 ,
		\u2_uk_K_r10_reg[37]/NET0131 ,
		_w7915_
	);
	LUT4 #(
		.INIT('hc963)
	) name2089 (
		decrypt_pad,
		\u2_R10_reg[31]/P0001 ,
		\u2_uk_K_r10_reg[0]/NET0131 ,
		\u2_uk_K_r10_reg[50]/NET0131 ,
		_w7916_
	);
	LUT4 #(
		.INIT('hc963)
	) name2090 (
		decrypt_pad,
		\u2_R10_reg[30]/NET0131 ,
		\u2_uk_K_r10_reg[43]/NET0131 ,
		\u2_uk_K_r10_reg[7]/NET0131 ,
		_w7917_
	);
	LUT4 #(
		.INIT('hc963)
	) name2091 (
		decrypt_pad,
		\u2_R10_reg[28]/NET0131 ,
		\u2_uk_K_r10_reg[15]/NET0131 ,
		\u2_uk_K_r10_reg[38]/NET0131 ,
		_w7918_
	);
	LUT4 #(
		.INIT('hc693)
	) name2092 (
		decrypt_pad,
		\u2_R10_reg[29]/NET0131 ,
		\u2_uk_K_r10_reg[37]/NET0131 ,
		\u2_uk_K_r10_reg[42]/NET0131 ,
		_w7919_
	);
	LUT2 #(
		.INIT('h2)
	) name2093 (
		_w7918_,
		_w7919_,
		_w7920_
	);
	LUT4 #(
		.INIT('hc693)
	) name2094 (
		decrypt_pad,
		\u2_R10_reg[1]/NET0131 ,
		\u2_uk_K_r10_reg[22]/NET0131 ,
		\u2_uk_K_r10_reg[31]/NET0131 ,
		_w7921_
	);
	LUT2 #(
		.INIT('h8)
	) name2095 (
		_w7918_,
		_w7921_,
		_w7922_
	);
	LUT4 #(
		.INIT('hdd2d)
	) name2096 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w7923_
	);
	LUT4 #(
		.INIT('h4000)
	) name2097 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w7924_
	);
	LUT3 #(
		.INIT('h01)
	) name2098 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7925_
	);
	LUT4 #(
		.INIT('h2031)
	) name2099 (
		_w7916_,
		_w7924_,
		_w7923_,
		_w7925_,
		_w7926_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		_w7915_,
		_w7926_,
		_w7927_
	);
	LUT2 #(
		.INIT('h1)
	) name2101 (
		_w7917_,
		_w7916_,
		_w7928_
	);
	LUT4 #(
		.INIT('h7b2a)
	) name2102 (
		_w7917_,
		_w7919_,
		_w7921_,
		_w7916_,
		_w7929_
	);
	LUT2 #(
		.INIT('h2)
	) name2103 (
		_w7918_,
		_w7929_,
		_w7930_
	);
	LUT4 #(
		.INIT('h0008)
	) name2104 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w7931_
	);
	LUT4 #(
		.INIT('hef00)
	) name2105 (
		_w7918_,
		_w7919_,
		_w7921_,
		_w7916_,
		_w7932_
	);
	LUT3 #(
		.INIT('h04)
	) name2106 (
		_w7918_,
		_w7917_,
		_w7921_,
		_w7933_
	);
	LUT2 #(
		.INIT('h8)
	) name2107 (
		_w7919_,
		_w7921_,
		_w7934_
	);
	LUT3 #(
		.INIT('h07)
	) name2108 (
		_w7919_,
		_w7921_,
		_w7916_,
		_w7935_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2109 (
		_w7931_,
		_w7932_,
		_w7933_,
		_w7935_,
		_w7936_
	);
	LUT3 #(
		.INIT('h0e)
	) name2110 (
		_w7930_,
		_w7936_,
		_w7915_,
		_w7937_
	);
	LUT4 #(
		.INIT('h0040)
	) name2111 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w7938_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name2112 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w7939_
	);
	LUT4 #(
		.INIT('h0400)
	) name2113 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w7940_
	);
	LUT4 #(
		.INIT('hf9be)
	) name2114 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w7941_
	);
	LUT2 #(
		.INIT('h2)
	) name2115 (
		_w7916_,
		_w7941_,
		_w7942_
	);
	LUT3 #(
		.INIT('h20)
	) name2116 (
		_w7917_,
		_w7916_,
		_w7915_,
		_w7943_
	);
	LUT3 #(
		.INIT('h08)
	) name2117 (
		_w7918_,
		_w7919_,
		_w7921_,
		_w7944_
	);
	LUT4 #(
		.INIT('h153f)
	) name2118 (
		_w7928_,
		_w7920_,
		_w7943_,
		_w7944_,
		_w7945_
	);
	LUT2 #(
		.INIT('h4)
	) name2119 (
		_w7942_,
		_w7945_,
		_w7946_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2120 (
		\u2_L10_reg[5]/NET0131 ,
		_w7937_,
		_w7927_,
		_w7946_,
		_w7947_
	);
	LUT4 #(
		.INIT('h1900)
	) name2121 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7948_
	);
	LUT4 #(
		.INIT('haa2a)
	) name2122 (
		_w7808_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7949_
	);
	LUT4 #(
		.INIT('h5545)
	) name2123 (
		_w7808_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7950_
	);
	LUT4 #(
		.INIT('h8acf)
	) name2124 (
		_w7901_,
		_w7948_,
		_w7949_,
		_w7950_,
		_w7951_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w7815_,
		_w7817_,
		_w7952_
	);
	LUT3 #(
		.INIT('h45)
	) name2126 (
		_w7807_,
		_w7951_,
		_w7952_,
		_w7953_
	);
	LUT4 #(
		.INIT('h6ee6)
	) name2127 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7954_
	);
	LUT3 #(
		.INIT('h45)
	) name2128 (
		_w7808_,
		_w7811_,
		_w7810_,
		_w7955_
	);
	LUT2 #(
		.INIT('h4)
	) name2129 (
		_w7954_,
		_w7955_,
		_w7956_
	);
	LUT3 #(
		.INIT('h04)
	) name2130 (
		_w7811_,
		_w7812_,
		_w7810_,
		_w7957_
	);
	LUT4 #(
		.INIT('heeae)
	) name2131 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7958_
	);
	LUT4 #(
		.INIT('ha010)
	) name2132 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7959_
	);
	LUT4 #(
		.INIT('h2000)
	) name2133 (
		_w7808_,
		_w7811_,
		_w7809_,
		_w7810_,
		_w7960_
	);
	LUT4 #(
		.INIT('h0032)
	) name2134 (
		_w7808_,
		_w7959_,
		_w7958_,
		_w7960_,
		_w7961_
	);
	LUT3 #(
		.INIT('hb6)
	) name2135 (
		_w7809_,
		_w7812_,
		_w7810_,
		_w7962_
	);
	LUT2 #(
		.INIT('h8)
	) name2136 (
		_w7808_,
		_w7811_,
		_w7963_
	);
	LUT2 #(
		.INIT('h4)
	) name2137 (
		_w7962_,
		_w7963_,
		_w7964_
	);
	LUT4 #(
		.INIT('h000d)
	) name2138 (
		_w7807_,
		_w7961_,
		_w7964_,
		_w7956_,
		_w7965_
	);
	LUT3 #(
		.INIT('h65)
	) name2139 (
		\u2_L10_reg[4]/NET0131 ,
		_w7953_,
		_w7965_,
		_w7966_
	);
	LUT4 #(
		.INIT('h1000)
	) name2140 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7967_
	);
	LUT2 #(
		.INIT('h2)
	) name2141 (
		_w7741_,
		_w7967_,
		_w7968_
	);
	LUT4 #(
		.INIT('hfb05)
	) name2142 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7969_
	);
	LUT3 #(
		.INIT('h80)
	) name2143 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7970_
	);
	LUT4 #(
		.INIT('h4401)
	) name2144 (
		_w7743_,
		_w7744_,
		_w7742_,
		_w7746_,
		_w7971_
	);
	LUT4 #(
		.INIT('h000d)
	) name2145 (
		_w7743_,
		_w7969_,
		_w7970_,
		_w7971_,
		_w7972_
	);
	LUT2 #(
		.INIT('h8)
	) name2146 (
		_w7968_,
		_w7972_,
		_w7973_
	);
	LUT4 #(
		.INIT('h3c9f)
	) name2147 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7974_
	);
	LUT2 #(
		.INIT('h2)
	) name2148 (
		_w7743_,
		_w7974_,
		_w7975_
	);
	LUT4 #(
		.INIT('hf3ec)
	) name2149 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w7976_
	);
	LUT2 #(
		.INIT('h1)
	) name2150 (
		_w7743_,
		_w7976_,
		_w7977_
	);
	LUT3 #(
		.INIT('h01)
	) name2151 (
		_w7765_,
		_w7741_,
		_w7749_,
		_w7978_
	);
	LUT3 #(
		.INIT('h10)
	) name2152 (
		_w7977_,
		_w7975_,
		_w7978_,
		_w7979_
	);
	LUT3 #(
		.INIT('ha9)
	) name2153 (
		\u2_L10_reg[17]/NET0131 ,
		_w7973_,
		_w7979_,
		_w7980_
	);
	LUT4 #(
		.INIT('h1001)
	) name2154 (
		_w7808_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7981_
	);
	LUT4 #(
		.INIT('h7343)
	) name2155 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7982_
	);
	LUT4 #(
		.INIT('h8000)
	) name2156 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7983_
	);
	LUT4 #(
		.INIT('h0031)
	) name2157 (
		_w7808_,
		_w7807_,
		_w7982_,
		_w7983_,
		_w7984_
	);
	LUT3 #(
		.INIT('h04)
	) name2158 (
		_w7808_,
		_w7809_,
		_w7812_,
		_w7985_
	);
	LUT4 #(
		.INIT('h0004)
	) name2159 (
		_w7823_,
		_w7807_,
		_w7957_,
		_w7985_,
		_w7986_
	);
	LUT4 #(
		.INIT('h2000)
	) name2160 (
		_w7808_,
		_w7811_,
		_w7809_,
		_w7812_,
		_w7987_
	);
	LUT4 #(
		.INIT('hdefd)
	) name2161 (
		_w7811_,
		_w7809_,
		_w7812_,
		_w7810_,
		_w7988_
	);
	LUT2 #(
		.INIT('h4)
	) name2162 (
		_w7987_,
		_w7988_,
		_w7989_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name2163 (
		_w7981_,
		_w7984_,
		_w7986_,
		_w7989_,
		_w7990_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name2164 (
		_w7811_,
		_w7812_,
		_w7831_,
		_w7817_,
		_w7991_
	);
	LUT3 #(
		.INIT('h65)
	) name2165 (
		\u2_L10_reg[19]/NET0131 ,
		_w7990_,
		_w7991_,
		_w7992_
	);
	LUT3 #(
		.INIT('h01)
	) name2166 (
		_w7838_,
		_w7842_,
		_w7837_,
		_w7993_
	);
	LUT3 #(
		.INIT('h02)
	) name2167 (
		_w7836_,
		_w7863_,
		_w7993_,
		_w7994_
	);
	LUT3 #(
		.INIT('h08)
	) name2168 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7995_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name2169 (
		_w7838_,
		_w7842_,
		_w7836_,
		_w7837_,
		_w7996_
	);
	LUT2 #(
		.INIT('h4)
	) name2170 (
		_w7995_,
		_w7996_,
		_w7997_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name2171 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w7998_
	);
	LUT4 #(
		.INIT('h0155)
	) name2172 (
		_w7835_,
		_w7994_,
		_w7997_,
		_w7998_,
		_w7999_
	);
	LUT4 #(
		.INIT('hbf2f)
	) name2173 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8000_
	);
	LUT4 #(
		.INIT('h2000)
	) name2174 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8001_
	);
	LUT4 #(
		.INIT('hdaff)
	) name2175 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8002_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2176 (
		_w7835_,
		_w7836_,
		_w8000_,
		_w8002_,
		_w8003_
	);
	LUT4 #(
		.INIT('h7bff)
	) name2177 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8004_
	);
	LUT4 #(
		.INIT('h6bff)
	) name2178 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8005_
	);
	LUT2 #(
		.INIT('h2)
	) name2179 (
		_w7836_,
		_w8005_,
		_w8006_
	);
	LUT2 #(
		.INIT('h4)
	) name2180 (
		_w7836_,
		_w8001_,
		_w8007_
	);
	LUT4 #(
		.INIT('hf3f1)
	) name2181 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8008_
	);
	LUT2 #(
		.INIT('h8)
	) name2182 (
		_w7835_,
		_w7836_,
		_w8009_
	);
	LUT4 #(
		.INIT('h7077)
	) name2183 (
		_w7837_,
		_w7850_,
		_w8008_,
		_w8009_,
		_w8010_
	);
	LUT4 #(
		.INIT('h0100)
	) name2184 (
		_w8006_,
		_w8007_,
		_w8003_,
		_w8010_,
		_w8011_
	);
	LUT3 #(
		.INIT('h65)
	) name2185 (
		\u2_L10_reg[1]/NET0131 ,
		_w7999_,
		_w8011_,
		_w8012_
	);
	LUT4 #(
		.INIT('h0004)
	) name2186 (
		_w7918_,
		_w7919_,
		_w7921_,
		_w7916_,
		_w8013_
	);
	LUT3 #(
		.INIT('hba)
	) name2187 (
		_w7917_,
		_w7919_,
		_w7916_,
		_w8014_
	);
	LUT4 #(
		.INIT('h1101)
	) name2188 (
		_w7931_,
		_w7915_,
		_w7922_,
		_w8014_,
		_w8015_
	);
	LUT4 #(
		.INIT('hf757)
	) name2189 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8016_
	);
	LUT4 #(
		.INIT('h0040)
	) name2190 (
		_w7918_,
		_w7917_,
		_w7921_,
		_w7916_,
		_w8017_
	);
	LUT4 #(
		.INIT('hbfbe)
	) name2191 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8018_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2192 (
		_w7916_,
		_w8016_,
		_w8017_,
		_w8018_,
		_w8019_
	);
	LUT3 #(
		.INIT('h40)
	) name2193 (
		_w8013_,
		_w8015_,
		_w8019_,
		_w8020_
	);
	LUT4 #(
		.INIT('hef00)
	) name2194 (
		_w7917_,
		_w7919_,
		_w7921_,
		_w7916_,
		_w8021_
	);
	LUT4 #(
		.INIT('h2f7f)
	) name2195 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8022_
	);
	LUT2 #(
		.INIT('h8)
	) name2196 (
		_w8021_,
		_w8022_,
		_w8023_
	);
	LUT3 #(
		.INIT('h02)
	) name2197 (
		_w7918_,
		_w7917_,
		_w7921_,
		_w8024_
	);
	LUT4 #(
		.INIT('h0800)
	) name2198 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8025_
	);
	LUT3 #(
		.INIT('h01)
	) name2199 (
		_w7916_,
		_w8025_,
		_w8024_,
		_w8026_
	);
	LUT4 #(
		.INIT('h0084)
	) name2200 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8027_
	);
	LUT4 #(
		.INIT('h0100)
	) name2201 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8028_
	);
	LUT3 #(
		.INIT('h02)
	) name2202 (
		_w7915_,
		_w8028_,
		_w8027_,
		_w8029_
	);
	LUT3 #(
		.INIT('he0)
	) name2203 (
		_w8023_,
		_w8026_,
		_w8029_,
		_w8030_
	);
	LUT4 #(
		.INIT('h0100)
	) name2204 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7916_,
		_w8031_
	);
	LUT3 #(
		.INIT('h02)
	) name2205 (
		_w7918_,
		_w7917_,
		_w7916_,
		_w8032_
	);
	LUT3 #(
		.INIT('h13)
	) name2206 (
		_w7934_,
		_w8031_,
		_w8032_,
		_w8033_
	);
	LUT4 #(
		.INIT('ha955)
	) name2207 (
		\u2_L10_reg[21]/NET0131 ,
		_w8020_,
		_w8030_,
		_w8033_,
		_w8034_
	);
	LUT4 #(
		.INIT('hfdc3)
	) name2208 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w8035_
	);
	LUT4 #(
		.INIT('heffb)
	) name2209 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w8036_
	);
	LUT4 #(
		.INIT('h0455)
	) name2210 (
		_w7743_,
		_w7741_,
		_w8035_,
		_w8036_,
		_w8037_
	);
	LUT4 #(
		.INIT('hdf3f)
	) name2211 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w8038_
	);
	LUT2 #(
		.INIT('h2)
	) name2212 (
		_w7743_,
		_w8038_,
		_w8039_
	);
	LUT3 #(
		.INIT('h07)
	) name2213 (
		_w7754_,
		_w7768_,
		_w7751_,
		_w8040_
	);
	LUT3 #(
		.INIT('h8a)
	) name2214 (
		_w7741_,
		_w8039_,
		_w8040_,
		_w8041_
	);
	LUT4 #(
		.INIT('hff47)
	) name2215 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w8042_
	);
	LUT2 #(
		.INIT('h2)
	) name2216 (
		_w7743_,
		_w8042_,
		_w8043_
	);
	LUT3 #(
		.INIT('h7e)
	) name2217 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w8044_
	);
	LUT3 #(
		.INIT('h40)
	) name2218 (
		_w7743_,
		_w7742_,
		_w7746_,
		_w8045_
	);
	LUT4 #(
		.INIT('h4000)
	) name2219 (
		_w7743_,
		_w7744_,
		_w7745_,
		_w7746_,
		_w8046_
	);
	LUT3 #(
		.INIT('h10)
	) name2220 (
		_w8045_,
		_w8046_,
		_w8044_,
		_w8047_
	);
	LUT4 #(
		.INIT('hbffd)
	) name2221 (
		_w7743_,
		_w7744_,
		_w7745_,
		_w7746_,
		_w8048_
	);
	LUT3 #(
		.INIT('h31)
	) name2222 (
		_w7742_,
		_w7769_,
		_w8048_,
		_w8049_
	);
	LUT4 #(
		.INIT('hba00)
	) name2223 (
		_w7741_,
		_w8043_,
		_w8047_,
		_w8049_,
		_w8050_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2224 (
		\u2_L10_reg[23]/NET0131 ,
		_w8041_,
		_w8037_,
		_w8050_,
		_w8051_
	);
	LUT4 #(
		.INIT('hc693)
	) name2225 (
		decrypt_pad,
		\u2_R10_reg[19]/NET0131 ,
		\u2_uk_K_r10_reg[2]/NET0131 ,
		\u2_uk_K_r10_reg[7]/NET0131 ,
		_w8052_
	);
	LUT4 #(
		.INIT('hc693)
	) name2226 (
		decrypt_pad,
		\u2_R10_reg[18]/NET0131 ,
		\u2_uk_K_r10_reg[15]/NET0131 ,
		\u2_uk_K_r10_reg[51]/NET0131 ,
		_w8053_
	);
	LUT4 #(
		.INIT('hc693)
	) name2227 (
		decrypt_pad,
		\u2_R10_reg[17]/NET0131 ,
		\u2_uk_K_r10_reg[21]/NET0131 ,
		\u2_uk_K_r10_reg[2]/NET0131 ,
		_w8054_
	);
	LUT4 #(
		.INIT('hc963)
	) name2228 (
		decrypt_pad,
		\u2_R10_reg[21]/NET0131 ,
		\u2_uk_K_r10_reg[23]/NET0131 ,
		\u2_uk_K_r10_reg[42]/NET0131 ,
		_w8055_
	);
	LUT4 #(
		.INIT('hc693)
	) name2229 (
		decrypt_pad,
		\u2_R10_reg[16]/NET0131 ,
		\u2_uk_K_r10_reg[30]/NET0131 ,
		\u2_uk_K_r10_reg[35]/NET0131 ,
		_w8056_
	);
	LUT3 #(
		.INIT('h80)
	) name2230 (
		_w8055_,
		_w8054_,
		_w8056_,
		_w8057_
	);
	LUT4 #(
		.INIT('h3ed0)
	) name2231 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8058_
	);
	LUT3 #(
		.INIT('h20)
	) name2232 (
		_w8055_,
		_w8054_,
		_w8056_,
		_w8059_
	);
	LUT4 #(
		.INIT('hf3af)
	) name2233 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8060_
	);
	LUT3 #(
		.INIT('h8b)
	) name2234 (
		_w8053_,
		_w8055_,
		_w8056_,
		_w8061_
	);
	LUT4 #(
		.INIT('h6040)
	) name2235 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8062_
	);
	LUT4 #(
		.INIT('h00e2)
	) name2236 (
		_w8060_,
		_w8052_,
		_w8058_,
		_w8062_,
		_w8063_
	);
	LUT4 #(
		.INIT('hc963)
	) name2237 (
		decrypt_pad,
		\u2_R10_reg[20]/NET0131 ,
		\u2_uk_K_r10_reg[22]/NET0131 ,
		\u2_uk_K_r10_reg[45]/P0001 ,
		_w8064_
	);
	LUT2 #(
		.INIT('h4)
	) name2238 (
		_w8063_,
		_w8064_,
		_w8065_
	);
	LUT4 #(
		.INIT('h2002)
	) name2239 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8066_
	);
	LUT4 #(
		.INIT('hdff9)
	) name2240 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8067_
	);
	LUT2 #(
		.INIT('h2)
	) name2241 (
		_w8052_,
		_w8067_,
		_w8068_
	);
	LUT4 #(
		.INIT('hfc5f)
	) name2242 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8069_
	);
	LUT2 #(
		.INIT('h4)
	) name2243 (
		_w8055_,
		_w8052_,
		_w8070_
	);
	LUT3 #(
		.INIT('hb0)
	) name2244 (
		_w8055_,
		_w8054_,
		_w8052_,
		_w8071_
	);
	LUT4 #(
		.INIT('h5501)
	) name2245 (
		_w8053_,
		_w8054_,
		_w8056_,
		_w8052_,
		_w8072_
	);
	LUT4 #(
		.INIT('he0ee)
	) name2246 (
		_w8069_,
		_w8070_,
		_w8071_,
		_w8072_,
		_w8073_
	);
	LUT4 #(
		.INIT('h4000)
	) name2247 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8074_
	);
	LUT2 #(
		.INIT('h2)
	) name2248 (
		_w8053_,
		_w8052_,
		_w8075_
	);
	LUT4 #(
		.INIT('h0020)
	) name2249 (
		_w8053_,
		_w8054_,
		_w8056_,
		_w8052_,
		_w8076_
	);
	LUT2 #(
		.INIT('h1)
	) name2250 (
		_w8074_,
		_w8076_,
		_w8077_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2251 (
		_w8064_,
		_w8073_,
		_w8068_,
		_w8077_,
		_w8078_
	);
	LUT3 #(
		.INIT('h65)
	) name2252 (
		\u2_L10_reg[25]/NET0131 ,
		_w8065_,
		_w8078_,
		_w8079_
	);
	LUT4 #(
		.INIT('h5551)
	) name2253 (
		_w7835_,
		_w7838_,
		_w7839_,
		_w7837_,
		_w8080_
	);
	LUT2 #(
		.INIT('h4)
	) name2254 (
		_w7845_,
		_w8080_,
		_w8081_
	);
	LUT3 #(
		.INIT('h0d)
	) name2255 (
		_w7854_,
		_w7843_,
		_w7848_,
		_w8082_
	);
	LUT2 #(
		.INIT('h8)
	) name2256 (
		_w8081_,
		_w8082_,
		_w8083_
	);
	LUT4 #(
		.INIT('h9b9f)
	) name2257 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7836_,
		_w8084_
	);
	LUT2 #(
		.INIT('h2)
	) name2258 (
		_w7837_,
		_w8084_,
		_w8085_
	);
	LUT4 #(
		.INIT('h77fb)
	) name2259 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8086_
	);
	LUT2 #(
		.INIT('h1)
	) name2260 (
		_w7836_,
		_w8086_,
		_w8087_
	);
	LUT4 #(
		.INIT('h0010)
	) name2261 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8088_
	);
	LUT3 #(
		.INIT('h02)
	) name2262 (
		_w7835_,
		_w7856_,
		_w8088_,
		_w8089_
	);
	LUT3 #(
		.INIT('h10)
	) name2263 (
		_w8087_,
		_w8085_,
		_w8089_,
		_w8090_
	);
	LUT4 #(
		.INIT('h0092)
	) name2264 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8091_
	);
	LUT4 #(
		.INIT('hf8fc)
	) name2265 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8092_
	);
	LUT4 #(
		.INIT('h0302)
	) name2266 (
		_w7835_,
		_w7836_,
		_w8091_,
		_w8092_,
		_w8093_
	);
	LUT3 #(
		.INIT('h02)
	) name2267 (
		_w7836_,
		_w7857_,
		_w7848_,
		_w8094_
	);
	LUT2 #(
		.INIT('h1)
	) name2268 (
		_w8093_,
		_w8094_,
		_w8095_
	);
	LUT4 #(
		.INIT('h55a9)
	) name2269 (
		\u2_L10_reg[26]/NET0131 ,
		_w8083_,
		_w8090_,
		_w8095_,
		_w8096_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name2270 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8097_
	);
	LUT2 #(
		.INIT('h2)
	) name2271 (
		_w7872_,
		_w8097_,
		_w8098_
	);
	LUT4 #(
		.INIT('hbfae)
	) name2272 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8099_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w7872_,
		_w8099_,
		_w8100_
	);
	LUT2 #(
		.INIT('h8)
	) name2274 (
		_w7872_,
		_w7874_,
		_w8101_
	);
	LUT4 #(
		.INIT('h7737)
	) name2275 (
		_w7872_,
		_w7874_,
		_w7875_,
		_w7873_,
		_w8102_
	);
	LUT4 #(
		.INIT('h0400)
	) name2276 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8103_
	);
	LUT3 #(
		.INIT('h0e)
	) name2277 (
		_w7876_,
		_w8102_,
		_w8103_,
		_w8104_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2278 (
		_w7871_,
		_w8100_,
		_w8098_,
		_w8104_,
		_w8105_
	);
	LUT4 #(
		.INIT('h2000)
	) name2279 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8106_
	);
	LUT4 #(
		.INIT('hdaff)
	) name2280 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8107_
	);
	LUT2 #(
		.INIT('h1)
	) name2281 (
		_w7872_,
		_w8107_,
		_w8108_
	);
	LUT4 #(
		.INIT('h2900)
	) name2282 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8109_
	);
	LUT4 #(
		.INIT('h5b59)
	) name2283 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8110_
	);
	LUT4 #(
		.INIT('h00e4)
	) name2284 (
		_w7872_,
		_w8110_,
		_w8099_,
		_w8109_,
		_w8111_
	);
	LUT3 #(
		.INIT('h32)
	) name2285 (
		_w7871_,
		_w8108_,
		_w8111_,
		_w8112_
	);
	LUT3 #(
		.INIT('h65)
	) name2286 (
		\u2_L10_reg[28]/NET0131 ,
		_w8105_,
		_w8112_,
		_w8113_
	);
	LUT4 #(
		.INIT('h0200)
	) name2287 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8114_
	);
	LUT2 #(
		.INIT('h1)
	) name2288 (
		_w8052_,
		_w8114_,
		_w8115_
	);
	LUT4 #(
		.INIT('h0008)
	) name2289 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8116_
	);
	LUT4 #(
		.INIT('h0040)
	) name2290 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8117_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2291 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8052_,
		_w8118_
	);
	LUT3 #(
		.INIT('h10)
	) name2292 (
		_w8116_,
		_w8117_,
		_w8118_,
		_w8119_
	);
	LUT2 #(
		.INIT('h1)
	) name2293 (
		_w8115_,
		_w8119_,
		_w8120_
	);
	LUT4 #(
		.INIT('hffd7)
	) name2294 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8121_
	);
	LUT4 #(
		.INIT('h0001)
	) name2295 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8122_
	);
	LUT4 #(
		.INIT('hf3fe)
	) name2296 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8123_
	);
	LUT2 #(
		.INIT('h1)
	) name2297 (
		_w8053_,
		_w8052_,
		_w8124_
	);
	LUT4 #(
		.INIT('hfb00)
	) name2298 (
		_w8053_,
		_w8056_,
		_w8052_,
		_w8064_,
		_w8125_
	);
	LUT4 #(
		.INIT('hd000)
	) name2299 (
		_w8052_,
		_w8123_,
		_w8121_,
		_w8125_,
		_w8126_
	);
	LUT4 #(
		.INIT('h0100)
	) name2300 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8127_
	);
	LUT4 #(
		.INIT('h00df)
	) name2301 (
		_w8055_,
		_w8054_,
		_w8056_,
		_w8052_,
		_w8128_
	);
	LUT3 #(
		.INIT('h04)
	) name2302 (
		_w8053_,
		_w8055_,
		_w8056_,
		_w8129_
	);
	LUT4 #(
		.INIT('hff3b)
	) name2303 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8130_
	);
	LUT4 #(
		.INIT('he2f3)
	) name2304 (
		_w8059_,
		_w8052_,
		_w8127_,
		_w8130_,
		_w8131_
	);
	LUT4 #(
		.INIT('h8000)
	) name2305 (
		_w8055_,
		_w8054_,
		_w8056_,
		_w8052_,
		_w8132_
	);
	LUT4 #(
		.INIT('h00fb)
	) name2306 (
		_w8053_,
		_w8054_,
		_w8056_,
		_w8064_,
		_w8133_
	);
	LUT3 #(
		.INIT('h10)
	) name2307 (
		_w8066_,
		_w8132_,
		_w8133_,
		_w8134_
	);
	LUT3 #(
		.INIT('h45)
	) name2308 (
		_w8126_,
		_w8131_,
		_w8134_,
		_w8135_
	);
	LUT3 #(
		.INIT('h56)
	) name2309 (
		\u2_L10_reg[8]/NET0131 ,
		_w8120_,
		_w8135_,
		_w8136_
	);
	LUT4 #(
		.INIT('hddbd)
	) name2310 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8137_
	);
	LUT4 #(
		.INIT('hefe7)
	) name2311 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8138_
	);
	LUT4 #(
		.INIT('hc480)
	) name2312 (
		_w7836_,
		_w8004_,
		_w8138_,
		_w8137_,
		_w8139_
	);
	LUT2 #(
		.INIT('h2)
	) name2313 (
		_w7835_,
		_w8139_,
		_w8140_
	);
	LUT4 #(
		.INIT('hcf21)
	) name2314 (
		_w7842_,
		_w7839_,
		_w7836_,
		_w7837_,
		_w8141_
	);
	LUT2 #(
		.INIT('h2)
	) name2315 (
		_w7838_,
		_w8141_,
		_w8142_
	);
	LUT4 #(
		.INIT('h0040)
	) name2316 (
		_w7838_,
		_w7842_,
		_w7836_,
		_w7837_,
		_w8143_
	);
	LUT3 #(
		.INIT('h02)
	) name2317 (
		_w7859_,
		_w7850_,
		_w8143_,
		_w8144_
	);
	LUT3 #(
		.INIT('h45)
	) name2318 (
		_w7835_,
		_w8142_,
		_w8144_,
		_w8145_
	);
	LUT4 #(
		.INIT('h7bfe)
	) name2319 (
		_w7838_,
		_w7842_,
		_w7839_,
		_w7837_,
		_w8146_
	);
	LUT2 #(
		.INIT('h1)
	) name2320 (
		_w7836_,
		_w8146_,
		_w8147_
	);
	LUT3 #(
		.INIT('h13)
	) name2321 (
		_w7844_,
		_w7855_,
		_w7867_,
		_w8148_
	);
	LUT2 #(
		.INIT('h4)
	) name2322 (
		_w8147_,
		_w8148_,
		_w8149_
	);
	LUT4 #(
		.INIT('h5655)
	) name2323 (
		\u2_L10_reg[10]/NET0131 ,
		_w8140_,
		_w8145_,
		_w8149_,
		_w8150_
	);
	LUT4 #(
		.INIT('h0010)
	) name2324 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8151_
	);
	LUT2 #(
		.INIT('h1)
	) name2325 (
		_w7773_,
		_w8151_,
		_w8152_
	);
	LUT4 #(
		.INIT('h0104)
	) name2326 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8153_
	);
	LUT3 #(
		.INIT('hc4)
	) name2327 (
		_w7777_,
		_w7774_,
		_w7778_,
		_w8154_
	);
	LUT3 #(
		.INIT('h31)
	) name2328 (
		_w7796_,
		_w8153_,
		_w8154_,
		_w8155_
	);
	LUT3 #(
		.INIT('h1d)
	) name2329 (
		_w7774_,
		_w7778_,
		_w7775_,
		_w8156_
	);
	LUT3 #(
		.INIT('h21)
	) name2330 (
		_w7777_,
		_w7774_,
		_w7778_,
		_w8157_
	);
	LUT3 #(
		.INIT('h0d)
	) name2331 (
		_w7785_,
		_w8156_,
		_w8157_,
		_w8158_
	);
	LUT3 #(
		.INIT('h80)
	) name2332 (
		_w8152_,
		_w8155_,
		_w8158_,
		_w8159_
	);
	LUT4 #(
		.INIT('h0020)
	) name2333 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8160_
	);
	LUT4 #(
		.INIT('h0002)
	) name2334 (
		_w7773_,
		_w7800_,
		_w7779_,
		_w8160_,
		_w8161_
	);
	LUT3 #(
		.INIT('h0e)
	) name2335 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w8162_
	);
	LUT4 #(
		.INIT('h888c)
	) name2336 (
		_w7776_,
		_w7774_,
		_w7778_,
		_w7775_,
		_w8163_
	);
	LUT3 #(
		.INIT('hb9)
	) name2337 (
		_w7777_,
		_w7776_,
		_w7774_,
		_w8164_
	);
	LUT4 #(
		.INIT('hcf45)
	) name2338 (
		_w7786_,
		_w8162_,
		_w8163_,
		_w8164_,
		_w8165_
	);
	LUT2 #(
		.INIT('h8)
	) name2339 (
		_w8161_,
		_w8165_,
		_w8166_
	);
	LUT3 #(
		.INIT('ha9)
	) name2340 (
		\u2_L10_reg[12]/NET0131 ,
		_w8159_,
		_w8166_,
		_w8167_
	);
	LUT4 #(
		.INIT('h9ed3)
	) name2341 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8168_
	);
	LUT4 #(
		.INIT('h77af)
	) name2342 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8169_
	);
	LUT4 #(
		.INIT('h77ac)
	) name2343 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8170_
	);
	LUT4 #(
		.INIT('h0810)
	) name2344 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8171_
	);
	LUT4 #(
		.INIT('h0d08)
	) name2345 (
		_w8052_,
		_w8170_,
		_w8171_,
		_w8168_,
		_w8172_
	);
	LUT2 #(
		.INIT('h1)
	) name2346 (
		_w8064_,
		_w8172_,
		_w8173_
	);
	LUT4 #(
		.INIT('h1000)
	) name2347 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8174_
	);
	LUT4 #(
		.INIT('hedff)
	) name2348 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8175_
	);
	LUT4 #(
		.INIT('h0400)
	) name2349 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8176_
	);
	LUT4 #(
		.INIT('h0700)
	) name2350 (
		_w8057_,
		_w8075_,
		_w8176_,
		_w8175_,
		_w8177_
	);
	LUT3 #(
		.INIT('hf6)
	) name2351 (
		_w8055_,
		_w8054_,
		_w8056_,
		_w8178_
	);
	LUT4 #(
		.INIT('hea00)
	) name2352 (
		_w8055_,
		_w8054_,
		_w8056_,
		_w8052_,
		_w8179_
	);
	LUT4 #(
		.INIT('h31f5)
	) name2353 (
		_w8124_,
		_w8169_,
		_w8178_,
		_w8179_,
		_w8180_
	);
	LUT4 #(
		.INIT('heffd)
	) name2354 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8181_
	);
	LUT3 #(
		.INIT('he4)
	) name2355 (
		_w8052_,
		_w8121_,
		_w8181_,
		_w8182_
	);
	LUT4 #(
		.INIT('hd500)
	) name2356 (
		_w8064_,
		_w8177_,
		_w8180_,
		_w8182_,
		_w8183_
	);
	LUT3 #(
		.INIT('h65)
	) name2357 (
		\u2_L10_reg[14]/NET0131 ,
		_w8173_,
		_w8183_,
		_w8184_
	);
	LUT3 #(
		.INIT('h01)
	) name2358 (
		_w7875_,
		_w7873_,
		_w7876_,
		_w8185_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2359 (
		_w7872_,
		_w7874_,
		_w7875_,
		_w7876_,
		_w8186_
	);
	LUT4 #(
		.INIT('h5515)
	) name2360 (
		_w7872_,
		_w7874_,
		_w7875_,
		_w7873_,
		_w8187_
	);
	LUT4 #(
		.INIT('h8acf)
	) name2361 (
		_w7890_,
		_w8185_,
		_w8186_,
		_w8187_,
		_w8188_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name2362 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8189_
	);
	LUT4 #(
		.INIT('h0010)
	) name2363 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8190_
	);
	LUT4 #(
		.INIT('h0010)
	) name2364 (
		_w7879_,
		_w7880_,
		_w8189_,
		_w8190_,
		_w8191_
	);
	LUT3 #(
		.INIT('h8a)
	) name2365 (
		_w7871_,
		_w8188_,
		_w8191_,
		_w8192_
	);
	LUT4 #(
		.INIT('hebed)
	) name2366 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8193_
	);
	LUT4 #(
		.INIT('h0313)
	) name2367 (
		_w7871_,
		_w7872_,
		_w8189_,
		_w8193_,
		_w8194_
	);
	LUT4 #(
		.INIT('hf6d6)
	) name2368 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8195_
	);
	LUT2 #(
		.INIT('h2)
	) name2369 (
		_w7872_,
		_w8195_,
		_w8196_
	);
	LUT3 #(
		.INIT('hb0)
	) name2370 (
		_w7875_,
		_w7873_,
		_w7876_,
		_w8197_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w7872_,
		_w7873_,
		_w8198_
	);
	LUT3 #(
		.INIT('h04)
	) name2372 (
		_w7874_,
		_w7875_,
		_w7876_,
		_w8199_
	);
	LUT4 #(
		.INIT('h7077)
	) name2373 (
		_w8101_,
		_w8197_,
		_w8198_,
		_w8199_,
		_w8200_
	);
	LUT4 #(
		.INIT('h2322)
	) name2374 (
		_w7871_,
		_w8194_,
		_w8196_,
		_w8200_,
		_w8201_
	);
	LUT3 #(
		.INIT('h9a)
	) name2375 (
		\u2_L10_reg[13]/NET0131 ,
		_w8192_,
		_w8201_,
		_w8202_
	);
	LUT4 #(
		.INIT('h5f4f)
	) name2376 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8203_
	);
	LUT4 #(
		.INIT('h5a4f)
	) name2377 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8204_
	);
	LUT4 #(
		.INIT('h0002)
	) name2378 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8205_
	);
	LUT4 #(
		.INIT('h3302)
	) name2379 (
		_w7916_,
		_w7915_,
		_w8204_,
		_w8205_,
		_w8206_
	);
	LUT3 #(
		.INIT('h4b)
	) name2380 (
		_w7917_,
		_w7919_,
		_w7921_,
		_w8207_
	);
	LUT4 #(
		.INIT('h1041)
	) name2381 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8208_
	);
	LUT4 #(
		.INIT('h00f7)
	) name2382 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7916_,
		_w8209_
	);
	LUT2 #(
		.INIT('h4)
	) name2383 (
		_w8208_,
		_w8209_,
		_w8210_
	);
	LUT3 #(
		.INIT('h02)
	) name2384 (
		_w7916_,
		_w7924_,
		_w8028_,
		_w8211_
	);
	LUT2 #(
		.INIT('h1)
	) name2385 (
		_w8210_,
		_w8211_,
		_w8212_
	);
	LUT3 #(
		.INIT('h20)
	) name2386 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w8213_
	);
	LUT4 #(
		.INIT('h0020)
	) name2387 (
		_w7917_,
		_w7919_,
		_w7921_,
		_w7916_,
		_w8214_
	);
	LUT3 #(
		.INIT('h01)
	) name2388 (
		_w8025_,
		_w8214_,
		_w8213_,
		_w8215_
	);
	LUT4 #(
		.INIT('h0100)
	) name2389 (
		_w7918_,
		_w7919_,
		_w7921_,
		_w7916_,
		_w8216_
	);
	LUT2 #(
		.INIT('h1)
	) name2390 (
		_w7938_,
		_w8216_,
		_w8217_
	);
	LUT4 #(
		.INIT('h0002)
	) name2391 (
		_w7918_,
		_w7919_,
		_w7916_,
		_w7915_,
		_w8218_
	);
	LUT4 #(
		.INIT('h00d5)
	) name2392 (
		_w7915_,
		_w8215_,
		_w8217_,
		_w8218_,
		_w8219_
	);
	LUT4 #(
		.INIT('h5655)
	) name2393 (
		\u2_L10_reg[15]/NET0131 ,
		_w8206_,
		_w8212_,
		_w8219_,
		_w8220_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2394 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7916_,
		_w8221_
	);
	LUT2 #(
		.INIT('h8)
	) name2395 (
		_w8207_,
		_w8221_,
		_w8222_
	);
	LUT4 #(
		.INIT('h0080)
	) name2396 (
		_w7918_,
		_w7917_,
		_w7921_,
		_w7916_,
		_w8223_
	);
	LUT3 #(
		.INIT('h01)
	) name2397 (
		_w7940_,
		_w8013_,
		_w8223_,
		_w8224_
	);
	LUT3 #(
		.INIT('h45)
	) name2398 (
		_w7915_,
		_w8222_,
		_w8224_,
		_w8225_
	);
	LUT4 #(
		.INIT('hae5e)
	) name2399 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8226_
	);
	LUT2 #(
		.INIT('h1)
	) name2400 (
		_w7916_,
		_w8226_,
		_w8227_
	);
	LUT3 #(
		.INIT('hd0)
	) name2401 (
		_w7918_,
		_w7921_,
		_w7916_,
		_w8228_
	);
	LUT4 #(
		.INIT('hbcf7)
	) name2402 (
		_w7918_,
		_w7917_,
		_w7919_,
		_w7921_,
		_w8229_
	);
	LUT3 #(
		.INIT('hb0)
	) name2403 (
		_w8203_,
		_w8228_,
		_w8229_,
		_w8230_
	);
	LUT3 #(
		.INIT('h8a)
	) name2404 (
		_w7915_,
		_w8227_,
		_w8230_,
		_w8231_
	);
	LUT2 #(
		.INIT('h1)
	) name2405 (
		_w7916_,
		_w7939_,
		_w8232_
	);
	LUT4 #(
		.INIT('h0200)
	) name2406 (
		_w7917_,
		_w7919_,
		_w7921_,
		_w7916_,
		_w8233_
	);
	LUT3 #(
		.INIT('h07)
	) name2407 (
		_w7928_,
		_w7944_,
		_w8233_,
		_w8234_
	);
	LUT2 #(
		.INIT('h4)
	) name2408 (
		_w8232_,
		_w8234_,
		_w8235_
	);
	LUT4 #(
		.INIT('h5655)
	) name2409 (
		\u2_L10_reg[27]/NET0131 ,
		_w8231_,
		_w8225_,
		_w8235_,
		_w8236_
	);
	LUT4 #(
		.INIT('h0006)
	) name2410 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8237_
	);
	LUT4 #(
		.INIT('h0800)
	) name2411 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8238_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2412 (
		_w7777_,
		_w7776_,
		_w7774_,
		_w7778_,
		_w8239_
	);
	LUT3 #(
		.INIT('h10)
	) name2413 (
		_w8237_,
		_w8238_,
		_w8239_,
		_w8240_
	);
	LUT4 #(
		.INIT('h01a1)
	) name2414 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8241_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name2415 (
		_w7777_,
		_w7776_,
		_w7774_,
		_w7775_,
		_w8242_
	);
	LUT2 #(
		.INIT('h4)
	) name2416 (
		_w8241_,
		_w8242_,
		_w8243_
	);
	LUT4 #(
		.INIT('h4000)
	) name2417 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8244_
	);
	LUT4 #(
		.INIT('haa02)
	) name2418 (
		_w7773_,
		_w8240_,
		_w8243_,
		_w8244_,
		_w8245_
	);
	LUT3 #(
		.INIT('h04)
	) name2419 (
		_w7777_,
		_w7776_,
		_w7775_,
		_w8246_
	);
	LUT2 #(
		.INIT('h2)
	) name2420 (
		_w8157_,
		_w8246_,
		_w8247_
	);
	LUT4 #(
		.INIT('h0240)
	) name2421 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8248_
	);
	LUT4 #(
		.INIT('h9000)
	) name2422 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8249_
	);
	LUT3 #(
		.INIT('hd8)
	) name2423 (
		_w7777_,
		_w7778_,
		_w7775_,
		_w8250_
	);
	LUT4 #(
		.INIT('h0301)
	) name2424 (
		_w7783_,
		_w8249_,
		_w8248_,
		_w8250_,
		_w8251_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2425 (
		_w7777_,
		_w7776_,
		_w7774_,
		_w7778_,
		_w8252_
	);
	LUT4 #(
		.INIT('h135f)
	) name2426 (
		_w7774_,
		_w7797_,
		_w7787_,
		_w8252_,
		_w8253_
	);
	LUT4 #(
		.INIT('hba00)
	) name2427 (
		_w7773_,
		_w8247_,
		_w8251_,
		_w8253_,
		_w8254_
	);
	LUT3 #(
		.INIT('h65)
	) name2428 (
		\u2_L10_reg[32]/NET0131 ,
		_w8245_,
		_w8254_,
		_w8255_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2429 (
		_w8055_,
		_w8054_,
		_w8056_,
		_w8052_,
		_w8256_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2430 (
		_w8061_,
		_w8128_,
		_w8129_,
		_w8256_,
		_w8257_
	);
	LUT4 #(
		.INIT('h080a)
	) name2431 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8258_
	);
	LUT2 #(
		.INIT('h1)
	) name2432 (
		_w8064_,
		_w8258_,
		_w8259_
	);
	LUT4 #(
		.INIT('hbbcf)
	) name2433 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8260_
	);
	LUT2 #(
		.INIT('h2)
	) name2434 (
		_w8052_,
		_w8260_,
		_w8261_
	);
	LUT4 #(
		.INIT('h0008)
	) name2435 (
		_w8055_,
		_w8054_,
		_w8056_,
		_w8052_,
		_w8262_
	);
	LUT4 #(
		.INIT('h0004)
	) name2436 (
		_w8074_,
		_w8064_,
		_w8114_,
		_w8262_,
		_w8263_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2437 (
		_w8257_,
		_w8259_,
		_w8261_,
		_w8263_,
		_w8264_
	);
	LUT3 #(
		.INIT('h02)
	) name2438 (
		_w8052_,
		_w8116_,
		_w8127_,
		_w8265_
	);
	LUT4 #(
		.INIT('h0800)
	) name2439 (
		_w8053_,
		_w8055_,
		_w8054_,
		_w8056_,
		_w8266_
	);
	LUT4 #(
		.INIT('h0001)
	) name2440 (
		_w8052_,
		_w8122_,
		_w8174_,
		_w8266_,
		_w8267_
	);
	LUT2 #(
		.INIT('h1)
	) name2441 (
		_w8265_,
		_w8267_,
		_w8268_
	);
	LUT3 #(
		.INIT('h56)
	) name2442 (
		\u2_L10_reg[3]/NET0131 ,
		_w8264_,
		_w8268_,
		_w8269_
	);
	LUT4 #(
		.INIT('hc693)
	) name2443 (
		decrypt_pad,
		\u2_R10_reg[10]/NET0131 ,
		\u2_uk_K_r10_reg[25]/NET0131 ,
		\u2_uk_K_r10_reg[34]/NET0131 ,
		_w8270_
	);
	LUT4 #(
		.INIT('hc693)
	) name2444 (
		decrypt_pad,
		\u2_R10_reg[9]/NET0131 ,
		\u2_uk_K_r10_reg[17]/NET0131 ,
		\u2_uk_K_r10_reg[26]/NET0131 ,
		_w8271_
	);
	LUT4 #(
		.INIT('hc693)
	) name2445 (
		decrypt_pad,
		\u2_R10_reg[13]/NET0131 ,
		\u2_uk_K_r10_reg[54]/NET0131 ,
		\u2_uk_K_r10_reg[6]/NET0131 ,
		_w8272_
	);
	LUT3 #(
		.INIT('h20)
	) name2446 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8273_
	);
	LUT4 #(
		.INIT('hc693)
	) name2447 (
		decrypt_pad,
		\u2_R10_reg[8]/NET0131 ,
		\u2_uk_K_r10_reg[20]/NET0131 ,
		\u2_uk_K_r10_reg[54]/NET0131 ,
		_w8274_
	);
	LUT2 #(
		.INIT('h1)
	) name2448 (
		_w8270_,
		_w8271_,
		_w8275_
	);
	LUT4 #(
		.INIT('h0001)
	) name2449 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8276_
	);
	LUT4 #(
		.INIT('hdfde)
	) name2450 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8277_
	);
	LUT4 #(
		.INIT('hc693)
	) name2451 (
		decrypt_pad,
		\u2_R10_reg[11]/NET0131 ,
		\u2_uk_K_r10_reg[26]/NET0131 ,
		\u2_uk_K_r10_reg[3]/NET0131 ,
		_w8278_
	);
	LUT2 #(
		.INIT('h4)
	) name2452 (
		_w8277_,
		_w8278_,
		_w8279_
	);
	LUT2 #(
		.INIT('h6)
	) name2453 (
		_w8272_,
		_w8274_,
		_w8280_
	);
	LUT4 #(
		.INIT('hc04c)
	) name2454 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8281_
	);
	LUT3 #(
		.INIT('he0)
	) name2455 (
		_w8271_,
		_w8272_,
		_w8278_,
		_w8282_
	);
	LUT2 #(
		.INIT('h4)
	) name2456 (
		_w8281_,
		_w8282_,
		_w8283_
	);
	LUT2 #(
		.INIT('h2)
	) name2457 (
		_w8270_,
		_w8274_,
		_w8284_
	);
	LUT4 #(
		.INIT('h3cbf)
	) name2458 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8285_
	);
	LUT4 #(
		.INIT('h0008)
	) name2459 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8286_
	);
	LUT4 #(
		.INIT('hc963)
	) name2460 (
		decrypt_pad,
		\u2_R10_reg[12]/NET0131 ,
		\u2_uk_K_r10_reg[18]/NET0131 ,
		\u2_uk_K_r10_reg[41]/NET0131 ,
		_w8287_
	);
	LUT4 #(
		.INIT('h3200)
	) name2461 (
		_w8278_,
		_w8286_,
		_w8285_,
		_w8287_,
		_w8288_
	);
	LUT2 #(
		.INIT('h4)
	) name2462 (
		_w8283_,
		_w8288_,
		_w8289_
	);
	LUT4 #(
		.INIT('h2002)
	) name2463 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8290_
	);
	LUT3 #(
		.INIT('h08)
	) name2464 (
		_w8271_,
		_w8272_,
		_w8278_,
		_w8291_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		_w8270_,
		_w8274_,
		_w8292_
	);
	LUT4 #(
		.INIT('h0800)
	) name2466 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8293_
	);
	LUT4 #(
		.INIT('h0013)
	) name2467 (
		_w8284_,
		_w8287_,
		_w8291_,
		_w8293_,
		_w8294_
	);
	LUT3 #(
		.INIT('h46)
	) name2468 (
		_w8272_,
		_w8274_,
		_w8278_,
		_w8295_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		_w8275_,
		_w8295_,
		_w8296_
	);
	LUT3 #(
		.INIT('heb)
	) name2470 (
		_w8270_,
		_w8271_,
		_w8295_,
		_w8297_
	);
	LUT3 #(
		.INIT('h40)
	) name2471 (
		_w8290_,
		_w8294_,
		_w8297_,
		_w8298_
	);
	LUT4 #(
		.INIT('h6665)
	) name2472 (
		\u2_L10_reg[6]/NET0131 ,
		_w8279_,
		_w8289_,
		_w8298_,
		_w8299_
	);
	LUT4 #(
		.INIT('h8b9c)
	) name2473 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8300_
	);
	LUT4 #(
		.INIT('h6800)
	) name2474 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8301_
	);
	LUT4 #(
		.INIT('h0098)
	) name2475 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8302_
	);
	LUT4 #(
		.INIT('h040e)
	) name2476 (
		_w7774_,
		_w8300_,
		_w8301_,
		_w8302_,
		_w8303_
	);
	LUT4 #(
		.INIT('h6899)
	) name2477 (
		_w7777_,
		_w7776_,
		_w7778_,
		_w7775_,
		_w8304_
	);
	LUT4 #(
		.INIT('h2301)
	) name2478 (
		_w7774_,
		_w7791_,
		_w8302_,
		_w8304_,
		_w8305_
	);
	LUT3 #(
		.INIT('h27)
	) name2479 (
		_w7774_,
		_w7791_,
		_w8301_,
		_w8306_
	);
	LUT4 #(
		.INIT('hd800)
	) name2480 (
		_w7773_,
		_w8303_,
		_w8305_,
		_w8306_,
		_w8307_
	);
	LUT2 #(
		.INIT('h9)
	) name2481 (
		\u2_L10_reg[7]/NET0131 ,
		_w8307_,
		_w8308_
	);
	LUT3 #(
		.INIT('hb7)
	) name2482 (
		_w7744_,
		_w7745_,
		_w7746_,
		_w8309_
	);
	LUT2 #(
		.INIT('h2)
	) name2483 (
		_w7757_,
		_w8309_,
		_w8310_
	);
	LUT4 #(
		.INIT('h8228)
	) name2484 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w8311_
	);
	LUT3 #(
		.INIT('he6)
	) name2485 (
		_w7745_,
		_w7742_,
		_w7746_,
		_w8312_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2486 (
		_w7741_,
		_w7759_,
		_w7967_,
		_w8312_,
		_w8313_
	);
	LUT4 #(
		.INIT('hd3c3)
	) name2487 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w8314_
	);
	LUT2 #(
		.INIT('h2)
	) name2488 (
		_w7743_,
		_w8314_,
		_w8315_
	);
	LUT4 #(
		.INIT('h0141)
	) name2489 (
		_w7743_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w8316_
	);
	LUT4 #(
		.INIT('h0802)
	) name2490 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w8317_
	);
	LUT4 #(
		.INIT('h4000)
	) name2491 (
		_w7744_,
		_w7745_,
		_w7742_,
		_w7746_,
		_w8318_
	);
	LUT4 #(
		.INIT('h0001)
	) name2492 (
		_w7741_,
		_w8318_,
		_w8317_,
		_w8316_,
		_w8319_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2493 (
		_w8311_,
		_w8313_,
		_w8315_,
		_w8319_,
		_w8320_
	);
	LUT3 #(
		.INIT('h56)
	) name2494 (
		\u2_L10_reg[9]/NET0131 ,
		_w8310_,
		_w8320_,
		_w8321_
	);
	LUT4 #(
		.INIT('h0a20)
	) name2495 (
		_w7872_,
		_w7874_,
		_w7875_,
		_w7873_,
		_w8322_
	);
	LUT4 #(
		.INIT('hfd75)
	) name2496 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8323_
	);
	LUT4 #(
		.INIT('h0032)
	) name2497 (
		_w7872_,
		_w7891_,
		_w8323_,
		_w8322_,
		_w8324_
	);
	LUT2 #(
		.INIT('h2)
	) name2498 (
		_w7871_,
		_w8324_,
		_w8325_
	);
	LUT4 #(
		.INIT('h8000)
	) name2499 (
		_w7872_,
		_w7874_,
		_w7875_,
		_w7873_,
		_w8326_
	);
	LUT3 #(
		.INIT('h01)
	) name2500 (
		_w7882_,
		_w8185_,
		_w8326_,
		_w8327_
	);
	LUT4 #(
		.INIT('h1003)
	) name2501 (
		_w7872_,
		_w7874_,
		_w7873_,
		_w7876_,
		_w8328_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		_w8106_,
		_w8328_,
		_w8329_
	);
	LUT4 #(
		.INIT('h1000)
	) name2503 (
		_w7872_,
		_w7874_,
		_w7875_,
		_w7873_,
		_w8330_
	);
	LUT4 #(
		.INIT('h77ef)
	) name2504 (
		_w7874_,
		_w7875_,
		_w7873_,
		_w7876_,
		_w8331_
	);
	LUT3 #(
		.INIT('h31)
	) name2505 (
		_w7872_,
		_w8330_,
		_w8331_,
		_w8332_
	);
	LUT4 #(
		.INIT('hea00)
	) name2506 (
		_w7871_,
		_w8327_,
		_w8329_,
		_w8332_,
		_w8333_
	);
	LUT3 #(
		.INIT('h65)
	) name2507 (
		\u2_L10_reg[18]/P0001 ,
		_w8325_,
		_w8333_,
		_w8334_
	);
	LUT4 #(
		.INIT('h1001)
	) name2508 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8335_
	);
	LUT4 #(
		.INIT('he35e)
	) name2509 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8336_
	);
	LUT3 #(
		.INIT('h32)
	) name2510 (
		_w8278_,
		_w8287_,
		_w8336_,
		_w8337_
	);
	LUT2 #(
		.INIT('h4)
	) name2511 (
		_w8270_,
		_w8278_,
		_w8338_
	);
	LUT3 #(
		.INIT('hae)
	) name2512 (
		_w8271_,
		_w8272_,
		_w8274_,
		_w8339_
	);
	LUT3 #(
		.INIT('ha2)
	) name2513 (
		_w8287_,
		_w8338_,
		_w8339_,
		_w8340_
	);
	LUT3 #(
		.INIT('he0)
	) name2514 (
		_w8272_,
		_w8274_,
		_w8278_,
		_w8341_
	);
	LUT3 #(
		.INIT('h8a)
	) name2515 (
		_w8270_,
		_w8271_,
		_w8274_,
		_w8342_
	);
	LUT3 #(
		.INIT('h0e)
	) name2516 (
		_w8270_,
		_w8271_,
		_w8278_,
		_w8343_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name2517 (
		_w8280_,
		_w8341_,
		_w8342_,
		_w8343_,
		_w8344_
	);
	LUT4 #(
		.INIT('h2333)
	) name2518 (
		_w8296_,
		_w8337_,
		_w8340_,
		_w8344_,
		_w8345_
	);
	LUT3 #(
		.INIT('h20)
	) name2519 (
		_w8270_,
		_w8271_,
		_w8274_,
		_w8346_
	);
	LUT4 #(
		.INIT('hdda1)
	) name2520 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8347_
	);
	LUT4 #(
		.INIT('h0200)
	) name2521 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8348_
	);
	LUT4 #(
		.INIT('h3302)
	) name2522 (
		_w8278_,
		_w8287_,
		_w8347_,
		_w8348_,
		_w8349_
	);
	LUT3 #(
		.INIT('h27)
	) name2523 (
		_w8271_,
		_w8272_,
		_w8274_,
		_w8350_
	);
	LUT4 #(
		.INIT('h1500)
	) name2524 (
		_w8270_,
		_w8272_,
		_w8274_,
		_w8278_,
		_w8351_
	);
	LUT4 #(
		.INIT('h7077)
	) name2525 (
		_w8291_,
		_w8292_,
		_w8350_,
		_w8351_,
		_w8352_
	);
	LUT2 #(
		.INIT('h4)
	) name2526 (
		_w8349_,
		_w8352_,
		_w8353_
	);
	LUT3 #(
		.INIT('h65)
	) name2527 (
		\u2_L10_reg[24]/NET0131 ,
		_w8345_,
		_w8353_,
		_w8354_
	);
	LUT4 #(
		.INIT('hfea5)
	) name2528 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8355_
	);
	LUT4 #(
		.INIT('h51f3)
	) name2529 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8356_
	);
	LUT3 #(
		.INIT('h08)
	) name2530 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8357_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name2531 (
		_w8287_,
		_w8357_,
		_w8355_,
		_w8356_,
		_w8358_
	);
	LUT2 #(
		.INIT('h2)
	) name2532 (
		_w8278_,
		_w8358_,
		_w8359_
	);
	LUT4 #(
		.INIT('h0888)
	) name2533 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8360_
	);
	LUT4 #(
		.INIT('h55f3)
	) name2534 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8361_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name2535 (
		_w8278_,
		_w8287_,
		_w8360_,
		_w8361_,
		_w8362_
	);
	LUT3 #(
		.INIT('h07)
	) name2536 (
		_w8270_,
		_w8274_,
		_w8278_,
		_w8363_
	);
	LUT4 #(
		.INIT('h4544)
	) name2537 (
		_w8287_,
		_w8335_,
		_w8350_,
		_w8363_,
		_w8364_
	);
	LUT4 #(
		.INIT('h0008)
	) name2538 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8278_,
		_w8365_
	);
	LUT3 #(
		.INIT('h8d)
	) name2539 (
		_w8274_,
		_w8278_,
		_w8287_,
		_w8366_
	);
	LUT3 #(
		.INIT('h13)
	) name2540 (
		_w8273_,
		_w8365_,
		_w8366_,
		_w8367_
	);
	LUT3 #(
		.INIT('h10)
	) name2541 (
		_w8362_,
		_w8364_,
		_w8367_,
		_w8368_
	);
	LUT3 #(
		.INIT('h9a)
	) name2542 (
		\u2_L10_reg[30]/NET0131 ,
		_w8359_,
		_w8368_,
		_w8369_
	);
	LUT4 #(
		.INIT('h696b)
	) name2543 (
		_w8271_,
		_w8272_,
		_w8274_,
		_w8278_,
		_w8370_
	);
	LUT4 #(
		.INIT('h0080)
	) name2544 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8371_
	);
	LUT4 #(
		.INIT('h0012)
	) name2545 (
		_w8270_,
		_w8272_,
		_w8274_,
		_w8278_,
		_w8372_
	);
	LUT4 #(
		.INIT('h0032)
	) name2546 (
		_w8270_,
		_w8371_,
		_w8370_,
		_w8372_,
		_w8373_
	);
	LUT2 #(
		.INIT('h2)
	) name2547 (
		_w8287_,
		_w8373_,
		_w8374_
	);
	LUT4 #(
		.INIT('h3fca)
	) name2548 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8375_
	);
	LUT4 #(
		.INIT('h5051)
	) name2549 (
		_w8278_,
		_w8287_,
		_w8346_,
		_w8375_,
		_w8376_
	);
	LUT4 #(
		.INIT('hf7fd)
	) name2550 (
		_w8270_,
		_w8271_,
		_w8272_,
		_w8274_,
		_w8377_
	);
	LUT2 #(
		.INIT('h2)
	) name2551 (
		_w8278_,
		_w8377_,
		_w8378_
	);
	LUT4 #(
		.INIT('h6800)
	) name2552 (
		_w8271_,
		_w8272_,
		_w8274_,
		_w8278_,
		_w8379_
	);
	LUT3 #(
		.INIT('h32)
	) name2553 (
		_w8276_,
		_w8287_,
		_w8379_,
		_w8380_
	);
	LUT3 #(
		.INIT('h01)
	) name2554 (
		_w8376_,
		_w8378_,
		_w8380_,
		_w8381_
	);
	LUT3 #(
		.INIT('h65)
	) name2555 (
		\u2_L10_reg[16]/NET0131 ,
		_w8374_,
		_w8381_,
		_w8382_
	);
	LUT4 #(
		.INIT('hc963)
	) name2556 (
		decrypt_pad,
		\u2_R9_reg[28]/NET0131 ,
		\u2_uk_K_r9_reg[31]/P0001 ,
		\u2_uk_K_r9_reg[50]/NET0131 ,
		_w8383_
	);
	LUT4 #(
		.INIT('hc963)
	) name2557 (
		decrypt_pad,
		\u2_R9_reg[27]/NET0131 ,
		\u2_uk_K_r9_reg[16]/NET0131 ,
		\u2_uk_K_r9_reg[8]/NET0131 ,
		_w8384_
	);
	LUT4 #(
		.INIT('hc693)
	) name2558 (
		decrypt_pad,
		\u2_R9_reg[26]/NET0131 ,
		\u2_uk_K_r9_reg[30]/NET0131 ,
		\u2_uk_K_r9_reg[7]/NET0131 ,
		_w8385_
	);
	LUT4 #(
		.INIT('hc693)
	) name2559 (
		decrypt_pad,
		\u2_R9_reg[24]/NET0131 ,
		\u2_uk_K_r9_reg[38]/NET0131 ,
		\u2_uk_K_r9_reg[42]/NET0131 ,
		_w8386_
	);
	LUT4 #(
		.INIT('hc693)
	) name2560 (
		decrypt_pad,
		\u2_R9_reg[25]/NET0131 ,
		\u2_uk_K_r9_reg[14]/NET0131 ,
		\u2_uk_K_r9_reg[22]/NET0131 ,
		_w8387_
	);
	LUT4 #(
		.INIT('hc693)
	) name2561 (
		decrypt_pad,
		\u2_R9_reg[29]/NET0131 ,
		\u2_uk_K_r9_reg[42]/NET0131 ,
		\u2_uk_K_r9_reg[50]/NET0131 ,
		_w8388_
	);
	LUT4 #(
		.INIT('h1000)
	) name2562 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8389_
	);
	LUT2 #(
		.INIT('h4)
	) name2563 (
		_w8386_,
		_w8388_,
		_w8390_
	);
	LUT4 #(
		.INIT('he3ff)
	) name2564 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8391_
	);
	LUT2 #(
		.INIT('h1)
	) name2565 (
		_w8384_,
		_w8391_,
		_w8392_
	);
	LUT2 #(
		.INIT('h6)
	) name2566 (
		_w8385_,
		_w8387_,
		_w8393_
	);
	LUT2 #(
		.INIT('h8)
	) name2567 (
		_w8384_,
		_w8386_,
		_w8394_
	);
	LUT4 #(
		.INIT('hc080)
	) name2568 (
		_w8385_,
		_w8384_,
		_w8386_,
		_w8388_,
		_w8395_
	);
	LUT4 #(
		.INIT('h0200)
	) name2569 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8396_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name2570 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8397_
	);
	LUT3 #(
		.INIT('h70)
	) name2571 (
		_w8393_,
		_w8395_,
		_w8397_,
		_w8398_
	);
	LUT3 #(
		.INIT('h8a)
	) name2572 (
		_w8383_,
		_w8392_,
		_w8398_,
		_w8399_
	);
	LUT2 #(
		.INIT('h6)
	) name2573 (
		_w8385_,
		_w8386_,
		_w8400_
	);
	LUT4 #(
		.INIT('h0002)
	) name2574 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8401_
	);
	LUT4 #(
		.INIT('h5a2d)
	) name2575 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8402_
	);
	LUT4 #(
		.INIT('h1000)
	) name2576 (
		_w8385_,
		_w8387_,
		_w8384_,
		_w8386_,
		_w8403_
	);
	LUT4 #(
		.INIT('h8400)
	) name2577 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8404_
	);
	LUT4 #(
		.INIT('h0302)
	) name2578 (
		_w8384_,
		_w8403_,
		_w8404_,
		_w8402_,
		_w8405_
	);
	LUT4 #(
		.INIT('h0008)
	) name2579 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8406_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name2580 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8407_
	);
	LUT4 #(
		.INIT('hfdc7)
	) name2581 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8408_
	);
	LUT4 #(
		.INIT('h0010)
	) name2582 (
		_w8385_,
		_w8387_,
		_w8384_,
		_w8388_,
		_w8409_
	);
	LUT4 #(
		.INIT('h0804)
	) name2583 (
		_w8385_,
		_w8387_,
		_w8384_,
		_w8386_,
		_w8410_
	);
	LUT4 #(
		.INIT('h0031)
	) name2584 (
		_w8384_,
		_w8409_,
		_w8408_,
		_w8410_,
		_w8411_
	);
	LUT3 #(
		.INIT('he0)
	) name2585 (
		_w8405_,
		_w8383_,
		_w8411_,
		_w8412_
	);
	LUT3 #(
		.INIT('h65)
	) name2586 (
		\u2_L9_reg[22]/NET0131 ,
		_w8399_,
		_w8412_,
		_w8413_
	);
	LUT4 #(
		.INIT('hc693)
	) name2587 (
		decrypt_pad,
		\u2_R9_reg[3]/NET0131 ,
		\u2_uk_K_r9_reg[41]/NET0131 ,
		\u2_uk_K_r9_reg[47]/NET0131 ,
		_w8414_
	);
	LUT4 #(
		.INIT('hc693)
	) name2588 (
		decrypt_pad,
		\u2_R9_reg[4]/NET0131 ,
		\u2_uk_K_r9_reg[19]/NET0131 ,
		\u2_uk_K_r9_reg[25]/NET0131 ,
		_w8415_
	);
	LUT4 #(
		.INIT('hc963)
	) name2589 (
		decrypt_pad,
		\u2_R9_reg[2]/NET0131 ,
		\u2_uk_K_r9_reg[13]/NET0131 ,
		\u2_uk_K_r9_reg[32]/NET0131 ,
		_w8416_
	);
	LUT4 #(
		.INIT('hc693)
	) name2590 (
		decrypt_pad,
		\u2_R9_reg[5]/NET0131 ,
		\u2_uk_K_r9_reg[47]/NET0131 ,
		\u2_uk_K_r9_reg[53]/NET0131 ,
		_w8417_
	);
	LUT4 #(
		.INIT('hc693)
	) name2591 (
		decrypt_pad,
		\u2_R9_reg[1]/NET0131 ,
		\u2_uk_K_r9_reg[17]/NET0131 ,
		\u2_uk_K_r9_reg[55]/NET0131 ,
		_w8418_
	);
	LUT4 #(
		.INIT('hc963)
	) name2592 (
		decrypt_pad,
		\u2_R9_reg[32]/NET0131 ,
		\u2_uk_K_r9_reg[34]/NET0131 ,
		\u2_uk_K_r9_reg[53]/NET0131 ,
		_w8419_
	);
	LUT4 #(
		.INIT('heff4)
	) name2593 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8420_
	);
	LUT3 #(
		.INIT('h80)
	) name2594 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8421_
	);
	LUT4 #(
		.INIT('h7dbd)
	) name2595 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8422_
	);
	LUT4 #(
		.INIT('h0155)
	) name2596 (
		_w8414_,
		_w8415_,
		_w8420_,
		_w8422_,
		_w8423_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name2597 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8424_
	);
	LUT2 #(
		.INIT('h2)
	) name2598 (
		_w8414_,
		_w8424_,
		_w8425_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name2599 (
		_w8414_,
		_w8418_,
		_w8417_,
		_w8416_,
		_w8426_
	);
	LUT2 #(
		.INIT('h4)
	) name2600 (
		_w8426_,
		_w8419_,
		_w8427_
	);
	LUT2 #(
		.INIT('h2)
	) name2601 (
		_w8414_,
		_w8416_,
		_w8428_
	);
	LUT3 #(
		.INIT('hc4)
	) name2602 (
		_w8414_,
		_w8418_,
		_w8416_,
		_w8429_
	);
	LUT3 #(
		.INIT('h0e)
	) name2603 (
		_w8417_,
		_w8416_,
		_w8419_,
		_w8430_
	);
	LUT3 #(
		.INIT('hb0)
	) name2604 (
		_w8429_,
		_w8430_,
		_w8415_,
		_w8431_
	);
	LUT3 #(
		.INIT('h10)
	) name2605 (
		_w8427_,
		_w8425_,
		_w8431_,
		_w8432_
	);
	LUT4 #(
		.INIT('hd3ff)
	) name2606 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8433_
	);
	LUT2 #(
		.INIT('h2)
	) name2607 (
		_w8414_,
		_w8433_,
		_w8434_
	);
	LUT2 #(
		.INIT('h8)
	) name2608 (
		_w8414_,
		_w8416_,
		_w8435_
	);
	LUT4 #(
		.INIT('h0080)
	) name2609 (
		_w8414_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8436_
	);
	LUT4 #(
		.INIT('hff7c)
	) name2610 (
		_w8414_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8437_
	);
	LUT4 #(
		.INIT('h0400)
	) name2611 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8438_
	);
	LUT4 #(
		.INIT('h0031)
	) name2612 (
		_w8418_,
		_w8415_,
		_w8437_,
		_w8438_,
		_w8439_
	);
	LUT2 #(
		.INIT('h4)
	) name2613 (
		_w8434_,
		_w8439_,
		_w8440_
	);
	LUT4 #(
		.INIT('h0200)
	) name2614 (
		_w8414_,
		_w8418_,
		_w8416_,
		_w8419_,
		_w8441_
	);
	LUT3 #(
		.INIT('h01)
	) name2615 (
		_w8418_,
		_w8417_,
		_w8419_,
		_w8442_
	);
	LUT3 #(
		.INIT('h13)
	) name2616 (
		_w8435_,
		_w8441_,
		_w8442_,
		_w8443_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2617 (
		_w8432_,
		_w8440_,
		_w8423_,
		_w8443_,
		_w8444_
	);
	LUT2 #(
		.INIT('h9)
	) name2618 (
		\u2_L9_reg[31]/NET0131 ,
		_w8444_,
		_w8445_
	);
	LUT4 #(
		.INIT('hc693)
	) name2619 (
		decrypt_pad,
		\u2_R9_reg[24]/NET0131 ,
		\u2_uk_K_r9_reg[43]/NET0131 ,
		\u2_uk_K_r9_reg[51]/NET0131 ,
		_w8446_
	);
	LUT4 #(
		.INIT('hc693)
	) name2620 (
		decrypt_pad,
		\u2_R9_reg[20]/NET0131 ,
		\u2_uk_K_r9_reg[22]/NET0131 ,
		\u2_uk_K_r9_reg[30]/NET0131 ,
		_w8447_
	);
	LUT4 #(
		.INIT('hc693)
	) name2621 (
		decrypt_pad,
		\u2_R9_reg[22]/NET0131 ,
		\u2_uk_K_r9_reg[28]/NET0131 ,
		\u2_uk_K_r9_reg[36]/NET0131 ,
		_w8448_
	);
	LUT4 #(
		.INIT('hc963)
	) name2622 (
		decrypt_pad,
		\u2_R9_reg[21]/NET0131 ,
		\u2_uk_K_r9_reg[14]/NET0131 ,
		\u2_uk_K_r9_reg[37]/NET0131 ,
		_w8449_
	);
	LUT4 #(
		.INIT('hc693)
	) name2623 (
		decrypt_pad,
		\u2_R9_reg[23]/NET0131 ,
		\u2_uk_K_r9_reg[45]/NET0131 ,
		\u2_uk_K_r9_reg[49]/NET0131 ,
		_w8450_
	);
	LUT4 #(
		.INIT('h4155)
	) name2624 (
		_w8450_,
		_w8447_,
		_w8448_,
		_w8449_,
		_w8451_
	);
	LUT4 #(
		.INIT('hc963)
	) name2625 (
		decrypt_pad,
		\u2_R9_reg[25]/NET0131 ,
		\u2_uk_K_r9_reg[15]/NET0131 ,
		\u2_uk_K_r9_reg[7]/NET0131 ,
		_w8452_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2626 (
		_w8450_,
		_w8447_,
		_w8452_,
		_w8449_,
		_w8453_
	);
	LUT3 #(
		.INIT('he6)
	) name2627 (
		_w8447_,
		_w8448_,
		_w8449_,
		_w8454_
	);
	LUT3 #(
		.INIT('h13)
	) name2628 (
		_w8453_,
		_w8451_,
		_w8454_,
		_w8455_
	);
	LUT4 #(
		.INIT('h0080)
	) name2629 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8456_
	);
	LUT2 #(
		.INIT('h2)
	) name2630 (
		_w8447_,
		_w8452_,
		_w8457_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w8450_,
		_w8448_,
		_w8458_
	);
	LUT3 #(
		.INIT('hce)
	) name2632 (
		_w8450_,
		_w8448_,
		_w8449_,
		_w8459_
	);
	LUT3 #(
		.INIT('h31)
	) name2633 (
		_w8457_,
		_w8456_,
		_w8459_,
		_w8460_
	);
	LUT3 #(
		.INIT('h45)
	) name2634 (
		_w8446_,
		_w8455_,
		_w8460_,
		_w8461_
	);
	LUT4 #(
		.INIT('h0002)
	) name2635 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8462_
	);
	LUT4 #(
		.INIT('h27fd)
	) name2636 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8463_
	);
	LUT2 #(
		.INIT('h2)
	) name2637 (
		_w8450_,
		_w8463_,
		_w8464_
	);
	LUT4 #(
		.INIT('h0415)
	) name2638 (
		_w8450_,
		_w8447_,
		_w8452_,
		_w8449_,
		_w8465_
	);
	LUT4 #(
		.INIT('h0b07)
	) name2639 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8466_
	);
	LUT3 #(
		.INIT('h0e)
	) name2640 (
		_w8458_,
		_w8465_,
		_w8466_,
		_w8467_
	);
	LUT3 #(
		.INIT('he0)
	) name2641 (
		_w8464_,
		_w8467_,
		_w8446_,
		_w8468_
	);
	LUT4 #(
		.INIT('h5155)
	) name2642 (
		_w8450_,
		_w8447_,
		_w8452_,
		_w8449_,
		_w8469_
	);
	LUT3 #(
		.INIT('h01)
	) name2643 (
		_w8448_,
		_w8469_,
		_w8453_,
		_w8470_
	);
	LUT4 #(
		.INIT('h7077)
	) name2644 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8471_
	);
	LUT4 #(
		.INIT('haa02)
	) name2645 (
		_w8450_,
		_w8447_,
		_w8452_,
		_w8448_,
		_w8472_
	);
	LUT3 #(
		.INIT('h01)
	) name2646 (
		_w8447_,
		_w8452_,
		_w8449_,
		_w8473_
	);
	LUT4 #(
		.INIT('h45cf)
	) name2647 (
		_w8458_,
		_w8471_,
		_w8472_,
		_w8473_,
		_w8474_
	);
	LUT2 #(
		.INIT('h4)
	) name2648 (
		_w8470_,
		_w8474_,
		_w8475_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2649 (
		\u2_L9_reg[11]/NET0131 ,
		_w8468_,
		_w8461_,
		_w8475_,
		_w8476_
	);
	LUT4 #(
		.INIT('hc963)
	) name2650 (
		decrypt_pad,
		\u2_R9_reg[13]/NET0131 ,
		\u2_uk_K_r9_reg[10]/NET0131 ,
		\u2_uk_K_r9_reg[4]/NET0131 ,
		_w8477_
	);
	LUT4 #(
		.INIT('hc693)
	) name2651 (
		decrypt_pad,
		\u2_R9_reg[12]/NET0131 ,
		\u2_uk_K_r9_reg[10]/NET0131 ,
		\u2_uk_K_r9_reg[48]/NET0131 ,
		_w8478_
	);
	LUT2 #(
		.INIT('h2)
	) name2652 (
		_w8477_,
		_w8478_,
		_w8479_
	);
	LUT2 #(
		.INIT('h9)
	) name2653 (
		_w8477_,
		_w8478_,
		_w8480_
	);
	LUT4 #(
		.INIT('hc963)
	) name2654 (
		decrypt_pad,
		\u2_R9_reg[14]/NET0131 ,
		\u2_uk_K_r9_reg[11]/NET0131 ,
		\u2_uk_K_r9_reg[5]/NET0131 ,
		_w8481_
	);
	LUT4 #(
		.INIT('hc693)
	) name2655 (
		decrypt_pad,
		\u2_R9_reg[15]/NET0131 ,
		\u2_uk_K_r9_reg[13]/NET0131 ,
		\u2_uk_K_r9_reg[19]/NET0131 ,
		_w8482_
	);
	LUT4 #(
		.INIT('h0012)
	) name2656 (
		_w8477_,
		_w8481_,
		_w8478_,
		_w8482_,
		_w8483_
	);
	LUT4 #(
		.INIT('hc693)
	) name2657 (
		decrypt_pad,
		\u2_R9_reg[17]/NET0131 ,
		\u2_uk_K_r9_reg[26]/NET0131 ,
		\u2_uk_K_r9_reg[32]/NET0131 ,
		_w8484_
	);
	LUT2 #(
		.INIT('h8)
	) name2658 (
		_w8477_,
		_w8482_,
		_w8485_
	);
	LUT4 #(
		.INIT('h2000)
	) name2659 (
		_w8477_,
		_w8484_,
		_w8478_,
		_w8482_,
		_w8486_
	);
	LUT2 #(
		.INIT('h4)
	) name2660 (
		_w8477_,
		_w8482_,
		_w8487_
	);
	LUT4 #(
		.INIT('h0400)
	) name2661 (
		_w8477_,
		_w8484_,
		_w8478_,
		_w8482_,
		_w8488_
	);
	LUT4 #(
		.INIT('hc963)
	) name2662 (
		decrypt_pad,
		\u2_R9_reg[16]/NET0131 ,
		\u2_uk_K_r9_reg[27]/NET0131 ,
		\u2_uk_K_r9_reg[46]/NET0131 ,
		_w8489_
	);
	LUT4 #(
		.INIT('h0100)
	) name2663 (
		_w8483_,
		_w8488_,
		_w8486_,
		_w8489_,
		_w8490_
	);
	LUT4 #(
		.INIT('h0008)
	) name2664 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8491_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name2665 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8492_
	);
	LUT3 #(
		.INIT('h01)
	) name2666 (
		_w8477_,
		_w8484_,
		_w8478_,
		_w8493_
	);
	LUT4 #(
		.INIT('h0001)
	) name2667 (
		_w8477_,
		_w8484_,
		_w8478_,
		_w8482_,
		_w8494_
	);
	LUT3 #(
		.INIT('h4c)
	) name2668 (
		_w8481_,
		_w8492_,
		_w8494_,
		_w8495_
	);
	LUT2 #(
		.INIT('h8)
	) name2669 (
		_w8490_,
		_w8495_,
		_w8496_
	);
	LUT2 #(
		.INIT('h1)
	) name2670 (
		_w8481_,
		_w8478_,
		_w8497_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2671 (
		_w8477_,
		_w8484_,
		_w8478_,
		_w8482_,
		_w8498_
	);
	LUT2 #(
		.INIT('h4)
	) name2672 (
		_w8497_,
		_w8498_,
		_w8499_
	);
	LUT4 #(
		.INIT('h0100)
	) name2673 (
		_w8477_,
		_w8484_,
		_w8478_,
		_w8482_,
		_w8500_
	);
	LUT4 #(
		.INIT('h0400)
	) name2674 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8501_
	);
	LUT3 #(
		.INIT('h01)
	) name2675 (
		_w8489_,
		_w8500_,
		_w8501_,
		_w8502_
	);
	LUT4 #(
		.INIT('hffde)
	) name2676 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8503_
	);
	LUT3 #(
		.INIT('h40)
	) name2677 (
		_w8484_,
		_w8481_,
		_w8478_,
		_w8504_
	);
	LUT4 #(
		.INIT('h8bbb)
	) name2678 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8505_
	);
	LUT3 #(
		.INIT('hc8)
	) name2679 (
		_w8482_,
		_w8503_,
		_w8505_,
		_w8506_
	);
	LUT3 #(
		.INIT('h40)
	) name2680 (
		_w8499_,
		_w8502_,
		_w8506_,
		_w8507_
	);
	LUT3 #(
		.INIT('hbe)
	) name2681 (
		_w8484_,
		_w8481_,
		_w8478_,
		_w8508_
	);
	LUT2 #(
		.INIT('h2)
	) name2682 (
		_w8487_,
		_w8508_,
		_w8509_
	);
	LUT3 #(
		.INIT('h02)
	) name2683 (
		_w8484_,
		_w8481_,
		_w8482_,
		_w8510_
	);
	LUT4 #(
		.INIT('h23af)
	) name2684 (
		_w8481_,
		_w8479_,
		_w8486_,
		_w8510_,
		_w8511_
	);
	LUT2 #(
		.INIT('h4)
	) name2685 (
		_w8509_,
		_w8511_,
		_w8512_
	);
	LUT4 #(
		.INIT('ha955)
	) name2686 (
		\u2_L9_reg[20]/NET0131 ,
		_w8496_,
		_w8507_,
		_w8512_,
		_w8513_
	);
	LUT4 #(
		.INIT('hc963)
	) name2687 (
		decrypt_pad,
		\u2_R9_reg[31]/P0001 ,
		\u2_uk_K_r9_reg[45]/NET0131 ,
		\u2_uk_K_r9_reg[9]/NET0131 ,
		_w8514_
	);
	LUT4 #(
		.INIT('hc693)
	) name2688 (
		decrypt_pad,
		\u2_R9_reg[1]/NET0131 ,
		\u2_uk_K_r9_reg[36]/NET0131 ,
		\u2_uk_K_r9_reg[44]/NET0131 ,
		_w8515_
	);
	LUT4 #(
		.INIT('hc693)
	) name2689 (
		decrypt_pad,
		\u2_R9_reg[30]/NET0131 ,
		\u2_uk_K_r9_reg[21]/NET0131 ,
		\u2_uk_K_r9_reg[29]/NET0131 ,
		_w8516_
	);
	LUT4 #(
		.INIT('hc963)
	) name2690 (
		decrypt_pad,
		\u2_R9_reg[28]/NET0131 ,
		\u2_uk_K_r9_reg[1]/NET0131 ,
		\u2_uk_K_r9_reg[52]/NET0131 ,
		_w8517_
	);
	LUT4 #(
		.INIT('hc963)
	) name2691 (
		decrypt_pad,
		\u2_R9_reg[29]/NET0131 ,
		\u2_uk_K_r9_reg[28]/NET0131 ,
		\u2_uk_K_r9_reg[51]/NET0131 ,
		_w8518_
	);
	LUT4 #(
		.INIT('h0020)
	) name2692 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8519_
	);
	LUT4 #(
		.INIT('heedf)
	) name2693 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8520_
	);
	LUT2 #(
		.INIT('h2)
	) name2694 (
		_w8514_,
		_w8520_,
		_w8521_
	);
	LUT2 #(
		.INIT('h1)
	) name2695 (
		_w8516_,
		_w8514_,
		_w8522_
	);
	LUT4 #(
		.INIT('h7d4c)
	) name2696 (
		_w8518_,
		_w8516_,
		_w8515_,
		_w8514_,
		_w8523_
	);
	LUT3 #(
		.INIT('h0b)
	) name2697 (
		_w8518_,
		_w8515_,
		_w8514_,
		_w8524_
	);
	LUT3 #(
		.INIT('hf4)
	) name2698 (
		_w8517_,
		_w8516_,
		_w8515_,
		_w8525_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name2699 (
		_w8517_,
		_w8523_,
		_w8524_,
		_w8525_,
		_w8526_
	);
	LUT4 #(
		.INIT('hc693)
	) name2700 (
		decrypt_pad,
		\u2_R9_reg[32]/NET0131 ,
		\u2_uk_K_r9_reg[15]/NET0131 ,
		\u2_uk_K_r9_reg[23]/NET0131 ,
		_w8527_
	);
	LUT3 #(
		.INIT('h0b)
	) name2701 (
		_w8521_,
		_w8526_,
		_w8527_,
		_w8528_
	);
	LUT3 #(
		.INIT('h20)
	) name2702 (
		_w8517_,
		_w8516_,
		_w8515_,
		_w8529_
	);
	LUT4 #(
		.INIT('hf539)
	) name2703 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8530_
	);
	LUT4 #(
		.INIT('h4000)
	) name2704 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8531_
	);
	LUT3 #(
		.INIT('h01)
	) name2705 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8532_
	);
	LUT4 #(
		.INIT('h2031)
	) name2706 (
		_w8514_,
		_w8531_,
		_w8530_,
		_w8532_,
		_w8533_
	);
	LUT4 #(
		.INIT('h0040)
	) name2707 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8534_
	);
	LUT4 #(
		.INIT('hffbe)
	) name2708 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8535_
	);
	LUT4 #(
		.INIT('h1000)
	) name2709 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8536_
	);
	LUT4 #(
		.INIT('hedbe)
	) name2710 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8537_
	);
	LUT2 #(
		.INIT('h2)
	) name2711 (
		_w8514_,
		_w8537_,
		_w8538_
	);
	LUT3 #(
		.INIT('h20)
	) name2712 (
		_w8517_,
		_w8518_,
		_w8527_,
		_w8539_
	);
	LUT3 #(
		.INIT('h08)
	) name2713 (
		_w8517_,
		_w8518_,
		_w8515_,
		_w8540_
	);
	LUT4 #(
		.INIT('hcedf)
	) name2714 (
		_w8516_,
		_w8514_,
		_w8539_,
		_w8540_,
		_w8541_
	);
	LUT4 #(
		.INIT('h3100)
	) name2715 (
		_w8527_,
		_w8538_,
		_w8533_,
		_w8541_,
		_w8542_
	);
	LUT3 #(
		.INIT('h9a)
	) name2716 (
		\u2_L9_reg[5]/NET0131 ,
		_w8528_,
		_w8542_,
		_w8543_
	);
	LUT4 #(
		.INIT('ha4f1)
	) name2717 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8482_,
		_w8544_
	);
	LUT2 #(
		.INIT('h2)
	) name2718 (
		_w8478_,
		_w8544_,
		_w8545_
	);
	LUT3 #(
		.INIT('h20)
	) name2719 (
		_w8484_,
		_w8481_,
		_w8482_,
		_w8546_
	);
	LUT4 #(
		.INIT('h0200)
	) name2720 (
		_w8484_,
		_w8481_,
		_w8478_,
		_w8482_,
		_w8547_
	);
	LUT3 #(
		.INIT('h04)
	) name2721 (
		_w8494_,
		_w8503_,
		_w8547_,
		_w8548_
	);
	LUT3 #(
		.INIT('h45)
	) name2722 (
		_w8489_,
		_w8545_,
		_w8548_,
		_w8549_
	);
	LUT4 #(
		.INIT('hcef7)
	) name2723 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8550_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name2724 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8551_
	);
	LUT4 #(
		.INIT('hfbdd)
	) name2725 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8552_
	);
	LUT4 #(
		.INIT('hc480)
	) name2726 (
		_w8482_,
		_w8551_,
		_w8552_,
		_w8550_,
		_w8553_
	);
	LUT4 #(
		.INIT('h7fbe)
	) name2727 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8554_
	);
	LUT3 #(
		.INIT('he3)
	) name2728 (
		_w8484_,
		_w8481_,
		_w8478_,
		_w8555_
	);
	LUT4 #(
		.INIT('hfc74)
	) name2729 (
		_w8477_,
		_w8482_,
		_w8554_,
		_w8555_,
		_w8556_
	);
	LUT3 #(
		.INIT('hd0)
	) name2730 (
		_w8489_,
		_w8553_,
		_w8556_,
		_w8557_
	);
	LUT3 #(
		.INIT('h65)
	) name2731 (
		\u2_L9_reg[10]/NET0131 ,
		_w8549_,
		_w8557_,
		_w8558_
	);
	LUT2 #(
		.INIT('h2)
	) name2732 (
		_w8383_,
		_w8406_,
		_w8559_
	);
	LUT3 #(
		.INIT('h0b)
	) name2733 (
		_w8384_,
		_w8396_,
		_w8389_,
		_w8560_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name2734 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8561_
	);
	LUT4 #(
		.INIT('h0420)
	) name2735 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8562_
	);
	LUT3 #(
		.INIT('h0d)
	) name2736 (
		_w8384_,
		_w8561_,
		_w8562_,
		_w8563_
	);
	LUT3 #(
		.INIT('h80)
	) name2737 (
		_w8559_,
		_w8560_,
		_w8563_,
		_w8564_
	);
	LUT4 #(
		.INIT('h0014)
	) name2738 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8565_
	);
	LUT4 #(
		.INIT('h2000)
	) name2739 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8566_
	);
	LUT3 #(
		.INIT('h20)
	) name2740 (
		_w8385_,
		_w8384_,
		_w8386_,
		_w8567_
	);
	LUT4 #(
		.INIT('h0001)
	) name2741 (
		_w8401_,
		_w8383_,
		_w8566_,
		_w8567_,
		_w8568_
	);
	LUT3 #(
		.INIT('h47)
	) name2742 (
		_w8385_,
		_w8387_,
		_w8384_,
		_w8569_
	);
	LUT3 #(
		.INIT('h21)
	) name2743 (
		_w8387_,
		_w8384_,
		_w8388_,
		_w8570_
	);
	LUT3 #(
		.INIT('h0d)
	) name2744 (
		_w8390_,
		_w8569_,
		_w8570_,
		_w8571_
	);
	LUT3 #(
		.INIT('h40)
	) name2745 (
		_w8565_,
		_w8568_,
		_w8571_,
		_w8572_
	);
	LUT3 #(
		.INIT('ha9)
	) name2746 (
		\u2_L9_reg[12]/NET0131 ,
		_w8564_,
		_w8572_,
		_w8573_
	);
	LUT4 #(
		.INIT('hc693)
	) name2747 (
		decrypt_pad,
		\u2_R9_reg[20]/NET0131 ,
		\u2_uk_K_r9_reg[0]/P0001 ,
		\u2_uk_K_r9_reg[8]/NET0131 ,
		_w8574_
	);
	LUT4 #(
		.INIT('hc693)
	) name2748 (
		decrypt_pad,
		\u2_R9_reg[18]/NET0131 ,
		\u2_uk_K_r9_reg[29]/NET0131 ,
		\u2_uk_K_r9_reg[37]/NET0131 ,
		_w8575_
	);
	LUT4 #(
		.INIT('hc693)
	) name2749 (
		decrypt_pad,
		\u2_R9_reg[17]/NET0131 ,
		\u2_uk_K_r9_reg[35]/NET0131 ,
		\u2_uk_K_r9_reg[43]/NET0131 ,
		_w8576_
	);
	LUT4 #(
		.INIT('hc963)
	) name2750 (
		decrypt_pad,
		\u2_R9_reg[16]/NET0131 ,
		\u2_uk_K_r9_reg[21]/NET0131 ,
		\u2_uk_K_r9_reg[44]/NET0131 ,
		_w8577_
	);
	LUT4 #(
		.INIT('hc693)
	) name2751 (
		decrypt_pad,
		\u2_R9_reg[21]/NET0131 ,
		\u2_uk_K_r9_reg[1]/NET0131 ,
		\u2_uk_K_r9_reg[9]/NET0131 ,
		_w8578_
	);
	LUT2 #(
		.INIT('h2)
	) name2752 (
		_w8577_,
		_w8578_,
		_w8579_
	);
	LUT4 #(
		.INIT('h2010)
	) name2753 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8580_
	);
	LUT3 #(
		.INIT('h10)
	) name2754 (
		_w8576_,
		_w8577_,
		_w8578_,
		_w8581_
	);
	LUT4 #(
		.INIT('hc693)
	) name2755 (
		decrypt_pad,
		\u2_R9_reg[19]/NET0131 ,
		\u2_uk_K_r9_reg[16]/NET0131 ,
		\u2_uk_K_r9_reg[52]/NET0131 ,
		_w8582_
	);
	LUT4 #(
		.INIT('h00f7)
	) name2756 (
		_w8576_,
		_w8575_,
		_w8578_,
		_w8582_,
		_w8583_
	);
	LUT3 #(
		.INIT('h10)
	) name2757 (
		_w8581_,
		_w8580_,
		_w8583_,
		_w8584_
	);
	LUT4 #(
		.INIT('hc005)
	) name2758 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8585_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2759 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8582_,
		_w8586_
	);
	LUT2 #(
		.INIT('h4)
	) name2760 (
		_w8585_,
		_w8586_,
		_w8587_
	);
	LUT4 #(
		.INIT('h4000)
	) name2761 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8588_
	);
	LUT4 #(
		.INIT('hbffd)
	) name2762 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8589_
	);
	LUT4 #(
		.INIT('h0155)
	) name2763 (
		_w8574_,
		_w8584_,
		_w8587_,
		_w8589_,
		_w8590_
	);
	LUT4 #(
		.INIT('hc25f)
	) name2764 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8591_
	);
	LUT2 #(
		.INIT('h4)
	) name2765 (
		_w8591_,
		_w8582_,
		_w8592_
	);
	LUT4 #(
		.INIT('h0021)
	) name2766 (
		_w8576_,
		_w8577_,
		_w8578_,
		_w8582_,
		_w8593_
	);
	LUT4 #(
		.INIT('h2313)
	) name2767 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8594_
	);
	LUT4 #(
		.INIT('h0080)
	) name2768 (
		_w8576_,
		_w8577_,
		_w8578_,
		_w8582_,
		_w8595_
	);
	LUT4 #(
		.INIT('hcc8c)
	) name2769 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8596_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2770 (
		_w8593_,
		_w8594_,
		_w8595_,
		_w8596_,
		_w8597_
	);
	LUT4 #(
		.INIT('h0400)
	) name2771 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8598_
	);
	LUT4 #(
		.INIT('h0408)
	) name2772 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8599_
	);
	LUT4 #(
		.INIT('hffdb)
	) name2773 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8600_
	);
	LUT3 #(
		.INIT('hb1)
	) name2774 (
		_w8582_,
		_w8599_,
		_w8600_,
		_w8601_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2775 (
		_w8592_,
		_w8597_,
		_w8574_,
		_w8601_,
		_w8602_
	);
	LUT3 #(
		.INIT('h65)
	) name2776 (
		\u2_L9_reg[14]/NET0131 ,
		_w8590_,
		_w8602_,
		_w8603_
	);
	LUT4 #(
		.INIT('h7773)
	) name2777 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8604_
	);
	LUT4 #(
		.INIT('h6673)
	) name2778 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8605_
	);
	LUT4 #(
		.INIT('h0002)
	) name2779 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8606_
	);
	LUT4 #(
		.INIT('h0301)
	) name2780 (
		_w8514_,
		_w8527_,
		_w8606_,
		_w8605_,
		_w8607_
	);
	LUT4 #(
		.INIT('h0040)
	) name2781 (
		_w8518_,
		_w8516_,
		_w8515_,
		_w8514_,
		_w8608_
	);
	LUT3 #(
		.INIT('h08)
	) name2782 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8609_
	);
	LUT4 #(
		.INIT('h0002)
	) name2783 (
		_w8527_,
		_w8534_,
		_w8608_,
		_w8609_,
		_w8610_
	);
	LUT4 #(
		.INIT('h0100)
	) name2784 (
		_w8517_,
		_w8518_,
		_w8515_,
		_w8514_,
		_w8611_
	);
	LUT4 #(
		.INIT('h2000)
	) name2785 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8612_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		_w8611_,
		_w8612_,
		_w8613_
	);
	LUT3 #(
		.INIT('h15)
	) name2787 (
		_w8607_,
		_w8610_,
		_w8613_,
		_w8614_
	);
	LUT4 #(
		.INIT('h00df)
	) name2788 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8514_,
		_w8615_
	);
	LUT4 #(
		.INIT('h0400)
	) name2789 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8616_
	);
	LUT3 #(
		.INIT('h02)
	) name2790 (
		_w8517_,
		_w8518_,
		_w8527_,
		_w8617_
	);
	LUT4 #(
		.INIT('h0200)
	) name2791 (
		_w8535_,
		_w8616_,
		_w8617_,
		_w8615_,
		_w8618_
	);
	LUT4 #(
		.INIT('h0100)
	) name2792 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8619_
	);
	LUT3 #(
		.INIT('h02)
	) name2793 (
		_w8514_,
		_w8531_,
		_w8619_,
		_w8620_
	);
	LUT2 #(
		.INIT('h1)
	) name2794 (
		_w8618_,
		_w8620_,
		_w8621_
	);
	LUT3 #(
		.INIT('h56)
	) name2795 (
		\u2_L9_reg[15]/NET0131 ,
		_w8614_,
		_w8621_,
		_w8622_
	);
	LUT4 #(
		.INIT('hfb05)
	) name2796 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8623_
	);
	LUT4 #(
		.INIT('h5001)
	) name2797 (
		_w8414_,
		_w8418_,
		_w8416_,
		_w8419_,
		_w8624_
	);
	LUT4 #(
		.INIT('h0200)
	) name2798 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8625_
	);
	LUT4 #(
		.INIT('h7d7f)
	) name2799 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8626_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2800 (
		_w8414_,
		_w8623_,
		_w8624_,
		_w8626_,
		_w8627_
	);
	LUT3 #(
		.INIT('hf9)
	) name2801 (
		_w8417_,
		_w8416_,
		_w8419_,
		_w8628_
	);
	LUT2 #(
		.INIT('h8)
	) name2802 (
		_w8414_,
		_w8418_,
		_w8629_
	);
	LUT2 #(
		.INIT('h4)
	) name2803 (
		_w8628_,
		_w8629_,
		_w8630_
	);
	LUT2 #(
		.INIT('h6)
	) name2804 (
		_w8417_,
		_w8419_,
		_w8631_
	);
	LUT4 #(
		.INIT('hbbec)
	) name2805 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8632_
	);
	LUT3 #(
		.INIT('h80)
	) name2806 (
		_w8418_,
		_w8417_,
		_w8419_,
		_w8633_
	);
	LUT3 #(
		.INIT('h6f)
	) name2807 (
		_w8418_,
		_w8417_,
		_w8419_,
		_w8634_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name2808 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8635_
	);
	LUT4 #(
		.INIT('he400)
	) name2809 (
		_w8414_,
		_w8632_,
		_w8634_,
		_w8635_,
		_w8636_
	);
	LUT4 #(
		.INIT('h3210)
	) name2810 (
		_w8415_,
		_w8630_,
		_w8636_,
		_w8627_,
		_w8637_
	);
	LUT2 #(
		.INIT('h9)
	) name2811 (
		\u2_L9_reg[17]/NET0131 ,
		_w8637_,
		_w8638_
	);
	LUT3 #(
		.INIT('h40)
	) name2812 (
		_w8477_,
		_w8484_,
		_w8478_,
		_w8639_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2813 (
		_w8484_,
		_w8481_,
		_w8478_,
		_w8482_,
		_w8640_
	);
	LUT4 #(
		.INIT('h1000)
	) name2814 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8641_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2815 (
		_w8484_,
		_w8481_,
		_w8478_,
		_w8482_,
		_w8642_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2816 (
		_w8639_,
		_w8640_,
		_w8641_,
		_w8642_,
		_w8643_
	);
	LUT4 #(
		.INIT('h7df7)
	) name2817 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8644_
	);
	LUT3 #(
		.INIT('h45)
	) name2818 (
		_w8489_,
		_w8643_,
		_w8644_,
		_w8645_
	);
	LUT3 #(
		.INIT('hc4)
	) name2819 (
		_w8484_,
		_w8481_,
		_w8478_,
		_w8646_
	);
	LUT2 #(
		.INIT('h2)
	) name2820 (
		_w8477_,
		_w8482_,
		_w8647_
	);
	LUT4 #(
		.INIT('h008a)
	) name2821 (
		_w8477_,
		_w8484_,
		_w8478_,
		_w8482_,
		_w8648_
	);
	LUT4 #(
		.INIT('hdfaf)
	) name2822 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8649_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2823 (
		_w8489_,
		_w8646_,
		_w8648_,
		_w8649_,
		_w8650_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name2824 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8651_
	);
	LUT2 #(
		.INIT('h2)
	) name2825 (
		_w8482_,
		_w8651_,
		_w8652_
	);
	LUT3 #(
		.INIT('h10)
	) name2826 (
		_w8477_,
		_w8481_,
		_w8478_,
		_w8653_
	);
	LUT4 #(
		.INIT('hbabb)
	) name2827 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8654_
	);
	LUT2 #(
		.INIT('h8)
	) name2828 (
		_w8482_,
		_w8489_,
		_w8655_
	);
	LUT2 #(
		.INIT('h4)
	) name2829 (
		_w8654_,
		_w8655_,
		_w8656_
	);
	LUT4 #(
		.INIT('h0777)
	) name2830 (
		_w8481_,
		_w8494_,
		_w8504_,
		_w8647_,
		_w8657_
	);
	LUT4 #(
		.INIT('h0100)
	) name2831 (
		_w8652_,
		_w8656_,
		_w8650_,
		_w8657_,
		_w8658_
	);
	LUT3 #(
		.INIT('h65)
	) name2832 (
		\u2_L9_reg[1]/NET0131 ,
		_w8645_,
		_w8658_,
		_w8659_
	);
	LUT4 #(
		.INIT('hdff5)
	) name2833 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8660_
	);
	LUT4 #(
		.INIT('h387f)
	) name2834 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8661_
	);
	LUT4 #(
		.INIT('hfe6f)
	) name2835 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8662_
	);
	LUT4 #(
		.INIT('hd800)
	) name2836 (
		_w8514_,
		_w8661_,
		_w8660_,
		_w8662_,
		_w8663_
	);
	LUT2 #(
		.INIT('h2)
	) name2837 (
		_w8527_,
		_w8663_,
		_w8664_
	);
	LUT4 #(
		.INIT('hdf57)
	) name2838 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8665_
	);
	LUT2 #(
		.INIT('h2)
	) name2839 (
		_w8514_,
		_w8665_,
		_w8666_
	);
	LUT4 #(
		.INIT('hbfbe)
	) name2840 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8667_
	);
	LUT4 #(
		.INIT('h0040)
	) name2841 (
		_w8517_,
		_w8516_,
		_w8515_,
		_w8514_,
		_w8668_
	);
	LUT2 #(
		.INIT('h2)
	) name2842 (
		_w8518_,
		_w8514_,
		_w8669_
	);
	LUT4 #(
		.INIT('h0004)
	) name2843 (
		_w8517_,
		_w8518_,
		_w8515_,
		_w8514_,
		_w8670_
	);
	LUT3 #(
		.INIT('h10)
	) name2844 (
		_w8668_,
		_w8670_,
		_w8667_,
		_w8671_
	);
	LUT2 #(
		.INIT('h4)
	) name2845 (
		_w8518_,
		_w8514_,
		_w8672_
	);
	LUT3 #(
		.INIT('h51)
	) name2846 (
		_w8519_,
		_w8529_,
		_w8672_,
		_w8673_
	);
	LUT4 #(
		.INIT('h4555)
	) name2847 (
		_w8527_,
		_w8666_,
		_w8671_,
		_w8673_,
		_w8674_
	);
	LUT4 #(
		.INIT('h0100)
	) name2848 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8514_,
		_w8675_
	);
	LUT3 #(
		.INIT('h07)
	) name2849 (
		_w8529_,
		_w8669_,
		_w8675_,
		_w8676_
	);
	LUT4 #(
		.INIT('h5655)
	) name2850 (
		\u2_L9_reg[21]/NET0131 ,
		_w8674_,
		_w8664_,
		_w8676_,
		_w8677_
	);
	LUT4 #(
		.INIT('h5ae2)
	) name2851 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8678_
	);
	LUT4 #(
		.INIT('hadfd)
	) name2852 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8679_
	);
	LUT4 #(
		.INIT('hdd7f)
	) name2853 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8680_
	);
	LUT4 #(
		.INIT('hd800)
	) name2854 (
		_w8582_,
		_w8678_,
		_w8679_,
		_w8680_,
		_w8681_
	);
	LUT4 #(
		.INIT('hf6a6)
	) name2855 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8682_
	);
	LUT3 #(
		.INIT('h8a)
	) name2856 (
		_w8575_,
		_w8577_,
		_w8578_,
		_w8683_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2857 (
		_w8576_,
		_w8575_,
		_w8578_,
		_w8582_,
		_w8684_
	);
	LUT4 #(
		.INIT('he0ee)
	) name2858 (
		_w8582_,
		_w8682_,
		_w8683_,
		_w8684_,
		_w8685_
	);
	LUT4 #(
		.INIT('hfe7b)
	) name2859 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8686_
	);
	LUT3 #(
		.INIT('h04)
	) name2860 (
		_w8576_,
		_w8575_,
		_w8582_,
		_w8687_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name2861 (
		_w8576_,
		_w8575_,
		_w8578_,
		_w8582_,
		_w8688_
	);
	LUT4 #(
		.INIT('hf351)
	) name2862 (
		_w8577_,
		_w8582_,
		_w8686_,
		_w8688_,
		_w8689_
	);
	LUT4 #(
		.INIT('he400)
	) name2863 (
		_w8574_,
		_w8685_,
		_w8681_,
		_w8689_,
		_w8690_
	);
	LUT2 #(
		.INIT('h9)
	) name2864 (
		\u2_L9_reg[25]/NET0131 ,
		_w8690_,
		_w8691_
	);
	LUT4 #(
		.INIT('hc693)
	) name2865 (
		decrypt_pad,
		\u2_R9_reg[5]/NET0131 ,
		\u2_uk_K_r9_reg[12]/NET0131 ,
		\u2_uk_K_r9_reg[18]/NET0131 ,
		_w8692_
	);
	LUT4 #(
		.INIT('hc693)
	) name2866 (
		decrypt_pad,
		\u2_R9_reg[4]/NET0131 ,
		\u2_uk_K_r9_reg[33]/NET0131 ,
		\u2_uk_K_r9_reg[39]/NET0131 ,
		_w8693_
	);
	LUT4 #(
		.INIT('hc693)
	) name2867 (
		decrypt_pad,
		\u2_R9_reg[9]/NET0131 ,
		\u2_uk_K_r9_reg[25]/NET0131 ,
		\u2_uk_K_r9_reg[6]/NET0131 ,
		_w8694_
	);
	LUT4 #(
		.INIT('hc693)
	) name2868 (
		decrypt_pad,
		\u2_R9_reg[6]/NET0131 ,
		\u2_uk_K_r9_reg[3]/NET0131 ,
		\u2_uk_K_r9_reg[41]/NET0131 ,
		_w8695_
	);
	LUT4 #(
		.INIT('hc038)
	) name2869 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8696_
	);
	LUT4 #(
		.INIT('hc963)
	) name2870 (
		decrypt_pad,
		\u2_R9_reg[7]/NET0131 ,
		\u2_uk_K_r9_reg[3]/NET0131 ,
		\u2_uk_K_r9_reg[54]/NET0131 ,
		_w8697_
	);
	LUT2 #(
		.INIT('h4)
	) name2871 (
		_w8696_,
		_w8697_,
		_w8698_
	);
	LUT4 #(
		.INIT('h0c05)
	) name2872 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8699_
	);
	LUT4 #(
		.INIT('h0080)
	) name2873 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8700_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2874 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8697_,
		_w8701_
	);
	LUT3 #(
		.INIT('h10)
	) name2875 (
		_w8699_,
		_w8700_,
		_w8701_,
		_w8702_
	);
	LUT3 #(
		.INIT('h40)
	) name2876 (
		_w8692_,
		_w8693_,
		_w8694_,
		_w8703_
	);
	LUT4 #(
		.INIT('h00bf)
	) name2877 (
		_w8692_,
		_w8693_,
		_w8694_,
		_w8697_,
		_w8704_
	);
	LUT2 #(
		.INIT('h4)
	) name2878 (
		_w8695_,
		_w8693_,
		_w8705_
	);
	LUT4 #(
		.INIT('h0200)
	) name2879 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8706_
	);
	LUT4 #(
		.INIT('hc693)
	) name2880 (
		decrypt_pad,
		\u2_R9_reg[8]/NET0131 ,
		\u2_uk_K_r9_reg[20]/NET0131 ,
		\u2_uk_K_r9_reg[26]/NET0131 ,
		_w8707_
	);
	LUT4 #(
		.INIT('h4500)
	) name2881 (
		_w8706_,
		_w8704_,
		_w8705_,
		_w8707_,
		_w8708_
	);
	LUT3 #(
		.INIT('he0)
	) name2882 (
		_w8698_,
		_w8702_,
		_w8708_,
		_w8709_
	);
	LUT2 #(
		.INIT('h2)
	) name2883 (
		_w8697_,
		_w8699_,
		_w8710_
	);
	LUT4 #(
		.INIT('h3c2f)
	) name2884 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8711_
	);
	LUT3 #(
		.INIT('h40)
	) name2885 (
		_w8700_,
		_w8701_,
		_w8711_,
		_w8712_
	);
	LUT4 #(
		.INIT('h2002)
	) name2886 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8713_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		_w8700_,
		_w8707_,
		_w8714_
	);
	LUT3 #(
		.INIT('h01)
	) name2888 (
		_w8700_,
		_w8707_,
		_w8713_,
		_w8715_
	);
	LUT3 #(
		.INIT('he0)
	) name2889 (
		_w8710_,
		_w8712_,
		_w8715_,
		_w8716_
	);
	LUT3 #(
		.INIT('ha9)
	) name2890 (
		\u2_L9_reg[28]/NET0131 ,
		_w8709_,
		_w8716_,
		_w8717_
	);
	LUT4 #(
		.INIT('h67dc)
	) name2891 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8718_
	);
	LUT4 #(
		.INIT('hd2f7)
	) name2892 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8719_
	);
	LUT4 #(
		.INIT('h0040)
	) name2893 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8720_
	);
	LUT4 #(
		.INIT('h00d8)
	) name2894 (
		_w8450_,
		_w8718_,
		_w8719_,
		_w8720_,
		_w8721_
	);
	LUT4 #(
		.INIT('h9aff)
	) name2895 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8722_
	);
	LUT4 #(
		.INIT('haa02)
	) name2896 (
		_w8450_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8723_
	);
	LUT4 #(
		.INIT('h9297)
	) name2897 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8724_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2898 (
		_w8450_,
		_w8722_,
		_w8723_,
		_w8724_,
		_w8725_
	);
	LUT4 #(
		.INIT('h0800)
	) name2899 (
		_w8450_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8726_
	);
	LUT2 #(
		.INIT('h1)
	) name2900 (
		_w8462_,
		_w8726_,
		_w8727_
	);
	LUT4 #(
		.INIT('hd800)
	) name2901 (
		_w8446_,
		_w8725_,
		_w8721_,
		_w8727_,
		_w8728_
	);
	LUT2 #(
		.INIT('h6)
	) name2902 (
		\u2_L9_reg[29]/NET0131 ,
		_w8728_,
		_w8729_
	);
	LUT4 #(
		.INIT('hd3d7)
	) name2903 (
		_w8477_,
		_w8484_,
		_w8478_,
		_w8482_,
		_w8730_
	);
	LUT2 #(
		.INIT('h2)
	) name2904 (
		_w8481_,
		_w8730_,
		_w8731_
	);
	LUT4 #(
		.INIT('h3ffb)
	) name2905 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8732_
	);
	LUT4 #(
		.INIT('h0002)
	) name2906 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8733_
	);
	LUT4 #(
		.INIT('h0702)
	) name2907 (
		_w8482_,
		_w8493_,
		_w8733_,
		_w8732_,
		_w8734_
	);
	LUT3 #(
		.INIT('h8a)
	) name2908 (
		_w8489_,
		_w8731_,
		_w8734_,
		_w8735_
	);
	LUT2 #(
		.INIT('h8)
	) name2909 (
		_w8485_,
		_w8646_,
		_w8736_
	);
	LUT3 #(
		.INIT('h01)
	) name2910 (
		_w8491_,
		_w8486_,
		_w8653_,
		_w8737_
	);
	LUT3 #(
		.INIT('h45)
	) name2911 (
		_w8489_,
		_w8736_,
		_w8737_,
		_w8738_
	);
	LUT2 #(
		.INIT('h4)
	) name2912 (
		_w8480_,
		_w8546_,
		_w8739_
	);
	LUT4 #(
		.INIT('heeae)
	) name2913 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8740_
	);
	LUT4 #(
		.INIT('h0902)
	) name2914 (
		_w8477_,
		_w8484_,
		_w8481_,
		_w8478_,
		_w8741_
	);
	LUT4 #(
		.INIT('h5501)
	) name2915 (
		_w8482_,
		_w8489_,
		_w8740_,
		_w8741_,
		_w8742_
	);
	LUT2 #(
		.INIT('h1)
	) name2916 (
		_w8739_,
		_w8742_,
		_w8743_
	);
	LUT4 #(
		.INIT('h5655)
	) name2917 (
		\u2_L9_reg[26]/NET0131 ,
		_w8735_,
		_w8738_,
		_w8743_,
		_w8744_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name2918 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8745_
	);
	LUT4 #(
		.INIT('h7f7c)
	) name2919 (
		_w8695_,
		_w8697_,
		_w8703_,
		_w8745_,
		_w8746_
	);
	LUT4 #(
		.INIT('h0144)
	) name2920 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8747_
	);
	LUT4 #(
		.INIT('h0800)
	) name2921 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8748_
	);
	LUT4 #(
		.INIT('h0010)
	) name2922 (
		_w8695_,
		_w8692_,
		_w8694_,
		_w8697_,
		_w8749_
	);
	LUT3 #(
		.INIT('h01)
	) name2923 (
		_w8747_,
		_w8748_,
		_w8749_,
		_w8750_
	);
	LUT3 #(
		.INIT('h15)
	) name2924 (
		_w8707_,
		_w8746_,
		_w8750_,
		_w8751_
	);
	LUT3 #(
		.INIT('h01)
	) name2925 (
		_w8695_,
		_w8692_,
		_w8694_,
		_w8752_
	);
	LUT4 #(
		.INIT('h0010)
	) name2926 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8753_
	);
	LUT4 #(
		.INIT('h9fe4)
	) name2927 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8754_
	);
	LUT4 #(
		.INIT('h0900)
	) name2928 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8755_
	);
	LUT4 #(
		.INIT('h0501)
	) name2929 (
		_w8697_,
		_w8707_,
		_w8755_,
		_w8754_,
		_w8756_
	);
	LUT3 #(
		.INIT('h2a)
	) name2930 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8757_
	);
	LUT4 #(
		.INIT('hae00)
	) name2931 (
		_w8692_,
		_w8693_,
		_w8694_,
		_w8707_,
		_w8758_
	);
	LUT4 #(
		.INIT('h0002)
	) name2932 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8759_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2933 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8697_,
		_w8760_
	);
	LUT4 #(
		.INIT('h4500)
	) name2934 (
		_w8759_,
		_w8757_,
		_w8758_,
		_w8760_,
		_w8761_
	);
	LUT2 #(
		.INIT('h1)
	) name2935 (
		_w8756_,
		_w8761_,
		_w8762_
	);
	LUT3 #(
		.INIT('h56)
	) name2936 (
		\u2_L9_reg[2]/NET0131 ,
		_w8751_,
		_w8762_,
		_w8763_
	);
	LUT4 #(
		.INIT('hd97b)
	) name2937 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8764_
	);
	LUT2 #(
		.INIT('h2)
	) name2938 (
		_w8450_,
		_w8764_,
		_w8765_
	);
	LUT4 #(
		.INIT('heebf)
	) name2939 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8766_
	);
	LUT4 #(
		.INIT('h0040)
	) name2940 (
		_w8450_,
		_w8447_,
		_w8452_,
		_w8448_,
		_w8767_
	);
	LUT4 #(
		.INIT('h0032)
	) name2941 (
		_w8450_,
		_w8462_,
		_w8766_,
		_w8767_,
		_w8768_
	);
	LUT3 #(
		.INIT('h45)
	) name2942 (
		_w8446_,
		_w8765_,
		_w8768_,
		_w8769_
	);
	LUT4 #(
		.INIT('h7c7f)
	) name2943 (
		_w8450_,
		_w8447_,
		_w8452_,
		_w8449_,
		_w8770_
	);
	LUT2 #(
		.INIT('h1)
	) name2944 (
		_w8448_,
		_w8770_,
		_w8771_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name2945 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8772_
	);
	LUT3 #(
		.INIT('h80)
	) name2946 (
		_w8452_,
		_w8448_,
		_w8449_,
		_w8773_
	);
	LUT3 #(
		.INIT('h0e)
	) name2947 (
		_w8450_,
		_w8772_,
		_w8773_,
		_w8774_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2948 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8775_
	);
	LUT4 #(
		.INIT('h5501)
	) name2949 (
		_w8450_,
		_w8447_,
		_w8452_,
		_w8448_,
		_w8776_
	);
	LUT3 #(
		.INIT('h9e)
	) name2950 (
		_w8447_,
		_w8452_,
		_w8449_,
		_w8777_
	);
	LUT2 #(
		.INIT('h8)
	) name2951 (
		_w8450_,
		_w8448_,
		_w8778_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2952 (
		_w8775_,
		_w8776_,
		_w8777_,
		_w8778_,
		_w8779_
	);
	LUT4 #(
		.INIT('h7500)
	) name2953 (
		_w8446_,
		_w8771_,
		_w8774_,
		_w8779_,
		_w8780_
	);
	LUT3 #(
		.INIT('h65)
	) name2954 (
		\u2_L9_reg[4]/NET0131 ,
		_w8769_,
		_w8780_,
		_w8781_
	);
	LUT3 #(
		.INIT('h02)
	) name2955 (
		_w8695_,
		_w8692_,
		_w8694_,
		_w8782_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2956 (
		_w8695_,
		_w8693_,
		_w8694_,
		_w8697_,
		_w8783_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2957 (
		_w8704_,
		_w8752_,
		_w8782_,
		_w8783_,
		_w8784_
	);
	LUT4 #(
		.INIT('h0004)
	) name2958 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8785_
	);
	LUT4 #(
		.INIT('h0002)
	) name2959 (
		_w8707_,
		_w8748_,
		_w8749_,
		_w8785_,
		_w8786_
	);
	LUT4 #(
		.INIT('h0600)
	) name2960 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8787_
	);
	LUT3 #(
		.INIT('h02)
	) name2961 (
		_w8692_,
		_w8693_,
		_w8694_,
		_w8788_
	);
	LUT2 #(
		.INIT('h1)
	) name2962 (
		_w8697_,
		_w8707_,
		_w8789_
	);
	LUT4 #(
		.INIT('h0100)
	) name2963 (
		_w8753_,
		_w8788_,
		_w8787_,
		_w8789_,
		_w8790_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name2964 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8791_
	);
	LUT4 #(
		.INIT('hf400)
	) name2965 (
		_w8784_,
		_w8786_,
		_w8790_,
		_w8791_,
		_w8792_
	);
	LUT4 #(
		.INIT('h1141)
	) name2966 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8793_
	);
	LUT4 #(
		.INIT('ha022)
	) name2967 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8794_
	);
	LUT4 #(
		.INIT('h0400)
	) name2968 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w8795_
	);
	LUT2 #(
		.INIT('h2)
	) name2969 (
		_w8697_,
		_w8707_,
		_w8796_
	);
	LUT4 #(
		.INIT('h0100)
	) name2970 (
		_w8794_,
		_w8795_,
		_w8793_,
		_w8796_,
		_w8797_
	);
	LUT3 #(
		.INIT('h56)
	) name2971 (
		\u2_L9_reg[13]/NET0131 ,
		_w8792_,
		_w8797_,
		_w8798_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name2972 (
		_w8450_,
		_w8447_,
		_w8452_,
		_w8448_,
		_w8799_
	);
	LUT4 #(
		.INIT('hef00)
	) name2973 (
		_w8452_,
		_w8448_,
		_w8449_,
		_w8446_,
		_w8800_
	);
	LUT3 #(
		.INIT('he0)
	) name2974 (
		_w8449_,
		_w8799_,
		_w8800_,
		_w8801_
	);
	LUT4 #(
		.INIT('h4010)
	) name2975 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8802_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name2976 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8803_
	);
	LUT3 #(
		.INIT('h31)
	) name2977 (
		_w8450_,
		_w8802_,
		_w8803_,
		_w8804_
	);
	LUT4 #(
		.INIT('h4e55)
	) name2978 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8805_
	);
	LUT2 #(
		.INIT('h2)
	) name2979 (
		_w8450_,
		_w8805_,
		_w8806_
	);
	LUT4 #(
		.INIT('h1001)
	) name2980 (
		_w8450_,
		_w8447_,
		_w8452_,
		_w8449_,
		_w8807_
	);
	LUT4 #(
		.INIT('h8000)
	) name2981 (
		_w8447_,
		_w8452_,
		_w8448_,
		_w8449_,
		_w8808_
	);
	LUT3 #(
		.INIT('h01)
	) name2982 (
		_w8446_,
		_w8808_,
		_w8807_,
		_w8809_
	);
	LUT4 #(
		.INIT('h7077)
	) name2983 (
		_w8801_,
		_w8804_,
		_w8806_,
		_w8809_,
		_w8810_
	);
	LUT2 #(
		.INIT('h4)
	) name2984 (
		_w8449_,
		_w8767_,
		_w8811_
	);
	LUT2 #(
		.INIT('h1)
	) name2985 (
		_w8470_,
		_w8811_,
		_w8812_
	);
	LUT3 #(
		.INIT('h65)
	) name2986 (
		\u2_L9_reg[19]/NET0131 ,
		_w8810_,
		_w8812_,
		_w8813_
	);
	LUT4 #(
		.INIT('h8088)
	) name2987 (
		_w8414_,
		_w8418_,
		_w8416_,
		_w8419_,
		_w8814_
	);
	LUT2 #(
		.INIT('h8)
	) name2988 (
		_w8631_,
		_w8814_,
		_w8815_
	);
	LUT4 #(
		.INIT('h020a)
	) name2989 (
		_w8415_,
		_w8435_,
		_w8438_,
		_w8442_,
		_w8816_
	);
	LUT4 #(
		.INIT('habbb)
	) name2990 (
		_w8414_,
		_w8418_,
		_w8417_,
		_w8416_,
		_w8817_
	);
	LUT2 #(
		.INIT('h2)
	) name2991 (
		_w8419_,
		_w8817_,
		_w8818_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2992 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8415_,
		_w8819_
	);
	LUT4 #(
		.INIT('h0008)
	) name2993 (
		_w8414_,
		_w8418_,
		_w8417_,
		_w8419_,
		_w8820_
	);
	LUT4 #(
		.INIT('h0100)
	) name2994 (
		_w8436_,
		_w8421_,
		_w8820_,
		_w8819_,
		_w8821_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2995 (
		_w8815_,
		_w8816_,
		_w8818_,
		_w8821_,
		_w8822_
	);
	LUT4 #(
		.INIT('hef99)
	) name2996 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8823_
	);
	LUT4 #(
		.INIT('hfdfb)
	) name2997 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8824_
	);
	LUT4 #(
		.INIT('h0455)
	) name2998 (
		_w8414_,
		_w8415_,
		_w8823_,
		_w8824_,
		_w8825_
	);
	LUT3 #(
		.INIT('had)
	) name2999 (
		_w8418_,
		_w8417_,
		_w8419_,
		_w8826_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name3000 (
		_w8414_,
		_w8416_,
		_w8633_,
		_w8826_,
		_w8827_
	);
	LUT2 #(
		.INIT('h4)
	) name3001 (
		_w8825_,
		_w8827_,
		_w8828_
	);
	LUT3 #(
		.INIT('h9a)
	) name3002 (
		\u2_L9_reg[23]/NET0131 ,
		_w8822_,
		_w8828_,
		_w8829_
	);
	LUT4 #(
		.INIT('hba76)
	) name3003 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8830_
	);
	LUT2 #(
		.INIT('h1)
	) name3004 (
		_w8514_,
		_w8830_,
		_w8831_
	);
	LUT3 #(
		.INIT('hd0)
	) name3005 (
		_w8517_,
		_w8515_,
		_w8514_,
		_w8832_
	);
	LUT4 #(
		.INIT('hbcdf)
	) name3006 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8833_
	);
	LUT3 #(
		.INIT('hb0)
	) name3007 (
		_w8604_,
		_w8832_,
		_w8833_,
		_w8834_
	);
	LUT3 #(
		.INIT('h8a)
	) name3008 (
		_w8527_,
		_w8831_,
		_w8834_,
		_w8835_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3009 (
		_w8518_,
		_w8516_,
		_w8515_,
		_w8514_,
		_w8836_
	);
	LUT4 #(
		.INIT('h0cbf)
	) name3010 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8837_
	);
	LUT2 #(
		.INIT('h8)
	) name3011 (
		_w8836_,
		_w8837_,
		_w8838_
	);
	LUT4 #(
		.INIT('h0080)
	) name3012 (
		_w8517_,
		_w8516_,
		_w8515_,
		_w8514_,
		_w8839_
	);
	LUT3 #(
		.INIT('h01)
	) name3013 (
		_w8536_,
		_w8670_,
		_w8839_,
		_w8840_
	);
	LUT3 #(
		.INIT('h45)
	) name3014 (
		_w8527_,
		_w8838_,
		_w8840_,
		_w8841_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name3015 (
		_w8517_,
		_w8518_,
		_w8516_,
		_w8515_,
		_w8842_
	);
	LUT2 #(
		.INIT('h1)
	) name3016 (
		_w8514_,
		_w8842_,
		_w8843_
	);
	LUT4 #(
		.INIT('h0400)
	) name3017 (
		_w8518_,
		_w8516_,
		_w8515_,
		_w8514_,
		_w8844_
	);
	LUT3 #(
		.INIT('h07)
	) name3018 (
		_w8522_,
		_w8540_,
		_w8844_,
		_w8845_
	);
	LUT2 #(
		.INIT('h4)
	) name3019 (
		_w8843_,
		_w8845_,
		_w8846_
	);
	LUT4 #(
		.INIT('h5655)
	) name3020 (
		\u2_L9_reg[27]/NET0131 ,
		_w8835_,
		_w8841_,
		_w8846_,
		_w8847_
	);
	LUT3 #(
		.INIT('hca)
	) name3021 (
		_w8385_,
		_w8387_,
		_w8388_,
		_w8848_
	);
	LUT4 #(
		.INIT('hbb50)
	) name3022 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8849_
	);
	LUT4 #(
		.INIT('hccc4)
	) name3023 (
		_w8387_,
		_w8384_,
		_w8386_,
		_w8388_,
		_w8850_
	);
	LUT2 #(
		.INIT('h4)
	) name3024 (
		_w8849_,
		_w8850_,
		_w8851_
	);
	LUT4 #(
		.INIT('h0080)
	) name3025 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8852_
	);
	LUT4 #(
		.INIT('hdee3)
	) name3026 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8853_
	);
	LUT3 #(
		.INIT('h32)
	) name3027 (
		_w8384_,
		_w8852_,
		_w8853_,
		_w8854_
	);
	LUT3 #(
		.INIT('h8a)
	) name3028 (
		_w8383_,
		_w8851_,
		_w8854_,
		_w8855_
	);
	LUT3 #(
		.INIT('h04)
	) name3029 (
		_w8385_,
		_w8386_,
		_w8388_,
		_w8856_
	);
	LUT2 #(
		.INIT('h2)
	) name3030 (
		_w8570_,
		_w8856_,
		_w8857_
	);
	LUT4 #(
		.INIT('h8040)
	) name3031 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8858_
	);
	LUT4 #(
		.INIT('h00c4)
	) name3032 (
		_w8394_,
		_w8407_,
		_w8848_,
		_w8858_,
		_w8859_
	);
	LUT4 #(
		.INIT('h0c08)
	) name3033 (
		_w8385_,
		_w8387_,
		_w8384_,
		_w8388_,
		_w8860_
	);
	LUT4 #(
		.INIT('h135f)
	) name3034 (
		_w8384_,
		_w8400_,
		_w8396_,
		_w8860_,
		_w8861_
	);
	LUT4 #(
		.INIT('hba00)
	) name3035 (
		_w8383_,
		_w8857_,
		_w8859_,
		_w8861_,
		_w8862_
	);
	LUT3 #(
		.INIT('h65)
	) name3036 (
		\u2_L9_reg[32]/NET0131 ,
		_w8855_,
		_w8862_,
		_w8863_
	);
	LUT4 #(
		.INIT('hc963)
	) name3037 (
		decrypt_pad,
		\u2_R9_reg[12]/NET0131 ,
		\u2_uk_K_r9_reg[4]/NET0131 ,
		\u2_uk_K_r9_reg[55]/NET0131 ,
		_w8864_
	);
	LUT4 #(
		.INIT('hc693)
	) name3038 (
		decrypt_pad,
		\u2_R9_reg[13]/NET0131 ,
		\u2_uk_K_r9_reg[11]/NET0131 ,
		\u2_uk_K_r9_reg[17]/NET0131 ,
		_w8865_
	);
	LUT4 #(
		.INIT('hc693)
	) name3039 (
		decrypt_pad,
		\u2_R9_reg[8]/NET0131 ,
		\u2_uk_K_r9_reg[34]/NET0131 ,
		\u2_uk_K_r9_reg[40]/NET0131 ,
		_w8866_
	);
	LUT2 #(
		.INIT('h6)
	) name3040 (
		_w8865_,
		_w8866_,
		_w8867_
	);
	LUT4 #(
		.INIT('hc963)
	) name3041 (
		decrypt_pad,
		\u2_R9_reg[9]/NET0131 ,
		\u2_uk_K_r9_reg[12]/NET0131 ,
		\u2_uk_K_r9_reg[6]/NET0131 ,
		_w8868_
	);
	LUT4 #(
		.INIT('hc963)
	) name3042 (
		decrypt_pad,
		\u2_R9_reg[10]/NET0131 ,
		\u2_uk_K_r9_reg[20]/NET0131 ,
		\u2_uk_K_r9_reg[39]/NET0131 ,
		_w8869_
	);
	LUT4 #(
		.INIT('h2100)
	) name3043 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8870_
	);
	LUT3 #(
		.INIT('h08)
	) name3044 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8871_
	);
	LUT4 #(
		.INIT('hc693)
	) name3045 (
		decrypt_pad,
		\u2_R9_reg[11]/NET0131 ,
		\u2_uk_K_r9_reg[40]/NET0131 ,
		\u2_uk_K_r9_reg[46]/NET0131 ,
		_w8872_
	);
	LUT2 #(
		.INIT('h2)
	) name3046 (
		_w8869_,
		_w8872_,
		_w8873_
	);
	LUT3 #(
		.INIT('h40)
	) name3047 (
		_w8865_,
		_w8868_,
		_w8869_,
		_w8874_
	);
	LUT4 #(
		.INIT('h4000)
	) name3048 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8875_
	);
	LUT4 #(
		.INIT('h0007)
	) name3049 (
		_w8871_,
		_w8873_,
		_w8875_,
		_w8870_,
		_w8876_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		_w8865_,
		_w8872_,
		_w8877_
	);
	LUT3 #(
		.INIT('h46)
	) name3051 (
		_w8865_,
		_w8866_,
		_w8872_,
		_w8878_
	);
	LUT2 #(
		.INIT('h1)
	) name3052 (
		_w8868_,
		_w8869_,
		_w8879_
	);
	LUT2 #(
		.INIT('h8)
	) name3053 (
		_w8879_,
		_w8878_,
		_w8880_
	);
	LUT3 #(
		.INIT('hed)
	) name3054 (
		_w8868_,
		_w8869_,
		_w8878_,
		_w8881_
	);
	LUT3 #(
		.INIT('h15)
	) name3055 (
		_w8864_,
		_w8876_,
		_w8881_,
		_w8882_
	);
	LUT4 #(
		.INIT('h959d)
	) name3056 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8883_
	);
	LUT4 #(
		.INIT('h0001)
	) name3057 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8884_
	);
	LUT4 #(
		.INIT('hddfe)
	) name3058 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8885_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3059 (
		_w8883_,
		_w8864_,
		_w8885_,
		_w8872_,
		_w8886_
	);
	LUT2 #(
		.INIT('h8)
	) name3060 (
		_w8869_,
		_w8864_,
		_w8887_
	);
	LUT3 #(
		.INIT('h04)
	) name3061 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8888_
	);
	LUT2 #(
		.INIT('h2)
	) name3062 (
		_w8864_,
		_w8872_,
		_w8889_
	);
	LUT3 #(
		.INIT('h80)
	) name3063 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8890_
	);
	LUT4 #(
		.INIT('h6f67)
	) name3064 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8891_
	);
	LUT4 #(
		.INIT('h7707)
	) name3065 (
		_w8887_,
		_w8888_,
		_w8889_,
		_w8891_,
		_w8892_
	);
	LUT2 #(
		.INIT('h4)
	) name3066 (
		_w8886_,
		_w8892_,
		_w8893_
	);
	LUT3 #(
		.INIT('h65)
	) name3067 (
		\u2_L9_reg[6]/NET0131 ,
		_w8882_,
		_w8893_,
		_w8894_
	);
	LUT4 #(
		.INIT('hf216)
	) name3068 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8895_
	);
	LUT4 #(
		.INIT('h2880)
	) name3069 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8896_
	);
	LUT4 #(
		.INIT('h5004)
	) name3070 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8897_
	);
	LUT4 #(
		.INIT('h1032)
	) name3071 (
		_w8384_,
		_w8896_,
		_w8895_,
		_w8897_,
		_w8898_
	);
	LUT2 #(
		.INIT('h2)
	) name3072 (
		_w8383_,
		_w8898_,
		_w8899_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name3073 (
		_w8384_,
		_w8401_,
		_w8383_,
		_w8897_,
		_w8900_
	);
	LUT2 #(
		.INIT('h4)
	) name3074 (
		_w8384_,
		_w8896_,
		_w8901_
	);
	LUT4 #(
		.INIT('h0880)
	) name3075 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8902_
	);
	LUT2 #(
		.INIT('h2)
	) name3076 (
		_w8384_,
		_w8902_,
		_w8903_
	);
	LUT4 #(
		.INIT('h7005)
	) name3077 (
		_w8385_,
		_w8387_,
		_w8386_,
		_w8388_,
		_w8904_
	);
	LUT3 #(
		.INIT('h0b)
	) name3078 (
		_w8401_,
		_w8383_,
		_w8904_,
		_w8905_
	);
	LUT4 #(
		.INIT('h0111)
	) name3079 (
		_w8901_,
		_w8900_,
		_w8903_,
		_w8905_,
		_w8906_
	);
	LUT3 #(
		.INIT('h65)
	) name3080 (
		\u2_L9_reg[7]/NET0131 ,
		_w8899_,
		_w8906_,
		_w8907_
	);
	LUT4 #(
		.INIT('h0010)
	) name3081 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8908_
	);
	LUT4 #(
		.INIT('h5fef)
	) name3082 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8909_
	);
	LUT4 #(
		.INIT('ha4ff)
	) name3083 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8910_
	);
	LUT4 #(
		.INIT('hfd79)
	) name3084 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8911_
	);
	LUT4 #(
		.INIT('hd800)
	) name3085 (
		_w8582_,
		_w8909_,
		_w8910_,
		_w8911_,
		_w8912_
	);
	LUT4 #(
		.INIT('haffe)
	) name3086 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8913_
	);
	LUT3 #(
		.INIT('h04)
	) name3087 (
		_w8575_,
		_w8577_,
		_w8582_,
		_w8914_
	);
	LUT4 #(
		.INIT('h0031)
	) name3088 (
		_w8582_,
		_w8599_,
		_w8913_,
		_w8914_,
		_w8915_
	);
	LUT4 #(
		.INIT('hf977)
	) name3089 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8916_
	);
	LUT4 #(
		.INIT('h5f13)
	) name3090 (
		_w8579_,
		_w8582_,
		_w8687_,
		_w8916_,
		_w8917_
	);
	LUT4 #(
		.INIT('he400)
	) name3091 (
		_w8574_,
		_w8912_,
		_w8915_,
		_w8917_,
		_w8918_
	);
	LUT2 #(
		.INIT('h9)
	) name3092 (
		\u2_L9_reg[8]/NET0131 ,
		_w8918_,
		_w8919_
	);
	LUT4 #(
		.INIT('hf700)
	) name3093 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8920_
	);
	LUT4 #(
		.INIT('h0400)
	) name3094 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8872_,
		_w8921_
	);
	LUT4 #(
		.INIT('h006d)
	) name3095 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8922_
	);
	LUT3 #(
		.INIT('h45)
	) name3096 (
		_w8920_,
		_w8921_,
		_w8922_,
		_w8923_
	);
	LUT4 #(
		.INIT('h0100)
	) name3097 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8924_
	);
	LUT3 #(
		.INIT('h14)
	) name3098 (
		_w8865_,
		_w8866_,
		_w8869_,
		_w8925_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3099 (
		_w8872_,
		_w8875_,
		_w8924_,
		_w8925_,
		_w8926_
	);
	LUT3 #(
		.INIT('ha8)
	) name3100 (
		_w8864_,
		_w8923_,
		_w8926_,
		_w8927_
	);
	LUT3 #(
		.INIT('h40)
	) name3101 (
		_w8868_,
		_w8866_,
		_w8869_,
		_w8928_
	);
	LUT4 #(
		.INIT('h00bf)
	) name3102 (
		_w8868_,
		_w8866_,
		_w8869_,
		_w8872_,
		_w8929_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3103 (
		_w8872_,
		_w8875_,
		_w8924_,
		_w8929_,
		_w8930_
	);
	LUT4 #(
		.INIT('h7d78)
	) name3104 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8931_
	);
	LUT3 #(
		.INIT('he0)
	) name3105 (
		_w8865_,
		_w8866_,
		_w8872_,
		_w8932_
	);
	LUT4 #(
		.INIT('h6800)
	) name3106 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8872_,
		_w8933_
	);
	LUT4 #(
		.INIT('h0504)
	) name3107 (
		_w8884_,
		_w8872_,
		_w8933_,
		_w8931_,
		_w8934_
	);
	LUT3 #(
		.INIT('h32)
	) name3108 (
		_w8864_,
		_w8930_,
		_w8934_,
		_w8935_
	);
	LUT3 #(
		.INIT('h65)
	) name3109 (
		\u2_L9_reg[16]/NET0131 ,
		_w8927_,
		_w8935_,
		_w8936_
	);
	LUT2 #(
		.INIT('h4)
	) name3110 (
		_w8869_,
		_w8872_,
		_w8937_
	);
	LUT3 #(
		.INIT('h31)
	) name3111 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8938_
	);
	LUT2 #(
		.INIT('h8)
	) name3112 (
		_w8937_,
		_w8938_,
		_w8939_
	);
	LUT3 #(
		.INIT('h0e)
	) name3113 (
		_w8868_,
		_w8869_,
		_w8872_,
		_w8940_
	);
	LUT3 #(
		.INIT('hb0)
	) name3114 (
		_w8868_,
		_w8866_,
		_w8869_,
		_w8941_
	);
	LUT4 #(
		.INIT('h23af)
	) name3115 (
		_w8867_,
		_w8932_,
		_w8940_,
		_w8941_,
		_w8942_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3116 (
		_w8864_,
		_w8880_,
		_w8939_,
		_w8942_,
		_w8943_
	);
	LUT4 #(
		.INIT('hcaf1)
	) name3117 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8944_
	);
	LUT4 #(
		.INIT('h1000)
	) name3118 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8945_
	);
	LUT4 #(
		.INIT('h5504)
	) name3119 (
		_w8864_,
		_w8872_,
		_w8944_,
		_w8945_,
		_w8946_
	);
	LUT4 #(
		.INIT('h0021)
	) name3120 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8947_
	);
	LUT4 #(
		.INIT('hb59e)
	) name3121 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8948_
	);
	LUT2 #(
		.INIT('h1)
	) name3122 (
		_w8864_,
		_w8872_,
		_w8949_
	);
	LUT2 #(
		.INIT('h4)
	) name3123 (
		_w8948_,
		_w8949_,
		_w8950_
	);
	LUT3 #(
		.INIT('he7)
	) name3124 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8951_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name3125 (
		_w8869_,
		_w8872_,
		_w8890_,
		_w8951_,
		_w8952_
	);
	LUT3 #(
		.INIT('h10)
	) name3126 (
		_w8946_,
		_w8950_,
		_w8952_,
		_w8953_
	);
	LUT3 #(
		.INIT('h65)
	) name3127 (
		\u2_L9_reg[24]/NET0131 ,
		_w8943_,
		_w8953_,
		_w8954_
	);
	LUT4 #(
		.INIT('hfae5)
	) name3128 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8955_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3129 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8956_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name3130 (
		_w8864_,
		_w8874_,
		_w8955_,
		_w8956_,
		_w8957_
	);
	LUT2 #(
		.INIT('h2)
	) name3131 (
		_w8872_,
		_w8957_,
		_w8958_
	);
	LUT4 #(
		.INIT('h0200)
	) name3132 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8959_
	);
	LUT3 #(
		.INIT('h0e)
	) name3133 (
		_w8868_,
		_w8866_,
		_w8872_,
		_w8960_
	);
	LUT4 #(
		.INIT('h0015)
	) name3134 (
		_w8947_,
		_w8956_,
		_w8960_,
		_w8959_,
		_w8961_
	);
	LUT2 #(
		.INIT('h1)
	) name3135 (
		_w8864_,
		_w8961_,
		_w8962_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name3136 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8869_,
		_w8963_
	);
	LUT2 #(
		.INIT('h2)
	) name3137 (
		_w8889_,
		_w8963_,
		_w8964_
	);
	LUT3 #(
		.INIT('h4c)
	) name3138 (
		_w8865_,
		_w8868_,
		_w8866_,
		_w8965_
	);
	LUT2 #(
		.INIT('h8)
	) name3139 (
		_w8887_,
		_w8965_,
		_w8966_
	);
	LUT4 #(
		.INIT('h0040)
	) name3140 (
		_w8865_,
		_w8868_,
		_w8869_,
		_w8872_,
		_w8967_
	);
	LUT3 #(
		.INIT('h07)
	) name3141 (
		_w8877_,
		_w8928_,
		_w8967_,
		_w8968_
	);
	LUT3 #(
		.INIT('h10)
	) name3142 (
		_w8964_,
		_w8966_,
		_w8968_,
		_w8969_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name3143 (
		\u2_L9_reg[30]/NET0131 ,
		_w8958_,
		_w8962_,
		_w8969_,
		_w8970_
	);
	LUT4 #(
		.INIT('h2a00)
	) name3144 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8971_
	);
	LUT4 #(
		.INIT('h0040)
	) name3145 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8972_
	);
	LUT3 #(
		.INIT('h02)
	) name3146 (
		_w8574_,
		_w8971_,
		_w8972_,
		_w8973_
	);
	LUT4 #(
		.INIT('h4404)
	) name3147 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8974_
	);
	LUT4 #(
		.INIT('h23f0)
	) name3148 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8975_
	);
	LUT3 #(
		.INIT('h10)
	) name3149 (
		_w8574_,
		_w8974_,
		_w8975_,
		_w8976_
	);
	LUT4 #(
		.INIT('hffde)
	) name3150 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8977_
	);
	LUT3 #(
		.INIT('h10)
	) name3151 (
		_w8582_,
		_w8588_,
		_w8977_,
		_w8978_
	);
	LUT3 #(
		.INIT('he0)
	) name3152 (
		_w8973_,
		_w8976_,
		_w8978_,
		_w8979_
	);
	LUT4 #(
		.INIT('hcff5)
	) name3153 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8980_
	);
	LUT3 #(
		.INIT('h20)
	) name3154 (
		_w8574_,
		_w8972_,
		_w8980_,
		_w8981_
	);
	LUT4 #(
		.INIT('hfc5f)
	) name3155 (
		_w8576_,
		_w8575_,
		_w8577_,
		_w8578_,
		_w8982_
	);
	LUT3 #(
		.INIT('h10)
	) name3156 (
		_w8574_,
		_w8974_,
		_w8982_,
		_w8983_
	);
	LUT3 #(
		.INIT('h02)
	) name3157 (
		_w8582_,
		_w8598_,
		_w8908_,
		_w8984_
	);
	LUT3 #(
		.INIT('he0)
	) name3158 (
		_w8981_,
		_w8983_,
		_w8984_,
		_w8985_
	);
	LUT3 #(
		.INIT('ha9)
	) name3159 (
		\u2_L9_reg[3]/NET0131 ,
		_w8979_,
		_w8985_,
		_w8986_
	);
	LUT4 #(
		.INIT('h9b99)
	) name3160 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8987_
	);
	LUT3 #(
		.INIT('h19)
	) name3161 (
		_w8418_,
		_w8417_,
		_w8419_,
		_w8988_
	);
	LUT4 #(
		.INIT('h4810)
	) name3162 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8989_
	);
	LUT4 #(
		.INIT('h0b01)
	) name3163 (
		_w8414_,
		_w8988_,
		_w8989_,
		_w8987_,
		_w8990_
	);
	LUT4 #(
		.INIT('hf77f)
	) name3164 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8991_
	);
	LUT2 #(
		.INIT('h1)
	) name3165 (
		_w8414_,
		_w8991_,
		_w8992_
	);
	LUT4 #(
		.INIT('h9060)
	) name3166 (
		_w8418_,
		_w8417_,
		_w8416_,
		_w8419_,
		_w8993_
	);
	LUT4 #(
		.INIT('h0013)
	) name3167 (
		_w8428_,
		_w8625_,
		_w8988_,
		_w8993_,
		_w8994_
	);
	LUT4 #(
		.INIT('h0e04)
	) name3168 (
		_w8415_,
		_w8990_,
		_w8992_,
		_w8994_,
		_w8995_
	);
	LUT2 #(
		.INIT('h9)
	) name3169 (
		\u2_L9_reg[9]/NET0131 ,
		_w8995_,
		_w8996_
	);
	LUT4 #(
		.INIT('h1a00)
	) name3170 (
		_w8692_,
		_w8693_,
		_w8694_,
		_w8697_,
		_w8997_
	);
	LUT2 #(
		.INIT('h8)
	) name3171 (
		_w8695_,
		_w8694_,
		_w8998_
	);
	LUT4 #(
		.INIT('h00c4)
	) name3172 (
		_w8692_,
		_w8693_,
		_w8694_,
		_w8697_,
		_w8999_
	);
	LUT4 #(
		.INIT('h2022)
	) name3173 (
		_w8707_,
		_w8759_,
		_w8998_,
		_w8999_,
		_w9000_
	);
	LUT2 #(
		.INIT('h2)
	) name3174 (
		_w8692_,
		_w8697_,
		_w9001_
	);
	LUT4 #(
		.INIT('he000)
	) name3175 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w9002_
	);
	LUT4 #(
		.INIT('h0109)
	) name3176 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8697_,
		_w9003_
	);
	LUT4 #(
		.INIT('h0405)
	) name3177 (
		_w8752_,
		_w9001_,
		_w9003_,
		_w9002_,
		_w9004_
	);
	LUT4 #(
		.INIT('h45cf)
	) name3178 (
		_w8714_,
		_w8997_,
		_w9000_,
		_w9004_,
		_w9005_
	);
	LUT4 #(
		.INIT('h0020)
	) name3179 (
		_w8692_,
		_w8693_,
		_w8694_,
		_w8697_,
		_w9006_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name3180 (
		_w8695_,
		_w8692_,
		_w8693_,
		_w8694_,
		_w9007_
	);
	LUT3 #(
		.INIT('h31)
	) name3181 (
		_w8697_,
		_w9006_,
		_w9007_,
		_w9008_
	);
	LUT3 #(
		.INIT('h65)
	) name3182 (
		\u2_L9_reg[18]/P0001 ,
		_w9005_,
		_w9008_,
		_w9009_
	);
	LUT4 #(
		.INIT('hc963)
	) name3183 (
		decrypt_pad,
		\u2_R8_reg[4]/NET0131 ,
		\u2_uk_K_r8_reg[11]/NET0131 ,
		\u2_uk_K_r8_reg[33]/NET0131 ,
		_w9010_
	);
	LUT4 #(
		.INIT('hc963)
	) name3184 (
		decrypt_pad,
		\u2_R8_reg[2]/NET0131 ,
		\u2_uk_K_r8_reg[24]/NET0131 ,
		\u2_uk_K_r8_reg[46]/NET0131 ,
		_w9011_
	);
	LUT4 #(
		.INIT('hc963)
	) name3185 (
		decrypt_pad,
		\u2_R8_reg[5]/NET0131 ,
		\u2_uk_K_r8_reg[39]/NET0131 ,
		\u2_uk_K_r8_reg[4]/NET0131 ,
		_w9012_
	);
	LUT2 #(
		.INIT('h6)
	) name3186 (
		_w9011_,
		_w9012_,
		_w9013_
	);
	LUT4 #(
		.INIT('hc963)
	) name3187 (
		decrypt_pad,
		\u2_R8_reg[3]/NET0131 ,
		\u2_uk_K_r8_reg[33]/NET0131 ,
		\u2_uk_K_r8_reg[55]/NET0131 ,
		_w9014_
	);
	LUT4 #(
		.INIT('hc693)
	) name3188 (
		decrypt_pad,
		\u2_R8_reg[32]/NET0131 ,
		\u2_uk_K_r8_reg[10]/NET0131 ,
		\u2_uk_K_r8_reg[20]/NET0131 ,
		_w9015_
	);
	LUT4 #(
		.INIT('hc963)
	) name3189 (
		decrypt_pad,
		\u2_R8_reg[1]/NET0131 ,
		\u2_uk_K_r8_reg[41]/NET0131 ,
		\u2_uk_K_r8_reg[6]/NET0131 ,
		_w9016_
	);
	LUT4 #(
		.INIT('h4044)
	) name3190 (
		_w9015_,
		_w9016_,
		_w9014_,
		_w9012_,
		_w9017_
	);
	LUT2 #(
		.INIT('h4)
	) name3191 (
		_w9013_,
		_w9017_,
		_w9018_
	);
	LUT4 #(
		.INIT('h0080)
	) name3192 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9019_
	);
	LUT2 #(
		.INIT('h2)
	) name3193 (
		_w9016_,
		_w9014_,
		_w9020_
	);
	LUT3 #(
		.INIT('h20)
	) name3194 (
		_w9015_,
		_w9011_,
		_w9012_,
		_w9021_
	);
	LUT4 #(
		.INIT('h223f)
	) name3195 (
		_w9016_,
		_w9014_,
		_w9019_,
		_w9021_,
		_w9022_
	);
	LUT2 #(
		.INIT('h4)
	) name3196 (
		_w9011_,
		_w9014_,
		_w9023_
	);
	LUT4 #(
		.INIT('h0200)
	) name3197 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9014_,
		_w9024_
	);
	LUT2 #(
		.INIT('h1)
	) name3198 (
		_w9016_,
		_w9012_,
		_w9025_
	);
	LUT3 #(
		.INIT('h40)
	) name3199 (
		_w9015_,
		_w9011_,
		_w9014_,
		_w9026_
	);
	LUT3 #(
		.INIT('h15)
	) name3200 (
		_w9024_,
		_w9025_,
		_w9026_,
		_w9027_
	);
	LUT4 #(
		.INIT('hba00)
	) name3201 (
		_w9010_,
		_w9018_,
		_w9022_,
		_w9027_,
		_w9028_
	);
	LUT4 #(
		.INIT('hfbda)
	) name3202 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9029_
	);
	LUT4 #(
		.INIT('h1000)
	) name3203 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9030_
	);
	LUT4 #(
		.INIT('h6ff3)
	) name3204 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9031_
	);
	LUT4 #(
		.INIT('h0155)
	) name3205 (
		_w9014_,
		_w9010_,
		_w9029_,
		_w9031_,
		_w9032_
	);
	LUT4 #(
		.INIT('h75c4)
	) name3206 (
		_w9016_,
		_w9011_,
		_w9014_,
		_w9012_,
		_w9033_
	);
	LUT2 #(
		.INIT('h1)
	) name3207 (
		_w9015_,
		_w9033_,
		_w9034_
	);
	LUT4 #(
		.INIT('h5011)
	) name3208 (
		_w9016_,
		_w9011_,
		_w9014_,
		_w9012_,
		_w9035_
	);
	LUT3 #(
		.INIT('ha2)
	) name3209 (
		_w9015_,
		_w9016_,
		_w9014_,
		_w9036_
	);
	LUT3 #(
		.INIT('h8a)
	) name3210 (
		_w9010_,
		_w9035_,
		_w9036_,
		_w9037_
	);
	LUT3 #(
		.INIT('h45)
	) name3211 (
		_w9032_,
		_w9034_,
		_w9037_,
		_w9038_
	);
	LUT3 #(
		.INIT('h95)
	) name3212 (
		\u2_L8_reg[31]/NET0131 ,
		_w9028_,
		_w9038_,
		_w9039_
	);
	LUT4 #(
		.INIT('hc693)
	) name3213 (
		decrypt_pad,
		\u2_R8_reg[24]/NET0131 ,
		\u2_uk_K_r8_reg[2]/NET0131 ,
		\u2_uk_K_r8_reg[37]/P0001 ,
		_w9040_
	);
	LUT4 #(
		.INIT('hc963)
	) name3214 (
		decrypt_pad,
		\u2_R8_reg[20]/NET0131 ,
		\u2_uk_K_r8_reg[16]/NET0131 ,
		\u2_uk_K_r8_reg[36]/NET0131 ,
		_w9041_
	);
	LUT4 #(
		.INIT('hc963)
	) name3215 (
		decrypt_pad,
		\u2_R8_reg[22]/NET0131 ,
		\u2_uk_K_r8_reg[22]/NET0131 ,
		\u2_uk_K_r8_reg[42]/NET0131 ,
		_w9042_
	);
	LUT4 #(
		.INIT('hc963)
	) name3216 (
		decrypt_pad,
		\u2_R8_reg[21]/NET0131 ,
		\u2_uk_K_r8_reg[0]/NET0131 ,
		\u2_uk_K_r8_reg[51]/NET0131 ,
		_w9043_
	);
	LUT4 #(
		.INIT('hc693)
	) name3217 (
		decrypt_pad,
		\u2_R8_reg[23]/NET0131 ,
		\u2_uk_K_r8_reg[0]/NET0131 ,
		\u2_uk_K_r8_reg[35]/NET0131 ,
		_w9044_
	);
	LUT4 #(
		.INIT('h4155)
	) name3218 (
		_w9044_,
		_w9041_,
		_w9042_,
		_w9043_,
		_w9045_
	);
	LUT4 #(
		.INIT('hc963)
	) name3219 (
		decrypt_pad,
		\u2_R8_reg[25]/NET0131 ,
		\u2_uk_K_r8_reg[1]/NET0131 ,
		\u2_uk_K_r8_reg[21]/NET0131 ,
		_w9046_
	);
	LUT4 #(
		.INIT('haa8a)
	) name3220 (
		_w9044_,
		_w9041_,
		_w9046_,
		_w9043_,
		_w9047_
	);
	LUT3 #(
		.INIT('he6)
	) name3221 (
		_w9041_,
		_w9042_,
		_w9043_,
		_w9048_
	);
	LUT3 #(
		.INIT('h13)
	) name3222 (
		_w9047_,
		_w9045_,
		_w9048_,
		_w9049_
	);
	LUT4 #(
		.INIT('h0080)
	) name3223 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9050_
	);
	LUT2 #(
		.INIT('h2)
	) name3224 (
		_w9041_,
		_w9046_,
		_w9051_
	);
	LUT2 #(
		.INIT('h1)
	) name3225 (
		_w9044_,
		_w9042_,
		_w9052_
	);
	LUT3 #(
		.INIT('hce)
	) name3226 (
		_w9044_,
		_w9042_,
		_w9043_,
		_w9053_
	);
	LUT3 #(
		.INIT('h31)
	) name3227 (
		_w9051_,
		_w9050_,
		_w9053_,
		_w9054_
	);
	LUT3 #(
		.INIT('h45)
	) name3228 (
		_w9040_,
		_w9049_,
		_w9054_,
		_w9055_
	);
	LUT4 #(
		.INIT('h0002)
	) name3229 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9056_
	);
	LUT4 #(
		.INIT('h27fd)
	) name3230 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9057_
	);
	LUT2 #(
		.INIT('h2)
	) name3231 (
		_w9044_,
		_w9057_,
		_w9058_
	);
	LUT4 #(
		.INIT('h0415)
	) name3232 (
		_w9044_,
		_w9041_,
		_w9046_,
		_w9043_,
		_w9059_
	);
	LUT4 #(
		.INIT('h0b07)
	) name3233 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9060_
	);
	LUT3 #(
		.INIT('h0e)
	) name3234 (
		_w9052_,
		_w9059_,
		_w9060_,
		_w9061_
	);
	LUT3 #(
		.INIT('he0)
	) name3235 (
		_w9058_,
		_w9061_,
		_w9040_,
		_w9062_
	);
	LUT4 #(
		.INIT('h5155)
	) name3236 (
		_w9044_,
		_w9041_,
		_w9046_,
		_w9043_,
		_w9063_
	);
	LUT3 #(
		.INIT('h01)
	) name3237 (
		_w9042_,
		_w9063_,
		_w9047_,
		_w9064_
	);
	LUT4 #(
		.INIT('h7077)
	) name3238 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9065_
	);
	LUT4 #(
		.INIT('haa02)
	) name3239 (
		_w9044_,
		_w9041_,
		_w9046_,
		_w9042_,
		_w9066_
	);
	LUT3 #(
		.INIT('h01)
	) name3240 (
		_w9041_,
		_w9046_,
		_w9043_,
		_w9067_
	);
	LUT4 #(
		.INIT('h45cf)
	) name3241 (
		_w9052_,
		_w9065_,
		_w9066_,
		_w9067_,
		_w9068_
	);
	LUT2 #(
		.INIT('h4)
	) name3242 (
		_w9064_,
		_w9068_,
		_w9069_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name3243 (
		\u2_L8_reg[11]/NET0131 ,
		_w9062_,
		_w9055_,
		_w9069_,
		_w9070_
	);
	LUT4 #(
		.INIT('hc693)
	) name3244 (
		decrypt_pad,
		\u2_R8_reg[27]/NET0131 ,
		\u2_uk_K_r8_reg[22]/NET0131 ,
		\u2_uk_K_r8_reg[2]/NET0131 ,
		_w9071_
	);
	LUT4 #(
		.INIT('hc963)
	) name3245 (
		decrypt_pad,
		\u2_R8_reg[24]/NET0131 ,
		\u2_uk_K_r8_reg[28]/NET0131 ,
		\u2_uk_K_r8_reg[52]/NET0131 ,
		_w9072_
	);
	LUT4 #(
		.INIT('hc693)
	) name3246 (
		decrypt_pad,
		\u2_R8_reg[25]/NET0131 ,
		\u2_uk_K_r8_reg[28]/NET0131 ,
		\u2_uk_K_r8_reg[8]/NET0131 ,
		_w9073_
	);
	LUT4 #(
		.INIT('hc693)
	) name3247 (
		decrypt_pad,
		\u2_R8_reg[29]/NET0131 ,
		\u2_uk_K_r8_reg[1]/NET0131 ,
		\u2_uk_K_r8_reg[36]/NET0131 ,
		_w9074_
	);
	LUT4 #(
		.INIT('hc963)
	) name3248 (
		decrypt_pad,
		\u2_R8_reg[28]/NET0131 ,
		\u2_uk_K_r8_reg[44]/NET0131 ,
		\u2_uk_K_r8_reg[9]/NET0131 ,
		_w9075_
	);
	LUT4 #(
		.INIT('hc693)
	) name3249 (
		decrypt_pad,
		\u2_R8_reg[26]/NET0131 ,
		\u2_uk_K_r8_reg[44]/NET0131 ,
		\u2_uk_K_r8_reg[52]/NET0131 ,
		_w9076_
	);
	LUT4 #(
		.INIT('h9afa)
	) name3250 (
		_w9073_,
		_w9076_,
		_w9074_,
		_w9075_,
		_w9077_
	);
	LUT4 #(
		.INIT('h0400)
	) name3251 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9078_
	);
	LUT3 #(
		.INIT('h02)
	) name3252 (
		_w9076_,
		_w9072_,
		_w9074_,
		_w9079_
	);
	LUT4 #(
		.INIT('h0008)
	) name3253 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9080_
	);
	LUT4 #(
		.INIT('hfbe6)
	) name3254 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9081_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3255 (
		_w9071_,
		_w9072_,
		_w9077_,
		_w9081_,
		_w9082_
	);
	LUT2 #(
		.INIT('h6)
	) name3256 (
		_w9076_,
		_w9072_,
		_w9083_
	);
	LUT4 #(
		.INIT('h0004)
	) name3257 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9084_
	);
	LUT4 #(
		.INIT('h3c5b)
	) name3258 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9085_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		_w9071_,
		_w9085_,
		_w9086_
	);
	LUT4 #(
		.INIT('h8200)
	) name3260 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9087_
	);
	LUT2 #(
		.INIT('h4)
	) name3261 (
		_w9071_,
		_w9074_,
		_w9088_
	);
	LUT3 #(
		.INIT('h10)
	) name3262 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9089_
	);
	LUT3 #(
		.INIT('h45)
	) name3263 (
		_w9087_,
		_w9088_,
		_w9089_,
		_w9090_
	);
	LUT3 #(
		.INIT('h0b)
	) name3264 (
		_w9086_,
		_w9090_,
		_w9075_,
		_w9091_
	);
	LUT4 #(
		.INIT('h4004)
	) name3265 (
		_w9071_,
		_w9073_,
		_w9076_,
		_w9072_,
		_w9092_
	);
	LUT4 #(
		.INIT('h1000)
	) name3266 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9093_
	);
	LUT4 #(
		.INIT('he5ff)
	) name3267 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9094_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name3268 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9095_
	);
	LUT4 #(
		.INIT('h04cc)
	) name3269 (
		_w9071_,
		_w9075_,
		_w9094_,
		_w9095_,
		_w9096_
	);
	LUT2 #(
		.INIT('h1)
	) name3270 (
		_w9092_,
		_w9096_,
		_w9097_
	);
	LUT4 #(
		.INIT('h5655)
	) name3271 (
		\u2_L8_reg[22]/NET0131 ,
		_w9091_,
		_w9082_,
		_w9097_,
		_w9098_
	);
	LUT4 #(
		.INIT('h0200)
	) name3272 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9099_
	);
	LUT4 #(
		.INIT('ha9ab)
	) name3273 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9100_
	);
	LUT2 #(
		.INIT('h2)
	) name3274 (
		_w9014_,
		_w9100_,
		_w9101_
	);
	LUT4 #(
		.INIT('h00a1)
	) name3275 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9014_,
		_w9102_
	);
	LUT4 #(
		.INIT('h0008)
	) name3276 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9103_
	);
	LUT3 #(
		.INIT('h80)
	) name3277 (
		_w9016_,
		_w9011_,
		_w9012_,
		_w9104_
	);
	LUT4 #(
		.INIT('h0002)
	) name3278 (
		_w9010_,
		_w9103_,
		_w9104_,
		_w9102_,
		_w9105_
	);
	LUT4 #(
		.INIT('h0440)
	) name3279 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9106_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3280 (
		_w9015_,
		_w9016_,
		_w9014_,
		_w9012_,
		_w9107_
	);
	LUT3 #(
		.INIT('h21)
	) name3281 (
		_w9015_,
		_w9016_,
		_w9012_,
		_w9108_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name3282 (
		_w9015_,
		_w9011_,
		_w9014_,
		_w9012_,
		_w9109_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3283 (
		_w9106_,
		_w9107_,
		_w9108_,
		_w9109_,
		_w9110_
	);
	LUT3 #(
		.INIT('h01)
	) name3284 (
		_w9010_,
		_w9019_,
		_w9030_,
		_w9111_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3285 (
		_w9101_,
		_w9105_,
		_w9110_,
		_w9111_,
		_w9112_
	);
	LUT2 #(
		.INIT('h6)
	) name3286 (
		\u2_L8_reg[17]/NET0131 ,
		_w9112_,
		_w9113_
	);
	LUT4 #(
		.INIT('hc693)
	) name3287 (
		decrypt_pad,
		\u2_R8_reg[15]/NET0131 ,
		\u2_uk_K_r8_reg[27]/NET0131 ,
		\u2_uk_K_r8_reg[5]/NET0131 ,
		_w9114_
	);
	LUT4 #(
		.INIT('hc693)
	) name3288 (
		decrypt_pad,
		\u2_R8_reg[13]/NET0131 ,
		\u2_uk_K_r8_reg[18]/NET0131 ,
		\u2_uk_K_r8_reg[53]/NET0131 ,
		_w9115_
	);
	LUT4 #(
		.INIT('hc693)
	) name3289 (
		decrypt_pad,
		\u2_R8_reg[12]/NET0131 ,
		\u2_uk_K_r8_reg[24]/NET0131 ,
		\u2_uk_K_r8_reg[34]/NET0131 ,
		_w9116_
	);
	LUT4 #(
		.INIT('hc963)
	) name3290 (
		decrypt_pad,
		\u2_R8_reg[17]/NET0131 ,
		\u2_uk_K_r8_reg[18]/NET0131 ,
		\u2_uk_K_r8_reg[40]/NET0131 ,
		_w9117_
	);
	LUT2 #(
		.INIT('h1)
	) name3291 (
		_w9116_,
		_w9117_,
		_w9118_
	);
	LUT4 #(
		.INIT('h4cc8)
	) name3292 (
		_w9115_,
		_w9114_,
		_w9116_,
		_w9117_,
		_w9119_
	);
	LUT4 #(
		.INIT('hc693)
	) name3293 (
		decrypt_pad,
		\u2_R8_reg[14]/NET0131 ,
		\u2_uk_K_r8_reg[19]/NET0131 ,
		\u2_uk_K_r8_reg[54]/NET0131 ,
		_w9120_
	);
	LUT3 #(
		.INIT('h20)
	) name3294 (
		_w9116_,
		_w9117_,
		_w9120_,
		_w9121_
	);
	LUT3 #(
		.INIT('h23)
	) name3295 (
		_w9115_,
		_w9114_,
		_w9117_,
		_w9122_
	);
	LUT3 #(
		.INIT('h23)
	) name3296 (
		_w9121_,
		_w9119_,
		_w9122_,
		_w9123_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name3297 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9124_
	);
	LUT3 #(
		.INIT('h04)
	) name3298 (
		_w9115_,
		_w9116_,
		_w9120_,
		_w9125_
	);
	LUT4 #(
		.INIT('h0040)
	) name3299 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9126_
	);
	LUT4 #(
		.INIT('hc963)
	) name3300 (
		decrypt_pad,
		\u2_R8_reg[16]/NET0131 ,
		\u2_uk_K_r8_reg[13]/P0001 ,
		\u2_uk_K_r8_reg[3]/NET0131 ,
		_w9127_
	);
	LUT3 #(
		.INIT('h80)
	) name3301 (
		_w9115_,
		_w9114_,
		_w9120_,
		_w9128_
	);
	LUT4 #(
		.INIT('h0800)
	) name3302 (
		_w9115_,
		_w9114_,
		_w9116_,
		_w9120_,
		_w9129_
	);
	LUT4 #(
		.INIT('h0100)
	) name3303 (
		_w9127_,
		_w9129_,
		_w9126_,
		_w9124_,
		_w9130_
	);
	LUT2 #(
		.INIT('h4)
	) name3304 (
		_w9123_,
		_w9130_,
		_w9131_
	);
	LUT4 #(
		.INIT('h0080)
	) name3305 (
		_w9115_,
		_w9114_,
		_w9116_,
		_w9117_,
		_w9132_
	);
	LUT2 #(
		.INIT('h4)
	) name3306 (
		_w9116_,
		_w9117_,
		_w9133_
	);
	LUT4 #(
		.INIT('h0020)
	) name3307 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9134_
	);
	LUT2 #(
		.INIT('h1)
	) name3308 (
		_w9132_,
		_w9134_,
		_w9135_
	);
	LUT4 #(
		.INIT('h0001)
	) name3309 (
		_w9115_,
		_w9114_,
		_w9116_,
		_w9117_,
		_w9136_
	);
	LUT4 #(
		.INIT('h8000)
	) name3310 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9137_
	);
	LUT4 #(
		.INIT('h004c)
	) name3311 (
		_w9120_,
		_w9127_,
		_w9136_,
		_w9137_,
		_w9138_
	);
	LUT4 #(
		.INIT('h0400)
	) name3312 (
		_w9115_,
		_w9114_,
		_w9116_,
		_w9117_,
		_w9139_
	);
	LUT4 #(
		.INIT('h0012)
	) name3313 (
		_w9115_,
		_w9114_,
		_w9116_,
		_w9120_,
		_w9140_
	);
	LUT2 #(
		.INIT('h1)
	) name3314 (
		_w9139_,
		_w9140_,
		_w9141_
	);
	LUT3 #(
		.INIT('h80)
	) name3315 (
		_w9135_,
		_w9138_,
		_w9141_,
		_w9142_
	);
	LUT2 #(
		.INIT('h4)
	) name3316 (
		_w9114_,
		_w9134_,
		_w9143_
	);
	LUT2 #(
		.INIT('h4)
	) name3317 (
		_w9115_,
		_w9114_,
		_w9144_
	);
	LUT3 #(
		.INIT('h01)
	) name3318 (
		_w9116_,
		_w9117_,
		_w9120_,
		_w9145_
	);
	LUT3 #(
		.INIT('hde)
	) name3319 (
		_w9116_,
		_w9117_,
		_w9120_,
		_w9146_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3320 (
		_w9144_,
		_w9120_,
		_w9146_,
		_w9132_,
		_w9147_
	);
	LUT2 #(
		.INIT('h4)
	) name3321 (
		_w9143_,
		_w9147_,
		_w9148_
	);
	LUT4 #(
		.INIT('ha955)
	) name3322 (
		\u2_L8_reg[20]/NET0131 ,
		_w9131_,
		_w9142_,
		_w9148_,
		_w9149_
	);
	LUT4 #(
		.INIT('hc963)
	) name3323 (
		decrypt_pad,
		\u2_R8_reg[9]/NET0131 ,
		\u2_uk_K_r8_reg[17]/NET0131 ,
		\u2_uk_K_r8_reg[39]/NET0131 ,
		_w9150_
	);
	LUT4 #(
		.INIT('hc963)
	) name3324 (
		decrypt_pad,
		\u2_R8_reg[4]/NET0131 ,
		\u2_uk_K_r8_reg[25]/NET0131 ,
		\u2_uk_K_r8_reg[47]/NET0131 ,
		_w9151_
	);
	LUT2 #(
		.INIT('h2)
	) name3325 (
		_w9150_,
		_w9151_,
		_w9152_
	);
	LUT2 #(
		.INIT('h9)
	) name3326 (
		_w9150_,
		_w9151_,
		_w9153_
	);
	LUT4 #(
		.INIT('hc693)
	) name3327 (
		decrypt_pad,
		\u2_R8_reg[5]/NET0131 ,
		\u2_uk_K_r8_reg[26]/NET0131 ,
		\u2_uk_K_r8_reg[4]/NET0131 ,
		_w9154_
	);
	LUT4 #(
		.INIT('hc693)
	) name3328 (
		decrypt_pad,
		\u2_R8_reg[6]/NET0131 ,
		\u2_uk_K_r8_reg[17]/NET0131 ,
		\u2_uk_K_r8_reg[27]/NET0131 ,
		_w9155_
	);
	LUT4 #(
		.INIT('hc693)
	) name3329 (
		decrypt_pad,
		\u2_R8_reg[7]/NET0131 ,
		\u2_uk_K_r8_reg[11]/NET0131 ,
		\u2_uk_K_r8_reg[46]/NET0131 ,
		_w9156_
	);
	LUT4 #(
		.INIT('h0071)
	) name3330 (
		_w9154_,
		_w9151_,
		_w9155_,
		_w9156_,
		_w9157_
	);
	LUT2 #(
		.INIT('h8)
	) name3331 (
		_w9153_,
		_w9157_,
		_w9158_
	);
	LUT4 #(
		.INIT('h0010)
	) name3332 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9159_
	);
	LUT4 #(
		.INIT('hc963)
	) name3333 (
		decrypt_pad,
		\u2_R8_reg[8]/NET0131 ,
		\u2_uk_K_r8_reg[12]/NET0131 ,
		\u2_uk_K_r8_reg[34]/NET0131 ,
		_w9160_
	);
	LUT4 #(
		.INIT('h0080)
	) name3334 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9161_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3335 (
		_w9154_,
		_w9151_,
		_w9155_,
		_w9156_,
		_w9162_
	);
	LUT4 #(
		.INIT('h0010)
	) name3336 (
		_w9159_,
		_w9161_,
		_w9160_,
		_w9162_,
		_w9163_
	);
	LUT2 #(
		.INIT('h2)
	) name3337 (
		_w9154_,
		_w9150_,
		_w9164_
	);
	LUT2 #(
		.INIT('h4)
	) name3338 (
		_w9154_,
		_w9150_,
		_w9165_
	);
	LUT4 #(
		.INIT('h0026)
	) name3339 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9166_
	);
	LUT3 #(
		.INIT('h80)
	) name3340 (
		_w9151_,
		_w9155_,
		_w9156_,
		_w9167_
	);
	LUT4 #(
		.INIT('h0105)
	) name3341 (
		_w9160_,
		_w9165_,
		_w9166_,
		_w9167_,
		_w9168_
	);
	LUT4 #(
		.INIT('hf700)
	) name3342 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9169_
	);
	LUT3 #(
		.INIT('h32)
	) name3343 (
		_w9154_,
		_w9155_,
		_w9156_,
		_w9170_
	);
	LUT4 #(
		.INIT('hf0f4)
	) name3344 (
		_w9154_,
		_w9150_,
		_w9155_,
		_w9156_,
		_w9171_
	);
	LUT4 #(
		.INIT('h4bfb)
	) name3345 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9172_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name3346 (
		_w9156_,
		_w9169_,
		_w9171_,
		_w9172_,
		_w9173_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3347 (
		_w9158_,
		_w9163_,
		_w9168_,
		_w9173_,
		_w9174_
	);
	LUT3 #(
		.INIT('h10)
	) name3348 (
		_w9154_,
		_w9151_,
		_w9155_,
		_w9175_
	);
	LUT4 #(
		.INIT('h0100)
	) name3349 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9176_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name3350 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9177_
	);
	LUT3 #(
		.INIT('hf2)
	) name3351 (
		_w9154_,
		_w9155_,
		_w9156_,
		_w9178_
	);
	LUT4 #(
		.INIT('h080c)
	) name3352 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9179_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3353 (
		_w9156_,
		_w9177_,
		_w9178_,
		_w9179_,
		_w9180_
	);
	LUT3 #(
		.INIT('h65)
	) name3354 (
		\u2_L8_reg[2]/NET0131 ,
		_w9174_,
		_w9180_,
		_w9181_
	);
	LUT4 #(
		.INIT('h67dc)
	) name3355 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9182_
	);
	LUT4 #(
		.INIT('hd2f7)
	) name3356 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9183_
	);
	LUT4 #(
		.INIT('h0040)
	) name3357 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9184_
	);
	LUT4 #(
		.INIT('h00d8)
	) name3358 (
		_w9044_,
		_w9182_,
		_w9183_,
		_w9184_,
		_w9185_
	);
	LUT4 #(
		.INIT('h9aff)
	) name3359 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9186_
	);
	LUT4 #(
		.INIT('haa02)
	) name3360 (
		_w9044_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9187_
	);
	LUT4 #(
		.INIT('h9297)
	) name3361 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9188_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3362 (
		_w9044_,
		_w9186_,
		_w9187_,
		_w9188_,
		_w9189_
	);
	LUT4 #(
		.INIT('h0800)
	) name3363 (
		_w9044_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9190_
	);
	LUT2 #(
		.INIT('h1)
	) name3364 (
		_w9056_,
		_w9190_,
		_w9191_
	);
	LUT4 #(
		.INIT('hd800)
	) name3365 (
		_w9040_,
		_w9189_,
		_w9185_,
		_w9191_,
		_w9192_
	);
	LUT2 #(
		.INIT('h6)
	) name3366 (
		\u2_L8_reg[29]/NET0131 ,
		_w9192_,
		_w9193_
	);
	LUT4 #(
		.INIT('hd97b)
	) name3367 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9194_
	);
	LUT2 #(
		.INIT('h2)
	) name3368 (
		_w9044_,
		_w9194_,
		_w9195_
	);
	LUT4 #(
		.INIT('heebf)
	) name3369 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9196_
	);
	LUT4 #(
		.INIT('h0040)
	) name3370 (
		_w9044_,
		_w9041_,
		_w9046_,
		_w9042_,
		_w9197_
	);
	LUT4 #(
		.INIT('h0032)
	) name3371 (
		_w9044_,
		_w9056_,
		_w9196_,
		_w9197_,
		_w9198_
	);
	LUT3 #(
		.INIT('h45)
	) name3372 (
		_w9040_,
		_w9195_,
		_w9198_,
		_w9199_
	);
	LUT4 #(
		.INIT('h7c7f)
	) name3373 (
		_w9044_,
		_w9041_,
		_w9046_,
		_w9043_,
		_w9200_
	);
	LUT2 #(
		.INIT('h1)
	) name3374 (
		_w9042_,
		_w9200_,
		_w9201_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name3375 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9202_
	);
	LUT3 #(
		.INIT('h80)
	) name3376 (
		_w9046_,
		_w9042_,
		_w9043_,
		_w9203_
	);
	LUT3 #(
		.INIT('h0e)
	) name3377 (
		_w9044_,
		_w9202_,
		_w9203_,
		_w9204_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3378 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9205_
	);
	LUT4 #(
		.INIT('h5501)
	) name3379 (
		_w9044_,
		_w9041_,
		_w9046_,
		_w9042_,
		_w9206_
	);
	LUT3 #(
		.INIT('h9e)
	) name3380 (
		_w9041_,
		_w9046_,
		_w9043_,
		_w9207_
	);
	LUT2 #(
		.INIT('h8)
	) name3381 (
		_w9044_,
		_w9042_,
		_w9208_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3382 (
		_w9205_,
		_w9206_,
		_w9207_,
		_w9208_,
		_w9209_
	);
	LUT4 #(
		.INIT('h7500)
	) name3383 (
		_w9040_,
		_w9201_,
		_w9204_,
		_w9209_,
		_w9210_
	);
	LUT3 #(
		.INIT('h65)
	) name3384 (
		\u2_L8_reg[4]/NET0131 ,
		_w9199_,
		_w9210_,
		_w9211_
	);
	LUT4 #(
		.INIT('hc693)
	) name3385 (
		decrypt_pad,
		\u2_R8_reg[32]/NET0131 ,
		\u2_uk_K_r8_reg[29]/NET0131 ,
		\u2_uk_K_r8_reg[9]/NET0131 ,
		_w9212_
	);
	LUT4 #(
		.INIT('hc693)
	) name3386 (
		decrypt_pad,
		\u2_R8_reg[31]/P0001 ,
		\u2_uk_K_r8_reg[23]/NET0131 ,
		\u2_uk_K_r8_reg[31]/NET0131 ,
		_w9213_
	);
	LUT4 #(
		.INIT('hc963)
	) name3387 (
		decrypt_pad,
		\u2_R8_reg[1]/NET0131 ,
		\u2_uk_K_r8_reg[30]/NET0131 ,
		\u2_uk_K_r8_reg[50]/NET0131 ,
		_w9214_
	);
	LUT4 #(
		.INIT('hc963)
	) name3388 (
		decrypt_pad,
		\u2_R8_reg[30]/NET0131 ,
		\u2_uk_K_r8_reg[15]/NET0131 ,
		\u2_uk_K_r8_reg[35]/NET0131 ,
		_w9215_
	);
	LUT4 #(
		.INIT('hc963)
	) name3389 (
		decrypt_pad,
		\u2_R8_reg[28]/NET0131 ,
		\u2_uk_K_r8_reg[42]/NET0131 ,
		\u2_uk_K_r8_reg[7]/NET0131 ,
		_w9216_
	);
	LUT4 #(
		.INIT('hc963)
	) name3390 (
		decrypt_pad,
		\u2_R8_reg[29]/NET0131 ,
		\u2_uk_K_r8_reg[14]/NET0131 ,
		\u2_uk_K_r8_reg[38]/NET0131 ,
		_w9217_
	);
	LUT4 #(
		.INIT('hfcf7)
	) name3391 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9218_
	);
	LUT2 #(
		.INIT('h2)
	) name3392 (
		_w9213_,
		_w9218_,
		_w9219_
	);
	LUT3 #(
		.INIT('h32)
	) name3393 (
		_w9215_,
		_w9213_,
		_w9214_,
		_w9220_
	);
	LUT3 #(
		.INIT('hc5)
	) name3394 (
		_w9216_,
		_w9217_,
		_w9214_,
		_w9221_
	);
	LUT2 #(
		.INIT('h8)
	) name3395 (
		_w9220_,
		_w9221_,
		_w9222_
	);
	LUT4 #(
		.INIT('h8000)
	) name3396 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9223_
	);
	LUT4 #(
		.INIT('h0040)
	) name3397 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9224_
	);
	LUT3 #(
		.INIT('h04)
	) name3398 (
		_w9215_,
		_w9216_,
		_w9213_,
		_w9225_
	);
	LUT3 #(
		.INIT('h01)
	) name3399 (
		_w9224_,
		_w9225_,
		_w9223_,
		_w9226_
	);
	LUT4 #(
		.INIT('h5455)
	) name3400 (
		_w9212_,
		_w9219_,
		_w9222_,
		_w9226_,
		_w9227_
	);
	LUT3 #(
		.INIT('h01)
	) name3401 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9228_
	);
	LUT4 #(
		.INIT('h44b4)
	) name3402 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9229_
	);
	LUT4 #(
		.INIT('h2000)
	) name3403 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9230_
	);
	LUT4 #(
		.INIT('h001d)
	) name3404 (
		_w9228_,
		_w9213_,
		_w9229_,
		_w9230_,
		_w9231_
	);
	LUT4 #(
		.INIT('h0001)
	) name3405 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9232_
	);
	LUT4 #(
		.INIT('h0200)
	) name3406 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9233_
	);
	LUT4 #(
		.INIT('hf9de)
	) name3407 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9234_
	);
	LUT2 #(
		.INIT('h2)
	) name3408 (
		_w9213_,
		_w9234_,
		_w9235_
	);
	LUT3 #(
		.INIT('h20)
	) name3409 (
		_w9216_,
		_w9217_,
		_w9212_,
		_w9236_
	);
	LUT4 #(
		.INIT('hcdcf)
	) name3410 (
		_w9215_,
		_w9213_,
		_w9224_,
		_w9236_,
		_w9237_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3411 (
		_w9231_,
		_w9212_,
		_w9235_,
		_w9237_,
		_w9238_
	);
	LUT3 #(
		.INIT('h9a)
	) name3412 (
		\u2_L8_reg[5]/NET0131 ,
		_w9227_,
		_w9238_,
		_w9239_
	);
	LUT4 #(
		.INIT('hfdbd)
	) name3413 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9240_
	);
	LUT4 #(
		.INIT('hf3db)
	) name3414 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9241_
	);
	LUT4 #(
		.INIT('h9000)
	) name3415 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9242_
	);
	LUT4 #(
		.INIT('h00e4)
	) name3416 (
		_w9114_,
		_w9241_,
		_w9240_,
		_w9242_,
		_w9243_
	);
	LUT2 #(
		.INIT('h2)
	) name3417 (
		_w9127_,
		_w9243_,
		_w9244_
	);
	LUT3 #(
		.INIT('h08)
	) name3418 (
		_w9115_,
		_w9116_,
		_w9120_,
		_w9245_
	);
	LUT4 #(
		.INIT('h0040)
	) name3419 (
		_w9114_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9246_
	);
	LUT3 #(
		.INIT('h01)
	) name3420 (
		_w9136_,
		_w9246_,
		_w9245_,
		_w9247_
	);
	LUT2 #(
		.INIT('h2)
	) name3421 (
		_w9117_,
		_w9120_,
		_w9248_
	);
	LUT3 #(
		.INIT('h40)
	) name3422 (
		_w9115_,
		_w9114_,
		_w9116_,
		_w9249_
	);
	LUT4 #(
		.INIT('h0020)
	) name3423 (
		_w9114_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9250_
	);
	LUT3 #(
		.INIT('h0b)
	) name3424 (
		_w9248_,
		_w9249_,
		_w9250_,
		_w9251_
	);
	LUT4 #(
		.INIT('h1555)
	) name3425 (
		_w9127_,
		_w9124_,
		_w9247_,
		_w9251_,
		_w9252_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name3426 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9253_
	);
	LUT2 #(
		.INIT('h1)
	) name3427 (
		_w9114_,
		_w9253_,
		_w9254_
	);
	LUT3 #(
		.INIT('h23)
	) name3428 (
		_w9120_,
		_w9129_,
		_w9132_,
		_w9255_
	);
	LUT2 #(
		.INIT('h4)
	) name3429 (
		_w9254_,
		_w9255_,
		_w9256_
	);
	LUT4 #(
		.INIT('h5655)
	) name3430 (
		\u2_L8_reg[10]/NET0131 ,
		_w9252_,
		_w9244_,
		_w9256_,
		_w9257_
	);
	LUT4 #(
		.INIT('h4000)
	) name3431 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9258_
	);
	LUT4 #(
		.INIT('hbfe9)
	) name3432 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9259_
	);
	LUT2 #(
		.INIT('h2)
	) name3433 (
		_w9071_,
		_w9075_,
		_w9260_
	);
	LUT4 #(
		.INIT('hff40)
	) name3434 (
		_w9071_,
		_w9076_,
		_w9072_,
		_w9075_,
		_w9261_
	);
	LUT2 #(
		.INIT('h1)
	) name3435 (
		_w9071_,
		_w9073_,
		_w9262_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3436 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9263_
	);
	LUT3 #(
		.INIT('h41)
	) name3437 (
		_w9071_,
		_w9073_,
		_w9074_,
		_w9264_
	);
	LUT4 #(
		.INIT('h000b)
	) name3438 (
		_w9262_,
		_w9263_,
		_w9264_,
		_w9261_,
		_w9265_
	);
	LUT2 #(
		.INIT('h8)
	) name3439 (
		_w9259_,
		_w9265_,
		_w9266_
	);
	LUT4 #(
		.INIT('h5f5e)
	) name3440 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9267_
	);
	LUT2 #(
		.INIT('h2)
	) name3441 (
		_w9071_,
		_w9267_,
		_w9268_
	);
	LUT3 #(
		.INIT('h02)
	) name3442 (
		_w9075_,
		_w9093_,
		_w9080_,
		_w9269_
	);
	LUT2 #(
		.INIT('h9)
	) name3443 (
		_w9072_,
		_w9074_,
		_w9270_
	);
	LUT4 #(
		.INIT('h3010)
	) name3444 (
		_w9071_,
		_w9073_,
		_w9076_,
		_w9072_,
		_w9271_
	);
	LUT4 #(
		.INIT('h0200)
	) name3445 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9272_
	);
	LUT3 #(
		.INIT('h0b)
	) name3446 (
		_w9270_,
		_w9271_,
		_w9272_,
		_w9273_
	);
	LUT3 #(
		.INIT('h40)
	) name3447 (
		_w9268_,
		_w9269_,
		_w9273_,
		_w9274_
	);
	LUT3 #(
		.INIT('ha9)
	) name3448 (
		\u2_L8_reg[12]/NET0131 ,
		_w9266_,
		_w9274_,
		_w9275_
	);
	LUT4 #(
		.INIT('h2000)
	) name3449 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9276_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name3450 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9277_
	);
	LUT4 #(
		.INIT('hf9ed)
	) name3451 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9278_
	);
	LUT4 #(
		.INIT('h0313)
	) name3452 (
		_w9160_,
		_w9156_,
		_w9277_,
		_w9278_,
		_w9279_
	);
	LUT4 #(
		.INIT('hae8e)
	) name3453 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9280_
	);
	LUT4 #(
		.INIT('hef00)
	) name3454 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9156_,
		_w9281_
	);
	LUT2 #(
		.INIT('h4)
	) name3455 (
		_w9280_,
		_w9281_,
		_w9282_
	);
	LUT2 #(
		.INIT('h8)
	) name3456 (
		_w9152_,
		_w9170_,
		_w9283_
	);
	LUT3 #(
		.INIT('h45)
	) name3457 (
		_w9160_,
		_w9164_,
		_w9167_,
		_w9284_
	);
	LUT3 #(
		.INIT('h10)
	) name3458 (
		_w9282_,
		_w9283_,
		_w9284_,
		_w9285_
	);
	LUT4 #(
		.INIT('h5140)
	) name3459 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9286_
	);
	LUT3 #(
		.INIT('h20)
	) name3460 (
		_w9150_,
		_w9151_,
		_w9155_,
		_w9287_
	);
	LUT3 #(
		.INIT('h01)
	) name3461 (
		_w9154_,
		_w9150_,
		_w9155_,
		_w9288_
	);
	LUT4 #(
		.INIT('heee4)
	) name3462 (
		_w9156_,
		_w9286_,
		_w9288_,
		_w9287_,
		_w9289_
	);
	LUT4 #(
		.INIT('h0002)
	) name3463 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9290_
	);
	LUT4 #(
		.INIT('h008a)
	) name3464 (
		_w9160_,
		_w9169_,
		_w9171_,
		_w9290_,
		_w9291_
	);
	LUT3 #(
		.INIT('h20)
	) name3465 (
		_w9277_,
		_w9289_,
		_w9291_,
		_w9292_
	);
	LUT4 #(
		.INIT('h999a)
	) name3466 (
		\u2_L8_reg[13]/NET0131 ,
		_w9279_,
		_w9285_,
		_w9292_,
		_w9293_
	);
	LUT4 #(
		.INIT('hc693)
	) name3467 (
		decrypt_pad,
		\u2_R8_reg[20]/NET0131 ,
		\u2_uk_K_r8_reg[14]/NET0131 ,
		\u2_uk_K_r8_reg[49]/NET0131 ,
		_w9294_
	);
	LUT4 #(
		.INIT('hc693)
	) name3468 (
		decrypt_pad,
		\u2_R8_reg[19]/NET0131 ,
		\u2_uk_K_r8_reg[30]/NET0131 ,
		\u2_uk_K_r8_reg[38]/NET0131 ,
		_w9295_
	);
	LUT4 #(
		.INIT('hc693)
	) name3469 (
		decrypt_pad,
		\u2_R8_reg[16]/NET0131 ,
		\u2_uk_K_r8_reg[31]/NET0131 ,
		\u2_uk_K_r8_reg[7]/NET0131 ,
		_w9296_
	);
	LUT4 #(
		.INIT('hc963)
	) name3470 (
		decrypt_pad,
		\u2_R8_reg[17]/NET0131 ,
		\u2_uk_K_r8_reg[29]/NET0131 ,
		\u2_uk_K_r8_reg[49]/NET0131 ,
		_w9297_
	);
	LUT4 #(
		.INIT('hc693)
	) name3471 (
		decrypt_pad,
		\u2_R8_reg[21]/NET0131 ,
		\u2_uk_K_r8_reg[15]/NET0131 ,
		\u2_uk_K_r8_reg[50]/NET0131 ,
		_w9298_
	);
	LUT4 #(
		.INIT('hc963)
	) name3472 (
		decrypt_pad,
		\u2_R8_reg[18]/NET0131 ,
		\u2_uk_K_r8_reg[23]/NET0131 ,
		\u2_uk_K_r8_reg[43]/NET0131 ,
		_w9299_
	);
	LUT4 #(
		.INIT('h0080)
	) name3473 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9300_
	);
	LUT4 #(
		.INIT('h0002)
	) name3474 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9301_
	);
	LUT4 #(
		.INIT('hcb79)
	) name3475 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9302_
	);
	LUT4 #(
		.INIT('h76ae)
	) name3476 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9303_
	);
	LUT4 #(
		.INIT('h0810)
	) name3477 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9304_
	);
	LUT4 #(
		.INIT('h00e4)
	) name3478 (
		_w9295_,
		_w9302_,
		_w9303_,
		_w9304_,
		_w9305_
	);
	LUT2 #(
		.INIT('h1)
	) name3479 (
		_w9294_,
		_w9305_,
		_w9306_
	);
	LUT4 #(
		.INIT('hdf9e)
	) name3480 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9295_,
		_w9307_
	);
	LUT2 #(
		.INIT('h1)
	) name3481 (
		_w9307_,
		_w9299_,
		_w9308_
	);
	LUT2 #(
		.INIT('h8)
	) name3482 (
		_w9296_,
		_w9298_,
		_w9309_
	);
	LUT2 #(
		.INIT('h4)
	) name3483 (
		_w9296_,
		_w9299_,
		_w9310_
	);
	LUT4 #(
		.INIT('h9b53)
	) name3484 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9311_
	);
	LUT2 #(
		.INIT('h2)
	) name3485 (
		_w9295_,
		_w9311_,
		_w9312_
	);
	LUT3 #(
		.INIT('hda)
	) name3486 (
		_w9297_,
		_w9295_,
		_w9299_,
		_w9313_
	);
	LUT4 #(
		.INIT('h0200)
	) name3487 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9314_
	);
	LUT3 #(
		.INIT('h0d)
	) name3488 (
		_w9309_,
		_w9313_,
		_w9314_,
		_w9315_
	);
	LUT4 #(
		.INIT('hef00)
	) name3489 (
		_w9308_,
		_w9312_,
		_w9315_,
		_w9294_,
		_w9316_
	);
	LUT4 #(
		.INIT('h0400)
	) name3490 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9317_
	);
	LUT4 #(
		.INIT('h1400)
	) name3491 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9318_
	);
	LUT4 #(
		.INIT('h0020)
	) name3492 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9319_
	);
	LUT4 #(
		.INIT('hfedf)
	) name3493 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9320_
	);
	LUT3 #(
		.INIT('hb1)
	) name3494 (
		_w9295_,
		_w9318_,
		_w9320_,
		_w9321_
	);
	LUT4 #(
		.INIT('h5655)
	) name3495 (
		\u2_L8_reg[14]/NET0131 ,
		_w9316_,
		_w9306_,
		_w9321_,
		_w9322_
	);
	LUT4 #(
		.INIT('h3c2f)
	) name3496 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9323_
	);
	LUT4 #(
		.INIT('h0004)
	) name3497 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9324_
	);
	LUT4 #(
		.INIT('h3302)
	) name3498 (
		_w9213_,
		_w9212_,
		_w9323_,
		_w9324_,
		_w9325_
	);
	LUT4 #(
		.INIT('h0010)
	) name3499 (
		_w9216_,
		_w9217_,
		_w9213_,
		_w9214_,
		_w9326_
	);
	LUT3 #(
		.INIT('h40)
	) name3500 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9327_
	);
	LUT4 #(
		.INIT('h0200)
	) name3501 (
		_w9215_,
		_w9217_,
		_w9213_,
		_w9214_,
		_w9328_
	);
	LUT4 #(
		.INIT('h0800)
	) name3502 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9329_
	);
	LUT4 #(
		.INIT('hf7df)
	) name3503 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9330_
	);
	LUT4 #(
		.INIT('h0100)
	) name3504 (
		_w9327_,
		_w9328_,
		_w9326_,
		_w9330_,
		_w9331_
	);
	LUT4 #(
		.INIT('h080c)
	) name3505 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9212_,
		_w9332_
	);
	LUT2 #(
		.INIT('h8)
	) name3506 (
		_w9217_,
		_w9214_,
		_w9333_
	);
	LUT4 #(
		.INIT('hefdf)
	) name3507 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9334_
	);
	LUT4 #(
		.INIT('h0100)
	) name3508 (
		_w9213_,
		_w9232_,
		_w9332_,
		_w9334_,
		_w9335_
	);
	LUT4 #(
		.INIT('h0100)
	) name3509 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9336_
	);
	LUT3 #(
		.INIT('h02)
	) name3510 (
		_w9213_,
		_w9230_,
		_w9336_,
		_w9337_
	);
	LUT4 #(
		.INIT('hddd0)
	) name3511 (
		_w9212_,
		_w9331_,
		_w9335_,
		_w9337_,
		_w9338_
	);
	LUT3 #(
		.INIT('h65)
	) name3512 (
		\u2_L8_reg[15]/NET0131 ,
		_w9325_,
		_w9338_,
		_w9339_
	);
	LUT4 #(
		.INIT('h404c)
	) name3513 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9340_
	);
	LUT4 #(
		.INIT('h0400)
	) name3514 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9341_
	);
	LUT4 #(
		.INIT('hfad8)
	) name3515 (
		_w9114_,
		_w9145_,
		_w9340_,
		_w9341_,
		_w9342_
	);
	LUT4 #(
		.INIT('h7fd7)
	) name3516 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9343_
	);
	LUT3 #(
		.INIT('h45)
	) name3517 (
		_w9127_,
		_w9342_,
		_w9343_,
		_w9344_
	);
	LUT4 #(
		.INIT('hafab)
	) name3518 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9345_
	);
	LUT4 #(
		.INIT('h6dff)
	) name3519 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9346_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3520 (
		_w9114_,
		_w9127_,
		_w9345_,
		_w9346_,
		_w9347_
	);
	LUT4 #(
		.INIT('hdf5d)
	) name3521 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9348_
	);
	LUT4 #(
		.INIT('h0800)
	) name3522 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9349_
	);
	LUT4 #(
		.INIT('he6ff)
	) name3523 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9350_
	);
	LUT4 #(
		.INIT('h04cc)
	) name3524 (
		_w9114_,
		_w9127_,
		_w9348_,
		_w9350_,
		_w9351_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name3525 (
		_w9114_,
		_w9120_,
		_w9136_,
		_w9349_,
		_w9352_
	);
	LUT3 #(
		.INIT('h10)
	) name3526 (
		_w9351_,
		_w9347_,
		_w9352_,
		_w9353_
	);
	LUT3 #(
		.INIT('h65)
	) name3527 (
		\u2_L8_reg[1]/NET0131 ,
		_w9344_,
		_w9353_,
		_w9354_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name3528 (
		_w9044_,
		_w9041_,
		_w9046_,
		_w9042_,
		_w9355_
	);
	LUT4 #(
		.INIT('hef00)
	) name3529 (
		_w9046_,
		_w9042_,
		_w9043_,
		_w9040_,
		_w9356_
	);
	LUT3 #(
		.INIT('he0)
	) name3530 (
		_w9043_,
		_w9355_,
		_w9356_,
		_w9357_
	);
	LUT4 #(
		.INIT('h4010)
	) name3531 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9358_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name3532 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9359_
	);
	LUT3 #(
		.INIT('h31)
	) name3533 (
		_w9044_,
		_w9358_,
		_w9359_,
		_w9360_
	);
	LUT4 #(
		.INIT('h4e55)
	) name3534 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9361_
	);
	LUT2 #(
		.INIT('h2)
	) name3535 (
		_w9044_,
		_w9361_,
		_w9362_
	);
	LUT4 #(
		.INIT('h1001)
	) name3536 (
		_w9044_,
		_w9041_,
		_w9046_,
		_w9043_,
		_w9363_
	);
	LUT4 #(
		.INIT('h8000)
	) name3537 (
		_w9041_,
		_w9046_,
		_w9042_,
		_w9043_,
		_w9364_
	);
	LUT3 #(
		.INIT('h01)
	) name3538 (
		_w9040_,
		_w9364_,
		_w9363_,
		_w9365_
	);
	LUT4 #(
		.INIT('h7077)
	) name3539 (
		_w9357_,
		_w9360_,
		_w9362_,
		_w9365_,
		_w9366_
	);
	LUT2 #(
		.INIT('h4)
	) name3540 (
		_w9043_,
		_w9197_,
		_w9367_
	);
	LUT2 #(
		.INIT('h1)
	) name3541 (
		_w9064_,
		_w9367_,
		_w9368_
	);
	LUT3 #(
		.INIT('h65)
	) name3542 (
		\u2_L8_reg[19]/NET0131 ,
		_w9366_,
		_w9368_,
		_w9369_
	);
	LUT2 #(
		.INIT('h1)
	) name3543 (
		_w9216_,
		_w9213_,
		_w9370_
	);
	LUT4 #(
		.INIT('hf0f4)
	) name3544 (
		_w9215_,
		_w9216_,
		_w9213_,
		_w9214_,
		_w9371_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name3545 (
		_w9216_,
		_w9217_,
		_w9213_,
		_w9214_,
		_w9372_
	);
	LUT4 #(
		.INIT('h7a7f)
	) name3546 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9373_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3547 (
		_w9329_,
		_w9371_,
		_w9372_,
		_w9373_,
		_w9374_
	);
	LUT4 #(
		.INIT('h0082)
	) name3548 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9375_
	);
	LUT3 #(
		.INIT('h02)
	) name3549 (
		_w9212_,
		_w9336_,
		_w9375_,
		_w9376_
	);
	LUT4 #(
		.INIT('hfff6)
	) name3550 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9377_
	);
	LUT3 #(
		.INIT('h53)
	) name3551 (
		_w9215_,
		_w9217_,
		_w9214_,
		_w9378_
	);
	LUT4 #(
		.INIT('h00df)
	) name3552 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9212_,
		_w9379_
	);
	LUT4 #(
		.INIT('hd000)
	) name3553 (
		_w9370_,
		_w9378_,
		_w9379_,
		_w9377_,
		_w9380_
	);
	LUT4 #(
		.INIT('hf737)
	) name3554 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9381_
	);
	LUT4 #(
		.INIT('hbfbb)
	) name3555 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9213_,
		_w9382_
	);
	LUT4 #(
		.INIT('hf531)
	) name3556 (
		_w9213_,
		_w9214_,
		_w9381_,
		_w9382_,
		_w9383_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3557 (
		_w9374_,
		_w9376_,
		_w9380_,
		_w9383_,
		_w9384_
	);
	LUT4 #(
		.INIT('h0100)
	) name3558 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9213_,
		_w9385_
	);
	LUT3 #(
		.INIT('h07)
	) name3559 (
		_w9225_,
		_w9333_,
		_w9385_,
		_w9386_
	);
	LUT3 #(
		.INIT('h65)
	) name3560 (
		\u2_L8_reg[21]/NET0131 ,
		_w9384_,
		_w9386_,
		_w9387_
	);
	LUT4 #(
		.INIT('ha888)
	) name3561 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9388_
	);
	LUT3 #(
		.INIT('h40)
	) name3562 (
		_w9015_,
		_w9011_,
		_w9012_,
		_w9389_
	);
	LUT3 #(
		.INIT('h04)
	) name3563 (
		_w9015_,
		_w9016_,
		_w9012_,
		_w9390_
	);
	LUT4 #(
		.INIT('hfad8)
	) name3564 (
		_w9014_,
		_w9390_,
		_w9388_,
		_w9389_,
		_w9391_
	);
	LUT4 #(
		.INIT('h070e)
	) name3565 (
		_w9016_,
		_w9011_,
		_w9010_,
		_w9012_,
		_w9392_
	);
	LUT4 #(
		.INIT('h4000)
	) name3566 (
		_w9015_,
		_w9016_,
		_w9014_,
		_w9012_,
		_w9393_
	);
	LUT3 #(
		.INIT('h02)
	) name3567 (
		_w9010_,
		_w9099_,
		_w9393_,
		_w9394_
	);
	LUT4 #(
		.INIT('h0777)
	) name3568 (
		_w9014_,
		_w9019_,
		_w9025_,
		_w9026_,
		_w9395_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3569 (
		_w9391_,
		_w9392_,
		_w9394_,
		_w9395_,
		_w9396_
	);
	LUT3 #(
		.INIT('hd9)
	) name3570 (
		_w9015_,
		_w9016_,
		_w9012_,
		_w9397_
	);
	LUT2 #(
		.INIT('h2)
	) name3571 (
		_w9023_,
		_w9397_,
		_w9398_
	);
	LUT4 #(
		.INIT('hee9b)
	) name3572 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9399_
	);
	LUT4 #(
		.INIT('h7ef7)
	) name3573 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9400_
	);
	LUT4 #(
		.INIT('h0455)
	) name3574 (
		_w9014_,
		_w9010_,
		_w9399_,
		_w9400_,
		_w9401_
	);
	LUT2 #(
		.INIT('h1)
	) name3575 (
		_w9398_,
		_w9401_,
		_w9402_
	);
	LUT3 #(
		.INIT('h9a)
	) name3576 (
		\u2_L8_reg[23]/NET0131 ,
		_w9396_,
		_w9402_,
		_w9403_
	);
	LUT3 #(
		.INIT('h80)
	) name3577 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9404_
	);
	LUT4 #(
		.INIT('h6a78)
	) name3578 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9405_
	);
	LUT4 #(
		.INIT('hf7a7)
	) name3579 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9406_
	);
	LUT4 #(
		.INIT('hdf3f)
	) name3580 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9407_
	);
	LUT4 #(
		.INIT('hd800)
	) name3581 (
		_w9295_,
		_w9405_,
		_w9406_,
		_w9407_,
		_w9408_
	);
	LUT2 #(
		.INIT('h2)
	) name3582 (
		_w9294_,
		_w9408_,
		_w9409_
	);
	LUT4 #(
		.INIT('h00f7)
	) name3583 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9295_,
		_w9410_
	);
	LUT3 #(
		.INIT('h04)
	) name3584 (
		_w9298_,
		_w9295_,
		_w9299_,
		_w9411_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name3585 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9412_
	);
	LUT4 #(
		.INIT('h0700)
	) name3586 (
		_w9310_,
		_w9410_,
		_w9411_,
		_w9412_,
		_w9413_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name3587 (
		_w9297_,
		_w9310_,
		_w9294_,
		_w9410_,
		_w9414_
	);
	LUT4 #(
		.INIT('hdefb)
	) name3588 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9415_
	);
	LUT4 #(
		.INIT('h0200)
	) name3589 (
		_w9296_,
		_w9297_,
		_w9295_,
		_w9299_,
		_w9416_
	);
	LUT4 #(
		.INIT('h0031)
	) name3590 (
		_w9295_,
		_w9300_,
		_w9415_,
		_w9416_,
		_w9417_
	);
	LUT3 #(
		.INIT('hb0)
	) name3591 (
		_w9413_,
		_w9414_,
		_w9417_,
		_w9418_
	);
	LUT3 #(
		.INIT('h65)
	) name3592 (
		\u2_L8_reg[25]/NET0131 ,
		_w9409_,
		_w9418_,
		_w9419_
	);
	LUT3 #(
		.INIT('hb1)
	) name3593 (
		_w9115_,
		_w9114_,
		_w9120_,
		_w9420_
	);
	LUT4 #(
		.INIT('h0c04)
	) name3594 (
		_w9118_,
		_w9127_,
		_w9349_,
		_w9420_,
		_w9421_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name3595 (
		_w9115_,
		_w9114_,
		_w9116_,
		_w9117_,
		_w9422_
	);
	LUT4 #(
		.INIT('h3f2f)
	) name3596 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9423_
	);
	LUT3 #(
		.INIT('h51)
	) name3597 (
		_w9114_,
		_w9116_,
		_w9120_,
		_w9424_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3598 (
		_w9120_,
		_w9422_,
		_w9423_,
		_w9424_,
		_w9425_
	);
	LUT3 #(
		.INIT('h51)
	) name3599 (
		_w9127_,
		_w9128_,
		_w9133_,
		_w9426_
	);
	LUT4 #(
		.INIT('h153f)
	) name3600 (
		_w9135_,
		_w9421_,
		_w9425_,
		_w9426_,
		_w9427_
	);
	LUT3 #(
		.INIT('he0)
	) name3601 (
		_w9114_,
		_w9117_,
		_w9127_,
		_w9428_
	);
	LUT2 #(
		.INIT('h2)
	) name3602 (
		_w9125_,
		_w9428_,
		_w9429_
	);
	LUT4 #(
		.INIT('heafa)
	) name3603 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9430_
	);
	LUT4 #(
		.INIT('h0082)
	) name3604 (
		_w9115_,
		_w9116_,
		_w9117_,
		_w9120_,
		_w9431_
	);
	LUT4 #(
		.INIT('h0054)
	) name3605 (
		_w9114_,
		_w9127_,
		_w9430_,
		_w9431_,
		_w9432_
	);
	LUT3 #(
		.INIT('h02)
	) name3606 (
		_w9114_,
		_w9126_,
		_w9134_,
		_w9433_
	);
	LUT3 #(
		.INIT('h54)
	) name3607 (
		_w9429_,
		_w9432_,
		_w9433_,
		_w9434_
	);
	LUT3 #(
		.INIT('h65)
	) name3608 (
		\u2_L8_reg[26]/NET0131 ,
		_w9427_,
		_w9434_,
		_w9435_
	);
	LUT3 #(
		.INIT('h0d)
	) name3609 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9436_
	);
	LUT4 #(
		.INIT('h92f0)
	) name3610 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9437_
	);
	LUT2 #(
		.INIT('h2)
	) name3611 (
		_w9156_,
		_w9437_,
		_w9438_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name3612 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9439_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3613 (
		_w9154_,
		_w9151_,
		_w9155_,
		_w9156_,
		_w9440_
	);
	LUT3 #(
		.INIT('h40)
	) name3614 (
		_w9276_,
		_w9440_,
		_w9439_,
		_w9441_
	);
	LUT4 #(
		.INIT('h0440)
	) name3615 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9442_
	);
	LUT2 #(
		.INIT('h2)
	) name3616 (
		_w9160_,
		_w9442_,
		_w9443_
	);
	LUT3 #(
		.INIT('he0)
	) name3617 (
		_w9438_,
		_w9441_,
		_w9443_,
		_w9444_
	);
	LUT4 #(
		.INIT('h5b4b)
	) name3618 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9445_
	);
	LUT4 #(
		.INIT('h4e5f)
	) name3619 (
		_w9156_,
		_w9175_,
		_w9439_,
		_w9445_,
		_w9446_
	);
	LUT4 #(
		.INIT('h4100)
	) name3620 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9447_
	);
	LUT3 #(
		.INIT('h01)
	) name3621 (
		_w9160_,
		_w9276_,
		_w9447_,
		_w9448_
	);
	LUT2 #(
		.INIT('h4)
	) name3622 (
		_w9446_,
		_w9448_,
		_w9449_
	);
	LUT3 #(
		.INIT('ha9)
	) name3623 (
		\u2_L8_reg[28]/NET0131 ,
		_w9444_,
		_w9449_,
		_w9450_
	);
	LUT3 #(
		.INIT('h02)
	) name3624 (
		_w9295_,
		_w9301_,
		_w9404_,
		_w9451_
	);
	LUT4 #(
		.INIT('h4044)
	) name3625 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9452_
	);
	LUT2 #(
		.INIT('h2)
	) name3626 (
		_w9410_,
		_w9452_,
		_w9453_
	);
	LUT4 #(
		.INIT('hdeaf)
	) name3627 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9454_
	);
	LUT4 #(
		.INIT('h0155)
	) name3628 (
		_w9294_,
		_w9451_,
		_w9453_,
		_w9454_,
		_w9455_
	);
	LUT4 #(
		.INIT('h0001)
	) name3629 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9456_
	);
	LUT4 #(
		.INIT('hf7f6)
	) name3630 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9457_
	);
	LUT3 #(
		.INIT('h02)
	) name3631 (
		_w9296_,
		_w9295_,
		_w9299_,
		_w9458_
	);
	LUT4 #(
		.INIT('h0031)
	) name3632 (
		_w9295_,
		_w9318_,
		_w9457_,
		_w9458_,
		_w9459_
	);
	LUT4 #(
		.INIT('hcbbf)
	) name3633 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9460_
	);
	LUT4 #(
		.INIT('haf23)
	) name3634 (
		_w9298_,
		_w9295_,
		_w9416_,
		_w9460_,
		_w9461_
	);
	LUT3 #(
		.INIT('hd0)
	) name3635 (
		_w9294_,
		_w9459_,
		_w9461_,
		_w9462_
	);
	LUT3 #(
		.INIT('h65)
	) name3636 (
		\u2_L8_reg[8]/NET0131 ,
		_w9455_,
		_w9462_,
		_w9463_
	);
	LUT4 #(
		.INIT('hc010)
	) name3637 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9464_
	);
	LUT3 #(
		.INIT('hb7)
	) name3638 (
		_w9216_,
		_w9217_,
		_w9214_,
		_w9465_
	);
	LUT4 #(
		.INIT('he2f3)
	) name3639 (
		_w9228_,
		_w9213_,
		_w9464_,
		_w9465_,
		_w9466_
	);
	LUT4 #(
		.INIT('hdaf7)
	) name3640 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9467_
	);
	LUT3 #(
		.INIT('h8a)
	) name3641 (
		_w9212_,
		_w9466_,
		_w9467_,
		_w9468_
	);
	LUT4 #(
		.INIT('h0203)
	) name3642 (
		_w9215_,
		_w9217_,
		_w9214_,
		_w9212_,
		_w9469_
	);
	LUT3 #(
		.INIT('h4a)
	) name3643 (
		_w9215_,
		_w9217_,
		_w9214_,
		_w9470_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3644 (
		_w9213_,
		_w9379_,
		_w9469_,
		_w9470_,
		_w9471_
	);
	LUT4 #(
		.INIT('h0004)
	) name3645 (
		_w9216_,
		_w9217_,
		_w9213_,
		_w9214_,
		_w9472_
	);
	LUT4 #(
		.INIT('h0800)
	) name3646 (
		_w9215_,
		_w9216_,
		_w9213_,
		_w9214_,
		_w9473_
	);
	LUT4 #(
		.INIT('h5554)
	) name3647 (
		_w9212_,
		_w9233_,
		_w9472_,
		_w9473_,
		_w9474_
	);
	LUT4 #(
		.INIT('hfb9f)
	) name3648 (
		_w9215_,
		_w9216_,
		_w9217_,
		_w9214_,
		_w9475_
	);
	LUT2 #(
		.INIT('h1)
	) name3649 (
		_w9213_,
		_w9475_,
		_w9476_
	);
	LUT3 #(
		.INIT('h01)
	) name3650 (
		_w9471_,
		_w9474_,
		_w9476_,
		_w9477_
	);
	LUT3 #(
		.INIT('h65)
	) name3651 (
		\u2_L8_reg[27]/NET0131 ,
		_w9468_,
		_w9477_,
		_w9478_
	);
	LUT4 #(
		.INIT('hb005)
	) name3652 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9479_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name3653 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9480_
	);
	LUT3 #(
		.INIT('h01)
	) name3654 (
		_w9071_,
		_w9479_,
		_w9480_,
		_w9481_
	);
	LUT3 #(
		.INIT('h08)
	) name3655 (
		_w9076_,
		_w9072_,
		_w9074_,
		_w9482_
	);
	LUT4 #(
		.INIT('hddfa)
	) name3656 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9483_
	);
	LUT4 #(
		.INIT('h1f15)
	) name3657 (
		_w9071_,
		_w9073_,
		_w9482_,
		_w9483_,
		_w9484_
	);
	LUT3 #(
		.INIT('h8a)
	) name3658 (
		_w9075_,
		_w9481_,
		_w9484_,
		_w9485_
	);
	LUT3 #(
		.INIT('h04)
	) name3659 (
		_w9076_,
		_w9072_,
		_w9074_,
		_w9486_
	);
	LUT4 #(
		.INIT('h8000)
	) name3660 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9487_
	);
	LUT4 #(
		.INIT('h7bd7)
	) name3661 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9488_
	);
	LUT3 #(
		.INIT('h40)
	) name3662 (
		_w9073_,
		_w9072_,
		_w9074_,
		_w9489_
	);
	LUT4 #(
		.INIT('h5153)
	) name3663 (
		_w9071_,
		_w9264_,
		_w9486_,
		_w9489_,
		_w9490_
	);
	LUT4 #(
		.INIT('h4404)
	) name3664 (
		_w9071_,
		_w9073_,
		_w9072_,
		_w9074_,
		_w9491_
	);
	LUT4 #(
		.INIT('h135f)
	) name3665 (
		_w9071_,
		_w9083_,
		_w9078_,
		_w9491_,
		_w9492_
	);
	LUT4 #(
		.INIT('hea00)
	) name3666 (
		_w9075_,
		_w9488_,
		_w9490_,
		_w9492_,
		_w9493_
	);
	LUT3 #(
		.INIT('h65)
	) name3667 (
		\u2_L8_reg[32]/NET0131 ,
		_w9485_,
		_w9493_,
		_w9494_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3668 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9495_
	);
	LUT4 #(
		.INIT('h22e6)
	) name3669 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9496_
	);
	LUT3 #(
		.INIT('h10)
	) name3670 (
		_w9294_,
		_w9495_,
		_w9496_,
		_w9497_
	);
	LUT4 #(
		.INIT('hbf3f)
	) name3671 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9498_
	);
	LUT3 #(
		.INIT('h40)
	) name3672 (
		_w9314_,
		_w9294_,
		_w9498_,
		_w9499_
	);
	LUT4 #(
		.INIT('h0800)
	) name3673 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9500_
	);
	LUT4 #(
		.INIT('h0001)
	) name3674 (
		_w9295_,
		_w9319_,
		_w9456_,
		_w9500_,
		_w9501_
	);
	LUT3 #(
		.INIT('he0)
	) name3675 (
		_w9497_,
		_w9499_,
		_w9501_,
		_w9502_
	);
	LUT4 #(
		.INIT('h1098)
	) name3676 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9503_
	);
	LUT3 #(
		.INIT('h04)
	) name3677 (
		_w9314_,
		_w9294_,
		_w9503_,
		_w9504_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name3678 (
		_w9296_,
		_w9298_,
		_w9297_,
		_w9299_,
		_w9505_
	);
	LUT3 #(
		.INIT('h10)
	) name3679 (
		_w9294_,
		_w9495_,
		_w9505_,
		_w9506_
	);
	LUT3 #(
		.INIT('h02)
	) name3680 (
		_w9295_,
		_w9301_,
		_w9317_,
		_w9507_
	);
	LUT3 #(
		.INIT('he0)
	) name3681 (
		_w9504_,
		_w9506_,
		_w9507_,
		_w9508_
	);
	LUT3 #(
		.INIT('ha9)
	) name3682 (
		\u2_L8_reg[3]/NET0131 ,
		_w9502_,
		_w9508_,
		_w9509_
	);
	LUT4 #(
		.INIT('hc693)
	) name3683 (
		decrypt_pad,
		\u2_R8_reg[13]/NET0131 ,
		\u2_uk_K_r8_reg[25]/NET0131 ,
		\u2_uk_K_r8_reg[3]/NET0131 ,
		_w9510_
	);
	LUT4 #(
		.INIT('hc693)
	) name3684 (
		decrypt_pad,
		\u2_R8_reg[9]/NET0131 ,
		\u2_uk_K_r8_reg[20]/NET0131 ,
		\u2_uk_K_r8_reg[55]/NET0131 ,
		_w9511_
	);
	LUT4 #(
		.INIT('hc963)
	) name3685 (
		decrypt_pad,
		\u2_R8_reg[11]/NET0131 ,
		\u2_uk_K_r8_reg[32]/NET0131 ,
		\u2_uk_K_r8_reg[54]/NET0131 ,
		_w9512_
	);
	LUT3 #(
		.INIT('h0b)
	) name3686 (
		_w9510_,
		_w9511_,
		_w9512_,
		_w9513_
	);
	LUT4 #(
		.INIT('hc693)
	) name3687 (
		decrypt_pad,
		\u2_R8_reg[10]/NET0131 ,
		\u2_uk_K_r8_reg[53]/NET0131 ,
		\u2_uk_K_r8_reg[6]/NET0131 ,
		_w9514_
	);
	LUT4 #(
		.INIT('hc963)
	) name3688 (
		decrypt_pad,
		\u2_R8_reg[8]/NET0131 ,
		\u2_uk_K_r8_reg[26]/NET0131 ,
		\u2_uk_K_r8_reg[48]/NET0131 ,
		_w9515_
	);
	LUT4 #(
		.INIT('h3b0b)
	) name3689 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9516_
	);
	LUT4 #(
		.INIT('h1000)
	) name3690 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9517_
	);
	LUT4 #(
		.INIT('hc693)
	) name3691 (
		decrypt_pad,
		\u2_R8_reg[12]/NET0131 ,
		\u2_uk_K_r8_reg[12]/NET0131 ,
		\u2_uk_K_r8_reg[47]/NET0131 ,
		_w9518_
	);
	LUT4 #(
		.INIT('h5100)
	) name3692 (
		_w9517_,
		_w9513_,
		_w9516_,
		_w9518_,
		_w9519_
	);
	LUT2 #(
		.INIT('h6)
	) name3693 (
		_w9510_,
		_w9515_,
		_w9520_
	);
	LUT4 #(
		.INIT('h9990)
	) name3694 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9521_
	);
	LUT4 #(
		.INIT('h0990)
	) name3695 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9522_
	);
	LUT4 #(
		.INIT('h4000)
	) name3696 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9523_
	);
	LUT4 #(
		.INIT('h0400)
	) name3697 (
		_w9515_,
		_w9511_,
		_w9514_,
		_w9512_,
		_w9524_
	);
	LUT3 #(
		.INIT('h01)
	) name3698 (
		_w9518_,
		_w9524_,
		_w9523_,
		_w9525_
	);
	LUT4 #(
		.INIT('h2000)
	) name3699 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9526_
	);
	LUT4 #(
		.INIT('h0203)
	) name3700 (
		_w9515_,
		_w9511_,
		_w9514_,
		_w9512_,
		_w9527_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3701 (
		_w9512_,
		_w9526_,
		_w9520_,
		_w9527_,
		_w9528_
	);
	LUT4 #(
		.INIT('h4555)
	) name3702 (
		_w9519_,
		_w9522_,
		_w9525_,
		_w9528_,
		_w9529_
	);
	LUT4 #(
		.INIT('h95b5)
	) name3703 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9530_
	);
	LUT4 #(
		.INIT('h0001)
	) name3704 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9531_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name3705 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9532_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3706 (
		_w9512_,
		_w9518_,
		_w9530_,
		_w9532_,
		_w9533_
	);
	LUT3 #(
		.INIT('h56)
	) name3707 (
		\u2_L8_reg[6]/NET0131 ,
		_w9529_,
		_w9533_,
		_w9534_
	);
	LUT4 #(
		.INIT('h0770)
	) name3708 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9535_
	);
	LUT4 #(
		.INIT('h3882)
	) name3709 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9074_,
		_w9536_
	);
	LUT2 #(
		.INIT('h4)
	) name3710 (
		_w9071_,
		_w9075_,
		_w9537_
	);
	LUT2 #(
		.INIT('h9)
	) name3711 (
		_w9071_,
		_w9075_,
		_w9538_
	);
	LUT3 #(
		.INIT('h10)
	) name3712 (
		_w9084_,
		_w9536_,
		_w9538_,
		_w9539_
	);
	LUT3 #(
		.INIT('h09)
	) name3713 (
		_w9073_,
		_w9076_,
		_w9072_,
		_w9540_
	);
	LUT3 #(
		.INIT('h28)
	) name3714 (
		_w9073_,
		_w9072_,
		_w9074_,
		_w9541_
	);
	LUT4 #(
		.INIT('h0004)
	) name3715 (
		_w9482_,
		_w9537_,
		_w9541_,
		_w9540_,
		_w9542_
	);
	LUT4 #(
		.INIT('h0004)
	) name3716 (
		_w9079_,
		_w9260_,
		_w9487_,
		_w9535_,
		_w9543_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3717 (
		_w9258_,
		_w9539_,
		_w9542_,
		_w9543_,
		_w9544_
	);
	LUT2 #(
		.INIT('h6)
	) name3718 (
		\u2_L8_reg[7]/NET0131 ,
		_w9544_,
		_w9545_
	);
	LUT3 #(
		.INIT('h9f)
	) name3719 (
		_w9015_,
		_w9011_,
		_w9012_,
		_w9546_
	);
	LUT2 #(
		.INIT('h2)
	) name3720 (
		_w9020_,
		_w9546_,
		_w9547_
	);
	LUT3 #(
		.INIT('h43)
	) name3721 (
		_w9015_,
		_w9016_,
		_w9012_,
		_w9548_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name3722 (
		_w9015_,
		_w9011_,
		_w9014_,
		_w9012_,
		_w9549_
	);
	LUT3 #(
		.INIT('h84)
	) name3723 (
		_w9016_,
		_w9014_,
		_w9012_,
		_w9550_
	);
	LUT3 #(
		.INIT('h0e)
	) name3724 (
		_w9548_,
		_w9549_,
		_w9550_,
		_w9551_
	);
	LUT4 #(
		.INIT('h2810)
	) name3725 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9552_
	);
	LUT2 #(
		.INIT('h1)
	) name3726 (
		_w9010_,
		_w9552_,
		_w9553_
	);
	LUT4 #(
		.INIT('h9060)
	) name3727 (
		_w9015_,
		_w9016_,
		_w9011_,
		_w9012_,
		_w9554_
	);
	LUT4 #(
		.INIT('h040c)
	) name3728 (
		_w9023_,
		_w9010_,
		_w9103_,
		_w9548_,
		_w9555_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3729 (
		_w9551_,
		_w9553_,
		_w9554_,
		_w9555_,
		_w9556_
	);
	LUT3 #(
		.INIT('h56)
	) name3730 (
		\u2_L8_reg[9]/NET0131 ,
		_w9547_,
		_w9556_,
		_w9557_
	);
	LUT4 #(
		.INIT('h6979)
	) name3731 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9512_,
		_w9558_
	);
	LUT3 #(
		.INIT('h07)
	) name3732 (
		_w9515_,
		_w9514_,
		_w9512_,
		_w9559_
	);
	LUT4 #(
		.INIT('h0014)
	) name3733 (
		_w9510_,
		_w9515_,
		_w9514_,
		_w9512_,
		_w9560_
	);
	LUT4 #(
		.INIT('h0032)
	) name3734 (
		_w9514_,
		_w9526_,
		_w9558_,
		_w9560_,
		_w9561_
	);
	LUT3 #(
		.INIT('he0)
	) name3735 (
		_w9510_,
		_w9515_,
		_w9512_,
		_w9562_
	);
	LUT4 #(
		.INIT('h6800)
	) name3736 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9512_,
		_w9563_
	);
	LUT3 #(
		.INIT('h0d)
	) name3737 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9564_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name3738 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9565_
	);
	LUT4 #(
		.INIT('h0f02)
	) name3739 (
		_w9512_,
		_w9531_,
		_w9563_,
		_w9565_,
		_w9566_
	);
	LUT3 #(
		.INIT('h08)
	) name3740 (
		_w9515_,
		_w9514_,
		_w9512_,
		_w9567_
	);
	LUT4 #(
		.INIT('h0020)
	) name3741 (
		_w9515_,
		_w9511_,
		_w9514_,
		_w9512_,
		_w9568_
	);
	LUT4 #(
		.INIT('hbeff)
	) name3742 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9569_
	);
	LUT3 #(
		.INIT('h31)
	) name3743 (
		_w9512_,
		_w9568_,
		_w9569_,
		_w9570_
	);
	LUT4 #(
		.INIT('hd800)
	) name3744 (
		_w9518_,
		_w9561_,
		_w9566_,
		_w9570_,
		_w9571_
	);
	LUT2 #(
		.INIT('h9)
	) name3745 (
		\u2_L8_reg[16]/NET0131 ,
		_w9571_,
		_w9572_
	);
	LUT4 #(
		.INIT('h2600)
	) name3746 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9156_,
		_w9573_
	);
	LUT4 #(
		.INIT('hef2f)
	) name3747 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9574_
	);
	LUT4 #(
		.INIT('h0032)
	) name3748 (
		_w9156_,
		_w9176_,
		_w9574_,
		_w9573_,
		_w9575_
	);
	LUT4 #(
		.INIT('h0121)
	) name3749 (
		_w9154_,
		_w9151_,
		_w9155_,
		_w9156_,
		_w9576_
	);
	LUT4 #(
		.INIT('h6000)
	) name3750 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9155_,
		_w9577_
	);
	LUT4 #(
		.INIT('h8000)
	) name3751 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9156_,
		_w9578_
	);
	LUT4 #(
		.INIT('h0001)
	) name3752 (
		_w9288_,
		_w9578_,
		_w9577_,
		_w9576_,
		_w9579_
	);
	LUT4 #(
		.INIT('h0008)
	) name3753 (
		_w9154_,
		_w9150_,
		_w9151_,
		_w9156_,
		_w9580_
	);
	LUT4 #(
		.INIT('h8300)
	) name3754 (
		_w9150_,
		_w9151_,
		_w9155_,
		_w9156_,
		_w9581_
	);
	LUT3 #(
		.INIT('h23)
	) name3755 (
		_w9436_,
		_w9580_,
		_w9581_,
		_w9582_
	);
	LUT4 #(
		.INIT('he400)
	) name3756 (
		_w9160_,
		_w9579_,
		_w9575_,
		_w9582_,
		_w9583_
	);
	LUT2 #(
		.INIT('h9)
	) name3757 (
		\u2_L8_reg[18]/P0001 ,
		_w9583_,
		_w9584_
	);
	LUT3 #(
		.INIT('hed)
	) name3758 (
		_w9510_,
		_w9515_,
		_w9514_,
		_w9585_
	);
	LUT3 #(
		.INIT('h20)
	) name3759 (
		_w9515_,
		_w9511_,
		_w9514_,
		_w9586_
	);
	LUT4 #(
		.INIT('hef00)
	) name3760 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9512_,
		_w9587_
	);
	LUT3 #(
		.INIT('h20)
	) name3761 (
		_w9585_,
		_w9586_,
		_w9587_,
		_w9588_
	);
	LUT4 #(
		.INIT('h0009)
	) name3762 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9589_
	);
	LUT4 #(
		.INIT('h6640)
	) name3763 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9590_
	);
	LUT3 #(
		.INIT('h01)
	) name3764 (
		_w9512_,
		_w9590_,
		_w9589_,
		_w9591_
	);
	LUT3 #(
		.INIT('h54)
	) name3765 (
		_w9518_,
		_w9588_,
		_w9591_,
		_w9592_
	);
	LUT2 #(
		.INIT('h4)
	) name3766 (
		_w9512_,
		_w9521_,
		_w9593_
	);
	LUT3 #(
		.INIT('h2a)
	) name3767 (
		_w9518_,
		_w9520_,
		_w9527_,
		_w9594_
	);
	LUT3 #(
		.INIT('hd0)
	) name3768 (
		_w9515_,
		_w9511_,
		_w9514_,
		_w9595_
	);
	LUT2 #(
		.INIT('h4)
	) name3769 (
		_w9514_,
		_w9512_,
		_w9596_
	);
	LUT4 #(
		.INIT('h153f)
	) name3770 (
		_w9562_,
		_w9564_,
		_w9596_,
		_w9595_,
		_w9597_
	);
	LUT3 #(
		.INIT('h40)
	) name3771 (
		_w9593_,
		_w9594_,
		_w9597_,
		_w9598_
	);
	LUT2 #(
		.INIT('h8)
	) name3772 (
		_w9510_,
		_w9511_,
		_w9599_
	);
	LUT3 #(
		.INIT('h53)
	) name3773 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9600_
	);
	LUT4 #(
		.INIT('h0700)
	) name3774 (
		_w9510_,
		_w9515_,
		_w9514_,
		_w9512_,
		_w9601_
	);
	LUT4 #(
		.INIT('h7077)
	) name3775 (
		_w9567_,
		_w9599_,
		_w9600_,
		_w9601_,
		_w9602_
	);
	LUT4 #(
		.INIT('ha955)
	) name3776 (
		\u2_L8_reg[24]/NET0131 ,
		_w9592_,
		_w9598_,
		_w9602_,
		_w9603_
	);
	LUT4 #(
		.INIT('h8c00)
	) name3777 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9604_
	);
	LUT4 #(
		.INIT('h00fb)
	) name3778 (
		_w9510_,
		_w9511_,
		_w9514_,
		_w9518_,
		_w9605_
	);
	LUT2 #(
		.INIT('h4)
	) name3779 (
		_w9604_,
		_w9605_,
		_w9606_
	);
	LUT4 #(
		.INIT('h0004)
	) name3780 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9607_
	);
	LUT4 #(
		.INIT('haa2a)
	) name3781 (
		_w9512_,
		_w9518_,
		_w9585_,
		_w9607_,
		_w9608_
	);
	LUT2 #(
		.INIT('h4)
	) name3782 (
		_w9606_,
		_w9608_,
		_w9609_
	);
	LUT4 #(
		.INIT('h23ef)
	) name3783 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9610_
	);
	LUT4 #(
		.INIT('h7000)
	) name3784 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9611_
	);
	LUT4 #(
		.INIT('h0c08)
	) name3785 (
		_w9512_,
		_w9518_,
		_w9611_,
		_w9610_,
		_w9612_
	);
	LUT2 #(
		.INIT('h1)
	) name3786 (
		_w9518_,
		_w9589_,
		_w9613_
	);
	LUT4 #(
		.INIT('h0200)
	) name3787 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9514_,
		_w9614_
	);
	LUT3 #(
		.INIT('h0d)
	) name3788 (
		_w9559_,
		_w9600_,
		_w9614_,
		_w9615_
	);
	LUT4 #(
		.INIT('hf700)
	) name3789 (
		_w9510_,
		_w9515_,
		_w9511_,
		_w9512_,
		_w9616_
	);
	LUT4 #(
		.INIT('hf040)
	) name3790 (
		_w9510_,
		_w9511_,
		_w9514_,
		_w9512_,
		_w9617_
	);
	LUT2 #(
		.INIT('h4)
	) name3791 (
		_w9616_,
		_w9617_,
		_w9618_
	);
	LUT4 #(
		.INIT('h00ea)
	) name3792 (
		_w9612_,
		_w9613_,
		_w9615_,
		_w9618_,
		_w9619_
	);
	LUT3 #(
		.INIT('h9a)
	) name3793 (
		\u2_L8_reg[30]/NET0131 ,
		_w9609_,
		_w9619_,
		_w9620_
	);
	LUT4 #(
		.INIT('hc693)
	) name3794 (
		decrypt_pad,
		\u2_R7_reg[26]/NET0131 ,
		\u2_uk_K_r7_reg[31]/NET0131 ,
		\u2_uk_K_r7_reg[38]/NET0131 ,
		_w9621_
	);
	LUT4 #(
		.INIT('hc693)
	) name3795 (
		decrypt_pad,
		\u2_R7_reg[25]/NET0131 ,
		\u2_uk_K_r7_reg[42]/NET0131 ,
		\u2_uk_K_r7_reg[49]/NET0131 ,
		_w9622_
	);
	LUT4 #(
		.INIT('hc963)
	) name3796 (
		decrypt_pad,
		\u2_R7_reg[24]/NET0131 ,
		\u2_uk_K_r7_reg[14]/NET0131 ,
		\u2_uk_K_r7_reg[7]/NET0131 ,
		_w9623_
	);
	LUT4 #(
		.INIT('hc693)
	) name3797 (
		decrypt_pad,
		\u2_R7_reg[29]/NET0131 ,
		\u2_uk_K_r7_reg[15]/NET0131 ,
		\u2_uk_K_r7_reg[22]/NET0131 ,
		_w9624_
	);
	LUT2 #(
		.INIT('h4)
	) name3798 (
		_w9623_,
		_w9624_,
		_w9625_
	);
	LUT4 #(
		.INIT('h0200)
	) name3799 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9626_
	);
	LUT4 #(
		.INIT('h0008)
	) name3800 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9627_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name3801 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9628_
	);
	LUT4 #(
		.INIT('hc693)
	) name3802 (
		decrypt_pad,
		\u2_R7_reg[28]/NET0131 ,
		\u2_uk_K_r7_reg[23]/P0001 ,
		\u2_uk_K_r7_reg[30]/P0001 ,
		_w9629_
	);
	LUT4 #(
		.INIT('h9cfc)
	) name3803 (
		_w9621_,
		_w9622_,
		_w9624_,
		_w9629_,
		_w9630_
	);
	LUT4 #(
		.INIT('hc693)
	) name3804 (
		decrypt_pad,
		\u2_R7_reg[27]/NET0131 ,
		\u2_uk_K_r7_reg[36]/NET0131 ,
		\u2_uk_K_r7_reg[43]/NET0131 ,
		_w9631_
	);
	LUT4 #(
		.INIT('h3b00)
	) name3805 (
		_w9623_,
		_w9628_,
		_w9630_,
		_w9631_,
		_w9632_
	);
	LUT2 #(
		.INIT('h4)
	) name3806 (
		_w9622_,
		_w9631_,
		_w9633_
	);
	LUT4 #(
		.INIT('heef2)
	) name3807 (
		_w9621_,
		_w9622_,
		_w9624_,
		_w9631_,
		_w9634_
	);
	LUT2 #(
		.INIT('h6)
	) name3808 (
		_w9621_,
		_w9623_,
		_w9635_
	);
	LUT4 #(
		.INIT('h0002)
	) name3809 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9636_
	);
	LUT4 #(
		.INIT('h5afd)
	) name3810 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9637_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name3811 (
		_w9623_,
		_w9633_,
		_w9634_,
		_w9637_,
		_w9638_
	);
	LUT4 #(
		.INIT('h1000)
	) name3812 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9639_
	);
	LUT4 #(
		.INIT('he3ff)
	) name3813 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9640_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name3814 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9641_
	);
	LUT3 #(
		.INIT('he0)
	) name3815 (
		_w9631_,
		_w9640_,
		_w9641_,
		_w9642_
	);
	LUT4 #(
		.INIT('h0100)
	) name3816 (
		_w9621_,
		_w9622_,
		_w9624_,
		_w9631_,
		_w9643_
	);
	LUT4 #(
		.INIT('h0084)
	) name3817 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9631_,
		_w9644_
	);
	LUT2 #(
		.INIT('h1)
	) name3818 (
		_w9643_,
		_w9644_,
		_w9645_
	);
	LUT4 #(
		.INIT('he400)
	) name3819 (
		_w9629_,
		_w9638_,
		_w9642_,
		_w9645_,
		_w9646_
	);
	LUT3 #(
		.INIT('h65)
	) name3820 (
		\u2_L7_reg[22]/NET0131 ,
		_w9632_,
		_w9646_,
		_w9647_
	);
	LUT4 #(
		.INIT('hc693)
	) name3821 (
		decrypt_pad,
		\u2_R7_reg[4]/NET0131 ,
		\u2_uk_K_r7_reg[47]/NET0131 ,
		\u2_uk_K_r7_reg[54]/NET0131 ,
		_w9648_
	);
	LUT4 #(
		.INIT('hc693)
	) name3822 (
		decrypt_pad,
		\u2_R7_reg[3]/NET0131 ,
		\u2_uk_K_r7_reg[12]/NET0131 ,
		\u2_uk_K_r7_reg[19]/NET0131 ,
		_w9649_
	);
	LUT4 #(
		.INIT('hc693)
	) name3823 (
		decrypt_pad,
		\u2_R7_reg[1]/NET0131 ,
		\u2_uk_K_r7_reg[20]/NET0131 ,
		\u2_uk_K_r7_reg[27]/NET0131 ,
		_w9650_
	);
	LUT4 #(
		.INIT('hc693)
	) name3824 (
		decrypt_pad,
		\u2_R7_reg[5]/NET0131 ,
		\u2_uk_K_r7_reg[18]/NET0131 ,
		\u2_uk_K_r7_reg[25]/NET0131 ,
		_w9651_
	);
	LUT4 #(
		.INIT('hc963)
	) name3825 (
		decrypt_pad,
		\u2_R7_reg[2]/NET0131 ,
		\u2_uk_K_r7_reg[10]/NET0131 ,
		\u2_uk_K_r7_reg[3]/NET0131 ,
		_w9652_
	);
	LUT4 #(
		.INIT('hc693)
	) name3826 (
		decrypt_pad,
		\u2_R7_reg[32]/NET0131 ,
		\u2_uk_K_r7_reg[24]/NET0131 ,
		\u2_uk_K_r7_reg[6]/NET0131 ,
		_w9653_
	);
	LUT3 #(
		.INIT('heb)
	) name3827 (
		_w9653_,
		_w9652_,
		_w9651_,
		_w9654_
	);
	LUT4 #(
		.INIT('hc8af)
	) name3828 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9655_
	);
	LUT2 #(
		.INIT('h4)
	) name3829 (
		_w9650_,
		_w9652_,
		_w9656_
	);
	LUT4 #(
		.INIT('h1908)
	) name3830 (
		_w9653_,
		_w9650_,
		_w9649_,
		_w9652_,
		_w9657_
	);
	LUT4 #(
		.INIT('h1102)
	) name3831 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9658_
	);
	LUT4 #(
		.INIT('h000d)
	) name3832 (
		_w9649_,
		_w9655_,
		_w9657_,
		_w9658_,
		_w9659_
	);
	LUT2 #(
		.INIT('h2)
	) name3833 (
		_w9648_,
		_w9659_,
		_w9660_
	);
	LUT4 #(
		.INIT('h5dbb)
	) name3834 (
		_w9653_,
		_w9650_,
		_w9649_,
		_w9651_,
		_w9661_
	);
	LUT2 #(
		.INIT('h1)
	) name3835 (
		_w9652_,
		_w9661_,
		_w9662_
	);
	LUT3 #(
		.INIT('h48)
	) name3836 (
		_w9653_,
		_w9650_,
		_w9651_,
		_w9663_
	);
	LUT2 #(
		.INIT('h1)
	) name3837 (
		_w9650_,
		_w9651_,
		_w9664_
	);
	LUT4 #(
		.INIT('hfbda)
	) name3838 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9665_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name3839 (
		_w9649_,
		_w9652_,
		_w9663_,
		_w9665_,
		_w9666_
	);
	LUT3 #(
		.INIT('h45)
	) name3840 (
		_w9648_,
		_w9662_,
		_w9666_,
		_w9667_
	);
	LUT4 #(
		.INIT('h1000)
	) name3841 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9668_
	);
	LUT4 #(
		.INIT('h6ff3)
	) name3842 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9669_
	);
	LUT2 #(
		.INIT('h1)
	) name3843 (
		_w9649_,
		_w9669_,
		_w9670_
	);
	LUT2 #(
		.INIT('h2)
	) name3844 (
		_w9649_,
		_w9652_,
		_w9671_
	);
	LUT4 #(
		.INIT('h0020)
	) name3845 (
		_w9653_,
		_w9650_,
		_w9649_,
		_w9652_,
		_w9672_
	);
	LUT3 #(
		.INIT('h04)
	) name3846 (
		_w9653_,
		_w9649_,
		_w9651_,
		_w9673_
	);
	LUT3 #(
		.INIT('h15)
	) name3847 (
		_w9672_,
		_w9656_,
		_w9673_,
		_w9674_
	);
	LUT2 #(
		.INIT('h4)
	) name3848 (
		_w9670_,
		_w9674_,
		_w9675_
	);
	LUT4 #(
		.INIT('h5655)
	) name3849 (
		\u2_L7_reg[31]/NET0131 ,
		_w9667_,
		_w9660_,
		_w9675_,
		_w9676_
	);
	LUT4 #(
		.INIT('hc693)
	) name3850 (
		decrypt_pad,
		\u2_R7_reg[24]/NET0131 ,
		\u2_uk_K_r7_reg[16]/NET0131 ,
		\u2_uk_K_r7_reg[23]/P0001 ,
		_w9677_
	);
	LUT4 #(
		.INIT('hc693)
	) name3851 (
		decrypt_pad,
		\u2_R7_reg[23]/NET0131 ,
		\u2_uk_K_r7_reg[14]/NET0131 ,
		\u2_uk_K_r7_reg[21]/NET0131 ,
		_w9678_
	);
	LUT4 #(
		.INIT('hc963)
	) name3852 (
		decrypt_pad,
		\u2_R7_reg[20]/NET0131 ,
		\u2_uk_K_r7_reg[2]/NET0131 ,
		\u2_uk_K_r7_reg[50]/NET0131 ,
		_w9679_
	);
	LUT4 #(
		.INIT('hc693)
	) name3853 (
		decrypt_pad,
		\u2_R7_reg[21]/NET0131 ,
		\u2_uk_K_r7_reg[38]/NET0131 ,
		\u2_uk_K_r7_reg[45]/NET0131 ,
		_w9680_
	);
	LUT4 #(
		.INIT('hc693)
	) name3854 (
		decrypt_pad,
		\u2_R7_reg[22]/NET0131 ,
		\u2_uk_K_r7_reg[1]/NET0131 ,
		\u2_uk_K_r7_reg[8]/NET0131 ,
		_w9681_
	);
	LUT4 #(
		.INIT('hc693)
	) name3855 (
		decrypt_pad,
		\u2_R7_reg[25]/NET0131 ,
		\u2_uk_K_r7_reg[35]/NET0131 ,
		\u2_uk_K_r7_reg[42]/NET0131 ,
		_w9682_
	);
	LUT4 #(
		.INIT('heb73)
	) name3856 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9683_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		_w9678_,
		_w9683_,
		_w9684_
	);
	LUT2 #(
		.INIT('h2)
	) name3858 (
		_w9679_,
		_w9682_,
		_w9685_
	);
	LUT4 #(
		.INIT('h0002)
	) name3859 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9686_
	);
	LUT4 #(
		.INIT('h1fbd)
	) name3860 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9687_
	);
	LUT2 #(
		.INIT('h1)
	) name3861 (
		_w9678_,
		_w9681_,
		_w9688_
	);
	LUT4 #(
		.INIT('h0400)
	) name3862 (
		_w9678_,
		_w9679_,
		_w9681_,
		_w9682_,
		_w9689_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3863 (
		_w9678_,
		_w9680_,
		_w9687_,
		_w9689_,
		_w9690_
	);
	LUT3 #(
		.INIT('h8a)
	) name3864 (
		_w9677_,
		_w9684_,
		_w9690_,
		_w9691_
	);
	LUT4 #(
		.INIT('h1682)
	) name3865 (
		_w9678_,
		_w9679_,
		_w9681_,
		_w9680_,
		_w9692_
	);
	LUT3 #(
		.INIT('hce)
	) name3866 (
		_w9678_,
		_w9681_,
		_w9680_,
		_w9693_
	);
	LUT4 #(
		.INIT('h0800)
	) name3867 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9694_
	);
	LUT4 #(
		.INIT('h0200)
	) name3868 (
		_w9678_,
		_w9679_,
		_w9680_,
		_w9682_,
		_w9695_
	);
	LUT4 #(
		.INIT('h1101)
	) name3869 (
		_w9694_,
		_w9695_,
		_w9685_,
		_w9693_,
		_w9696_
	);
	LUT3 #(
		.INIT('h45)
	) name3870 (
		_w9677_,
		_w9692_,
		_w9696_,
		_w9697_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name3871 (
		_w9678_,
		_w9679_,
		_w9680_,
		_w9682_,
		_w9698_
	);
	LUT2 #(
		.INIT('h1)
	) name3872 (
		_w9681_,
		_w9698_,
		_w9699_
	);
	LUT4 #(
		.INIT('h3323)
	) name3873 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9700_
	);
	LUT4 #(
		.INIT('h8a0a)
	) name3874 (
		_w9678_,
		_w9679_,
		_w9681_,
		_w9682_,
		_w9701_
	);
	LUT3 #(
		.INIT('h01)
	) name3875 (
		_w9679_,
		_w9680_,
		_w9682_,
		_w9702_
	);
	LUT4 #(
		.INIT('h45cf)
	) name3876 (
		_w9688_,
		_w9700_,
		_w9701_,
		_w9702_,
		_w9703_
	);
	LUT2 #(
		.INIT('h4)
	) name3877 (
		_w9699_,
		_w9703_,
		_w9704_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name3878 (
		\u2_L7_reg[11]/NET0131 ,
		_w9697_,
		_w9691_,
		_w9704_,
		_w9705_
	);
	LUT4 #(
		.INIT('hc963)
	) name3879 (
		decrypt_pad,
		\u2_R7_reg[17]/NET0131 ,
		\u2_uk_K_r7_reg[4]/NET0131 ,
		\u2_uk_K_r7_reg[54]/NET0131 ,
		_w9706_
	);
	LUT4 #(
		.INIT('hc693)
	) name3880 (
		decrypt_pad,
		\u2_R7_reg[12]/NET0131 ,
		\u2_uk_K_r7_reg[13]/NET0131 ,
		\u2_uk_K_r7_reg[20]/NET0131 ,
		_w9707_
	);
	LUT2 #(
		.INIT('h4)
	) name3881 (
		_w9706_,
		_w9707_,
		_w9708_
	);
	LUT4 #(
		.INIT('hc693)
	) name3882 (
		decrypt_pad,
		\u2_R7_reg[14]/NET0131 ,
		\u2_uk_K_r7_reg[33]/NET0131 ,
		\u2_uk_K_r7_reg[40]/NET0131 ,
		_w9709_
	);
	LUT4 #(
		.INIT('hc693)
	) name3883 (
		decrypt_pad,
		\u2_R7_reg[13]/NET0131 ,
		\u2_uk_K_r7_reg[32]/NET0131 ,
		\u2_uk_K_r7_reg[39]/NET0131 ,
		_w9710_
	);
	LUT4 #(
		.INIT('hc693)
	) name3884 (
		decrypt_pad,
		\u2_R7_reg[15]/NET0131 ,
		\u2_uk_K_r7_reg[41]/NET0131 ,
		\u2_uk_K_r7_reg[48]/NET0131 ,
		_w9711_
	);
	LUT4 #(
		.INIT('hc080)
	) name3885 (
		_w9707_,
		_w9710_,
		_w9711_,
		_w9709_,
		_w9712_
	);
	LUT4 #(
		.INIT('h0001)
	) name3886 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9713_
	);
	LUT4 #(
		.INIT('hc693)
	) name3887 (
		decrypt_pad,
		\u2_R7_reg[16]/NET0131 ,
		\u2_uk_K_r7_reg[17]/NET0131 ,
		\u2_uk_K_r7_reg[24]/NET0131 ,
		_w9714_
	);
	LUT4 #(
		.INIT('h000b)
	) name3888 (
		_w9708_,
		_w9712_,
		_w9713_,
		_w9714_,
		_w9715_
	);
	LUT3 #(
		.INIT('h15)
	) name3889 (
		_w9706_,
		_w9707_,
		_w9709_,
		_w9716_
	);
	LUT3 #(
		.INIT('h07)
	) name3890 (
		_w9706_,
		_w9710_,
		_w9711_,
		_w9717_
	);
	LUT4 #(
		.INIT('h1000)
	) name3891 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9718_
	);
	LUT3 #(
		.INIT('h0b)
	) name3892 (
		_w9716_,
		_w9717_,
		_w9718_,
		_w9719_
	);
	LUT4 #(
		.INIT('h0008)
	) name3893 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9720_
	);
	LUT2 #(
		.INIT('h1)
	) name3894 (
		_w9706_,
		_w9710_,
		_w9721_
	);
	LUT4 #(
		.INIT('h0100)
	) name3895 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9711_,
		_w9722_
	);
	LUT2 #(
		.INIT('h1)
	) name3896 (
		_w9720_,
		_w9722_,
		_w9723_
	);
	LUT3 #(
		.INIT('h80)
	) name3897 (
		_w9715_,
		_w9719_,
		_w9723_,
		_w9724_
	);
	LUT3 #(
		.INIT('h06)
	) name3898 (
		_w9707_,
		_w9710_,
		_w9709_,
		_w9725_
	);
	LUT3 #(
		.INIT('h10)
	) name3899 (
		_w9707_,
		_w9710_,
		_w9709_,
		_w9726_
	);
	LUT4 #(
		.INIT('h0100)
	) name3900 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9727_
	);
	LUT4 #(
		.INIT('hfec3)
	) name3901 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9728_
	);
	LUT2 #(
		.INIT('h1)
	) name3902 (
		_w9711_,
		_w9728_,
		_w9729_
	);
	LUT3 #(
		.INIT('h40)
	) name3903 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9730_
	);
	LUT4 #(
		.INIT('h4000)
	) name3904 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9711_,
		_w9731_
	);
	LUT2 #(
		.INIT('h6)
	) name3905 (
		_w9707_,
		_w9709_,
		_w9732_
	);
	LUT4 #(
		.INIT('h8020)
	) name3906 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9733_
	);
	LUT4 #(
		.INIT('h0200)
	) name3907 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9711_,
		_w9734_
	);
	LUT4 #(
		.INIT('h0004)
	) name3908 (
		_w9731_,
		_w9714_,
		_w9733_,
		_w9734_,
		_w9735_
	);
	LUT2 #(
		.INIT('h4)
	) name3909 (
		_w9729_,
		_w9735_,
		_w9736_
	);
	LUT4 #(
		.INIT('hbfdf)
	) name3910 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9711_,
		_w9737_
	);
	LUT3 #(
		.INIT('h84)
	) name3911 (
		_w9707_,
		_w9711_,
		_w9709_,
		_w9738_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3912 (
		_w9737_,
		_w9709_,
		_w9721_,
		_w9738_,
		_w9739_
	);
	LUT4 #(
		.INIT('ha955)
	) name3913 (
		\u2_L7_reg[20]/NET0131 ,
		_w9724_,
		_w9736_,
		_w9739_,
		_w9740_
	);
	LUT4 #(
		.INIT('hc693)
	) name3914 (
		decrypt_pad,
		\u2_R7_reg[28]/NET0131 ,
		\u2_uk_K_r7_reg[21]/NET0131 ,
		\u2_uk_K_r7_reg[28]/NET0131 ,
		_w9741_
	);
	LUT4 #(
		.INIT('hc963)
	) name3915 (
		decrypt_pad,
		\u2_R7_reg[1]/NET0131 ,
		\u2_uk_K_r7_reg[16]/NET0131 ,
		\u2_uk_K_r7_reg[9]/NET0131 ,
		_w9742_
	);
	LUT4 #(
		.INIT('hc963)
	) name3916 (
		decrypt_pad,
		\u2_R7_reg[29]/NET0131 ,
		\u2_uk_K_r7_reg[0]/NET0131 ,
		\u2_uk_K_r7_reg[52]/NET0131 ,
		_w9743_
	);
	LUT4 #(
		.INIT('hc963)
	) name3917 (
		decrypt_pad,
		\u2_R7_reg[30]/NET0131 ,
		\u2_uk_K_r7_reg[1]/NET0131 ,
		\u2_uk_K_r7_reg[49]/NET0131 ,
		_w9744_
	);
	LUT4 #(
		.INIT('h0200)
	) name3918 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9745_
	);
	LUT4 #(
		.INIT('hf9fb)
	) name3919 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9746_
	);
	LUT4 #(
		.INIT('hc693)
	) name3920 (
		decrypt_pad,
		\u2_R7_reg[31]/P0001 ,
		\u2_uk_K_r7_reg[37]/NET0131 ,
		\u2_uk_K_r7_reg[44]/NET0131 ,
		_w9747_
	);
	LUT2 #(
		.INIT('h4)
	) name3921 (
		_w9746_,
		_w9747_,
		_w9748_
	);
	LUT3 #(
		.INIT('h0d)
	) name3922 (
		_w9741_,
		_w9742_,
		_w9747_,
		_w9749_
	);
	LUT2 #(
		.INIT('h2)
	) name3923 (
		_w9742_,
		_w9743_,
		_w9750_
	);
	LUT3 #(
		.INIT('hd8)
	) name3924 (
		_w9742_,
		_w9743_,
		_w9744_,
		_w9751_
	);
	LUT2 #(
		.INIT('h8)
	) name3925 (
		_w9749_,
		_w9751_,
		_w9752_
	);
	LUT4 #(
		.INIT('h0020)
	) name3926 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9753_
	);
	LUT4 #(
		.INIT('h8000)
	) name3927 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9754_
	);
	LUT3 #(
		.INIT('h02)
	) name3928 (
		_w9741_,
		_w9744_,
		_w9747_,
		_w9755_
	);
	LUT3 #(
		.INIT('h01)
	) name3929 (
		_w9754_,
		_w9755_,
		_w9753_,
		_w9756_
	);
	LUT4 #(
		.INIT('hc693)
	) name3930 (
		decrypt_pad,
		\u2_R7_reg[32]/NET0131 ,
		\u2_uk_K_r7_reg[43]/NET0131 ,
		\u2_uk_K_r7_reg[50]/NET0131 ,
		_w9757_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3931 (
		_w9748_,
		_w9752_,
		_w9756_,
		_w9757_,
		_w9758_
	);
	LUT4 #(
		.INIT('hcf45)
	) name3932 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9759_
	);
	LUT3 #(
		.INIT('h02)
	) name3933 (
		_w9747_,
		_w9753_,
		_w9759_,
		_w9760_
	);
	LUT4 #(
		.INIT('h0001)
	) name3934 (
		_w9741_,
		_w9743_,
		_w9744_,
		_w9747_,
		_w9761_
	);
	LUT4 #(
		.INIT('h4000)
	) name3935 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9762_
	);
	LUT2 #(
		.INIT('h1)
	) name3936 (
		_w9761_,
		_w9762_,
		_w9763_
	);
	LUT3 #(
		.INIT('h8a)
	) name3937 (
		_w9757_,
		_w9760_,
		_w9763_,
		_w9764_
	);
	LUT4 #(
		.INIT('h0400)
	) name3938 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9765_
	);
	LUT4 #(
		.INIT('h0001)
	) name3939 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9766_
	);
	LUT4 #(
		.INIT('h1008)
	) name3940 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9767_
	);
	LUT4 #(
		.INIT('hebf6)
	) name3941 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9768_
	);
	LUT2 #(
		.INIT('h2)
	) name3942 (
		_w9747_,
		_w9768_,
		_w9769_
	);
	LUT2 #(
		.INIT('h2)
	) name3943 (
		_w9741_,
		_w9743_,
		_w9770_
	);
	LUT3 #(
		.INIT('h20)
	) name3944 (
		_w9744_,
		_w9747_,
		_w9757_,
		_w9771_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3945 (
		_w9747_,
		_w9753_,
		_w9770_,
		_w9771_,
		_w9772_
	);
	LUT2 #(
		.INIT('h4)
	) name3946 (
		_w9769_,
		_w9772_,
		_w9773_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name3947 (
		\u2_L7_reg[5]/NET0131 ,
		_w9758_,
		_w9764_,
		_w9773_,
		_w9774_
	);
	LUT4 #(
		.INIT('h0020)
	) name3948 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9775_
	);
	LUT4 #(
		.INIT('hbbdb)
	) name3949 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9776_
	);
	LUT4 #(
		.INIT('h8200)
	) name3950 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9777_
	);
	LUT4 #(
		.INIT('hefe7)
	) name3951 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9778_
	);
	LUT4 #(
		.INIT('h3120)
	) name3952 (
		_w9711_,
		_w9777_,
		_w9778_,
		_w9776_,
		_w9779_
	);
	LUT2 #(
		.INIT('h2)
	) name3953 (
		_w9714_,
		_w9779_,
		_w9780_
	);
	LUT2 #(
		.INIT('h8)
	) name3954 (
		_w9711_,
		_w9709_,
		_w9781_
	);
	LUT4 #(
		.INIT('hdcfe)
	) name3955 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9711_,
		_w9782_
	);
	LUT2 #(
		.INIT('h1)
	) name3956 (
		_w9781_,
		_w9782_,
		_w9783_
	);
	LUT2 #(
		.INIT('h4)
	) name3957 (
		_w9710_,
		_w9711_,
		_w9784_
	);
	LUT3 #(
		.INIT('h8a)
	) name3958 (
		_w9707_,
		_w9710_,
		_w9711_,
		_w9785_
	);
	LUT3 #(
		.INIT('h0e)
	) name3959 (
		_w9706_,
		_w9710_,
		_w9709_,
		_w9786_
	);
	LUT2 #(
		.INIT('h8)
	) name3960 (
		_w9785_,
		_w9786_,
		_w9787_
	);
	LUT3 #(
		.INIT('h3b)
	) name3961 (
		_w9706_,
		_w9707_,
		_w9709_,
		_w9788_
	);
	LUT3 #(
		.INIT('h51)
	) name3962 (
		_w9718_,
		_w9784_,
		_w9788_,
		_w9789_
	);
	LUT4 #(
		.INIT('h5455)
	) name3963 (
		_w9714_,
		_w9783_,
		_w9787_,
		_w9789_,
		_w9790_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name3964 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9791_
	);
	LUT3 #(
		.INIT('hc8)
	) name3965 (
		_w9706_,
		_w9707_,
		_w9709_,
		_w9792_
	);
	LUT4 #(
		.INIT('hfa32)
	) name3966 (
		_w9711_,
		_w9712_,
		_w9791_,
		_w9792_,
		_w9793_
	);
	LUT4 #(
		.INIT('h5655)
	) name3967 (
		\u2_L7_reg[10]/NET0131 ,
		_w9790_,
		_w9780_,
		_w9793_,
		_w9794_
	);
	LUT4 #(
		.INIT('h2006)
	) name3968 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9795_
	);
	LUT4 #(
		.INIT('h134c)
	) name3969 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9796_
	);
	LUT2 #(
		.INIT('h1)
	) name3970 (
		_w9631_,
		_w9796_,
		_w9797_
	);
	LUT3 #(
		.INIT('h47)
	) name3971 (
		_w9621_,
		_w9622_,
		_w9631_,
		_w9798_
	);
	LUT4 #(
		.INIT('h0010)
	) name3972 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9799_
	);
	LUT4 #(
		.INIT('h0301)
	) name3973 (
		_w9625_,
		_w9629_,
		_w9799_,
		_w9798_,
		_w9800_
	);
	LUT3 #(
		.INIT('h10)
	) name3974 (
		_w9797_,
		_w9795_,
		_w9800_,
		_w9801_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name3975 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9802_
	);
	LUT2 #(
		.INIT('h2)
	) name3976 (
		_w9631_,
		_w9802_,
		_w9803_
	);
	LUT3 #(
		.INIT('h04)
	) name3977 (
		_w9627_,
		_w9629_,
		_w9639_,
		_w9804_
	);
	LUT4 #(
		.INIT('h0420)
	) name3978 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w9805_
	);
	LUT3 #(
		.INIT('h0d)
	) name3979 (
		_w9626_,
		_w9631_,
		_w9805_,
		_w9806_
	);
	LUT3 #(
		.INIT('h40)
	) name3980 (
		_w9803_,
		_w9804_,
		_w9806_,
		_w9807_
	);
	LUT3 #(
		.INIT('ha9)
	) name3981 (
		\u2_L7_reg[12]/NET0131 ,
		_w9801_,
		_w9807_,
		_w9808_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name3982 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9809_
	);
	LUT4 #(
		.INIT('h5b4b)
	) name3983 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9810_
	);
	LUT4 #(
		.INIT('h0002)
	) name3984 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9811_
	);
	LUT4 #(
		.INIT('h3302)
	) name3985 (
		_w9747_,
		_w9757_,
		_w9810_,
		_w9811_,
		_w9812_
	);
	LUT3 #(
		.INIT('h73)
	) name3986 (
		_w9741_,
		_w9744_,
		_w9747_,
		_w9813_
	);
	LUT4 #(
		.INIT('h0100)
	) name3987 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9747_,
		_w9814_
	);
	LUT3 #(
		.INIT('h08)
	) name3988 (
		_w9741_,
		_w9743_,
		_w9744_,
		_w9815_
	);
	LUT4 #(
		.INIT('h1000)
	) name3989 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9816_
	);
	LUT4 #(
		.INIT('hef5f)
	) name3990 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9817_
	);
	LUT4 #(
		.INIT('h3100)
	) name3991 (
		_w9750_,
		_w9814_,
		_w9813_,
		_w9817_,
		_w9818_
	);
	LUT2 #(
		.INIT('h2)
	) name3992 (
		_w9757_,
		_w9818_,
		_w9819_
	);
	LUT4 #(
		.INIT('h0040)
	) name3993 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9820_
	);
	LUT4 #(
		.INIT('h2022)
	) name3994 (
		_w9741_,
		_w9743_,
		_w9744_,
		_w9757_,
		_w9821_
	);
	LUT4 #(
		.INIT('h0001)
	) name3995 (
		_w9747_,
		_w9816_,
		_w9820_,
		_w9821_,
		_w9822_
	);
	LUT4 #(
		.INIT('h0004)
	) name3996 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9823_
	);
	LUT3 #(
		.INIT('h02)
	) name3997 (
		_w9747_,
		_w9762_,
		_w9823_,
		_w9824_
	);
	LUT3 #(
		.INIT('h0b)
	) name3998 (
		_w9766_,
		_w9822_,
		_w9824_,
		_w9825_
	);
	LUT4 #(
		.INIT('h5556)
	) name3999 (
		\u2_L7_reg[15]/NET0131 ,
		_w9812_,
		_w9819_,
		_w9825_,
		_w9826_
	);
	LUT4 #(
		.INIT('h0200)
	) name4000 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9827_
	);
	LUT4 #(
		.INIT('ha9ab)
	) name4001 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9828_
	);
	LUT2 #(
		.INIT('h2)
	) name4002 (
		_w9649_,
		_w9828_,
		_w9829_
	);
	LUT4 #(
		.INIT('h0008)
	) name4003 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9830_
	);
	LUT4 #(
		.INIT('h0a01)
	) name4004 (
		_w9653_,
		_w9650_,
		_w9649_,
		_w9652_,
		_w9831_
	);
	LUT3 #(
		.INIT('h80)
	) name4005 (
		_w9650_,
		_w9652_,
		_w9651_,
		_w9832_
	);
	LUT4 #(
		.INIT('h0002)
	) name4006 (
		_w9648_,
		_w9830_,
		_w9831_,
		_w9832_,
		_w9833_
	);
	LUT4 #(
		.INIT('hddea)
	) name4007 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9834_
	);
	LUT2 #(
		.INIT('h1)
	) name4008 (
		_w9649_,
		_w9834_,
		_w9835_
	);
	LUT3 #(
		.INIT('h31)
	) name4009 (
		_w9650_,
		_w9649_,
		_w9651_,
		_w9836_
	);
	LUT4 #(
		.INIT('h88a2)
	) name4010 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w9837_
	);
	LUT4 #(
		.INIT('h1011)
	) name4011 (
		_w9648_,
		_w9668_,
		_w9836_,
		_w9837_,
		_w9838_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4012 (
		_w9829_,
		_w9833_,
		_w9835_,
		_w9838_,
		_w9839_
	);
	LUT2 #(
		.INIT('h8)
	) name4013 (
		_w9650_,
		_w9649_,
		_w9840_
	);
	LUT2 #(
		.INIT('h4)
	) name4014 (
		_w9654_,
		_w9840_,
		_w9841_
	);
	LUT3 #(
		.INIT('h56)
	) name4015 (
		\u2_L7_reg[17]/NET0131 ,
		_w9839_,
		_w9841_,
		_w9842_
	);
	LUT4 #(
		.INIT('hc693)
	) name4016 (
		decrypt_pad,
		\u2_R7_reg[19]/NET0131 ,
		\u2_uk_K_r7_reg[44]/NET0131 ,
		\u2_uk_K_r7_reg[51]/NET0131 ,
		_w9843_
	);
	LUT4 #(
		.INIT('hc693)
	) name4017 (
		decrypt_pad,
		\u2_R7_reg[18]/NET0131 ,
		\u2_uk_K_r7_reg[2]/NET0131 ,
		\u2_uk_K_r7_reg[9]/NET0131 ,
		_w9844_
	);
	LUT4 #(
		.INIT('hc963)
	) name4018 (
		decrypt_pad,
		\u2_R7_reg[17]/NET0131 ,
		\u2_uk_K_r7_reg[15]/NET0131 ,
		\u2_uk_K_r7_reg[8]/NET0131 ,
		_w9845_
	);
	LUT4 #(
		.INIT('hc693)
	) name4019 (
		decrypt_pad,
		\u2_R7_reg[16]/NET0131 ,
		\u2_uk_K_r7_reg[45]/NET0131 ,
		\u2_uk_K_r7_reg[52]/NET0131 ,
		_w9846_
	);
	LUT4 #(
		.INIT('hc693)
	) name4020 (
		decrypt_pad,
		\u2_R7_reg[21]/NET0131 ,
		\u2_uk_K_r7_reg[29]/NET0131 ,
		\u2_uk_K_r7_reg[36]/NET0131 ,
		_w9847_
	);
	LUT3 #(
		.INIT('h04)
	) name4021 (
		_w9845_,
		_w9846_,
		_w9847_,
		_w9848_
	);
	LUT4 #(
		.INIT('h0010)
	) name4022 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9849_
	);
	LUT4 #(
		.INIT('h4000)
	) name4023 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9850_
	);
	LUT4 #(
		.INIT('hbc67)
	) name4024 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9851_
	);
	LUT4 #(
		.INIT('h5bf8)
	) name4025 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9852_
	);
	LUT4 #(
		.INIT('h2004)
	) name4026 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9853_
	);
	LUT4 #(
		.INIT('h00d8)
	) name4027 (
		_w9843_,
		_w9852_,
		_w9851_,
		_w9853_,
		_w9854_
	);
	LUT4 #(
		.INIT('hc693)
	) name4028 (
		decrypt_pad,
		\u2_R7_reg[20]/NET0131 ,
		\u2_uk_K_r7_reg[28]/NET0131 ,
		\u2_uk_K_r7_reg[35]/NET0131 ,
		_w9855_
	);
	LUT2 #(
		.INIT('h1)
	) name4029 (
		_w9854_,
		_w9855_,
		_w9856_
	);
	LUT4 #(
		.INIT('ha43f)
	) name4030 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9857_
	);
	LUT2 #(
		.INIT('h2)
	) name4031 (
		_w9843_,
		_w9857_,
		_w9858_
	);
	LUT3 #(
		.INIT('hde)
	) name4032 (
		_w9845_,
		_w9846_,
		_w9847_,
		_w9859_
	);
	LUT2 #(
		.INIT('h1)
	) name4033 (
		_w9843_,
		_w9844_,
		_w9860_
	);
	LUT2 #(
		.INIT('h4)
	) name4034 (
		_w9859_,
		_w9860_,
		_w9861_
	);
	LUT2 #(
		.INIT('h9)
	) name4035 (
		_w9844_,
		_w9845_,
		_w9862_
	);
	LUT4 #(
		.INIT('h0060)
	) name4036 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9863_
	);
	LUT4 #(
		.INIT('h7000)
	) name4037 (
		_w9843_,
		_w9844_,
		_w9846_,
		_w9847_,
		_w9864_
	);
	LUT3 #(
		.INIT('h13)
	) name4038 (
		_w9862_,
		_w9863_,
		_w9864_,
		_w9865_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4039 (
		_w9855_,
		_w9858_,
		_w9861_,
		_w9865_,
		_w9866_
	);
	LUT4 #(
		.INIT('h0040)
	) name4040 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9867_
	);
	LUT4 #(
		.INIT('hffbd)
	) name4041 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9868_
	);
	LUT4 #(
		.INIT('h0200)
	) name4042 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9869_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name4043 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9870_
	);
	LUT3 #(
		.INIT('hd8)
	) name4044 (
		_w9843_,
		_w9868_,
		_w9870_,
		_w9871_
	);
	LUT4 #(
		.INIT('h5655)
	) name4045 (
		\u2_L7_reg[14]/NET0131 ,
		_w9856_,
		_w9866_,
		_w9871_,
		_w9872_
	);
	LUT3 #(
		.INIT('hea)
	) name4046 (
		_w9706_,
		_w9710_,
		_w9709_,
		_w9873_
	);
	LUT2 #(
		.INIT('h2)
	) name4047 (
		_w9738_,
		_w9873_,
		_w9874_
	);
	LUT3 #(
		.INIT('hd8)
	) name4048 (
		_w9706_,
		_w9710_,
		_w9709_,
		_w9875_
	);
	LUT4 #(
		.INIT('h1101)
	) name4049 (
		_w9714_,
		_w9733_,
		_w9785_,
		_w9875_,
		_w9876_
	);
	LUT4 #(
		.INIT('hdf0f)
	) name4050 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9877_
	);
	LUT3 #(
		.INIT('h0b)
	) name4051 (
		_w9706_,
		_w9707_,
		_w9711_,
		_w9878_
	);
	LUT2 #(
		.INIT('h4)
	) name4052 (
		_w9877_,
		_w9878_,
		_w9879_
	);
	LUT4 #(
		.INIT('h4000)
	) name4053 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9880_
	);
	LUT3 #(
		.INIT('h02)
	) name4054 (
		_w9714_,
		_w9726_,
		_w9880_,
		_w9881_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4055 (
		_w9874_,
		_w9876_,
		_w9879_,
		_w9881_,
		_w9882_
	);
	LUT3 #(
		.INIT('h01)
	) name4056 (
		_w9711_,
		_w9727_,
		_w9880_,
		_w9883_
	);
	LUT4 #(
		.INIT('hf5f1)
	) name4057 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9884_
	);
	LUT2 #(
		.INIT('h2)
	) name4058 (
		_w9714_,
		_w9884_,
		_w9885_
	);
	LUT3 #(
		.INIT('h02)
	) name4059 (
		_w9711_,
		_w9718_,
		_w9777_,
		_w9886_
	);
	LUT3 #(
		.INIT('h45)
	) name4060 (
		_w9883_,
		_w9885_,
		_w9886_,
		_w9887_
	);
	LUT3 #(
		.INIT('h56)
	) name4061 (
		\u2_L7_reg[1]/NET0131 ,
		_w9882_,
		_w9887_,
		_w9888_
	);
	LUT4 #(
		.INIT('h0010)
	) name4062 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9747_,
		_w9889_
	);
	LUT3 #(
		.INIT('h01)
	) name4063 (
		_w9745_,
		_w9757_,
		_w9889_,
		_w9890_
	);
	LUT3 #(
		.INIT('h8b)
	) name4064 (
		_w9742_,
		_w9743_,
		_w9744_,
		_w9891_
	);
	LUT2 #(
		.INIT('h8)
	) name4065 (
		_w9741_,
		_w9747_,
		_w9892_
	);
	LUT3 #(
		.INIT('h45)
	) name4066 (
		_w9766_,
		_w9891_,
		_w9892_,
		_w9893_
	);
	LUT4 #(
		.INIT('hf7f5)
	) name4067 (
		_w9741_,
		_w9743_,
		_w9744_,
		_w9747_,
		_w9894_
	);
	LUT4 #(
		.INIT('h3f1f)
	) name4068 (
		_w9742_,
		_w9743_,
		_w9744_,
		_w9747_,
		_w9895_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name4069 (
		_w9741_,
		_w9742_,
		_w9894_,
		_w9895_,
		_w9896_
	);
	LUT3 #(
		.INIT('h80)
	) name4070 (
		_w9890_,
		_w9893_,
		_w9896_,
		_w9897_
	);
	LUT4 #(
		.INIT('h2100)
	) name4071 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w9898_
	);
	LUT3 #(
		.INIT('h02)
	) name4072 (
		_w9757_,
		_w9823_,
		_w9898_,
		_w9899_
	);
	LUT3 #(
		.INIT('hb0)
	) name4073 (
		_w9743_,
		_w9744_,
		_w9747_,
		_w9900_
	);
	LUT3 #(
		.INIT('hec)
	) name4074 (
		_w9741_,
		_w9742_,
		_w9744_,
		_w9901_
	);
	LUT3 #(
		.INIT('h40)
	) name4075 (
		_w9815_,
		_w9900_,
		_w9901_,
		_w9902_
	);
	LUT3 #(
		.INIT('hda)
	) name4076 (
		_w9742_,
		_w9743_,
		_w9744_,
		_w9903_
	);
	LUT2 #(
		.INIT('h2)
	) name4077 (
		_w9741_,
		_w9747_,
		_w9904_
	);
	LUT2 #(
		.INIT('h4)
	) name4078 (
		_w9903_,
		_w9904_,
		_w9905_
	);
	LUT3 #(
		.INIT('h10)
	) name4079 (
		_w9902_,
		_w9905_,
		_w9899_,
		_w9906_
	);
	LUT3 #(
		.INIT('h07)
	) name4080 (
		_w9741_,
		_w9742_,
		_w9747_,
		_w9907_
	);
	LUT4 #(
		.INIT('h010d)
	) name4081 (
		_w9741_,
		_w9743_,
		_w9744_,
		_w9747_,
		_w9908_
	);
	LUT2 #(
		.INIT('h4)
	) name4082 (
		_w9907_,
		_w9908_,
		_w9909_
	);
	LUT4 #(
		.INIT('h55a9)
	) name4083 (
		\u2_L7_reg[21]/NET0131 ,
		_w9897_,
		_w9906_,
		_w9909_,
		_w9910_
	);
	LUT4 #(
		.INIT('h3ce4)
	) name4084 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9911_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name4085 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9912_
	);
	LUT4 #(
		.INIT('hbb7f)
	) name4086 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9913_
	);
	LUT4 #(
		.INIT('hd800)
	) name4087 (
		_w9843_,
		_w9911_,
		_w9912_,
		_w9913_,
		_w9914_
	);
	LUT2 #(
		.INIT('h2)
	) name4088 (
		_w9855_,
		_w9914_,
		_w9915_
	);
	LUT4 #(
		.INIT('hfe7d)
	) name4089 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9916_
	);
	LUT2 #(
		.INIT('h2)
	) name4090 (
		_w9843_,
		_w9916_,
		_w9917_
	);
	LUT3 #(
		.INIT('ha2)
	) name4091 (
		_w9843_,
		_w9845_,
		_w9847_,
		_w9918_
	);
	LUT4 #(
		.INIT('h2223)
	) name4092 (
		_w9843_,
		_w9844_,
		_w9845_,
		_w9846_,
		_w9919_
	);
	LUT2 #(
		.INIT('h4)
	) name4093 (
		_w9918_,
		_w9919_,
		_w9920_
	);
	LUT4 #(
		.INIT('h0010)
	) name4094 (
		_w9843_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w9921_
	);
	LUT2 #(
		.INIT('h2)
	) name4095 (
		_w9843_,
		_w9847_,
		_w9922_
	);
	LUT3 #(
		.INIT('h08)
	) name4096 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9923_
	);
	LUT3 #(
		.INIT('h45)
	) name4097 (
		_w9921_,
		_w9922_,
		_w9923_,
		_w9924_
	);
	LUT4 #(
		.INIT('h0400)
	) name4098 (
		_w9843_,
		_w9844_,
		_w9845_,
		_w9846_,
		_w9925_
	);
	LUT2 #(
		.INIT('h1)
	) name4099 (
		_w9850_,
		_w9925_,
		_w9926_
	);
	LUT4 #(
		.INIT('hba00)
	) name4100 (
		_w9855_,
		_w9920_,
		_w9924_,
		_w9926_,
		_w9927_
	);
	LUT4 #(
		.INIT('h5655)
	) name4101 (
		\u2_L7_reg[25]/NET0131 ,
		_w9915_,
		_w9917_,
		_w9927_,
		_w9928_
	);
	LUT4 #(
		.INIT('h008a)
	) name4102 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9711_,
		_w9929_
	);
	LUT4 #(
		.INIT('h0010)
	) name4103 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9930_
	);
	LUT4 #(
		.INIT('h0203)
	) name4104 (
		_w9732_,
		_w9722_,
		_w9930_,
		_w9929_,
		_w9931_
	);
	LUT4 #(
		.INIT('hdddf)
	) name4105 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9711_,
		_w9932_
	);
	LUT4 #(
		.INIT('h7030)
	) name4106 (
		_w9730_,
		_w9709_,
		_w9714_,
		_w9932_,
		_w9933_
	);
	LUT2 #(
		.INIT('h8)
	) name4107 (
		_w9931_,
		_w9933_,
		_w9934_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name4108 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9709_,
		_w9935_
	);
	LUT2 #(
		.INIT('h1)
	) name4109 (
		_w9711_,
		_w9935_,
		_w9936_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4110 (
		_w9707_,
		_w9710_,
		_w9709_,
		_w9714_,
		_w9937_
	);
	LUT2 #(
		.INIT('h4)
	) name4111 (
		_w9731_,
		_w9937_,
		_w9938_
	);
	LUT3 #(
		.INIT('hd0)
	) name4112 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9939_
	);
	LUT3 #(
		.INIT('h13)
	) name4113 (
		_w9781_,
		_w9775_,
		_w9939_,
		_w9940_
	);
	LUT3 #(
		.INIT('h40)
	) name4114 (
		_w9936_,
		_w9938_,
		_w9940_,
		_w9941_
	);
	LUT3 #(
		.INIT('h2b)
	) name4115 (
		_w9706_,
		_w9707_,
		_w9710_,
		_w9942_
	);
	LUT2 #(
		.INIT('h1)
	) name4116 (
		_w9711_,
		_w9709_,
		_w9943_
	);
	LUT3 #(
		.INIT('h10)
	) name4117 (
		_w9730_,
		_w9942_,
		_w9943_,
		_w9944_
	);
	LUT2 #(
		.INIT('h8)
	) name4118 (
		_w9706_,
		_w9711_,
		_w9945_
	);
	LUT2 #(
		.INIT('h8)
	) name4119 (
		_w9725_,
		_w9945_,
		_w9946_
	);
	LUT2 #(
		.INIT('h1)
	) name4120 (
		_w9944_,
		_w9946_,
		_w9947_
	);
	LUT4 #(
		.INIT('ha955)
	) name4121 (
		\u2_L7_reg[26]/NET0131 ,
		_w9934_,
		_w9941_,
		_w9947_,
		_w9948_
	);
	LUT4 #(
		.INIT('hc693)
	) name4122 (
		decrypt_pad,
		\u2_R7_reg[8]/NET0131 ,
		\u2_uk_K_r7_reg[48]/NET0131 ,
		\u2_uk_K_r7_reg[55]/P0001 ,
		_w9949_
	);
	LUT4 #(
		.INIT('hc693)
	) name4123 (
		decrypt_pad,
		\u2_R7_reg[7]/NET0131 ,
		\u2_uk_K_r7_reg[25]/NET0131 ,
		\u2_uk_K_r7_reg[32]/NET0131 ,
		_w9950_
	);
	LUT4 #(
		.INIT('hc963)
	) name4124 (
		decrypt_pad,
		\u2_R7_reg[6]/NET0131 ,
		\u2_uk_K_r7_reg[13]/NET0131 ,
		\u2_uk_K_r7_reg[6]/NET0131 ,
		_w9951_
	);
	LUT4 #(
		.INIT('hc963)
	) name4125 (
		decrypt_pad,
		\u2_R7_reg[4]/NET0131 ,
		\u2_uk_K_r7_reg[11]/NET0131 ,
		\u2_uk_K_r7_reg[4]/NET0131 ,
		_w9952_
	);
	LUT4 #(
		.INIT('hc963)
	) name4126 (
		decrypt_pad,
		\u2_R7_reg[9]/NET0131 ,
		\u2_uk_K_r7_reg[3]/NET0131 ,
		\u2_uk_K_r7_reg[53]/NET0131 ,
		_w9953_
	);
	LUT4 #(
		.INIT('hc693)
	) name4127 (
		decrypt_pad,
		\u2_R7_reg[5]/NET0131 ,
		\u2_uk_K_r7_reg[40]/NET0131 ,
		\u2_uk_K_r7_reg[47]/NET0131 ,
		_w9954_
	);
	LUT4 #(
		.INIT('h5a4f)
	) name4128 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9955_
	);
	LUT4 #(
		.INIT('hf5fc)
	) name4129 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9956_
	);
	LUT4 #(
		.INIT('hbf7b)
	) name4130 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9957_
	);
	LUT4 #(
		.INIT('hd800)
	) name4131 (
		_w9950_,
		_w9956_,
		_w9955_,
		_w9957_,
		_w9958_
	);
	LUT2 #(
		.INIT('h1)
	) name4132 (
		_w9949_,
		_w9958_,
		_w9959_
	);
	LUT4 #(
		.INIT('hfb7b)
	) name4133 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9960_
	);
	LUT2 #(
		.INIT('h1)
	) name4134 (
		_w9960_,
		_w9950_,
		_w9961_
	);
	LUT3 #(
		.INIT('h02)
	) name4135 (
		_w9954_,
		_w9952_,
		_w9953_,
		_w9962_
	);
	LUT4 #(
		.INIT('h5fa7)
	) name4136 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9963_
	);
	LUT2 #(
		.INIT('h2)
	) name4137 (
		_w9950_,
		_w9963_,
		_w9964_
	);
	LUT2 #(
		.INIT('h1)
	) name4138 (
		_w9950_,
		_w9956_,
		_w9965_
	);
	LUT4 #(
		.INIT('h0400)
	) name4139 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9966_
	);
	LUT3 #(
		.INIT('h0b)
	) name4140 (
		_w9954_,
		_w9953_,
		_w9950_,
		_w9967_
	);
	LUT2 #(
		.INIT('h4)
	) name4141 (
		_w9951_,
		_w9952_,
		_w9968_
	);
	LUT3 #(
		.INIT('h45)
	) name4142 (
		_w9966_,
		_w9967_,
		_w9968_,
		_w9969_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4143 (
		_w9949_,
		_w9964_,
		_w9965_,
		_w9969_,
		_w9970_
	);
	LUT4 #(
		.INIT('h5556)
	) name4144 (
		\u2_L7_reg[28]/NET0131 ,
		_w9961_,
		_w9970_,
		_w9959_,
		_w9971_
	);
	LUT4 #(
		.INIT('hcd6f)
	) name4145 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9972_
	);
	LUT2 #(
		.INIT('h1)
	) name4146 (
		_w9678_,
		_w9972_,
		_w9973_
	);
	LUT4 #(
		.INIT('h5fb4)
	) name4147 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9974_
	);
	LUT4 #(
		.INIT('h0400)
	) name4148 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9975_
	);
	LUT4 #(
		.INIT('h0051)
	) name4149 (
		_w9677_,
		_w9678_,
		_w9974_,
		_w9975_,
		_w9976_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name4150 (
		_w9678_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9977_
	);
	LUT4 #(
		.INIT('h8967)
	) name4151 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9978_
	);
	LUT2 #(
		.INIT('h4)
	) name4152 (
		_w9977_,
		_w9978_,
		_w9979_
	);
	LUT4 #(
		.INIT('haf6f)
	) name4153 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9980_
	);
	LUT3 #(
		.INIT('ha2)
	) name4154 (
		_w9677_,
		_w9678_,
		_w9980_,
		_w9981_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4155 (
		_w9973_,
		_w9976_,
		_w9979_,
		_w9981_,
		_w9982_
	);
	LUT4 #(
		.INIT('h2000)
	) name4156 (
		_w9678_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w9983_
	);
	LUT2 #(
		.INIT('h1)
	) name4157 (
		_w9686_,
		_w9983_,
		_w9984_
	);
	LUT3 #(
		.INIT('h9a)
	) name4158 (
		\u2_L7_reg[29]/NET0131 ,
		_w9982_,
		_w9984_,
		_w9985_
	);
	LUT4 #(
		.INIT('h0122)
	) name4159 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9986_
	);
	LUT4 #(
		.INIT('h0800)
	) name4160 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9987_
	);
	LUT4 #(
		.INIT('h0010)
	) name4161 (
		_w9954_,
		_w9951_,
		_w9953_,
		_w9950_,
		_w9988_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name4162 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9989_
	);
	LUT4 #(
		.INIT('h00bf)
	) name4163 (
		_w9954_,
		_w9952_,
		_w9953_,
		_w9950_,
		_w9990_
	);
	LUT4 #(
		.INIT('h1011)
	) name4164 (
		_w9987_,
		_w9988_,
		_w9989_,
		_w9990_,
		_w9991_
	);
	LUT3 #(
		.INIT('h45)
	) name4165 (
		_w9949_,
		_w9986_,
		_w9991_,
		_w9992_
	);
	LUT4 #(
		.INIT('h2010)
	) name4166 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9993_
	);
	LUT4 #(
		.INIT('ha200)
	) name4167 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9950_,
		_w9994_
	);
	LUT3 #(
		.INIT('ha8)
	) name4168 (
		_w9949_,
		_w9993_,
		_w9994_,
		_w9995_
	);
	LUT3 #(
		.INIT('h04)
	) name4169 (
		_w9954_,
		_w9951_,
		_w9953_,
		_w9996_
	);
	LUT4 #(
		.INIT('h0004)
	) name4170 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9997_
	);
	LUT4 #(
		.INIT('h4000)
	) name4171 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w9998_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4172 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9950_,
		_w9999_
	);
	LUT4 #(
		.INIT('h0b00)
	) name4173 (
		_w9949_,
		_w9998_,
		_w9997_,
		_w9999_,
		_w10000_
	);
	LUT4 #(
		.INIT('hbff2)
	) name4174 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10001_
	);
	LUT4 #(
		.INIT('h0900)
	) name4175 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10002_
	);
	LUT4 #(
		.INIT('h0051)
	) name4176 (
		_w9950_,
		_w9949_,
		_w10001_,
		_w10002_,
		_w10003_
	);
	LUT3 #(
		.INIT('h54)
	) name4177 (
		_w9995_,
		_w10000_,
		_w10003_,
		_w10004_
	);
	LUT3 #(
		.INIT('h65)
	) name4178 (
		\u2_L7_reg[2]/NET0131 ,
		_w9992_,
		_w10004_,
		_w10005_
	);
	LUT4 #(
		.INIT('hc010)
	) name4179 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w10006_
	);
	LUT4 #(
		.INIT('h0800)
	) name4180 (
		_w9678_,
		_w9679_,
		_w9681_,
		_w9682_,
		_w10007_
	);
	LUT3 #(
		.INIT('h02)
	) name4181 (
		_w9677_,
		_w10006_,
		_w10007_,
		_w10008_
	);
	LUT4 #(
		.INIT('he65f)
	) name4182 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w10009_
	);
	LUT2 #(
		.INIT('h2)
	) name4183 (
		_w9678_,
		_w10009_,
		_w10010_
	);
	LUT3 #(
		.INIT('h01)
	) name4184 (
		_w9677_,
		_w9686_,
		_w9689_,
		_w10011_
	);
	LUT3 #(
		.INIT('h45)
	) name4185 (
		_w10008_,
		_w10010_,
		_w10011_,
		_w10012_
	);
	LUT4 #(
		.INIT('hfbaf)
	) name4186 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w10013_
	);
	LUT3 #(
		.INIT('h01)
	) name4187 (
		_w9679_,
		_w9681_,
		_w9682_,
		_w10014_
	);
	LUT3 #(
		.INIT('h04)
	) name4188 (
		_w9681_,
		_w9680_,
		_w9682_,
		_w10015_
	);
	LUT4 #(
		.INIT('heece)
	) name4189 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w10016_
	);
	LUT4 #(
		.INIT('h3210)
	) name4190 (
		_w9677_,
		_w10014_,
		_w10013_,
		_w10016_,
		_w10017_
	);
	LUT4 #(
		.INIT('h1551)
	) name4191 (
		_w9678_,
		_w9679_,
		_w9680_,
		_w9682_,
		_w10018_
	);
	LUT3 #(
		.INIT('hbe)
	) name4192 (
		_w9679_,
		_w9680_,
		_w9682_,
		_w10019_
	);
	LUT4 #(
		.INIT('h8a28)
	) name4193 (
		_w9678_,
		_w9679_,
		_w9680_,
		_w9682_,
		_w10020_
	);
	LUT3 #(
		.INIT('h02)
	) name4194 (
		_w9681_,
		_w10020_,
		_w10018_,
		_w10021_
	);
	LUT3 #(
		.INIT('h0e)
	) name4195 (
		_w9678_,
		_w10017_,
		_w10021_,
		_w10022_
	);
	LUT3 #(
		.INIT('h65)
	) name4196 (
		\u2_L7_reg[4]/NET0131 ,
		_w10012_,
		_w10022_,
		_w10023_
	);
	LUT3 #(
		.INIT('h01)
	) name4197 (
		_w9954_,
		_w9951_,
		_w9953_,
		_w10024_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4198 (
		_w9951_,
		_w9952_,
		_w9953_,
		_w9950_,
		_w10025_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4199 (
		_w9996_,
		_w9990_,
		_w10024_,
		_w10025_,
		_w10026_
	);
	LUT4 #(
		.INIT('h0002)
	) name4200 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10027_
	);
	LUT4 #(
		.INIT('h0002)
	) name4201 (
		_w9949_,
		_w9987_,
		_w9988_,
		_w10027_,
		_w10028_
	);
	LUT4 #(
		.INIT('h0600)
	) name4202 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10029_
	);
	LUT4 #(
		.INIT('h0010)
	) name4203 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10030_
	);
	LUT2 #(
		.INIT('h1)
	) name4204 (
		_w9950_,
		_w9949_,
		_w10031_
	);
	LUT4 #(
		.INIT('h0100)
	) name4205 (
		_w9962_,
		_w10030_,
		_w10029_,
		_w10031_,
		_w10032_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name4206 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10033_
	);
	LUT4 #(
		.INIT('hf400)
	) name4207 (
		_w10026_,
		_w10028_,
		_w10032_,
		_w10033_,
		_w10034_
	);
	LUT4 #(
		.INIT('h1321)
	) name4208 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10035_
	);
	LUT4 #(
		.INIT('hc044)
	) name4209 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10036_
	);
	LUT2 #(
		.INIT('h2)
	) name4210 (
		_w9950_,
		_w9949_,
		_w10037_
	);
	LUT3 #(
		.INIT('h10)
	) name4211 (
		_w10035_,
		_w10036_,
		_w10037_,
		_w10038_
	);
	LUT3 #(
		.INIT('h56)
	) name4212 (
		\u2_L7_reg[13]/NET0131 ,
		_w10034_,
		_w10038_,
		_w10039_
	);
	LUT4 #(
		.INIT('h7525)
	) name4213 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w10040_
	);
	LUT4 #(
		.INIT('h8000)
	) name4214 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w10041_
	);
	LUT4 #(
		.INIT('h0e04)
	) name4215 (
		_w9678_,
		_w10019_,
		_w10041_,
		_w10040_,
		_w10042_
	);
	LUT2 #(
		.INIT('h1)
	) name4216 (
		_w9677_,
		_w10042_,
		_w10043_
	);
	LUT4 #(
		.INIT('hdadf)
	) name4217 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w10044_
	);
	LUT3 #(
		.INIT('h31)
	) name4218 (
		_w9678_,
		_w10015_,
		_w10044_,
		_w10045_
	);
	LUT4 #(
		.INIT('hb8bb)
	) name4219 (
		_w9678_,
		_w9679_,
		_w9681_,
		_w9682_,
		_w10046_
	);
	LUT4 #(
		.INIT('h4004)
	) name4220 (
		_w9679_,
		_w9681_,
		_w9680_,
		_w9682_,
		_w10047_
	);
	LUT3 #(
		.INIT('h0e)
	) name4221 (
		_w9680_,
		_w10046_,
		_w10047_,
		_w10048_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name4222 (
		_w9681_,
		_w9680_,
		_w9698_,
		_w9689_,
		_w10049_
	);
	LUT4 #(
		.INIT('hd500)
	) name4223 (
		_w9677_,
		_w10045_,
		_w10048_,
		_w10049_,
		_w10050_
	);
	LUT3 #(
		.INIT('h65)
	) name4224 (
		\u2_L7_reg[19]/NET0131 ,
		_w10043_,
		_w10050_,
		_w10051_
	);
	LUT4 #(
		.INIT('hee9b)
	) name4225 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w10052_
	);
	LUT4 #(
		.INIT('h7ef7)
	) name4226 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w10053_
	);
	LUT4 #(
		.INIT('h0455)
	) name4227 (
		_w9649_,
		_w9648_,
		_w10052_,
		_w10053_,
		_w10054_
	);
	LUT3 #(
		.INIT('hc4)
	) name4228 (
		_w9653_,
		_w9649_,
		_w9652_,
		_w10055_
	);
	LUT2 #(
		.INIT('h8)
	) name4229 (
		_w9663_,
		_w10055_,
		_w10056_
	);
	LUT3 #(
		.INIT('h07)
	) name4230 (
		_w9656_,
		_w9673_,
		_w9827_,
		_w10057_
	);
	LUT3 #(
		.INIT('h8a)
	) name4231 (
		_w9648_,
		_w10056_,
		_w10057_,
		_w10058_
	);
	LUT4 #(
		.INIT('h0a08)
	) name4232 (
		_w9653_,
		_w9650_,
		_w9649_,
		_w9652_,
		_w10059_
	);
	LUT3 #(
		.INIT('h54)
	) name4233 (
		_w9664_,
		_w9673_,
		_w10059_,
		_w10060_
	);
	LUT4 #(
		.INIT('h4000)
	) name4234 (
		_w9653_,
		_w9649_,
		_w9652_,
		_w9651_,
		_w10061_
	);
	LUT3 #(
		.INIT('h7e)
	) name4235 (
		_w9650_,
		_w9652_,
		_w9651_,
		_w10062_
	);
	LUT2 #(
		.INIT('h4)
	) name4236 (
		_w10061_,
		_w10062_,
		_w10063_
	);
	LUT3 #(
		.INIT('hd9)
	) name4237 (
		_w9653_,
		_w9650_,
		_w9651_,
		_w10064_
	);
	LUT2 #(
		.INIT('h2)
	) name4238 (
		_w9671_,
		_w10064_,
		_w10065_
	);
	LUT4 #(
		.INIT('h00ba)
	) name4239 (
		_w9648_,
		_w10060_,
		_w10063_,
		_w10065_,
		_w10066_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name4240 (
		\u2_L7_reg[23]/NET0131 ,
		_w10058_,
		_w10054_,
		_w10066_,
		_w10067_
	);
	LUT4 #(
		.INIT('h9f9a)
	) name4241 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w10068_
	);
	LUT2 #(
		.INIT('h1)
	) name4242 (
		_w9747_,
		_w10068_,
		_w10069_
	);
	LUT3 #(
		.INIT('hd0)
	) name4243 (
		_w9741_,
		_w9742_,
		_w9747_,
		_w10070_
	);
	LUT4 #(
		.INIT('hbdf3)
	) name4244 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w10071_
	);
	LUT3 #(
		.INIT('h70)
	) name4245 (
		_w9809_,
		_w10070_,
		_w10071_,
		_w10072_
	);
	LUT3 #(
		.INIT('h8a)
	) name4246 (
		_w9757_,
		_w10069_,
		_w10072_,
		_w10073_
	);
	LUT3 #(
		.INIT('ha2)
	) name4247 (
		_w9742_,
		_w9743_,
		_w9744_,
		_w10074_
	);
	LUT4 #(
		.INIT('h1030)
	) name4248 (
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_,
		_w10075_
	);
	LUT3 #(
		.INIT('h02)
	) name4249 (
		_w9747_,
		_w10075_,
		_w10074_,
		_w10076_
	);
	LUT4 #(
		.INIT('h0080)
	) name4250 (
		_w9741_,
		_w9742_,
		_w9744_,
		_w9747_,
		_w10077_
	);
	LUT3 #(
		.INIT('h01)
	) name4251 (
		_w9765_,
		_w9889_,
		_w10077_,
		_w10078_
	);
	LUT4 #(
		.INIT('h1000)
	) name4252 (
		_w9742_,
		_w9743_,
		_w9744_,
		_w9747_,
		_w10079_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4253 (
		_w9747_,
		_w9753_,
		_w9767_,
		_w10079_,
		_w10080_
	);
	LUT4 #(
		.INIT('hba00)
	) name4254 (
		_w9757_,
		_w10076_,
		_w10078_,
		_w10080_,
		_w10081_
	);
	LUT3 #(
		.INIT('h65)
	) name4255 (
		\u2_L7_reg[27]/NET0131 ,
		_w10073_,
		_w10081_,
		_w10082_
	);
	LUT3 #(
		.INIT('h40)
	) name4256 (
		_w9622_,
		_w9623_,
		_w9624_,
		_w10083_
	);
	LUT4 #(
		.INIT('hdee3)
	) name4257 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w10084_
	);
	LUT2 #(
		.INIT('h1)
	) name4258 (
		_w9631_,
		_w10084_,
		_w10085_
	);
	LUT3 #(
		.INIT('h08)
	) name4259 (
		_w9621_,
		_w9623_,
		_w9624_,
		_w10086_
	);
	LUT4 #(
		.INIT('hbbfc)
	) name4260 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w10087_
	);
	LUT4 #(
		.INIT('h1f13)
	) name4261 (
		_w9622_,
		_w9631_,
		_w10086_,
		_w10087_,
		_w10088_
	);
	LUT3 #(
		.INIT('h8a)
	) name4262 (
		_w9629_,
		_w10085_,
		_w10088_,
		_w10089_
	);
	LUT3 #(
		.INIT('h04)
	) name4263 (
		_w9621_,
		_w9623_,
		_w9624_,
		_w10090_
	);
	LUT2 #(
		.INIT('h6)
	) name4264 (
		_w9622_,
		_w9624_,
		_w10091_
	);
	LUT4 #(
		.INIT('hab89)
	) name4265 (
		_w9631_,
		_w10090_,
		_w10091_,
		_w10083_,
		_w10092_
	);
	LUT4 #(
		.INIT('h7db7)
	) name4266 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w10093_
	);
	LUT4 #(
		.INIT('h00a2)
	) name4267 (
		_w9622_,
		_w9623_,
		_w9624_,
		_w9631_,
		_w10094_
	);
	LUT4 #(
		.INIT('h0777)
	) name4268 (
		_w9626_,
		_w9631_,
		_w9635_,
		_w10094_,
		_w10095_
	);
	LUT4 #(
		.INIT('hba00)
	) name4269 (
		_w9629_,
		_w10092_,
		_w10093_,
		_w10095_,
		_w10096_
	);
	LUT3 #(
		.INIT('h65)
	) name4270 (
		\u2_L7_reg[32]/NET0131 ,
		_w10089_,
		_w10096_,
		_w10097_
	);
	LUT4 #(
		.INIT('hc693)
	) name4271 (
		decrypt_pad,
		\u2_R7_reg[12]/NET0131 ,
		\u2_uk_K_r7_reg[26]/NET0131 ,
		\u2_uk_K_r7_reg[33]/NET0131 ,
		_w10098_
	);
	LUT4 #(
		.INIT('hc693)
	) name4272 (
		decrypt_pad,
		\u2_R7_reg[11]/NET0131 ,
		\u2_uk_K_r7_reg[11]/NET0131 ,
		\u2_uk_K_r7_reg[18]/NET0131 ,
		_w10099_
	);
	LUT4 #(
		.INIT('hc693)
	) name4273 (
		decrypt_pad,
		\u2_R7_reg[9]/NET0131 ,
		\u2_uk_K_r7_reg[34]/NET0131 ,
		\u2_uk_K_r7_reg[41]/NET0131 ,
		_w10100_
	);
	LUT4 #(
		.INIT('hc693)
	) name4274 (
		decrypt_pad,
		\u2_R7_reg[10]/NET0131 ,
		\u2_uk_K_r7_reg[10]/NET0131 ,
		\u2_uk_K_r7_reg[17]/NET0131 ,
		_w10101_
	);
	LUT4 #(
		.INIT('hc963)
	) name4275 (
		decrypt_pad,
		\u2_R7_reg[8]/NET0131 ,
		\u2_uk_K_r7_reg[12]/NET0131 ,
		\u2_uk_K_r7_reg[5]/NET0131 ,
		_w10102_
	);
	LUT4 #(
		.INIT('hc693)
	) name4276 (
		decrypt_pad,
		\u2_R7_reg[13]/NET0131 ,
		\u2_uk_K_r7_reg[39]/NET0131 ,
		\u2_uk_K_r7_reg[46]/NET0131 ,
		_w10103_
	);
	LUT4 #(
		.INIT('h4000)
	) name4277 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10104_
	);
	LUT2 #(
		.INIT('h4)
	) name4278 (
		_w10099_,
		_w10104_,
		_w10105_
	);
	LUT2 #(
		.INIT('h6)
	) name4279 (
		_w10102_,
		_w10103_,
		_w10106_
	);
	LUT4 #(
		.INIT('h9990)
	) name4280 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10107_
	);
	LUT4 #(
		.INIT('h0990)
	) name4281 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10108_
	);
	LUT2 #(
		.INIT('h4)
	) name4282 (
		_w10102_,
		_w10099_,
		_w10109_
	);
	LUT4 #(
		.INIT('h000b)
	) name4283 (
		_w10102_,
		_w10099_,
		_w10100_,
		_w10101_,
		_w10110_
	);
	LUT2 #(
		.INIT('h2)
	) name4284 (
		_w10099_,
		_w10101_,
		_w10111_
	);
	LUT4 #(
		.INIT('h0040)
	) name4285 (
		_w10102_,
		_w10099_,
		_w10100_,
		_w10101_,
		_w10112_
	);
	LUT4 #(
		.INIT('h2000)
	) name4286 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10113_
	);
	LUT4 #(
		.INIT('h0007)
	) name4287 (
		_w10106_,
		_w10110_,
		_w10112_,
		_w10113_,
		_w10114_
	);
	LUT4 #(
		.INIT('h5455)
	) name4288 (
		_w10098_,
		_w10108_,
		_w10105_,
		_w10114_,
		_w10115_
	);
	LUT2 #(
		.INIT('h8)
	) name4289 (
		_w10098_,
		_w10101_,
		_w10116_
	);
	LUT3 #(
		.INIT('h10)
	) name4290 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10117_
	);
	LUT4 #(
		.INIT('h93d3)
	) name4291 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10118_
	);
	LUT2 #(
		.INIT('h8)
	) name4292 (
		_w10098_,
		_w10099_,
		_w10119_
	);
	LUT4 #(
		.INIT('h7077)
	) name4293 (
		_w10116_,
		_w10117_,
		_w10118_,
		_w10119_,
		_w10120_
	);
	LUT4 #(
		.INIT('h0001)
	) name4294 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10121_
	);
	LUT4 #(
		.INIT('hf3fe)
	) name4295 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10122_
	);
	LUT2 #(
		.INIT('h2)
	) name4296 (
		_w10098_,
		_w10099_,
		_w10123_
	);
	LUT3 #(
		.INIT('h80)
	) name4297 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10124_
	);
	LUT3 #(
		.INIT('h08)
	) name4298 (
		_w10103_,
		_w10100_,
		_w10101_,
		_w10125_
	);
	LUT2 #(
		.INIT('h2)
	) name4299 (
		_w10102_,
		_w10100_,
		_w10126_
	);
	LUT3 #(
		.INIT('h02)
	) name4300 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10127_
	);
	LUT4 #(
		.INIT('h7d3d)
	) name4301 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10128_
	);
	LUT4 #(
		.INIT('hf3d1)
	) name4302 (
		_w10098_,
		_w10099_,
		_w10122_,
		_w10128_,
		_w10129_
	);
	LUT2 #(
		.INIT('h8)
	) name4303 (
		_w10120_,
		_w10129_,
		_w10130_
	);
	LUT3 #(
		.INIT('h65)
	) name4304 (
		\u2_L7_reg[6]/NET0131 ,
		_w10115_,
		_w10130_,
		_w10131_
	);
	LUT3 #(
		.INIT('h28)
	) name4305 (
		_w9622_,
		_w9623_,
		_w9624_,
		_w10132_
	);
	LUT4 #(
		.INIT('h2880)
	) name4306 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w10133_
	);
	LUT4 #(
		.INIT('h5004)
	) name4307 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w10134_
	);
	LUT2 #(
		.INIT('h2)
	) name4308 (
		_w9631_,
		_w10134_,
		_w10135_
	);
	LUT3 #(
		.INIT('h09)
	) name4309 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w10136_
	);
	LUT4 #(
		.INIT('h00f7)
	) name4310 (
		_w9621_,
		_w9623_,
		_w9624_,
		_w9631_,
		_w10137_
	);
	LUT3 #(
		.INIT('h10)
	) name4311 (
		_w10132_,
		_w10136_,
		_w10137_,
		_w10138_
	);
	LUT4 #(
		.INIT('h888a)
	) name4312 (
		_w9629_,
		_w10133_,
		_w10135_,
		_w10138_,
		_w10139_
	);
	LUT4 #(
		.INIT('h5150)
	) name4313 (
		_w9629_,
		_w9631_,
		_w9636_,
		_w10134_,
		_w10140_
	);
	LUT4 #(
		.INIT('h7885)
	) name4314 (
		_w9621_,
		_w9622_,
		_w9623_,
		_w9624_,
		_w10141_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4315 (
		_w9629_,
		_w9631_,
		_w9636_,
		_w10141_,
		_w10142_
	);
	LUT2 #(
		.INIT('h4)
	) name4316 (
		_w9631_,
		_w10133_,
		_w10143_
	);
	LUT3 #(
		.INIT('h01)
	) name4317 (
		_w10142_,
		_w10143_,
		_w10140_,
		_w10144_
	);
	LUT3 #(
		.INIT('h65)
	) name4318 (
		\u2_L7_reg[7]/NET0131 ,
		_w10139_,
		_w10144_,
		_w10145_
	);
	LUT4 #(
		.INIT('h3fef)
	) name4319 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10146_
	);
	LUT4 #(
		.INIT('hc2ff)
	) name4320 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10147_
	);
	LUT4 #(
		.INIT('hfb79)
	) name4321 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10148_
	);
	LUT4 #(
		.INIT('hd800)
	) name4322 (
		_w9843_,
		_w10146_,
		_w10147_,
		_w10148_,
		_w10149_
	);
	LUT4 #(
		.INIT('h0001)
	) name4323 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10150_
	);
	LUT4 #(
		.INIT('hcffe)
	) name4324 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10151_
	);
	LUT3 #(
		.INIT('h10)
	) name4325 (
		_w9843_,
		_w9844_,
		_w9846_,
		_w10152_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4326 (
		_w9843_,
		_w9870_,
		_w10151_,
		_w10152_,
		_w10153_
	);
	LUT4 #(
		.INIT('hf977)
	) name4327 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10154_
	);
	LUT4 #(
		.INIT('hbf15)
	) name4328 (
		_w9843_,
		_w9844_,
		_w9848_,
		_w10154_,
		_w10155_
	);
	LUT4 #(
		.INIT('hd800)
	) name4329 (
		_w9855_,
		_w10153_,
		_w10149_,
		_w10155_,
		_w10156_
	);
	LUT2 #(
		.INIT('h9)
	) name4330 (
		\u2_L7_reg[8]/NET0131 ,
		_w10156_,
		_w10157_
	);
	LUT3 #(
		.INIT('h84)
	) name4331 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10158_
	);
	LUT4 #(
		.INIT('h5ba5)
	) name4332 (
		_w10102_,
		_w10099_,
		_w10103_,
		_w10100_,
		_w10159_
	);
	LUT2 #(
		.INIT('h1)
	) name4333 (
		_w10101_,
		_w10159_,
		_w10160_
	);
	LUT4 #(
		.INIT('h0102)
	) name4334 (
		_w10102_,
		_w10099_,
		_w10103_,
		_w10101_,
		_w10161_
	);
	LUT3 #(
		.INIT('h02)
	) name4335 (
		_w10098_,
		_w10104_,
		_w10161_,
		_w10162_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name4336 (
		_w10102_,
		_w10099_,
		_w10103_,
		_w10100_,
		_w10163_
	);
	LUT3 #(
		.INIT('h70)
	) name4337 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10164_
	);
	LUT4 #(
		.INIT('h844c)
	) name4338 (
		_w10102_,
		_w10099_,
		_w10103_,
		_w10100_,
		_w10165_
	);
	LUT4 #(
		.INIT('h3332)
	) name4339 (
		_w10102_,
		_w10099_,
		_w10103_,
		_w10101_,
		_w10166_
	);
	LUT3 #(
		.INIT('h23)
	) name4340 (
		_w10158_,
		_w10165_,
		_w10166_,
		_w10167_
	);
	LUT2 #(
		.INIT('h1)
	) name4341 (
		_w10098_,
		_w10121_,
		_w10168_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4342 (
		_w10160_,
		_w10162_,
		_w10167_,
		_w10168_,
		_w10169_
	);
	LUT4 #(
		.INIT('hdeff)
	) name4343 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10170_
	);
	LUT4 #(
		.INIT('h0200)
	) name4344 (
		_w10102_,
		_w10099_,
		_w10100_,
		_w10101_,
		_w10171_
	);
	LUT3 #(
		.INIT('h0d)
	) name4345 (
		_w10099_,
		_w10170_,
		_w10171_,
		_w10172_
	);
	LUT3 #(
		.INIT('h65)
	) name4346 (
		\u2_L7_reg[16]/NET0131 ,
		_w10169_,
		_w10172_,
		_w10173_
	);
	LUT4 #(
		.INIT('h0009)
	) name4347 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10174_
	);
	LUT4 #(
		.INIT('h9bd6)
	) name4348 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10175_
	);
	LUT3 #(
		.INIT('h54)
	) name4349 (
		_w10098_,
		_w10099_,
		_w10175_,
		_w10176_
	);
	LUT2 #(
		.INIT('h4)
	) name4350 (
		_w10099_,
		_w10107_,
		_w10177_
	);
	LUT3 #(
		.INIT('h2a)
	) name4351 (
		_w10098_,
		_w10106_,
		_w10110_,
		_w10178_
	);
	LUT3 #(
		.INIT('h0b)
	) name4352 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10179_
	);
	LUT4 #(
		.INIT('hc800)
	) name4353 (
		_w10102_,
		_w10099_,
		_w10103_,
		_w10101_,
		_w10180_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name4354 (
		_w10111_,
		_w10126_,
		_w10179_,
		_w10180_,
		_w10181_
	);
	LUT4 #(
		.INIT('h4555)
	) name4355 (
		_w10176_,
		_w10177_,
		_w10178_,
		_w10181_,
		_w10182_
	);
	LUT4 #(
		.INIT('he4ab)
	) name4356 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10183_
	);
	LUT4 #(
		.INIT('h0200)
	) name4357 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10184_
	);
	LUT4 #(
		.INIT('h5504)
	) name4358 (
		_w10098_,
		_w10099_,
		_w10183_,
		_w10184_,
		_w10185_
	);
	LUT2 #(
		.INIT('h8)
	) name4359 (
		_w10109_,
		_w10125_,
		_w10186_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name4360 (
		_w10099_,
		_w10101_,
		_w10127_,
		_w10124_,
		_w10187_
	);
	LUT3 #(
		.INIT('h10)
	) name4361 (
		_w10185_,
		_w10186_,
		_w10187_,
		_w10188_
	);
	LUT3 #(
		.INIT('h65)
	) name4362 (
		\u2_L7_reg[24]/NET0131 ,
		_w10182_,
		_w10188_,
		_w10189_
	);
	LUT4 #(
		.INIT('h75cf)
	) name4363 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10190_
	);
	LUT2 #(
		.INIT('h2)
	) name4364 (
		_w10099_,
		_w10190_,
		_w10191_
	);
	LUT4 #(
		.INIT('h0400)
	) name4365 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10192_
	);
	LUT3 #(
		.INIT('hb1)
	) name4366 (
		_w10102_,
		_w10100_,
		_w10101_,
		_w10193_
	);
	LUT3 #(
		.INIT('h45)
	) name4367 (
		_w10099_,
		_w10103_,
		_w10100_,
		_w10194_
	);
	LUT4 #(
		.INIT('h0045)
	) name4368 (
		_w10174_,
		_w10193_,
		_w10194_,
		_w10192_,
		_w10195_
	);
	LUT3 #(
		.INIT('h45)
	) name4369 (
		_w10098_,
		_w10191_,
		_w10195_,
		_w10196_
	);
	LUT4 #(
		.INIT('h0440)
	) name4370 (
		_w10102_,
		_w10099_,
		_w10103_,
		_w10101_,
		_w10197_
	);
	LUT4 #(
		.INIT('haa80)
	) name4371 (
		_w10098_,
		_w10111_,
		_w10127_,
		_w10197_,
		_w10198_
	);
	LUT4 #(
		.INIT('hba00)
	) name4372 (
		_w10099_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10199_
	);
	LUT2 #(
		.INIT('h4)
	) name4373 (
		_w10163_,
		_w10199_,
		_w10200_
	);
	LUT4 #(
		.INIT('h45ef)
	) name4374 (
		_w10102_,
		_w10103_,
		_w10100_,
		_w10101_,
		_w10201_
	);
	LUT4 #(
		.INIT('h5f13)
	) name4375 (
		_w10116_,
		_w10123_,
		_w10164_,
		_w10201_,
		_w10202_
	);
	LUT3 #(
		.INIT('h10)
	) name4376 (
		_w10198_,
		_w10200_,
		_w10202_,
		_w10203_
	);
	LUT3 #(
		.INIT('h9a)
	) name4377 (
		\u2_L7_reg[30]/NET0131 ,
		_w10196_,
		_w10203_,
		_w10204_
	);
	LUT4 #(
		.INIT('hfa3f)
	) name4378 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10205_
	);
	LUT2 #(
		.INIT('h2)
	) name4379 (
		_w9843_,
		_w10205_,
		_w10206_
	);
	LUT3 #(
		.INIT('ha2)
	) name4380 (
		_w9843_,
		_w9844_,
		_w9845_,
		_w10207_
	);
	LUT4 #(
		.INIT('h45f0)
	) name4381 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10208_
	);
	LUT3 #(
		.INIT('h54)
	) name4382 (
		_w9855_,
		_w10207_,
		_w10208_,
		_w10209_
	);
	LUT3 #(
		.INIT('h8c)
	) name4383 (
		_w9844_,
		_w9846_,
		_w9847_,
		_w10210_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4384 (
		_w9843_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10211_
	);
	LUT2 #(
		.INIT('h4)
	) name4385 (
		_w10210_,
		_w10211_,
		_w10212_
	);
	LUT4 #(
		.INIT('h0400)
	) name4386 (
		_w9843_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10213_
	);
	LUT4 #(
		.INIT('h0020)
	) name4387 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10214_
	);
	LUT4 #(
		.INIT('h0004)
	) name4388 (
		_w9850_,
		_w9855_,
		_w10214_,
		_w10213_,
		_w10215_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4389 (
		_w10206_,
		_w10209_,
		_w10212_,
		_w10215_,
		_w10216_
	);
	LUT4 #(
		.INIT('h2000)
	) name4390 (
		_w9844_,
		_w9845_,
		_w9846_,
		_w9847_,
		_w10217_
	);
	LUT4 #(
		.INIT('h0001)
	) name4391 (
		_w9843_,
		_w9867_,
		_w10150_,
		_w10217_,
		_w10218_
	);
	LUT3 #(
		.INIT('h02)
	) name4392 (
		_w9843_,
		_w9849_,
		_w9869_,
		_w10219_
	);
	LUT2 #(
		.INIT('h1)
	) name4393 (
		_w10218_,
		_w10219_,
		_w10220_
	);
	LUT3 #(
		.INIT('h56)
	) name4394 (
		\u2_L7_reg[3]/NET0131 ,
		_w10216_,
		_w10220_,
		_w10221_
	);
	LUT3 #(
		.INIT('h08)
	) name4395 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w10222_
	);
	LUT4 #(
		.INIT('h0800)
	) name4396 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w10223_
	);
	LUT4 #(
		.INIT('h2010)
	) name4397 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w10224_
	);
	LUT3 #(
		.INIT('h01)
	) name4398 (
		_w9648_,
		_w10224_,
		_w10223_,
		_w10225_
	);
	LUT3 #(
		.INIT('h43)
	) name4399 (
		_w9653_,
		_w9650_,
		_w9651_,
		_w10226_
	);
	LUT4 #(
		.INIT('h0403)
	) name4400 (
		_w9653_,
		_w9650_,
		_w9649_,
		_w9651_,
		_w10227_
	);
	LUT3 #(
		.INIT('h48)
	) name4401 (
		_w9650_,
		_w9649_,
		_w9651_,
		_w10228_
	);
	LUT3 #(
		.INIT('h45)
	) name4402 (
		_w10227_,
		_w10222_,
		_w10228_,
		_w10229_
	);
	LUT4 #(
		.INIT('h9060)
	) name4403 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w10230_
	);
	LUT4 #(
		.INIT('h040c)
	) name4404 (
		_w9671_,
		_w9648_,
		_w9830_,
		_w10226_,
		_w10231_
	);
	LUT4 #(
		.INIT('h7077)
	) name4405 (
		_w10225_,
		_w10229_,
		_w10230_,
		_w10231_,
		_w10232_
	);
	LUT3 #(
		.INIT('h13)
	) name4406 (
		_w9653_,
		_w9649_,
		_w9652_,
		_w10233_
	);
	LUT4 #(
		.INIT('hc800)
	) name4407 (
		_w9653_,
		_w9650_,
		_w9652_,
		_w9651_,
		_w10234_
	);
	LUT2 #(
		.INIT('h8)
	) name4408 (
		_w10233_,
		_w10234_,
		_w10235_
	);
	LUT3 #(
		.INIT('h56)
	) name4409 (
		\u2_L7_reg[9]/NET0131 ,
		_w10232_,
		_w10235_,
		_w10236_
	);
	LUT4 #(
		.INIT('h1a00)
	) name4410 (
		_w9954_,
		_w9952_,
		_w9953_,
		_w9950_,
		_w10237_
	);
	LUT4 #(
		.INIT('hcfaf)
	) name4411 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10238_
	);
	LUT4 #(
		.INIT('h0032)
	) name4412 (
		_w9950_,
		_w9997_,
		_w10238_,
		_w10237_,
		_w10239_
	);
	LUT4 #(
		.INIT('hbf6e)
	) name4413 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10240_
	);
	LUT4 #(
		.INIT('h8000)
	) name4414 (
		_w9954_,
		_w9952_,
		_w9953_,
		_w9950_,
		_w10241_
	);
	LUT4 #(
		.INIT('h0109)
	) name4415 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9950_,
		_w10242_
	);
	LUT3 #(
		.INIT('h10)
	) name4416 (
		_w10241_,
		_w10242_,
		_w10240_,
		_w10243_
	);
	LUT4 #(
		.INIT('h0020)
	) name4417 (
		_w9954_,
		_w9952_,
		_w9953_,
		_w9950_,
		_w10244_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name4418 (
		_w9954_,
		_w9951_,
		_w9952_,
		_w9953_,
		_w10245_
	);
	LUT3 #(
		.INIT('h31)
	) name4419 (
		_w9950_,
		_w10244_,
		_w10245_,
		_w10246_
	);
	LUT4 #(
		.INIT('hd800)
	) name4420 (
		_w9949_,
		_w10239_,
		_w10243_,
		_w10246_,
		_w10247_
	);
	LUT2 #(
		.INIT('h9)
	) name4421 (
		\u2_L7_reg[18]/P0001 ,
		_w10247_,
		_w10248_
	);
	LUT4 #(
		.INIT('hc963)
	) name4422 (
		decrypt_pad,
		\u2_R6_reg[4]/NET0131 ,
		\u2_uk_K_r6_reg[47]/NET0131 ,
		\u2_uk_K_r6_reg[54]/NET0131 ,
		_w10249_
	);
	LUT4 #(
		.INIT('hc963)
	) name4423 (
		decrypt_pad,
		\u2_R6_reg[3]/NET0131 ,
		\u2_uk_K_r6_reg[12]/NET0131 ,
		\u2_uk_K_r6_reg[19]/NET0131 ,
		_w10250_
	);
	LUT4 #(
		.INIT('hc693)
	) name4424 (
		decrypt_pad,
		\u2_R6_reg[2]/NET0131 ,
		\u2_uk_K_r6_reg[10]/NET0131 ,
		\u2_uk_K_r6_reg[3]/NET0131 ,
		_w10251_
	);
	LUT4 #(
		.INIT('hc963)
	) name4425 (
		decrypt_pad,
		\u2_R6_reg[5]/NET0131 ,
		\u2_uk_K_r6_reg[18]/NET0131 ,
		\u2_uk_K_r6_reg[25]/NET0131 ,
		_w10252_
	);
	LUT4 #(
		.INIT('hc963)
	) name4426 (
		decrypt_pad,
		\u2_R6_reg[1]/NET0131 ,
		\u2_uk_K_r6_reg[20]/NET0131 ,
		\u2_uk_K_r6_reg[27]/NET0131 ,
		_w10253_
	);
	LUT4 #(
		.INIT('hc963)
	) name4427 (
		decrypt_pad,
		\u2_R6_reg[32]/NET0131 ,
		\u2_uk_K_r6_reg[24]/NET0131 ,
		\u2_uk_K_r6_reg[6]/NET0131 ,
		_w10254_
	);
	LUT4 #(
		.INIT('hfdba)
	) name4428 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10255_
	);
	LUT2 #(
		.INIT('h1)
	) name4429 (
		_w10250_,
		_w10255_,
		_w10256_
	);
	LUT4 #(
		.INIT('h0800)
	) name4430 (
		_w10251_,
		_w10252_,
		_w10254_,
		_w10250_,
		_w10257_
	);
	LUT4 #(
		.INIT('hf6fe)
	) name4431 (
		_w10251_,
		_w10252_,
		_w10254_,
		_w10250_,
		_w10258_
	);
	LUT2 #(
		.INIT('h2)
	) name4432 (
		_w10253_,
		_w10258_,
		_w10259_
	);
	LUT4 #(
		.INIT('h0800)
	) name4433 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10260_
	);
	LUT2 #(
		.INIT('h8)
	) name4434 (
		_w10252_,
		_w10254_,
		_w10261_
	);
	LUT2 #(
		.INIT('h4)
	) name4435 (
		_w10251_,
		_w10250_,
		_w10262_
	);
	LUT3 #(
		.INIT('hae)
	) name4436 (
		_w10251_,
		_w10253_,
		_w10250_,
		_w10263_
	);
	LUT4 #(
		.INIT('h7707)
	) name4437 (
		_w10260_,
		_w10250_,
		_w10261_,
		_w10263_,
		_w10264_
	);
	LUT4 #(
		.INIT('h5455)
	) name4438 (
		_w10249_,
		_w10256_,
		_w10259_,
		_w10264_,
		_w10265_
	);
	LUT4 #(
		.INIT('h0132)
	) name4439 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10266_
	);
	LUT3 #(
		.INIT('h02)
	) name4440 (
		_w10251_,
		_w10252_,
		_w10254_,
		_w10267_
	);
	LUT4 #(
		.INIT('hcfc5)
	) name4441 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10268_
	);
	LUT4 #(
		.INIT('h0400)
	) name4442 (
		_w10251_,
		_w10252_,
		_w10254_,
		_w10250_,
		_w10269_
	);
	LUT3 #(
		.INIT('h08)
	) name4443 (
		_w10253_,
		_w10254_,
		_w10250_,
		_w10270_
	);
	LUT4 #(
		.INIT('h0031)
	) name4444 (
		_w10250_,
		_w10269_,
		_w10268_,
		_w10270_,
		_w10271_
	);
	LUT2 #(
		.INIT('h4)
	) name4445 (
		_w10253_,
		_w10250_,
		_w10272_
	);
	LUT3 #(
		.INIT('had)
	) name4446 (
		_w10251_,
		_w10252_,
		_w10254_,
		_w10273_
	);
	LUT4 #(
		.INIT('h7bdb)
	) name4447 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10274_
	);
	LUT4 #(
		.INIT('hfbc8)
	) name4448 (
		_w10253_,
		_w10250_,
		_w10273_,
		_w10274_,
		_w10275_
	);
	LUT4 #(
		.INIT('h7500)
	) name4449 (
		_w10249_,
		_w10266_,
		_w10271_,
		_w10275_,
		_w10276_
	);
	LUT3 #(
		.INIT('h65)
	) name4450 (
		\u2_L6_reg[31]/NET0131 ,
		_w10265_,
		_w10276_,
		_w10277_
	);
	LUT4 #(
		.INIT('hc963)
	) name4451 (
		decrypt_pad,
		\u2_R6_reg[23]/NET0131 ,
		\u2_uk_K_r6_reg[14]/NET0131 ,
		\u2_uk_K_r6_reg[21]/NET0131 ,
		_w10278_
	);
	LUT4 #(
		.INIT('hc963)
	) name4452 (
		decrypt_pad,
		\u2_R6_reg[22]/NET0131 ,
		\u2_uk_K_r6_reg[1]/NET0131 ,
		\u2_uk_K_r6_reg[8]/NET0131 ,
		_w10279_
	);
	LUT4 #(
		.INIT('hc693)
	) name4453 (
		decrypt_pad,
		\u2_R6_reg[20]/NET0131 ,
		\u2_uk_K_r6_reg[2]/NET0131 ,
		\u2_uk_K_r6_reg[50]/NET0131 ,
		_w10280_
	);
	LUT4 #(
		.INIT('hc963)
	) name4454 (
		decrypt_pad,
		\u2_R6_reg[25]/NET0131 ,
		\u2_uk_K_r6_reg[35]/NET0131 ,
		\u2_uk_K_r6_reg[42]/NET0131 ,
		_w10281_
	);
	LUT4 #(
		.INIT('hc963)
	) name4455 (
		decrypt_pad,
		\u2_R6_reg[21]/NET0131 ,
		\u2_uk_K_r6_reg[38]/NET0131 ,
		\u2_uk_K_r6_reg[45]/NET0131 ,
		_w10282_
	);
	LUT3 #(
		.INIT('h20)
	) name4456 (
		_w10280_,
		_w10282_,
		_w10281_,
		_w10283_
	);
	LUT4 #(
		.INIT('h168a)
	) name4457 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10284_
	);
	LUT2 #(
		.INIT('h1)
	) name4458 (
		_w10278_,
		_w10284_,
		_w10285_
	);
	LUT4 #(
		.INIT('hc963)
	) name4459 (
		decrypt_pad,
		\u2_R6_reg[24]/NET0131 ,
		\u2_uk_K_r6_reg[16]/NET0131 ,
		\u2_uk_K_r6_reg[23]/P0001 ,
		_w10286_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4460 (
		_w10278_,
		_w10279_,
		_w10280_,
		_w10282_,
		_w10287_
	);
	LUT4 #(
		.INIT('h0004)
	) name4461 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10288_
	);
	LUT4 #(
		.INIT('h3ffb)
	) name4462 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10289_
	);
	LUT3 #(
		.INIT('h2a)
	) name4463 (
		_w10286_,
		_w10287_,
		_w10289_,
		_w10290_
	);
	LUT2 #(
		.INIT('h4)
	) name4464 (
		_w10285_,
		_w10290_,
		_w10291_
	);
	LUT4 #(
		.INIT('h0040)
	) name4465 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10292_
	);
	LUT4 #(
		.INIT('h0800)
	) name4466 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10293_
	);
	LUT4 #(
		.INIT('h0200)
	) name4467 (
		_w10278_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10294_
	);
	LUT3 #(
		.INIT('h01)
	) name4468 (
		_w10293_,
		_w10294_,
		_w10292_,
		_w10295_
	);
	LUT4 #(
		.INIT('h1400)
	) name4469 (
		_w10278_,
		_w10279_,
		_w10280_,
		_w10282_,
		_w10296_
	);
	LUT2 #(
		.INIT('h8)
	) name4470 (
		_w10278_,
		_w10279_,
		_w10297_
	);
	LUT4 #(
		.INIT('h0080)
	) name4471 (
		_w10278_,
		_w10279_,
		_w10280_,
		_w10282_,
		_w10298_
	);
	LUT4 #(
		.INIT('h0010)
	) name4472 (
		_w10278_,
		_w10279_,
		_w10280_,
		_w10281_,
		_w10299_
	);
	LUT4 #(
		.INIT('hfded)
	) name4473 (
		_w10278_,
		_w10279_,
		_w10280_,
		_w10281_,
		_w10300_
	);
	LUT3 #(
		.INIT('h10)
	) name4474 (
		_w10296_,
		_w10298_,
		_w10300_,
		_w10301_
	);
	LUT3 #(
		.INIT('h15)
	) name4475 (
		_w10286_,
		_w10295_,
		_w10301_,
		_w10302_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name4476 (
		_w10278_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10303_
	);
	LUT2 #(
		.INIT('h1)
	) name4477 (
		_w10279_,
		_w10303_,
		_w10304_
	);
	LUT4 #(
		.INIT('h0010)
	) name4478 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10305_
	);
	LUT4 #(
		.INIT('h77ef)
	) name4479 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10306_
	);
	LUT3 #(
		.INIT('h01)
	) name4480 (
		_w10280_,
		_w10282_,
		_w10281_,
		_w10307_
	);
	LUT4 #(
		.INIT('he4f5)
	) name4481 (
		_w10278_,
		_w10279_,
		_w10306_,
		_w10307_,
		_w10308_
	);
	LUT2 #(
		.INIT('h4)
	) name4482 (
		_w10304_,
		_w10308_,
		_w10309_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name4483 (
		\u2_L6_reg[11]/NET0131 ,
		_w10302_,
		_w10291_,
		_w10309_,
		_w10310_
	);
	LUT4 #(
		.INIT('hc693)
	) name4484 (
		decrypt_pad,
		\u2_R6_reg[24]/NET0131 ,
		\u2_uk_K_r6_reg[14]/NET0131 ,
		\u2_uk_K_r6_reg[7]/NET0131 ,
		_w10311_
	);
	LUT4 #(
		.INIT('hc963)
	) name4485 (
		decrypt_pad,
		\u2_R6_reg[27]/NET0131 ,
		\u2_uk_K_r6_reg[36]/NET0131 ,
		\u2_uk_K_r6_reg[43]/NET0131 ,
		_w10312_
	);
	LUT2 #(
		.INIT('h2)
	) name4486 (
		_w10311_,
		_w10312_,
		_w10313_
	);
	LUT4 #(
		.INIT('hc963)
	) name4487 (
		decrypt_pad,
		\u2_R6_reg[25]/NET0131 ,
		\u2_uk_K_r6_reg[42]/NET0131 ,
		\u2_uk_K_r6_reg[49]/NET0131 ,
		_w10314_
	);
	LUT4 #(
		.INIT('hc963)
	) name4488 (
		decrypt_pad,
		\u2_R6_reg[26]/NET0131 ,
		\u2_uk_K_r6_reg[31]/NET0131 ,
		\u2_uk_K_r6_reg[38]/NET0131 ,
		_w10315_
	);
	LUT4 #(
		.INIT('hc963)
	) name4489 (
		decrypt_pad,
		\u2_R6_reg[29]/NET0131 ,
		\u2_uk_K_r6_reg[15]/NET0131 ,
		\u2_uk_K_r6_reg[22]/NET0131 ,
		_w10316_
	);
	LUT2 #(
		.INIT('h2)
	) name4490 (
		_w10315_,
		_w10316_,
		_w10317_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4491 (
		_w10311_,
		_w10315_,
		_w10316_,
		_w10312_,
		_w10318_
	);
	LUT3 #(
		.INIT('h32)
	) name4492 (
		_w10314_,
		_w10313_,
		_w10318_,
		_w10319_
	);
	LUT4 #(
		.INIT('hc963)
	) name4493 (
		decrypt_pad,
		\u2_R6_reg[28]/NET0131 ,
		\u2_uk_K_r6_reg[23]/P0001 ,
		\u2_uk_K_r6_reg[30]/P0001 ,
		_w10320_
	);
	LUT3 #(
		.INIT('h8b)
	) name4494 (
		_w10314_,
		_w10315_,
		_w10316_,
		_w10321_
	);
	LUT3 #(
		.INIT('h51)
	) name4495 (
		_w10320_,
		_w10313_,
		_w10321_,
		_w10322_
	);
	LUT2 #(
		.INIT('h4)
	) name4496 (
		_w10319_,
		_w10322_,
		_w10323_
	);
	LUT3 #(
		.INIT('h9b)
	) name4497 (
		_w10314_,
		_w10315_,
		_w10316_,
		_w10324_
	);
	LUT2 #(
		.INIT('h8)
	) name4498 (
		_w10311_,
		_w10312_,
		_w10325_
	);
	LUT2 #(
		.INIT('h4)
	) name4499 (
		_w10324_,
		_w10325_,
		_w10326_
	);
	LUT4 #(
		.INIT('h1001)
	) name4500 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10327_
	);
	LUT2 #(
		.INIT('h6)
	) name4501 (
		_w10314_,
		_w10311_,
		_w10328_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4502 (
		_w10314_,
		_w10315_,
		_w10316_,
		_w10312_,
		_w10329_
	);
	LUT3 #(
		.INIT('h15)
	) name4503 (
		_w10327_,
		_w10328_,
		_w10329_,
		_w10330_
	);
	LUT3 #(
		.INIT('h8a)
	) name4504 (
		_w10320_,
		_w10326_,
		_w10330_,
		_w10331_
	);
	LUT4 #(
		.INIT('h2010)
	) name4505 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10332_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name4506 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10333_
	);
	LUT3 #(
		.INIT('h02)
	) name4507 (
		_w10312_,
		_w10333_,
		_w10332_,
		_w10334_
	);
	LUT4 #(
		.INIT('haf23)
	) name4508 (
		_w10320_,
		_w10314_,
		_w10316_,
		_w10312_,
		_w10335_
	);
	LUT2 #(
		.INIT('h9)
	) name4509 (
		_w10311_,
		_w10315_,
		_w10336_
	);
	LUT4 #(
		.INIT('h82c3)
	) name4510 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10312_,
		_w10337_
	);
	LUT2 #(
		.INIT('h4)
	) name4511 (
		_w10335_,
		_w10337_,
		_w10338_
	);
	LUT2 #(
		.INIT('h1)
	) name4512 (
		_w10334_,
		_w10338_,
		_w10339_
	);
	LUT4 #(
		.INIT('h5655)
	) name4513 (
		\u2_L6_reg[22]/NET0131 ,
		_w10331_,
		_w10323_,
		_w10339_,
		_w10340_
	);
	LUT4 #(
		.INIT('hcff8)
	) name4514 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10341_
	);
	LUT3 #(
		.INIT('h6f)
	) name4515 (
		_w10253_,
		_w10252_,
		_w10254_,
		_w10342_
	);
	LUT4 #(
		.INIT('hf7df)
	) name4516 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10343_
	);
	LUT4 #(
		.INIT('he400)
	) name4517 (
		_w10250_,
		_w10341_,
		_w10342_,
		_w10343_,
		_w10344_
	);
	LUT4 #(
		.INIT('hffb7)
	) name4518 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10345_
	);
	LUT2 #(
		.INIT('h2)
	) name4519 (
		_w10250_,
		_w10345_,
		_w10346_
	);
	LUT4 #(
		.INIT('h1000)
	) name4520 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10347_
	);
	LUT4 #(
		.INIT('hef11)
	) name4521 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10348_
	);
	LUT4 #(
		.INIT('h00a1)
	) name4522 (
		_w10251_,
		_w10253_,
		_w10254_,
		_w10250_,
		_w10349_
	);
	LUT4 #(
		.INIT('h0400)
	) name4523 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10350_
	);
	LUT4 #(
		.INIT('h7b7f)
	) name4524 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10351_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4525 (
		_w10250_,
		_w10348_,
		_w10349_,
		_w10351_,
		_w10352_
	);
	LUT4 #(
		.INIT('h3120)
	) name4526 (
		_w10249_,
		_w10346_,
		_w10352_,
		_w10344_,
		_w10353_
	);
	LUT2 #(
		.INIT('h9)
	) name4527 (
		\u2_L6_reg[17]/NET0131 ,
		_w10353_,
		_w10354_
	);
	LUT4 #(
		.INIT('hc963)
	) name4528 (
		decrypt_pad,
		\u2_R6_reg[15]/NET0131 ,
		\u2_uk_K_r6_reg[41]/NET0131 ,
		\u2_uk_K_r6_reg[48]/NET0131 ,
		_w10355_
	);
	LUT4 #(
		.INIT('hc963)
	) name4529 (
		decrypt_pad,
		\u2_R6_reg[14]/NET0131 ,
		\u2_uk_K_r6_reg[33]/NET0131 ,
		\u2_uk_K_r6_reg[40]/NET0131 ,
		_w10356_
	);
	LUT4 #(
		.INIT('hc963)
	) name4530 (
		decrypt_pad,
		\u2_R6_reg[12]/NET0131 ,
		\u2_uk_K_r6_reg[13]/NET0131 ,
		\u2_uk_K_r6_reg[20]/NET0131 ,
		_w10357_
	);
	LUT4 #(
		.INIT('hc963)
	) name4531 (
		decrypt_pad,
		\u2_R6_reg[13]/NET0131 ,
		\u2_uk_K_r6_reg[32]/NET0131 ,
		\u2_uk_K_r6_reg[39]/NET0131 ,
		_w10358_
	);
	LUT4 #(
		.INIT('h0012)
	) name4532 (
		_w10357_,
		_w10355_,
		_w10358_,
		_w10356_,
		_w10359_
	);
	LUT4 #(
		.INIT('hc693)
	) name4533 (
		decrypt_pad,
		\u2_R6_reg[17]/NET0131 ,
		\u2_uk_K_r6_reg[4]/NET0131 ,
		\u2_uk_K_r6_reg[54]/NET0131 ,
		_w10360_
	);
	LUT4 #(
		.INIT('h0020)
	) name4534 (
		_w10360_,
		_w10357_,
		_w10355_,
		_w10358_,
		_w10361_
	);
	LUT2 #(
		.INIT('h8)
	) name4535 (
		_w10357_,
		_w10355_,
		_w10362_
	);
	LUT4 #(
		.INIT('h4000)
	) name4536 (
		_w10360_,
		_w10357_,
		_w10355_,
		_w10358_,
		_w10363_
	);
	LUT4 #(
		.INIT('hc963)
	) name4537 (
		decrypt_pad,
		\u2_R6_reg[16]/NET0131 ,
		\u2_uk_K_r6_reg[17]/NET0131 ,
		\u2_uk_K_r6_reg[24]/NET0131 ,
		_w10364_
	);
	LUT4 #(
		.INIT('h0100)
	) name4538 (
		_w10361_,
		_w10363_,
		_w10359_,
		_w10364_,
		_w10365_
	);
	LUT4 #(
		.INIT('h0020)
	) name4539 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10366_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name4540 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10367_
	);
	LUT3 #(
		.INIT('h10)
	) name4541 (
		_w10357_,
		_w10358_,
		_w10356_,
		_w10368_
	);
	LUT4 #(
		.INIT('h0100)
	) name4542 (
		_w10357_,
		_w10355_,
		_w10358_,
		_w10356_,
		_w10369_
	);
	LUT3 #(
		.INIT('h8c)
	) name4543 (
		_w10360_,
		_w10367_,
		_w10369_,
		_w10370_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name4544 (
		_w10360_,
		_w10357_,
		_w10355_,
		_w10358_,
		_w10371_
	);
	LUT4 #(
		.INIT('h70e0)
	) name4545 (
		_w10360_,
		_w10357_,
		_w10355_,
		_w10358_,
		_w10372_
	);
	LUT3 #(
		.INIT('h40)
	) name4546 (
		_w10360_,
		_w10357_,
		_w10356_,
		_w10373_
	);
	LUT3 #(
		.INIT('h31)
	) name4547 (
		_w10360_,
		_w10355_,
		_w10358_,
		_w10374_
	);
	LUT3 #(
		.INIT('h45)
	) name4548 (
		_w10372_,
		_w10373_,
		_w10374_,
		_w10375_
	);
	LUT2 #(
		.INIT('h8)
	) name4549 (
		_w10355_,
		_w10356_,
		_w10376_
	);
	LUT4 #(
		.INIT('h4000)
	) name4550 (
		_w10357_,
		_w10355_,
		_w10358_,
		_w10356_,
		_w10377_
	);
	LUT4 #(
		.INIT('h0001)
	) name4551 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10378_
	);
	LUT4 #(
		.INIT('h1000)
	) name4552 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10379_
	);
	LUT4 #(
		.INIT('heff7)
	) name4553 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10380_
	);
	LUT4 #(
		.INIT('h0100)
	) name4554 (
		_w10364_,
		_w10378_,
		_w10377_,
		_w10380_,
		_w10381_
	);
	LUT4 #(
		.INIT('h7077)
	) name4555 (
		_w10365_,
		_w10370_,
		_w10375_,
		_w10381_,
		_w10382_
	);
	LUT4 #(
		.INIT('h0400)
	) name4556 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10383_
	);
	LUT4 #(
		.INIT('hffbe)
	) name4557 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10384_
	);
	LUT4 #(
		.INIT('he4ee)
	) name4558 (
		_w10355_,
		_w10366_,
		_w10383_,
		_w10384_,
		_w10385_
	);
	LUT3 #(
		.INIT('h56)
	) name4559 (
		\u2_L6_reg[20]/NET0131 ,
		_w10382_,
		_w10385_,
		_w10386_
	);
	LUT4 #(
		.INIT('h3fd2)
	) name4560 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10387_
	);
	LUT4 #(
		.INIT('hab6f)
	) name4561 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10388_
	);
	LUT4 #(
		.INIT('h0200)
	) name4562 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10389_
	);
	LUT4 #(
		.INIT('h00e4)
	) name4563 (
		_w10278_,
		_w10388_,
		_w10387_,
		_w10389_,
		_w10390_
	);
	LUT2 #(
		.INIT('h1)
	) name4564 (
		_w10286_,
		_w10390_,
		_w10391_
	);
	LUT4 #(
		.INIT('hcf6f)
	) name4565 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10392_
	);
	LUT2 #(
		.INIT('h2)
	) name4566 (
		_w10278_,
		_w10392_,
		_w10393_
	);
	LUT4 #(
		.INIT('h0102)
	) name4567 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10394_
	);
	LUT4 #(
		.INIT('h77dc)
	) name4568 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10395_
	);
	LUT4 #(
		.INIT('h0302)
	) name4569 (
		_w10278_,
		_w10299_,
		_w10293_,
		_w10395_,
		_w10396_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4570 (
		_w10286_,
		_w10393_,
		_w10394_,
		_w10396_,
		_w10397_
	);
	LUT4 #(
		.INIT('h2000)
	) name4571 (
		_w10278_,
		_w10279_,
		_w10282_,
		_w10281_,
		_w10398_
	);
	LUT2 #(
		.INIT('h1)
	) name4572 (
		_w10288_,
		_w10398_,
		_w10399_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name4573 (
		\u2_L6_reg[29]/NET0131 ,
		_w10397_,
		_w10391_,
		_w10399_,
		_w10400_
	);
	LUT4 #(
		.INIT('hc963)
	) name4574 (
		decrypt_pad,
		\u2_R6_reg[8]/NET0131 ,
		\u2_uk_K_r6_reg[48]/NET0131 ,
		\u2_uk_K_r6_reg[55]/P0001 ,
		_w10401_
	);
	LUT4 #(
		.INIT('hc963)
	) name4575 (
		decrypt_pad,
		\u2_R6_reg[5]/NET0131 ,
		\u2_uk_K_r6_reg[40]/NET0131 ,
		\u2_uk_K_r6_reg[47]/NET0131 ,
		_w10402_
	);
	LUT4 #(
		.INIT('hc693)
	) name4576 (
		decrypt_pad,
		\u2_R6_reg[9]/NET0131 ,
		\u2_uk_K_r6_reg[3]/NET0131 ,
		\u2_uk_K_r6_reg[53]/NET0131 ,
		_w10403_
	);
	LUT4 #(
		.INIT('hc693)
	) name4577 (
		decrypt_pad,
		\u2_R6_reg[4]/NET0131 ,
		\u2_uk_K_r6_reg[11]/NET0131 ,
		\u2_uk_K_r6_reg[4]/NET0131 ,
		_w10404_
	);
	LUT3 #(
		.INIT('h04)
	) name4578 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10405_
	);
	LUT3 #(
		.INIT('hd9)
	) name4579 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10406_
	);
	LUT4 #(
		.INIT('hc693)
	) name4580 (
		decrypt_pad,
		\u2_R6_reg[6]/NET0131 ,
		\u2_uk_K_r6_reg[13]/NET0131 ,
		\u2_uk_K_r6_reg[6]/NET0131 ,
		_w10407_
	);
	LUT4 #(
		.INIT('h0026)
	) name4581 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10408_
	);
	LUT4 #(
		.INIT('hc963)
	) name4582 (
		decrypt_pad,
		\u2_R6_reg[7]/NET0131 ,
		\u2_uk_K_r6_reg[25]/NET0131 ,
		\u2_uk_K_r6_reg[32]/NET0131 ,
		_w10409_
	);
	LUT4 #(
		.INIT('h4000)
	) name4583 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10410_
	);
	LUT3 #(
		.INIT('h15)
	) name4584 (
		_w10408_,
		_w10409_,
		_w10410_,
		_w10411_
	);
	LUT2 #(
		.INIT('h8)
	) name4585 (
		_w10404_,
		_w10407_,
		_w10412_
	);
	LUT4 #(
		.INIT('h4bfb)
	) name4586 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10413_
	);
	LUT3 #(
		.INIT('hcd)
	) name4587 (
		_w10402_,
		_w10407_,
		_w10409_,
		_w10414_
	);
	LUT2 #(
		.INIT('h2)
	) name4588 (
		_w10403_,
		_w10404_,
		_w10415_
	);
	LUT4 #(
		.INIT('h084c)
	) name4589 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10416_
	);
	LUT4 #(
		.INIT('h0eee)
	) name4590 (
		_w10409_,
		_w10413_,
		_w10414_,
		_w10416_,
		_w10417_
	);
	LUT3 #(
		.INIT('h15)
	) name4591 (
		_w10401_,
		_w10411_,
		_w10417_,
		_w10418_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name4592 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10419_
	);
	LUT4 #(
		.INIT('h080c)
	) name4593 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10420_
	);
	LUT3 #(
		.INIT('h0d)
	) name4594 (
		_w10402_,
		_w10407_,
		_w10409_,
		_w10421_
	);
	LUT4 #(
		.INIT('hf200)
	) name4595 (
		_w10401_,
		_w10419_,
		_w10420_,
		_w10421_,
		_w10422_
	);
	LUT4 #(
		.INIT('h0080)
	) name4596 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10423_
	);
	LUT4 #(
		.INIT('h0010)
	) name4597 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10424_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4598 (
		_w10402_,
		_w10404_,
		_w10407_,
		_w10409_,
		_w10425_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4599 (
		_w10401_,
		_w10424_,
		_w10425_,
		_w10423_,
		_w10426_
	);
	LUT4 #(
		.INIT('hfc54)
	) name4600 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10427_
	);
	LUT4 #(
		.INIT('hdc00)
	) name4601 (
		_w10402_,
		_w10404_,
		_w10407_,
		_w10409_,
		_w10428_
	);
	LUT2 #(
		.INIT('h4)
	) name4602 (
		_w10427_,
		_w10428_,
		_w10429_
	);
	LUT3 #(
		.INIT('h01)
	) name4603 (
		_w10426_,
		_w10429_,
		_w10422_,
		_w10430_
	);
	LUT3 #(
		.INIT('h65)
	) name4604 (
		\u2_L6_reg[2]/NET0131 ,
		_w10418_,
		_w10430_,
		_w10431_
	);
	LUT4 #(
		.INIT('he63f)
	) name4605 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10432_
	);
	LUT2 #(
		.INIT('h2)
	) name4606 (
		_w10278_,
		_w10432_,
		_w10433_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name4607 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10434_
	);
	LUT4 #(
		.INIT('h1000)
	) name4608 (
		_w10278_,
		_w10279_,
		_w10280_,
		_w10281_,
		_w10435_
	);
	LUT4 #(
		.INIT('h0032)
	) name4609 (
		_w10278_,
		_w10288_,
		_w10434_,
		_w10435_,
		_w10436_
	);
	LUT3 #(
		.INIT('h45)
	) name4610 (
		_w10286_,
		_w10433_,
		_w10436_,
		_w10437_
	);
	LUT4 #(
		.INIT('heeae)
	) name4611 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10438_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		_w10278_,
		_w10438_,
		_w10439_
	);
	LUT3 #(
		.INIT('h80)
	) name4613 (
		_w10279_,
		_w10282_,
		_w10281_,
		_w10440_
	);
	LUT4 #(
		.INIT('h2000)
	) name4614 (
		_w10278_,
		_w10279_,
		_w10280_,
		_w10281_,
		_w10441_
	);
	LUT3 #(
		.INIT('h01)
	) name4615 (
		_w10305_,
		_w10440_,
		_w10441_,
		_w10442_
	);
	LUT3 #(
		.INIT('hb6)
	) name4616 (
		_w10280_,
		_w10282_,
		_w10281_,
		_w10443_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name4617 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10444_
	);
	LUT4 #(
		.INIT('h4445)
	) name4618 (
		_w10278_,
		_w10279_,
		_w10280_,
		_w10281_,
		_w10445_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name4619 (
		_w10297_,
		_w10443_,
		_w10444_,
		_w10445_,
		_w10446_
	);
	LUT4 #(
		.INIT('h7500)
	) name4620 (
		_w10286_,
		_w10439_,
		_w10442_,
		_w10446_,
		_w10447_
	);
	LUT3 #(
		.INIT('h65)
	) name4621 (
		\u2_L6_reg[4]/NET0131 ,
		_w10437_,
		_w10447_,
		_w10448_
	);
	LUT4 #(
		.INIT('hc963)
	) name4622 (
		decrypt_pad,
		\u2_R6_reg[32]/NET0131 ,
		\u2_uk_K_r6_reg[43]/NET0131 ,
		\u2_uk_K_r6_reg[50]/NET0131 ,
		_w10449_
	);
	LUT4 #(
		.INIT('hc963)
	) name4623 (
		decrypt_pad,
		\u2_R6_reg[31]/P0001 ,
		\u2_uk_K_r6_reg[37]/NET0131 ,
		\u2_uk_K_r6_reg[44]/NET0131 ,
		_w10450_
	);
	LUT4 #(
		.INIT('hc693)
	) name4624 (
		decrypt_pad,
		\u2_R6_reg[30]/NET0131 ,
		\u2_uk_K_r6_reg[1]/NET0131 ,
		\u2_uk_K_r6_reg[49]/NET0131 ,
		_w10451_
	);
	LUT4 #(
		.INIT('hc963)
	) name4625 (
		decrypt_pad,
		\u2_R6_reg[28]/NET0131 ,
		\u2_uk_K_r6_reg[21]/NET0131 ,
		\u2_uk_K_r6_reg[28]/NET0131 ,
		_w10452_
	);
	LUT4 #(
		.INIT('hc693)
	) name4626 (
		decrypt_pad,
		\u2_R6_reg[29]/NET0131 ,
		\u2_uk_K_r6_reg[0]/NET0131 ,
		\u2_uk_K_r6_reg[52]/NET0131 ,
		_w10453_
	);
	LUT4 #(
		.INIT('hc693)
	) name4627 (
		decrypt_pad,
		\u2_R6_reg[1]/NET0131 ,
		\u2_uk_K_r6_reg[16]/NET0131 ,
		\u2_uk_K_r6_reg[9]/NET0131 ,
		_w10454_
	);
	LUT4 #(
		.INIT('h23a5)
	) name4628 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10455_
	);
	LUT3 #(
		.INIT('h02)
	) name4629 (
		_w10451_,
		_w10453_,
		_w10454_,
		_w10456_
	);
	LUT4 #(
		.INIT('h0020)
	) name4630 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10457_
	);
	LUT4 #(
		.INIT('hfcdf)
	) name4631 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10458_
	);
	LUT4 #(
		.INIT('h0040)
	) name4632 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10459_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name4633 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10460_
	);
	LUT4 #(
		.INIT('hb800)
	) name4634 (
		_w10458_,
		_w10450_,
		_w10455_,
		_w10460_,
		_w10461_
	);
	LUT2 #(
		.INIT('h1)
	) name4635 (
		_w10449_,
		_w10461_,
		_w10462_
	);
	LUT4 #(
		.INIT('haf23)
	) name4636 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10463_
	);
	LUT4 #(
		.INIT('h0001)
	) name4637 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10464_
	);
	LUT4 #(
		.INIT('h0008)
	) name4638 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10465_
	);
	LUT4 #(
		.INIT('hfff6)
	) name4639 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10466_
	);
	LUT4 #(
		.INIT('hedf6)
	) name4640 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10467_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4641 (
		_w10449_,
		_w10459_,
		_w10463_,
		_w10467_,
		_w10468_
	);
	LUT4 #(
		.INIT('h0800)
	) name4642 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10469_
	);
	LUT4 #(
		.INIT('h0021)
	) name4643 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10450_,
		_w10470_
	);
	LUT3 #(
		.INIT('ha8)
	) name4644 (
		_w10449_,
		_w10469_,
		_w10470_,
		_w10471_
	);
	LUT4 #(
		.INIT('h0b01)
	) name4645 (
		_w10450_,
		_w10459_,
		_w10471_,
		_w10468_,
		_w10472_
	);
	LUT3 #(
		.INIT('h9a)
	) name4646 (
		\u2_L6_reg[5]/NET0131 ,
		_w10462_,
		_w10472_,
		_w10473_
	);
	LUT4 #(
		.INIT('hefe7)
	) name4647 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10474_
	);
	LUT2 #(
		.INIT('h2)
	) name4648 (
		_w10355_,
		_w10474_,
		_w10475_
	);
	LUT4 #(
		.INIT('h7dff)
	) name4649 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10476_
	);
	LUT4 #(
		.INIT('hbb1b)
	) name4650 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10477_
	);
	LUT3 #(
		.INIT('h08)
	) name4651 (
		_w10357_,
		_w10358_,
		_w10356_,
		_w10478_
	);
	LUT4 #(
		.INIT('h3313)
	) name4652 (
		_w10357_,
		_w10355_,
		_w10358_,
		_w10356_,
		_w10479_
	);
	LUT3 #(
		.INIT('h8a)
	) name4653 (
		_w10476_,
		_w10477_,
		_w10479_,
		_w10480_
	);
	LUT3 #(
		.INIT('h8a)
	) name4654 (
		_w10364_,
		_w10475_,
		_w10480_,
		_w10481_
	);
	LUT4 #(
		.INIT('hdfce)
	) name4655 (
		_w10360_,
		_w10357_,
		_w10355_,
		_w10358_,
		_w10482_
	);
	LUT2 #(
		.INIT('h1)
	) name4656 (
		_w10376_,
		_w10482_,
		_w10483_
	);
	LUT3 #(
		.INIT('hce)
	) name4657 (
		_w10360_,
		_w10358_,
		_w10356_,
		_w10484_
	);
	LUT2 #(
		.INIT('h2)
	) name4658 (
		_w10362_,
		_w10484_,
		_w10485_
	);
	LUT4 #(
		.INIT('h0008)
	) name4659 (
		_w10360_,
		_w10357_,
		_w10355_,
		_w10356_,
		_w10486_
	);
	LUT3 #(
		.INIT('h01)
	) name4660 (
		_w10379_,
		_w10478_,
		_w10486_,
		_w10487_
	);
	LUT4 #(
		.INIT('h5455)
	) name4661 (
		_w10364_,
		_w10483_,
		_w10485_,
		_w10487_,
		_w10488_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name4662 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10489_
	);
	LUT2 #(
		.INIT('h1)
	) name4663 (
		_w10355_,
		_w10489_,
		_w10490_
	);
	LUT3 #(
		.INIT('h0b)
	) name4664 (
		_w10356_,
		_w10363_,
		_w10377_,
		_w10491_
	);
	LUT2 #(
		.INIT('h4)
	) name4665 (
		_w10490_,
		_w10491_,
		_w10492_
	);
	LUT4 #(
		.INIT('h5655)
	) name4666 (
		\u2_L6_reg[10]/NET0131 ,
		_w10488_,
		_w10481_,
		_w10492_,
		_w10493_
	);
	LUT2 #(
		.INIT('h4)
	) name4667 (
		_w10311_,
		_w10316_,
		_w10494_
	);
	LUT4 #(
		.INIT('hab00)
	) name4668 (
		_w10311_,
		_w10315_,
		_w10316_,
		_w10312_,
		_w10495_
	);
	LUT2 #(
		.INIT('h4)
	) name4669 (
		_w10328_,
		_w10495_,
		_w10496_
	);
	LUT4 #(
		.INIT('h0660)
	) name4670 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10497_
	);
	LUT4 #(
		.INIT('h1000)
	) name4671 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10498_
	);
	LUT4 #(
		.INIT('h008a)
	) name4672 (
		_w10320_,
		_w10312_,
		_w10498_,
		_w10497_,
		_w10499_
	);
	LUT2 #(
		.INIT('h4)
	) name4673 (
		_w10496_,
		_w10499_,
		_w10500_
	);
	LUT4 #(
		.INIT('h4012)
	) name4674 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10501_
	);
	LUT3 #(
		.INIT('h32)
	) name4675 (
		_w10314_,
		_w10315_,
		_w10316_,
		_w10502_
	);
	LUT3 #(
		.INIT('h2a)
	) name4676 (
		_w10311_,
		_w10315_,
		_w10312_,
		_w10503_
	);
	LUT3 #(
		.INIT('h45)
	) name4677 (
		_w10320_,
		_w10502_,
		_w10503_,
		_w10504_
	);
	LUT3 #(
		.INIT('h27)
	) name4678 (
		_w10314_,
		_w10315_,
		_w10312_,
		_w10505_
	);
	LUT3 #(
		.INIT('h09)
	) name4679 (
		_w10314_,
		_w10316_,
		_w10312_,
		_w10506_
	);
	LUT3 #(
		.INIT('h0d)
	) name4680 (
		_w10494_,
		_w10505_,
		_w10506_,
		_w10507_
	);
	LUT3 #(
		.INIT('h40)
	) name4681 (
		_w10501_,
		_w10504_,
		_w10507_,
		_w10508_
	);
	LUT3 #(
		.INIT('ha9)
	) name4682 (
		\u2_L6_reg[12]/NET0131 ,
		_w10500_,
		_w10508_,
		_w10509_
	);
	LUT4 #(
		.INIT('h2000)
	) name4683 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10510_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name4684 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10511_
	);
	LUT4 #(
		.INIT('h0400)
	) name4685 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10512_
	);
	LUT4 #(
		.INIT('hf9ed)
	) name4686 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10513_
	);
	LUT4 #(
		.INIT('h0313)
	) name4687 (
		_w10401_,
		_w10409_,
		_w10511_,
		_w10513_,
		_w10514_
	);
	LUT3 #(
		.INIT('h8e)
	) name4688 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10515_
	);
	LUT4 #(
		.INIT('h3010)
	) name4689 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10516_
	);
	LUT3 #(
		.INIT('h02)
	) name4690 (
		_w10409_,
		_w10515_,
		_w10516_,
		_w10517_
	);
	LUT3 #(
		.INIT('hd0)
	) name4691 (
		_w10402_,
		_w10403_,
		_w10409_,
		_w10518_
	);
	LUT2 #(
		.INIT('h8)
	) name4692 (
		_w10412_,
		_w10518_,
		_w10519_
	);
	LUT3 #(
		.INIT('h51)
	) name4693 (
		_w10401_,
		_w10415_,
		_w10414_,
		_w10520_
	);
	LUT3 #(
		.INIT('h10)
	) name4694 (
		_w10519_,
		_w10517_,
		_w10520_,
		_w10521_
	);
	LUT4 #(
		.INIT('h0002)
	) name4695 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10522_
	);
	LUT4 #(
		.INIT('h002a)
	) name4696 (
		_w10401_,
		_w10414_,
		_w10416_,
		_w10522_,
		_w10523_
	);
	LUT4 #(
		.INIT('h5140)
	) name4697 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10524_
	);
	LUT3 #(
		.INIT('h01)
	) name4698 (
		_w10402_,
		_w10403_,
		_w10407_,
		_w10525_
	);
	LUT4 #(
		.INIT('hf3ee)
	) name4699 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10526_
	);
	LUT4 #(
		.INIT('h80c4)
	) name4700 (
		_w10409_,
		_w10511_,
		_w10526_,
		_w10524_,
		_w10527_
	);
	LUT2 #(
		.INIT('h8)
	) name4701 (
		_w10523_,
		_w10527_,
		_w10528_
	);
	LUT4 #(
		.INIT('h999a)
	) name4702 (
		\u2_L6_reg[13]/NET0131 ,
		_w10514_,
		_w10521_,
		_w10528_,
		_w10529_
	);
	LUT4 #(
		.INIT('hc963)
	) name4703 (
		decrypt_pad,
		\u2_R6_reg[20]/NET0131 ,
		\u2_uk_K_r6_reg[28]/NET0131 ,
		\u2_uk_K_r6_reg[35]/NET0131 ,
		_w10530_
	);
	LUT4 #(
		.INIT('hc963)
	) name4704 (
		decrypt_pad,
		\u2_R6_reg[19]/NET0131 ,
		\u2_uk_K_r6_reg[44]/NET0131 ,
		\u2_uk_K_r6_reg[51]/NET0131 ,
		_w10531_
	);
	LUT4 #(
		.INIT('hc963)
	) name4705 (
		decrypt_pad,
		\u2_R6_reg[16]/NET0131 ,
		\u2_uk_K_r6_reg[45]/NET0131 ,
		\u2_uk_K_r6_reg[52]/NET0131 ,
		_w10532_
	);
	LUT4 #(
		.INIT('hc693)
	) name4706 (
		decrypt_pad,
		\u2_R6_reg[17]/NET0131 ,
		\u2_uk_K_r6_reg[15]/NET0131 ,
		\u2_uk_K_r6_reg[8]/NET0131 ,
		_w10533_
	);
	LUT4 #(
		.INIT('hc963)
	) name4707 (
		decrypt_pad,
		\u2_R6_reg[21]/NET0131 ,
		\u2_uk_K_r6_reg[29]/NET0131 ,
		\u2_uk_K_r6_reg[36]/NET0131 ,
		_w10534_
	);
	LUT4 #(
		.INIT('hc963)
	) name4708 (
		decrypt_pad,
		\u2_R6_reg[18]/NET0131 ,
		\u2_uk_K_r6_reg[2]/NET0131 ,
		\u2_uk_K_r6_reg[9]/NET0131 ,
		_w10535_
	);
	LUT4 #(
		.INIT('h0080)
	) name4709 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10536_
	);
	LUT4 #(
		.INIT('h0002)
	) name4710 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10537_
	);
	LUT4 #(
		.INIT('hcb79)
	) name4711 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10538_
	);
	LUT4 #(
		.INIT('h76ae)
	) name4712 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10539_
	);
	LUT4 #(
		.INIT('h0810)
	) name4713 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10540_
	);
	LUT4 #(
		.INIT('h00e4)
	) name4714 (
		_w10531_,
		_w10538_,
		_w10539_,
		_w10540_,
		_w10541_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w10530_,
		_w10541_,
		_w10542_
	);
	LUT4 #(
		.INIT('hdf9e)
	) name4716 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10531_,
		_w10543_
	);
	LUT2 #(
		.INIT('h1)
	) name4717 (
		_w10543_,
		_w10535_,
		_w10544_
	);
	LUT2 #(
		.INIT('h8)
	) name4718 (
		_w10532_,
		_w10534_,
		_w10545_
	);
	LUT2 #(
		.INIT('h4)
	) name4719 (
		_w10532_,
		_w10535_,
		_w10546_
	);
	LUT4 #(
		.INIT('h9b53)
	) name4720 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10547_
	);
	LUT2 #(
		.INIT('h2)
	) name4721 (
		_w10531_,
		_w10547_,
		_w10548_
	);
	LUT3 #(
		.INIT('hda)
	) name4722 (
		_w10533_,
		_w10531_,
		_w10535_,
		_w10549_
	);
	LUT4 #(
		.INIT('h0200)
	) name4723 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10550_
	);
	LUT3 #(
		.INIT('h0d)
	) name4724 (
		_w10545_,
		_w10549_,
		_w10550_,
		_w10551_
	);
	LUT4 #(
		.INIT('hef00)
	) name4725 (
		_w10544_,
		_w10548_,
		_w10551_,
		_w10530_,
		_w10552_
	);
	LUT4 #(
		.INIT('h0400)
	) name4726 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10553_
	);
	LUT4 #(
		.INIT('h1400)
	) name4727 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10554_
	);
	LUT4 #(
		.INIT('h0020)
	) name4728 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10555_
	);
	LUT4 #(
		.INIT('hfedf)
	) name4729 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10556_
	);
	LUT3 #(
		.INIT('hb1)
	) name4730 (
		_w10531_,
		_w10554_,
		_w10556_,
		_w10557_
	);
	LUT4 #(
		.INIT('h5655)
	) name4731 (
		\u2_L6_reg[14]/NET0131 ,
		_w10552_,
		_w10542_,
		_w10557_,
		_w10558_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name4732 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10559_
	);
	LUT4 #(
		.INIT('h3c3b)
	) name4733 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10560_
	);
	LUT4 #(
		.INIT('h0010)
	) name4734 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10561_
	);
	LUT4 #(
		.INIT('h5504)
	) name4735 (
		_w10449_,
		_w10450_,
		_w10560_,
		_w10561_,
		_w10562_
	);
	LUT3 #(
		.INIT('h40)
	) name4736 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10563_
	);
	LUT4 #(
		.INIT('h0020)
	) name4737 (
		_w10451_,
		_w10453_,
		_w10454_,
		_w10450_,
		_w10564_
	);
	LUT3 #(
		.INIT('h01)
	) name4738 (
		_w10465_,
		_w10563_,
		_w10564_,
		_w10565_
	);
	LUT4 #(
		.INIT('h0100)
	) name4739 (
		_w10453_,
		_w10452_,
		_w10454_,
		_w10450_,
		_w10566_
	);
	LUT4 #(
		.INIT('h2000)
	) name4740 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10567_
	);
	LUT2 #(
		.INIT('h1)
	) name4741 (
		_w10566_,
		_w10567_,
		_w10568_
	);
	LUT3 #(
		.INIT('h2a)
	) name4742 (
		_w10449_,
		_w10565_,
		_w10568_,
		_w10569_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4743 (
		_w10449_,
		_w10451_,
		_w10453_,
		_w10452_,
		_w10570_
	);
	LUT4 #(
		.INIT('h0400)
	) name4744 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10571_
	);
	LUT4 #(
		.INIT('h0004)
	) name4745 (
		_w10450_,
		_w10466_,
		_w10571_,
		_w10570_,
		_w10572_
	);
	LUT4 #(
		.INIT('h0100)
	) name4746 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10573_
	);
	LUT3 #(
		.INIT('h02)
	) name4747 (
		_w10450_,
		_w10469_,
		_w10573_,
		_w10574_
	);
	LUT2 #(
		.INIT('h1)
	) name4748 (
		_w10572_,
		_w10574_,
		_w10575_
	);
	LUT4 #(
		.INIT('h5556)
	) name4749 (
		\u2_L6_reg[15]/NET0131 ,
		_w10562_,
		_w10569_,
		_w10575_,
		_w10576_
	);
	LUT4 #(
		.INIT('h7343)
	) name4750 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10577_
	);
	LUT2 #(
		.INIT('h2)
	) name4751 (
		_w10278_,
		_w10577_,
		_w10578_
	);
	LUT4 #(
		.INIT('h1001)
	) name4752 (
		_w10278_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10579_
	);
	LUT4 #(
		.INIT('h8000)
	) name4753 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10580_
	);
	LUT3 #(
		.INIT('h01)
	) name4754 (
		_w10286_,
		_w10580_,
		_w10579_,
		_w10581_
	);
	LUT4 #(
		.INIT('h2000)
	) name4755 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10582_
	);
	LUT3 #(
		.INIT('h04)
	) name4756 (
		_w10278_,
		_w10280_,
		_w10282_,
		_w10583_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4757 (
		_w10286_,
		_w10279_,
		_w10282_,
		_w10281_,
		_w10584_
	);
	LUT3 #(
		.INIT('h10)
	) name4758 (
		_w10582_,
		_w10583_,
		_w10584_,
		_w10585_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name4759 (
		_w10279_,
		_w10280_,
		_w10282_,
		_w10281_,
		_w10586_
	);
	LUT3 #(
		.INIT('h31)
	) name4760 (
		_w10278_,
		_w10394_,
		_w10586_,
		_w10587_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name4761 (
		_w10578_,
		_w10581_,
		_w10585_,
		_w10587_,
		_w10588_
	);
	LUT4 #(
		.INIT('hefcc)
	) name4762 (
		_w10278_,
		_w10279_,
		_w10283_,
		_w10303_,
		_w10589_
	);
	LUT3 #(
		.INIT('h65)
	) name4763 (
		\u2_L6_reg[19]/NET0131 ,
		_w10588_,
		_w10589_,
		_w10590_
	);
	LUT4 #(
		.INIT('h084c)
	) name4764 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10591_
	);
	LUT3 #(
		.INIT('h01)
	) name4765 (
		_w10360_,
		_w10357_,
		_w10356_,
		_w10592_
	);
	LUT4 #(
		.INIT('hfad8)
	) name4766 (
		_w10355_,
		_w10383_,
		_w10591_,
		_w10592_,
		_w10593_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name4767 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10594_
	);
	LUT3 #(
		.INIT('h45)
	) name4768 (
		_w10364_,
		_w10593_,
		_w10594_,
		_w10595_
	);
	LUT4 #(
		.INIT('hdf4f)
	) name4769 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10596_
	);
	LUT4 #(
		.INIT('h4000)
	) name4770 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10597_
	);
	LUT4 #(
		.INIT('hbcff)
	) name4771 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10598_
	);
	LUT4 #(
		.INIT('h04cc)
	) name4772 (
		_w10355_,
		_w10364_,
		_w10596_,
		_w10598_,
		_w10599_
	);
	LUT4 #(
		.INIT('h6dff)
	) name4773 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10600_
	);
	LUT2 #(
		.INIT('h2)
	) name4774 (
		_w10355_,
		_w10600_,
		_w10601_
	);
	LUT4 #(
		.INIT('hf5f1)
	) name4775 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10602_
	);
	LUT2 #(
		.INIT('h8)
	) name4776 (
		_w10355_,
		_w10364_,
		_w10603_
	);
	LUT2 #(
		.INIT('h4)
	) name4777 (
		_w10602_,
		_w10603_,
		_w10604_
	);
	LUT4 #(
		.INIT('hccef)
	) name4778 (
		_w10360_,
		_w10355_,
		_w10368_,
		_w10597_,
		_w10605_
	);
	LUT4 #(
		.INIT('h0100)
	) name4779 (
		_w10601_,
		_w10604_,
		_w10599_,
		_w10605_,
		_w10606_
	);
	LUT3 #(
		.INIT('h65)
	) name4780 (
		\u2_L6_reg[1]/NET0131 ,
		_w10595_,
		_w10606_,
		_w10607_
	);
	LUT4 #(
		.INIT('h4050)
	) name4781 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10608_
	);
	LUT3 #(
		.INIT('h01)
	) name4782 (
		_w10450_,
		_w10567_,
		_w10608_,
		_w10609_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4783 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10450_,
		_w10610_
	);
	LUT4 #(
		.INIT('h627f)
	) name4784 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10611_
	);
	LUT2 #(
		.INIT('h8)
	) name4785 (
		_w10610_,
		_w10611_,
		_w10612_
	);
	LUT4 #(
		.INIT('h0082)
	) name4786 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10613_
	);
	LUT3 #(
		.INIT('h02)
	) name4787 (
		_w10449_,
		_w10573_,
		_w10613_,
		_w10614_
	);
	LUT3 #(
		.INIT('he0)
	) name4788 (
		_w10609_,
		_w10612_,
		_w10614_,
		_w10615_
	);
	LUT4 #(
		.INIT('h009f)
	) name4789 (
		_w10451_,
		_w10452_,
		_w10454_,
		_w10450_,
		_w10616_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name4790 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10617_
	);
	LUT3 #(
		.INIT('h13)
	) name4791 (
		_w10610_,
		_w10616_,
		_w10617_,
		_w10618_
	);
	LUT4 #(
		.INIT('h0002)
	) name4792 (
		_w10453_,
		_w10452_,
		_w10454_,
		_w10450_,
		_w10619_
	);
	LUT2 #(
		.INIT('h1)
	) name4793 (
		_w10457_,
		_w10619_,
		_w10620_
	);
	LUT4 #(
		.INIT('h4000)
	) name4794 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10621_
	);
	LUT4 #(
		.INIT('h5515)
	) name4795 (
		_w10449_,
		_w10451_,
		_w10453_,
		_w10452_,
		_w10622_
	);
	LUT3 #(
		.INIT('h04)
	) name4796 (
		_w10464_,
		_w10622_,
		_w10621_,
		_w10623_
	);
	LUT3 #(
		.INIT('h40)
	) name4797 (
		_w10618_,
		_w10620_,
		_w10623_,
		_w10624_
	);
	LUT3 #(
		.INIT('ha9)
	) name4798 (
		\u2_L6_reg[21]/NET0131 ,
		_w10615_,
		_w10624_,
		_w10625_
	);
	LUT4 #(
		.INIT('hfdc3)
	) name4799 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10626_
	);
	LUT4 #(
		.INIT('h7bef)
	) name4800 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10627_
	);
	LUT4 #(
		.INIT('h0233)
	) name4801 (
		_w10249_,
		_w10250_,
		_w10626_,
		_w10627_,
		_w10628_
	);
	LUT4 #(
		.INIT('hf73f)
	) name4802 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10629_
	);
	LUT2 #(
		.INIT('h2)
	) name4803 (
		_w10250_,
		_w10629_,
		_w10630_
	);
	LUT3 #(
		.INIT('h07)
	) name4804 (
		_w10267_,
		_w10272_,
		_w10347_,
		_w10631_
	);
	LUT3 #(
		.INIT('h8a)
	) name4805 (
		_w10249_,
		_w10630_,
		_w10631_,
		_w10632_
	);
	LUT3 #(
		.INIT('had)
	) name4806 (
		_w10253_,
		_w10252_,
		_w10254_,
		_w10633_
	);
	LUT2 #(
		.INIT('h2)
	) name4807 (
		_w10262_,
		_w10633_,
		_w10634_
	);
	LUT4 #(
		.INIT('h0080)
	) name4808 (
		_w10251_,
		_w10252_,
		_w10254_,
		_w10250_,
		_w10635_
	);
	LUT3 #(
		.INIT('h7e)
	) name4809 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10636_
	);
	LUT2 #(
		.INIT('h4)
	) name4810 (
		_w10635_,
		_w10636_,
		_w10637_
	);
	LUT4 #(
		.INIT('h0200)
	) name4811 (
		_w10253_,
		_w10252_,
		_w10254_,
		_w10250_,
		_w10638_
	);
	LUT3 #(
		.INIT('h01)
	) name4812 (
		_w10257_,
		_w10270_,
		_w10638_,
		_w10639_
	);
	LUT4 #(
		.INIT('h3222)
	) name4813 (
		_w10249_,
		_w10634_,
		_w10637_,
		_w10639_,
		_w10640_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name4814 (
		\u2_L6_reg[23]/NET0131 ,
		_w10628_,
		_w10632_,
		_w10640_,
		_w10641_
	);
	LUT3 #(
		.INIT('h80)
	) name4815 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10642_
	);
	LUT4 #(
		.INIT('h6a78)
	) name4816 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10643_
	);
	LUT4 #(
		.INIT('hf7a7)
	) name4817 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10644_
	);
	LUT4 #(
		.INIT('hdf3f)
	) name4818 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10645_
	);
	LUT4 #(
		.INIT('hd800)
	) name4819 (
		_w10531_,
		_w10643_,
		_w10644_,
		_w10645_,
		_w10646_
	);
	LUT2 #(
		.INIT('h2)
	) name4820 (
		_w10530_,
		_w10646_,
		_w10647_
	);
	LUT4 #(
		.INIT('h00f7)
	) name4821 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10531_,
		_w10648_
	);
	LUT3 #(
		.INIT('h04)
	) name4822 (
		_w10534_,
		_w10531_,
		_w10535_,
		_w10649_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name4823 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10650_
	);
	LUT4 #(
		.INIT('h0700)
	) name4824 (
		_w10546_,
		_w10648_,
		_w10649_,
		_w10650_,
		_w10651_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name4825 (
		_w10533_,
		_w10546_,
		_w10530_,
		_w10648_,
		_w10652_
	);
	LUT4 #(
		.INIT('hdefb)
	) name4826 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10653_
	);
	LUT4 #(
		.INIT('h0200)
	) name4827 (
		_w10532_,
		_w10533_,
		_w10531_,
		_w10535_,
		_w10654_
	);
	LUT4 #(
		.INIT('h0031)
	) name4828 (
		_w10531_,
		_w10536_,
		_w10653_,
		_w10654_,
		_w10655_
	);
	LUT3 #(
		.INIT('hb0)
	) name4829 (
		_w10651_,
		_w10652_,
		_w10655_,
		_w10656_
	);
	LUT3 #(
		.INIT('h65)
	) name4830 (
		\u2_L6_reg[25]/NET0131 ,
		_w10647_,
		_w10656_,
		_w10657_
	);
	LUT4 #(
		.INIT('h0002)
	) name4831 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10658_
	);
	LUT4 #(
		.INIT('h070f)
	) name4832 (
		_w10360_,
		_w10357_,
		_w10355_,
		_w10356_,
		_w10659_
	);
	LUT3 #(
		.INIT('h45)
	) name4833 (
		_w10371_,
		_w10658_,
		_w10659_,
		_w10660_
	);
	LUT4 #(
		.INIT('hdddf)
	) name4834 (
		_w10360_,
		_w10357_,
		_w10355_,
		_w10358_,
		_w10661_
	);
	LUT2 #(
		.INIT('h2)
	) name4835 (
		_w10356_,
		_w10661_,
		_w10662_
	);
	LUT4 #(
		.INIT('h0010)
	) name4836 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10663_
	);
	LUT3 #(
		.INIT('h02)
	) name4837 (
		_w10364_,
		_w10597_,
		_w10663_,
		_w10664_
	);
	LUT3 #(
		.INIT('h10)
	) name4838 (
		_w10660_,
		_w10662_,
		_w10664_,
		_w10665_
	);
	LUT3 #(
		.INIT('h01)
	) name4839 (
		_w10360_,
		_w10355_,
		_w10358_,
		_w10666_
	);
	LUT3 #(
		.INIT('h01)
	) name4840 (
		_w10363_,
		_w10364_,
		_w10666_,
		_w10667_
	);
	LUT3 #(
		.INIT('hd0)
	) name4841 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10668_
	);
	LUT4 #(
		.INIT('h0111)
	) name4842 (
		_w10366_,
		_w10369_,
		_w10376_,
		_w10668_,
		_w10669_
	);
	LUT2 #(
		.INIT('h8)
	) name4843 (
		_w10667_,
		_w10669_,
		_w10670_
	);
	LUT3 #(
		.INIT('h02)
	) name4844 (
		_w10357_,
		_w10358_,
		_w10364_,
		_w10671_
	);
	LUT4 #(
		.INIT('h0904)
	) name4845 (
		_w10360_,
		_w10357_,
		_w10355_,
		_w10358_,
		_w10672_
	);
	LUT3 #(
		.INIT('h54)
	) name4846 (
		_w10356_,
		_w10671_,
		_w10672_,
		_w10673_
	);
	LUT4 #(
		.INIT('hffd7)
	) name4847 (
		_w10360_,
		_w10357_,
		_w10358_,
		_w10356_,
		_w10674_
	);
	LUT2 #(
		.INIT('h2)
	) name4848 (
		_w10355_,
		_w10674_,
		_w10675_
	);
	LUT2 #(
		.INIT('h1)
	) name4849 (
		_w10673_,
		_w10675_,
		_w10676_
	);
	LUT4 #(
		.INIT('ha955)
	) name4850 (
		\u2_L6_reg[26]/NET0131 ,
		_w10665_,
		_w10670_,
		_w10676_,
		_w10677_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name4851 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10678_
	);
	LUT2 #(
		.INIT('h8)
	) name4852 (
		_w10409_,
		_w10678_,
		_w10679_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name4853 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10680_
	);
	LUT3 #(
		.INIT('h10)
	) name4854 (
		_w10402_,
		_w10404_,
		_w10407_,
		_w10681_
	);
	LUT4 #(
		.INIT('h0001)
	) name4855 (
		_w10405_,
		_w10409_,
		_w10510_,
		_w10681_,
		_w10682_
	);
	LUT4 #(
		.INIT('h6100)
	) name4856 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10683_
	);
	LUT2 #(
		.INIT('h1)
	) name4857 (
		_w10401_,
		_w10683_,
		_w10684_
	);
	LUT4 #(
		.INIT('hba00)
	) name4858 (
		_w10679_,
		_w10680_,
		_w10682_,
		_w10684_,
		_w10685_
	);
	LUT4 #(
		.INIT('h0010)
	) name4859 (
		_w10409_,
		_w10510_,
		_w10678_,
		_w10681_,
		_w10686_
	);
	LUT4 #(
		.INIT('h8280)
	) name4860 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10687_
	);
	LUT4 #(
		.INIT('hef00)
	) name4861 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10409_,
		_w10688_
	);
	LUT2 #(
		.INIT('h4)
	) name4862 (
		_w10687_,
		_w10688_,
		_w10689_
	);
	LUT3 #(
		.INIT('h0b)
	) name4863 (
		_w10402_,
		_w10403_,
		_w10409_,
		_w10690_
	);
	LUT2 #(
		.INIT('h2)
	) name4864 (
		_w10404_,
		_w10407_,
		_w10691_
	);
	LUT4 #(
		.INIT('h2022)
	) name4865 (
		_w10401_,
		_w10512_,
		_w10690_,
		_w10691_,
		_w10692_
	);
	LUT3 #(
		.INIT('he0)
	) name4866 (
		_w10686_,
		_w10689_,
		_w10692_,
		_w10693_
	);
	LUT3 #(
		.INIT('ha9)
	) name4867 (
		\u2_L6_reg[28]/NET0131 ,
		_w10685_,
		_w10693_,
		_w10694_
	);
	LUT3 #(
		.INIT('h02)
	) name4868 (
		_w10531_,
		_w10537_,
		_w10642_,
		_w10695_
	);
	LUT4 #(
		.INIT('h4044)
	) name4869 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10696_
	);
	LUT2 #(
		.INIT('h2)
	) name4870 (
		_w10648_,
		_w10696_,
		_w10697_
	);
	LUT4 #(
		.INIT('hdeaf)
	) name4871 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10698_
	);
	LUT4 #(
		.INIT('h0155)
	) name4872 (
		_w10530_,
		_w10695_,
		_w10697_,
		_w10698_,
		_w10699_
	);
	LUT4 #(
		.INIT('h0001)
	) name4873 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10700_
	);
	LUT4 #(
		.INIT('hf7f6)
	) name4874 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10701_
	);
	LUT3 #(
		.INIT('h02)
	) name4875 (
		_w10532_,
		_w10531_,
		_w10535_,
		_w10702_
	);
	LUT4 #(
		.INIT('h0031)
	) name4876 (
		_w10531_,
		_w10554_,
		_w10701_,
		_w10702_,
		_w10703_
	);
	LUT4 #(
		.INIT('hcbbf)
	) name4877 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10704_
	);
	LUT4 #(
		.INIT('haf23)
	) name4878 (
		_w10534_,
		_w10531_,
		_w10654_,
		_w10704_,
		_w10705_
	);
	LUT3 #(
		.INIT('hd0)
	) name4879 (
		_w10530_,
		_w10703_,
		_w10705_,
		_w10706_
	);
	LUT3 #(
		.INIT('h65)
	) name4880 (
		\u2_L6_reg[8]/NET0131 ,
		_w10699_,
		_w10706_,
		_w10707_
	);
	LUT4 #(
		.INIT('hf23e)
	) name4881 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10708_
	);
	LUT2 #(
		.INIT('h1)
	) name4882 (
		_w10450_,
		_w10708_,
		_w10709_
	);
	LUT3 #(
		.INIT('hd0)
	) name4883 (
		_w10452_,
		_w10454_,
		_w10450_,
		_w10710_
	);
	LUT4 #(
		.INIT('he6df)
	) name4884 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10711_
	);
	LUT3 #(
		.INIT('h70)
	) name4885 (
		_w10559_,
		_w10710_,
		_w10711_,
		_w10712_
	);
	LUT3 #(
		.INIT('h8a)
	) name4886 (
		_w10449_,
		_w10709_,
		_w10712_,
		_w10713_
	);
	LUT3 #(
		.INIT('h4b)
	) name4887 (
		_w10451_,
		_w10453_,
		_w10454_,
		_w10714_
	);
	LUT4 #(
		.INIT('hc888)
	) name4888 (
		_w10456_,
		_w10450_,
		_w10622_,
		_w10714_,
		_w10715_
	);
	LUT4 #(
		.INIT('h0200)
	) name4889 (
		_w10451_,
		_w10453_,
		_w10452_,
		_w10454_,
		_w10716_
	);
	LUT4 #(
		.INIT('h0080)
	) name4890 (
		_w10451_,
		_w10452_,
		_w10454_,
		_w10450_,
		_w10717_
	);
	LUT4 #(
		.INIT('h5554)
	) name4891 (
		_w10449_,
		_w10619_,
		_w10717_,
		_w10716_,
		_w10718_
	);
	LUT3 #(
		.INIT('hb5)
	) name4892 (
		_w10453_,
		_w10452_,
		_w10454_,
		_w10719_
	);
	LUT3 #(
		.INIT('h06)
	) name4893 (
		_w10451_,
		_w10452_,
		_w10450_,
		_w10720_
	);
	LUT2 #(
		.INIT('h4)
	) name4894 (
		_w10719_,
		_w10720_,
		_w10721_
	);
	LUT3 #(
		.INIT('h01)
	) name4895 (
		_w10715_,
		_w10718_,
		_w10721_,
		_w10722_
	);
	LUT3 #(
		.INIT('h65)
	) name4896 (
		\u2_L6_reg[27]/NET0131 ,
		_w10713_,
		_w10722_,
		_w10723_
	);
	LUT4 #(
		.INIT('hbed9)
	) name4897 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10724_
	);
	LUT2 #(
		.INIT('h1)
	) name4898 (
		_w10312_,
		_w10724_,
		_w10725_
	);
	LUT3 #(
		.INIT('hc8)
	) name4899 (
		_w10314_,
		_w10311_,
		_w10312_,
		_w10726_
	);
	LUT4 #(
		.INIT('hf5ee)
	) name4900 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10727_
	);
	LUT4 #(
		.INIT('h5f13)
	) name4901 (
		_w10317_,
		_w10312_,
		_w10726_,
		_w10727_,
		_w10728_
	);
	LUT3 #(
		.INIT('h8a)
	) name4902 (
		_w10320_,
		_w10725_,
		_w10728_,
		_w10729_
	);
	LUT3 #(
		.INIT('h02)
	) name4903 (
		_w10311_,
		_w10315_,
		_w10316_,
		_w10730_
	);
	LUT2 #(
		.INIT('h2)
	) name4904 (
		_w10506_,
		_w10730_,
		_w10731_
	);
	LUT4 #(
		.INIT('h8020)
	) name4905 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10732_
	);
	LUT3 #(
		.INIT('h53)
	) name4906 (
		_w10314_,
		_w10315_,
		_w10316_,
		_w10733_
	);
	LUT3 #(
		.INIT('h13)
	) name4907 (
		_w10726_,
		_w10732_,
		_w10733_,
		_w10734_
	);
	LUT2 #(
		.INIT('h2)
	) name4908 (
		_w10320_,
		_w10312_,
		_w10735_
	);
	LUT4 #(
		.INIT('h00a2)
	) name4909 (
		_w10314_,
		_w10311_,
		_w10316_,
		_w10312_,
		_w10736_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name4910 (
		_w10336_,
		_w10498_,
		_w10735_,
		_w10736_,
		_w10737_
	);
	LUT4 #(
		.INIT('hba00)
	) name4911 (
		_w10320_,
		_w10731_,
		_w10734_,
		_w10737_,
		_w10738_
	);
	LUT3 #(
		.INIT('h65)
	) name4912 (
		\u2_L6_reg[32]/NET0131 ,
		_w10729_,
		_w10738_,
		_w10739_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4913 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10740_
	);
	LUT4 #(
		.INIT('h22e6)
	) name4914 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10741_
	);
	LUT3 #(
		.INIT('h10)
	) name4915 (
		_w10530_,
		_w10740_,
		_w10741_,
		_w10742_
	);
	LUT4 #(
		.INIT('hbf3f)
	) name4916 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10743_
	);
	LUT3 #(
		.INIT('h40)
	) name4917 (
		_w10550_,
		_w10530_,
		_w10743_,
		_w10744_
	);
	LUT4 #(
		.INIT('h0800)
	) name4918 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10745_
	);
	LUT4 #(
		.INIT('h0001)
	) name4919 (
		_w10531_,
		_w10555_,
		_w10700_,
		_w10745_,
		_w10746_
	);
	LUT3 #(
		.INIT('he0)
	) name4920 (
		_w10742_,
		_w10744_,
		_w10746_,
		_w10747_
	);
	LUT4 #(
		.INIT('h1098)
	) name4921 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10748_
	);
	LUT3 #(
		.INIT('h04)
	) name4922 (
		_w10550_,
		_w10530_,
		_w10748_,
		_w10749_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name4923 (
		_w10532_,
		_w10534_,
		_w10533_,
		_w10535_,
		_w10750_
	);
	LUT3 #(
		.INIT('h10)
	) name4924 (
		_w10530_,
		_w10740_,
		_w10750_,
		_w10751_
	);
	LUT3 #(
		.INIT('h02)
	) name4925 (
		_w10531_,
		_w10537_,
		_w10553_,
		_w10752_
	);
	LUT3 #(
		.INIT('he0)
	) name4926 (
		_w10749_,
		_w10751_,
		_w10752_,
		_w10753_
	);
	LUT3 #(
		.INIT('ha9)
	) name4927 (
		\u2_L6_reg[3]/NET0131 ,
		_w10747_,
		_w10753_,
		_w10754_
	);
	LUT4 #(
		.INIT('hc963)
	) name4928 (
		decrypt_pad,
		\u2_R6_reg[13]/NET0131 ,
		\u2_uk_K_r6_reg[39]/NET0131 ,
		\u2_uk_K_r6_reg[46]/NET0131 ,
		_w10755_
	);
	LUT4 #(
		.INIT('hc963)
	) name4929 (
		decrypt_pad,
		\u2_R6_reg[9]/NET0131 ,
		\u2_uk_K_r6_reg[34]/NET0131 ,
		\u2_uk_K_r6_reg[41]/NET0131 ,
		_w10756_
	);
	LUT4 #(
		.INIT('hc963)
	) name4930 (
		decrypt_pad,
		\u2_R6_reg[11]/NET0131 ,
		\u2_uk_K_r6_reg[11]/NET0131 ,
		\u2_uk_K_r6_reg[18]/NET0131 ,
		_w10757_
	);
	LUT3 #(
		.INIT('h0b)
	) name4931 (
		_w10755_,
		_w10756_,
		_w10757_,
		_w10758_
	);
	LUT4 #(
		.INIT('hc963)
	) name4932 (
		decrypt_pad,
		\u2_R6_reg[10]/NET0131 ,
		\u2_uk_K_r6_reg[10]/NET0131 ,
		\u2_uk_K_r6_reg[17]/NET0131 ,
		_w10759_
	);
	LUT4 #(
		.INIT('hc693)
	) name4933 (
		decrypt_pad,
		\u2_R6_reg[8]/NET0131 ,
		\u2_uk_K_r6_reg[12]/NET0131 ,
		\u2_uk_K_r6_reg[5]/NET0131 ,
		_w10760_
	);
	LUT4 #(
		.INIT('h3b0b)
	) name4934 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10761_
	);
	LUT4 #(
		.INIT('h1000)
	) name4935 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10762_
	);
	LUT4 #(
		.INIT('hc963)
	) name4936 (
		decrypt_pad,
		\u2_R6_reg[12]/NET0131 ,
		\u2_uk_K_r6_reg[26]/NET0131 ,
		\u2_uk_K_r6_reg[33]/NET0131 ,
		_w10763_
	);
	LUT4 #(
		.INIT('h5100)
	) name4937 (
		_w10762_,
		_w10758_,
		_w10761_,
		_w10763_,
		_w10764_
	);
	LUT2 #(
		.INIT('h6)
	) name4938 (
		_w10755_,
		_w10760_,
		_w10765_
	);
	LUT4 #(
		.INIT('h9990)
	) name4939 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10766_
	);
	LUT4 #(
		.INIT('h0990)
	) name4940 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10767_
	);
	LUT4 #(
		.INIT('h4000)
	) name4941 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10768_
	);
	LUT4 #(
		.INIT('h0400)
	) name4942 (
		_w10760_,
		_w10756_,
		_w10759_,
		_w10757_,
		_w10769_
	);
	LUT3 #(
		.INIT('h01)
	) name4943 (
		_w10763_,
		_w10769_,
		_w10768_,
		_w10770_
	);
	LUT4 #(
		.INIT('h2000)
	) name4944 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10771_
	);
	LUT4 #(
		.INIT('h0203)
	) name4945 (
		_w10760_,
		_w10756_,
		_w10759_,
		_w10757_,
		_w10772_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name4946 (
		_w10757_,
		_w10771_,
		_w10765_,
		_w10772_,
		_w10773_
	);
	LUT4 #(
		.INIT('h4555)
	) name4947 (
		_w10764_,
		_w10767_,
		_w10770_,
		_w10773_,
		_w10774_
	);
	LUT4 #(
		.INIT('h95b5)
	) name4948 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10775_
	);
	LUT4 #(
		.INIT('h0001)
	) name4949 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10776_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name4950 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10777_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4951 (
		_w10757_,
		_w10763_,
		_w10775_,
		_w10777_,
		_w10778_
	);
	LUT3 #(
		.INIT('h56)
	) name4952 (
		\u2_L6_reg[6]/NET0131 ,
		_w10774_,
		_w10778_,
		_w10779_
	);
	LUT4 #(
		.INIT('h135c)
	) name4953 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10780_
	);
	LUT2 #(
		.INIT('h4)
	) name4954 (
		_w10320_,
		_w10312_,
		_w10781_
	);
	LUT3 #(
		.INIT('h04)
	) name4955 (
		_w10732_,
		_w10781_,
		_w10780_,
		_w10782_
	);
	LUT4 #(
		.INIT('h6c82)
	) name4956 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10783_
	);
	LUT2 #(
		.INIT('h9)
	) name4957 (
		_w10320_,
		_w10312_,
		_w10784_
	);
	LUT2 #(
		.INIT('h4)
	) name4958 (
		_w10783_,
		_w10784_,
		_w10785_
	);
	LUT4 #(
		.INIT('h0010)
	) name4959 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10786_
	);
	LUT4 #(
		.INIT('h22a8)
	) name4960 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10316_,
		_w10787_
	);
	LUT3 #(
		.INIT('h41)
	) name4961 (
		_w10314_,
		_w10311_,
		_w10315_,
		_w10788_
	);
	LUT3 #(
		.INIT('h02)
	) name4962 (
		_w10735_,
		_w10787_,
		_w10788_,
		_w10789_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4963 (
		_w10782_,
		_w10785_,
		_w10786_,
		_w10789_,
		_w10790_
	);
	LUT2 #(
		.INIT('h6)
	) name4964 (
		\u2_L6_reg[7]/NET0131 ,
		_w10790_,
		_w10791_
	);
	LUT4 #(
		.INIT('h8228)
	) name4965 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10792_
	);
	LUT3 #(
		.INIT('h19)
	) name4966 (
		_w10253_,
		_w10252_,
		_w10254_,
		_w10793_
	);
	LUT4 #(
		.INIT('h0013)
	) name4967 (
		_w10262_,
		_w10350_,
		_w10793_,
		_w10792_,
		_w10794_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name4968 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10795_
	);
	LUT2 #(
		.INIT('h1)
	) name4969 (
		_w10250_,
		_w10795_,
		_w10796_
	);
	LUT4 #(
		.INIT('hc7c3)
	) name4970 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10797_
	);
	LUT4 #(
		.INIT('h9ffd)
	) name4971 (
		_w10251_,
		_w10253_,
		_w10252_,
		_w10254_,
		_w10798_
	);
	LUT4 #(
		.INIT('h8d00)
	) name4972 (
		_w10250_,
		_w10797_,
		_w10793_,
		_w10798_,
		_w10799_
	);
	LUT4 #(
		.INIT('h3210)
	) name4973 (
		_w10249_,
		_w10796_,
		_w10799_,
		_w10794_,
		_w10800_
	);
	LUT2 #(
		.INIT('h9)
	) name4974 (
		\u2_L6_reg[9]/NET0131 ,
		_w10800_,
		_w10801_
	);
	LUT4 #(
		.INIT('h6979)
	) name4975 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10757_,
		_w10802_
	);
	LUT3 #(
		.INIT('h07)
	) name4976 (
		_w10760_,
		_w10759_,
		_w10757_,
		_w10803_
	);
	LUT4 #(
		.INIT('h0014)
	) name4977 (
		_w10755_,
		_w10760_,
		_w10759_,
		_w10757_,
		_w10804_
	);
	LUT4 #(
		.INIT('h0032)
	) name4978 (
		_w10759_,
		_w10771_,
		_w10802_,
		_w10804_,
		_w10805_
	);
	LUT3 #(
		.INIT('he0)
	) name4979 (
		_w10755_,
		_w10760_,
		_w10757_,
		_w10806_
	);
	LUT4 #(
		.INIT('h6800)
	) name4980 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10757_,
		_w10807_
	);
	LUT3 #(
		.INIT('h0d)
	) name4981 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10808_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name4982 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10809_
	);
	LUT4 #(
		.INIT('h0f02)
	) name4983 (
		_w10757_,
		_w10776_,
		_w10807_,
		_w10809_,
		_w10810_
	);
	LUT3 #(
		.INIT('h08)
	) name4984 (
		_w10760_,
		_w10759_,
		_w10757_,
		_w10811_
	);
	LUT4 #(
		.INIT('h0020)
	) name4985 (
		_w10760_,
		_w10756_,
		_w10759_,
		_w10757_,
		_w10812_
	);
	LUT4 #(
		.INIT('hbeff)
	) name4986 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10813_
	);
	LUT3 #(
		.INIT('h31)
	) name4987 (
		_w10757_,
		_w10812_,
		_w10813_,
		_w10814_
	);
	LUT4 #(
		.INIT('hd800)
	) name4988 (
		_w10763_,
		_w10805_,
		_w10810_,
		_w10814_,
		_w10815_
	);
	LUT2 #(
		.INIT('h9)
	) name4989 (
		\u2_L6_reg[16]/NET0131 ,
		_w10815_,
		_w10816_
	);
	LUT4 #(
		.INIT('hef2f)
	) name4990 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10817_
	);
	LUT4 #(
		.INIT('h0100)
	) name4991 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10818_
	);
	LUT4 #(
		.INIT('h0b08)
	) name4992 (
		_w10406_,
		_w10409_,
		_w10818_,
		_w10817_,
		_w10819_
	);
	LUT4 #(
		.INIT('h0121)
	) name4993 (
		_w10402_,
		_w10404_,
		_w10407_,
		_w10409_,
		_w10820_
	);
	LUT4 #(
		.INIT('h9fff)
	) name4994 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10821_
	);
	LUT4 #(
		.INIT('h8000)
	) name4995 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10409_,
		_w10822_
	);
	LUT4 #(
		.INIT('h0100)
	) name4996 (
		_w10525_,
		_w10822_,
		_w10820_,
		_w10821_,
		_w10823_
	);
	LUT4 #(
		.INIT('h0008)
	) name4997 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10409_,
		_w10824_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name4998 (
		_w10402_,
		_w10403_,
		_w10404_,
		_w10407_,
		_w10825_
	);
	LUT3 #(
		.INIT('h31)
	) name4999 (
		_w10409_,
		_w10824_,
		_w10825_,
		_w10826_
	);
	LUT4 #(
		.INIT('hd800)
	) name5000 (
		_w10401_,
		_w10819_,
		_w10823_,
		_w10826_,
		_w10827_
	);
	LUT2 #(
		.INIT('h9)
	) name5001 (
		\u2_L6_reg[18]/P0001 ,
		_w10827_,
		_w10828_
	);
	LUT3 #(
		.INIT('hed)
	) name5002 (
		_w10755_,
		_w10760_,
		_w10759_,
		_w10829_
	);
	LUT3 #(
		.INIT('h20)
	) name5003 (
		_w10760_,
		_w10756_,
		_w10759_,
		_w10830_
	);
	LUT4 #(
		.INIT('hef00)
	) name5004 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10757_,
		_w10831_
	);
	LUT3 #(
		.INIT('h20)
	) name5005 (
		_w10829_,
		_w10830_,
		_w10831_,
		_w10832_
	);
	LUT4 #(
		.INIT('h0009)
	) name5006 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10833_
	);
	LUT4 #(
		.INIT('h6640)
	) name5007 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10834_
	);
	LUT3 #(
		.INIT('h01)
	) name5008 (
		_w10757_,
		_w10834_,
		_w10833_,
		_w10835_
	);
	LUT3 #(
		.INIT('h54)
	) name5009 (
		_w10763_,
		_w10832_,
		_w10835_,
		_w10836_
	);
	LUT2 #(
		.INIT('h4)
	) name5010 (
		_w10757_,
		_w10766_,
		_w10837_
	);
	LUT3 #(
		.INIT('h2a)
	) name5011 (
		_w10763_,
		_w10765_,
		_w10772_,
		_w10838_
	);
	LUT3 #(
		.INIT('hd0)
	) name5012 (
		_w10760_,
		_w10756_,
		_w10759_,
		_w10839_
	);
	LUT2 #(
		.INIT('h4)
	) name5013 (
		_w10759_,
		_w10757_,
		_w10840_
	);
	LUT4 #(
		.INIT('h153f)
	) name5014 (
		_w10806_,
		_w10808_,
		_w10840_,
		_w10839_,
		_w10841_
	);
	LUT3 #(
		.INIT('h40)
	) name5015 (
		_w10837_,
		_w10838_,
		_w10841_,
		_w10842_
	);
	LUT2 #(
		.INIT('h8)
	) name5016 (
		_w10755_,
		_w10756_,
		_w10843_
	);
	LUT3 #(
		.INIT('h53)
	) name5017 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10844_
	);
	LUT4 #(
		.INIT('h0700)
	) name5018 (
		_w10755_,
		_w10760_,
		_w10759_,
		_w10757_,
		_w10845_
	);
	LUT4 #(
		.INIT('h7077)
	) name5019 (
		_w10811_,
		_w10843_,
		_w10844_,
		_w10845_,
		_w10846_
	);
	LUT4 #(
		.INIT('ha955)
	) name5020 (
		\u2_L6_reg[24]/NET0131 ,
		_w10836_,
		_w10842_,
		_w10846_,
		_w10847_
	);
	LUT4 #(
		.INIT('h8c00)
	) name5021 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10848_
	);
	LUT4 #(
		.INIT('h00fb)
	) name5022 (
		_w10755_,
		_w10756_,
		_w10759_,
		_w10763_,
		_w10849_
	);
	LUT2 #(
		.INIT('h4)
	) name5023 (
		_w10848_,
		_w10849_,
		_w10850_
	);
	LUT4 #(
		.INIT('h0004)
	) name5024 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10851_
	);
	LUT4 #(
		.INIT('haa2a)
	) name5025 (
		_w10757_,
		_w10763_,
		_w10829_,
		_w10851_,
		_w10852_
	);
	LUT2 #(
		.INIT('h4)
	) name5026 (
		_w10850_,
		_w10852_,
		_w10853_
	);
	LUT4 #(
		.INIT('h23ef)
	) name5027 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10854_
	);
	LUT4 #(
		.INIT('h7000)
	) name5028 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10855_
	);
	LUT4 #(
		.INIT('h0c08)
	) name5029 (
		_w10757_,
		_w10763_,
		_w10855_,
		_w10854_,
		_w10856_
	);
	LUT2 #(
		.INIT('h1)
	) name5030 (
		_w10763_,
		_w10833_,
		_w10857_
	);
	LUT4 #(
		.INIT('h0200)
	) name5031 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10759_,
		_w10858_
	);
	LUT3 #(
		.INIT('h0d)
	) name5032 (
		_w10803_,
		_w10844_,
		_w10858_,
		_w10859_
	);
	LUT4 #(
		.INIT('hf700)
	) name5033 (
		_w10755_,
		_w10760_,
		_w10756_,
		_w10757_,
		_w10860_
	);
	LUT4 #(
		.INIT('hf040)
	) name5034 (
		_w10755_,
		_w10756_,
		_w10759_,
		_w10757_,
		_w10861_
	);
	LUT2 #(
		.INIT('h4)
	) name5035 (
		_w10860_,
		_w10861_,
		_w10862_
	);
	LUT4 #(
		.INIT('h00ea)
	) name5036 (
		_w10856_,
		_w10857_,
		_w10859_,
		_w10862_,
		_w10863_
	);
	LUT3 #(
		.INIT('h9a)
	) name5037 (
		\u2_L6_reg[30]/NET0131 ,
		_w10853_,
		_w10863_,
		_w10864_
	);
	LUT4 #(
		.INIT('hc693)
	) name5038 (
		decrypt_pad,
		\u2_R5_reg[28]/NET0131 ,
		\u2_uk_K_r5_reg[44]/NET0131 ,
		\u2_uk_K_r5_reg[9]/P0001 ,
		_w10865_
	);
	LUT4 #(
		.INIT('hc963)
	) name5039 (
		decrypt_pad,
		\u2_R5_reg[27]/NET0131 ,
		\u2_uk_K_r5_reg[22]/NET0131 ,
		\u2_uk_K_r5_reg[2]/NET0131 ,
		_w10866_
	);
	LUT4 #(
		.INIT('hc963)
	) name5040 (
		decrypt_pad,
		\u2_R5_reg[26]/NET0131 ,
		\u2_uk_K_r5_reg[44]/NET0131 ,
		\u2_uk_K_r5_reg[52]/NET0131 ,
		_w10867_
	);
	LUT4 #(
		.INIT('hc693)
	) name5041 (
		decrypt_pad,
		\u2_R5_reg[24]/NET0131 ,
		\u2_uk_K_r5_reg[28]/NET0131 ,
		\u2_uk_K_r5_reg[52]/NET0131 ,
		_w10868_
	);
	LUT4 #(
		.INIT('hc963)
	) name5042 (
		decrypt_pad,
		\u2_R5_reg[29]/NET0131 ,
		\u2_uk_K_r5_reg[1]/NET0131 ,
		\u2_uk_K_r5_reg[36]/NET0131 ,
		_w10869_
	);
	LUT4 #(
		.INIT('hc963)
	) name5043 (
		decrypt_pad,
		\u2_R5_reg[25]/NET0131 ,
		\u2_uk_K_r5_reg[28]/NET0131 ,
		\u2_uk_K_r5_reg[8]/NET0131 ,
		_w10870_
	);
	LUT4 #(
		.INIT('h5f67)
	) name5044 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w10871_
	);
	LUT2 #(
		.INIT('h1)
	) name5045 (
		_w10866_,
		_w10871_,
		_w10872_
	);
	LUT2 #(
		.INIT('h8)
	) name5046 (
		_w10868_,
		_w10866_,
		_w10873_
	);
	LUT4 #(
		.INIT('hddaf)
	) name5047 (
		_w10868_,
		_w10870_,
		_w10869_,
		_w10866_,
		_w10874_
	);
	LUT3 #(
		.INIT('h7b)
	) name5048 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10875_
	);
	LUT3 #(
		.INIT('h02)
	) name5049 (
		_w10868_,
		_w10867_,
		_w10869_,
		_w10876_
	);
	LUT4 #(
		.INIT('h0002)
	) name5050 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w10877_
	);
	LUT4 #(
		.INIT('h7bfd)
	) name5051 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w10878_
	);
	LUT3 #(
		.INIT('he0)
	) name5052 (
		_w10867_,
		_w10874_,
		_w10878_,
		_w10879_
	);
	LUT3 #(
		.INIT('h45)
	) name5053 (
		_w10865_,
		_w10872_,
		_w10879_,
		_w10880_
	);
	LUT3 #(
		.INIT('h9b)
	) name5054 (
		_w10870_,
		_w10867_,
		_w10869_,
		_w10881_
	);
	LUT4 #(
		.INIT('h1000)
	) name5055 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w10882_
	);
	LUT4 #(
		.INIT('heffe)
	) name5056 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w10883_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5057 (
		_w10865_,
		_w10873_,
		_w10881_,
		_w10883_,
		_w10884_
	);
	LUT4 #(
		.INIT('h0200)
	) name5058 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w10885_
	);
	LUT4 #(
		.INIT('hb9ff)
	) name5059 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w10886_
	);
	LUT4 #(
		.INIT('h005d)
	) name5060 (
		_w10875_,
		_w10865_,
		_w10886_,
		_w10866_,
		_w10887_
	);
	LUT4 #(
		.INIT('h0040)
	) name5061 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w10888_
	);
	LUT4 #(
		.INIT('hef9c)
	) name5062 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w10889_
	);
	LUT2 #(
		.INIT('h2)
	) name5063 (
		_w10866_,
		_w10889_,
		_w10890_
	);
	LUT3 #(
		.INIT('h01)
	) name5064 (
		_w10887_,
		_w10890_,
		_w10884_,
		_w10891_
	);
	LUT3 #(
		.INIT('h65)
	) name5065 (
		\u2_L5_reg[22]/NET0131 ,
		_w10880_,
		_w10891_,
		_w10892_
	);
	LUT4 #(
		.INIT('hc693)
	) name5066 (
		decrypt_pad,
		\u2_R5_reg[4]/NET0131 ,
		\u2_uk_K_r5_reg[11]/NET0131 ,
		\u2_uk_K_r5_reg[33]/NET0131 ,
		_w10893_
	);
	LUT4 #(
		.INIT('hc693)
	) name5067 (
		decrypt_pad,
		\u2_R5_reg[3]/NET0131 ,
		\u2_uk_K_r5_reg[33]/NET0131 ,
		\u2_uk_K_r5_reg[55]/NET0131 ,
		_w10894_
	);
	LUT4 #(
		.INIT('hc693)
	) name5068 (
		decrypt_pad,
		\u2_R5_reg[1]/NET0131 ,
		\u2_uk_K_r5_reg[41]/NET0131 ,
		\u2_uk_K_r5_reg[6]/NET0131 ,
		_w10895_
	);
	LUT4 #(
		.INIT('hc693)
	) name5069 (
		decrypt_pad,
		\u2_R5_reg[5]/NET0131 ,
		\u2_uk_K_r5_reg[39]/NET0131 ,
		\u2_uk_K_r5_reg[4]/NET0131 ,
		_w10896_
	);
	LUT4 #(
		.INIT('hc693)
	) name5070 (
		decrypt_pad,
		\u2_R5_reg[2]/NET0131 ,
		\u2_uk_K_r5_reg[24]/NET0131 ,
		\u2_uk_K_r5_reg[46]/NET0131 ,
		_w10897_
	);
	LUT4 #(
		.INIT('hc963)
	) name5071 (
		decrypt_pad,
		\u2_R5_reg[32]/NET0131 ,
		\u2_uk_K_r5_reg[10]/NET0131 ,
		\u2_uk_K_r5_reg[20]/NET0131 ,
		_w10898_
	);
	LUT4 #(
		.INIT('hcfc5)
	) name5072 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w10899_
	);
	LUT2 #(
		.INIT('h2)
	) name5073 (
		_w10894_,
		_w10899_,
		_w10900_
	);
	LUT2 #(
		.INIT('h2)
	) name5074 (
		_w10896_,
		_w10898_,
		_w10901_
	);
	LUT2 #(
		.INIT('h2)
	) name5075 (
		_w10894_,
		_w10897_,
		_w10902_
	);
	LUT3 #(
		.INIT('hd0)
	) name5076 (
		_w10894_,
		_w10897_,
		_w10895_,
		_w10903_
	);
	LUT4 #(
		.INIT('h500c)
	) name5077 (
		_w10894_,
		_w10897_,
		_w10895_,
		_w10898_,
		_w10904_
	);
	LUT2 #(
		.INIT('h1)
	) name5078 (
		_w10895_,
		_w10896_,
		_w10905_
	);
	LUT4 #(
		.INIT('h0100)
	) name5079 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w10906_
	);
	LUT4 #(
		.INIT('h0031)
	) name5080 (
		_w10901_,
		_w10904_,
		_w10903_,
		_w10906_,
		_w10907_
	);
	LUT3 #(
		.INIT('h8a)
	) name5081 (
		_w10893_,
		_w10900_,
		_w10907_,
		_w10908_
	);
	LUT4 #(
		.INIT('h4703)
	) name5082 (
		_w10894_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w10909_
	);
	LUT3 #(
		.INIT('h41)
	) name5083 (
		_w10897_,
		_w10896_,
		_w10898_,
		_w10910_
	);
	LUT2 #(
		.INIT('h4)
	) name5084 (
		_w10909_,
		_w10910_,
		_w10911_
	);
	LUT3 #(
		.INIT('h28)
	) name5085 (
		_w10895_,
		_w10896_,
		_w10898_,
		_w10912_
	);
	LUT2 #(
		.INIT('h2)
	) name5086 (
		_w10897_,
		_w10895_,
		_w10913_
	);
	LUT4 #(
		.INIT('hfdba)
	) name5087 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w10914_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name5088 (
		_w10894_,
		_w10897_,
		_w10912_,
		_w10914_,
		_w10915_
	);
	LUT3 #(
		.INIT('h45)
	) name5089 (
		_w10893_,
		_w10911_,
		_w10915_,
		_w10916_
	);
	LUT3 #(
		.INIT('h80)
	) name5090 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10917_
	);
	LUT4 #(
		.INIT('h7bdb)
	) name5091 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w10918_
	);
	LUT2 #(
		.INIT('h1)
	) name5092 (
		_w10894_,
		_w10918_,
		_w10919_
	);
	LUT4 #(
		.INIT('h0200)
	) name5093 (
		_w10894_,
		_w10897_,
		_w10895_,
		_w10898_,
		_w10920_
	);
	LUT3 #(
		.INIT('h02)
	) name5094 (
		_w10894_,
		_w10896_,
		_w10898_,
		_w10921_
	);
	LUT3 #(
		.INIT('h13)
	) name5095 (
		_w10913_,
		_w10920_,
		_w10921_,
		_w10922_
	);
	LUT2 #(
		.INIT('h4)
	) name5096 (
		_w10919_,
		_w10922_,
		_w10923_
	);
	LUT4 #(
		.INIT('h5655)
	) name5097 (
		\u2_L5_reg[31]/NET0131 ,
		_w10916_,
		_w10908_,
		_w10923_,
		_w10924_
	);
	LUT4 #(
		.INIT('hc963)
	) name5098 (
		decrypt_pad,
		\u2_R5_reg[24]/NET0131 ,
		\u2_uk_K_r5_reg[2]/NET0131 ,
		\u2_uk_K_r5_reg[37]/P0001 ,
		_w10925_
	);
	LUT4 #(
		.INIT('hc693)
	) name5099 (
		decrypt_pad,
		\u2_R5_reg[20]/NET0131 ,
		\u2_uk_K_r5_reg[16]/NET0131 ,
		\u2_uk_K_r5_reg[36]/NET0131 ,
		_w10926_
	);
	LUT4 #(
		.INIT('hc693)
	) name5100 (
		decrypt_pad,
		\u2_R5_reg[22]/NET0131 ,
		\u2_uk_K_r5_reg[22]/NET0131 ,
		\u2_uk_K_r5_reg[42]/NET0131 ,
		_w10927_
	);
	LUT4 #(
		.INIT('hc693)
	) name5101 (
		decrypt_pad,
		\u2_R5_reg[21]/NET0131 ,
		\u2_uk_K_r5_reg[0]/NET0131 ,
		\u2_uk_K_r5_reg[51]/NET0131 ,
		_w10928_
	);
	LUT4 #(
		.INIT('hc963)
	) name5102 (
		decrypt_pad,
		\u2_R5_reg[23]/NET0131 ,
		\u2_uk_K_r5_reg[0]/NET0131 ,
		\u2_uk_K_r5_reg[35]/NET0131 ,
		_w10929_
	);
	LUT4 #(
		.INIT('h4155)
	) name5103 (
		_w10929_,
		_w10926_,
		_w10927_,
		_w10928_,
		_w10930_
	);
	LUT4 #(
		.INIT('hc693)
	) name5104 (
		decrypt_pad,
		\u2_R5_reg[25]/NET0131 ,
		\u2_uk_K_r5_reg[1]/NET0131 ,
		\u2_uk_K_r5_reg[21]/NET0131 ,
		_w10931_
	);
	LUT4 #(
		.INIT('haa8a)
	) name5105 (
		_w10929_,
		_w10926_,
		_w10931_,
		_w10928_,
		_w10932_
	);
	LUT3 #(
		.INIT('he6)
	) name5106 (
		_w10926_,
		_w10927_,
		_w10928_,
		_w10933_
	);
	LUT3 #(
		.INIT('h13)
	) name5107 (
		_w10932_,
		_w10930_,
		_w10933_,
		_w10934_
	);
	LUT4 #(
		.INIT('h0080)
	) name5108 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w10935_
	);
	LUT2 #(
		.INIT('h2)
	) name5109 (
		_w10926_,
		_w10931_,
		_w10936_
	);
	LUT2 #(
		.INIT('h1)
	) name5110 (
		_w10929_,
		_w10927_,
		_w10937_
	);
	LUT3 #(
		.INIT('hce)
	) name5111 (
		_w10929_,
		_w10927_,
		_w10928_,
		_w10938_
	);
	LUT3 #(
		.INIT('h31)
	) name5112 (
		_w10936_,
		_w10935_,
		_w10938_,
		_w10939_
	);
	LUT3 #(
		.INIT('h45)
	) name5113 (
		_w10925_,
		_w10934_,
		_w10939_,
		_w10940_
	);
	LUT4 #(
		.INIT('h0002)
	) name5114 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w10941_
	);
	LUT4 #(
		.INIT('h27fd)
	) name5115 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w10942_
	);
	LUT2 #(
		.INIT('h2)
	) name5116 (
		_w10929_,
		_w10942_,
		_w10943_
	);
	LUT4 #(
		.INIT('h0415)
	) name5117 (
		_w10929_,
		_w10926_,
		_w10931_,
		_w10928_,
		_w10944_
	);
	LUT4 #(
		.INIT('h0b07)
	) name5118 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w10945_
	);
	LUT3 #(
		.INIT('h0e)
	) name5119 (
		_w10937_,
		_w10944_,
		_w10945_,
		_w10946_
	);
	LUT3 #(
		.INIT('he0)
	) name5120 (
		_w10943_,
		_w10946_,
		_w10925_,
		_w10947_
	);
	LUT4 #(
		.INIT('h5155)
	) name5121 (
		_w10929_,
		_w10926_,
		_w10931_,
		_w10928_,
		_w10948_
	);
	LUT3 #(
		.INIT('h01)
	) name5122 (
		_w10927_,
		_w10948_,
		_w10932_,
		_w10949_
	);
	LUT4 #(
		.INIT('h7077)
	) name5123 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w10950_
	);
	LUT4 #(
		.INIT('haa02)
	) name5124 (
		_w10929_,
		_w10926_,
		_w10931_,
		_w10927_,
		_w10951_
	);
	LUT3 #(
		.INIT('h01)
	) name5125 (
		_w10926_,
		_w10931_,
		_w10928_,
		_w10952_
	);
	LUT4 #(
		.INIT('h45cf)
	) name5126 (
		_w10937_,
		_w10950_,
		_w10951_,
		_w10952_,
		_w10953_
	);
	LUT2 #(
		.INIT('h4)
	) name5127 (
		_w10949_,
		_w10953_,
		_w10954_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5128 (
		\u2_L5_reg[11]/NET0131 ,
		_w10947_,
		_w10940_,
		_w10954_,
		_w10955_
	);
	LUT4 #(
		.INIT('hc963)
	) name5129 (
		decrypt_pad,
		\u2_R5_reg[14]/NET0131 ,
		\u2_uk_K_r5_reg[19]/NET0131 ,
		\u2_uk_K_r5_reg[54]/NET0131 ,
		_w10956_
	);
	LUT4 #(
		.INIT('hc963)
	) name5130 (
		decrypt_pad,
		\u2_R5_reg[12]/NET0131 ,
		\u2_uk_K_r5_reg[24]/NET0131 ,
		\u2_uk_K_r5_reg[34]/NET0131 ,
		_w10957_
	);
	LUT4 #(
		.INIT('hc693)
	) name5131 (
		decrypt_pad,
		\u2_R5_reg[17]/NET0131 ,
		\u2_uk_K_r5_reg[18]/NET0131 ,
		\u2_uk_K_r5_reg[40]/NET0131 ,
		_w10958_
	);
	LUT3 #(
		.INIT('h08)
	) name5132 (
		_w10957_,
		_w10956_,
		_w10958_,
		_w10959_
	);
	LUT4 #(
		.INIT('hc963)
	) name5133 (
		decrypt_pad,
		\u2_R5_reg[15]/NET0131 ,
		\u2_uk_K_r5_reg[27]/NET0131 ,
		\u2_uk_K_r5_reg[5]/NET0131 ,
		_w10960_
	);
	LUT4 #(
		.INIT('hc963)
	) name5134 (
		decrypt_pad,
		\u2_R5_reg[13]/NET0131 ,
		\u2_uk_K_r5_reg[18]/NET0131 ,
		\u2_uk_K_r5_reg[53]/NET0131 ,
		_w10961_
	);
	LUT3 #(
		.INIT('h0b)
	) name5135 (
		_w10961_,
		_w10958_,
		_w10960_,
		_w10962_
	);
	LUT4 #(
		.INIT('h7e00)
	) name5136 (
		_w10961_,
		_w10957_,
		_w10958_,
		_w10960_,
		_w10963_
	);
	LUT3 #(
		.INIT('h0b)
	) name5137 (
		_w10959_,
		_w10962_,
		_w10963_,
		_w10964_
	);
	LUT3 #(
		.INIT('h04)
	) name5138 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10965_
	);
	LUT4 #(
		.INIT('h0400)
	) name5139 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w10966_
	);
	LUT4 #(
		.INIT('hc693)
	) name5140 (
		decrypt_pad,
		\u2_R5_reg[16]/NET0131 ,
		\u2_uk_K_r5_reg[13]/P0001 ,
		\u2_uk_K_r5_reg[3]/NET0131 ,
		_w10967_
	);
	LUT2 #(
		.INIT('h1)
	) name5141 (
		_w10966_,
		_w10967_,
		_w10968_
	);
	LUT4 #(
		.INIT('h0001)
	) name5142 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w10969_
	);
	LUT2 #(
		.INIT('h8)
	) name5143 (
		_w10956_,
		_w10960_,
		_w10970_
	);
	LUT3 #(
		.INIT('h80)
	) name5144 (
		_w10961_,
		_w10956_,
		_w10960_,
		_w10971_
	);
	LUT4 #(
		.INIT('h2000)
	) name5145 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10960_,
		_w10972_
	);
	LUT4 #(
		.INIT('h0020)
	) name5146 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w10973_
	);
	LUT3 #(
		.INIT('h01)
	) name5147 (
		_w10972_,
		_w10973_,
		_w10969_,
		_w10974_
	);
	LUT3 #(
		.INIT('h40)
	) name5148 (
		_w10964_,
		_w10968_,
		_w10974_,
		_w10975_
	);
	LUT2 #(
		.INIT('h9)
	) name5149 (
		_w10961_,
		_w10957_,
		_w10976_
	);
	LUT4 #(
		.INIT('h0010)
	) name5150 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w10977_
	);
	LUT4 #(
		.INIT('hf9e9)
	) name5151 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w10978_
	);
	LUT2 #(
		.INIT('h1)
	) name5152 (
		_w10960_,
		_w10978_,
		_w10979_
	);
	LUT2 #(
		.INIT('h4)
	) name5153 (
		_w10957_,
		_w10958_,
		_w10980_
	);
	LUT4 #(
		.INIT('h0200)
	) name5154 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w10981_
	);
	LUT4 #(
		.INIT('h7dff)
	) name5155 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w10982_
	);
	LUT4 #(
		.INIT('h1000)
	) name5156 (
		_w10961_,
		_w10957_,
		_w10958_,
		_w10960_,
		_w10983_
	);
	LUT4 #(
		.INIT('h0800)
	) name5157 (
		_w10961_,
		_w10957_,
		_w10958_,
		_w10960_,
		_w10984_
	);
	LUT4 #(
		.INIT('h0008)
	) name5158 (
		_w10967_,
		_w10982_,
		_w10984_,
		_w10983_,
		_w10985_
	);
	LUT2 #(
		.INIT('h4)
	) name5159 (
		_w10979_,
		_w10985_,
		_w10986_
	);
	LUT4 #(
		.INIT('hffb6)
	) name5160 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w10987_
	);
	LUT3 #(
		.INIT('hb1)
	) name5161 (
		_w10960_,
		_w10981_,
		_w10987_,
		_w10988_
	);
	LUT4 #(
		.INIT('ha955)
	) name5162 (
		\u2_L5_reg[20]/NET0131 ,
		_w10975_,
		_w10986_,
		_w10988_,
		_w10989_
	);
	LUT4 #(
		.INIT('hc963)
	) name5163 (
		decrypt_pad,
		\u2_R5_reg[32]/NET0131 ,
		\u2_uk_K_r5_reg[29]/NET0131 ,
		\u2_uk_K_r5_reg[9]/P0001 ,
		_w10990_
	);
	LUT4 #(
		.INIT('hc693)
	) name5164 (
		decrypt_pad,
		\u2_R5_reg[28]/NET0131 ,
		\u2_uk_K_r5_reg[42]/NET0131 ,
		\u2_uk_K_r5_reg[7]/NET0131 ,
		_w10991_
	);
	LUT4 #(
		.INIT('hc693)
	) name5165 (
		decrypt_pad,
		\u2_R5_reg[30]/NET0131 ,
		\u2_uk_K_r5_reg[15]/NET0131 ,
		\u2_uk_K_r5_reg[35]/NET0131 ,
		_w10992_
	);
	LUT4 #(
		.INIT('hc693)
	) name5166 (
		decrypt_pad,
		\u2_R5_reg[29]/NET0131 ,
		\u2_uk_K_r5_reg[14]/NET0131 ,
		\u2_uk_K_r5_reg[38]/NET0131 ,
		_w10993_
	);
	LUT4 #(
		.INIT('hc693)
	) name5167 (
		decrypt_pad,
		\u2_R5_reg[1]/NET0131 ,
		\u2_uk_K_r5_reg[30]/NET0131 ,
		\u2_uk_K_r5_reg[50]/NET0131 ,
		_w10994_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name5168 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w10995_
	);
	LUT4 #(
		.INIT('hc963)
	) name5169 (
		decrypt_pad,
		\u2_R5_reg[31]/P0001 ,
		\u2_uk_K_r5_reg[23]/NET0131 ,
		\u2_uk_K_r5_reg[31]/NET0131 ,
		_w10996_
	);
	LUT4 #(
		.INIT('h0020)
	) name5170 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w10997_
	);
	LUT3 #(
		.INIT('h02)
	) name5171 (
		_w10996_,
		_w10997_,
		_w10995_,
		_w10998_
	);
	LUT4 #(
		.INIT('h0041)
	) name5172 (
		_w10996_,
		_w10991_,
		_w10992_,
		_w10993_,
		_w10999_
	);
	LUT4 #(
		.INIT('h4000)
	) name5173 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11000_
	);
	LUT2 #(
		.INIT('h1)
	) name5174 (
		_w10999_,
		_w11000_,
		_w11001_
	);
	LUT3 #(
		.INIT('h8a)
	) name5175 (
		_w10990_,
		_w10998_,
		_w11001_,
		_w11002_
	);
	LUT4 #(
		.INIT('h0d99)
	) name5176 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11003_
	);
	LUT4 #(
		.INIT('h8020)
	) name5177 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11004_
	);
	LUT4 #(
		.INIT('hfaf7)
	) name5178 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11005_
	);
	LUT4 #(
		.INIT('h3120)
	) name5179 (
		_w10996_,
		_w11004_,
		_w11005_,
		_w11003_,
		_w11006_
	);
	LUT4 #(
		.INIT('h0240)
	) name5180 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11007_
	);
	LUT4 #(
		.INIT('h0001)
	) name5181 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11008_
	);
	LUT4 #(
		.INIT('h0400)
	) name5182 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11009_
	);
	LUT4 #(
		.INIT('hf9be)
	) name5183 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11010_
	);
	LUT3 #(
		.INIT('hb1)
	) name5184 (
		_w10996_,
		_w10997_,
		_w11010_,
		_w11011_
	);
	LUT3 #(
		.INIT('he0)
	) name5185 (
		_w10990_,
		_w11006_,
		_w11011_,
		_w11012_
	);
	LUT3 #(
		.INIT('h9a)
	) name5186 (
		\u2_L5_reg[5]/NET0131 ,
		_w11002_,
		_w11012_,
		_w11013_
	);
	LUT4 #(
		.INIT('hfbdd)
	) name5187 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11014_
	);
	LUT4 #(
		.INIT('h6fff)
	) name5188 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11015_
	);
	LUT4 #(
		.INIT('hfd3b)
	) name5189 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11016_
	);
	LUT4 #(
		.INIT('hc840)
	) name5190 (
		_w10960_,
		_w11015_,
		_w11016_,
		_w11014_,
		_w11017_
	);
	LUT2 #(
		.INIT('h2)
	) name5191 (
		_w10967_,
		_w11017_,
		_w11018_
	);
	LUT3 #(
		.INIT('h40)
	) name5192 (
		_w10956_,
		_w10958_,
		_w10960_,
		_w11019_
	);
	LUT4 #(
		.INIT('h98cd)
	) name5193 (
		_w10961_,
		_w10956_,
		_w10958_,
		_w10960_,
		_w11020_
	);
	LUT2 #(
		.INIT('h2)
	) name5194 (
		_w10957_,
		_w11020_,
		_w11021_
	);
	LUT4 #(
		.INIT('hcefe)
	) name5195 (
		_w10961_,
		_w10957_,
		_w10958_,
		_w10960_,
		_w11022_
	);
	LUT3 #(
		.INIT('h32)
	) name5196 (
		_w10970_,
		_w10973_,
		_w11022_,
		_w11023_
	);
	LUT3 #(
		.INIT('h45)
	) name5197 (
		_w10967_,
		_w11021_,
		_w11023_,
		_w11024_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name5198 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11025_
	);
	LUT2 #(
		.INIT('h1)
	) name5199 (
		_w10960_,
		_w11025_,
		_w11026_
	);
	LUT3 #(
		.INIT('h23)
	) name5200 (
		_w10956_,
		_w10972_,
		_w10984_,
		_w11027_
	);
	LUT2 #(
		.INIT('h4)
	) name5201 (
		_w11026_,
		_w11027_,
		_w11028_
	);
	LUT4 #(
		.INIT('h5655)
	) name5202 (
		\u2_L5_reg[10]/NET0131 ,
		_w11018_,
		_w11024_,
		_w11028_,
		_w11029_
	);
	LUT4 #(
		.INIT('h0400)
	) name5203 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11030_
	);
	LUT4 #(
		.INIT('h000b)
	) name5204 (
		_w10866_,
		_w10882_,
		_w10888_,
		_w11030_,
		_w11031_
	);
	LUT4 #(
		.INIT('h7776)
	) name5205 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11032_
	);
	LUT2 #(
		.INIT('h2)
	) name5206 (
		_w10866_,
		_w11032_,
		_w11033_
	);
	LUT4 #(
		.INIT('h0020)
	) name5207 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11034_
	);
	LUT3 #(
		.INIT('h02)
	) name5208 (
		_w10865_,
		_w10885_,
		_w11034_,
		_w11035_
	);
	LUT3 #(
		.INIT('h40)
	) name5209 (
		_w11033_,
		_w11035_,
		_w11031_,
		_w11036_
	);
	LUT4 #(
		.INIT('hde54)
	) name5210 (
		_w10868_,
		_w10870_,
		_w10869_,
		_w10866_,
		_w11037_
	);
	LUT2 #(
		.INIT('h2)
	) name5211 (
		_w10867_,
		_w11037_,
		_w11038_
	);
	LUT4 #(
		.INIT('h0004)
	) name5212 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11039_
	);
	LUT3 #(
		.INIT('h01)
	) name5213 (
		_w10865_,
		_w10877_,
		_w11039_,
		_w11040_
	);
	LUT3 #(
		.INIT('h51)
	) name5214 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w11041_
	);
	LUT3 #(
		.INIT('hc8)
	) name5215 (
		_w10870_,
		_w10869_,
		_w10866_,
		_w11042_
	);
	LUT3 #(
		.INIT('h09)
	) name5216 (
		_w10870_,
		_w10869_,
		_w10866_,
		_w11043_
	);
	LUT3 #(
		.INIT('h07)
	) name5217 (
		_w11041_,
		_w11042_,
		_w11043_,
		_w11044_
	);
	LUT3 #(
		.INIT('h40)
	) name5218 (
		_w11038_,
		_w11040_,
		_w11044_,
		_w11045_
	);
	LUT3 #(
		.INIT('ha9)
	) name5219 (
		\u2_L5_reg[12]/NET0131 ,
		_w11036_,
		_w11045_,
		_w11046_
	);
	LUT4 #(
		.INIT('hc963)
	) name5220 (
		decrypt_pad,
		\u2_R5_reg[19]/NET0131 ,
		\u2_uk_K_r5_reg[30]/NET0131 ,
		\u2_uk_K_r5_reg[38]/NET0131 ,
		_w11047_
	);
	LUT4 #(
		.INIT('hc693)
	) name5221 (
		decrypt_pad,
		\u2_R5_reg[18]/NET0131 ,
		\u2_uk_K_r5_reg[23]/NET0131 ,
		\u2_uk_K_r5_reg[43]/NET0131 ,
		_w11048_
	);
	LUT4 #(
		.INIT('hc693)
	) name5222 (
		decrypt_pad,
		\u2_R5_reg[17]/NET0131 ,
		\u2_uk_K_r5_reg[29]/NET0131 ,
		\u2_uk_K_r5_reg[49]/NET0131 ,
		_w11049_
	);
	LUT4 #(
		.INIT('hc963)
	) name5223 (
		decrypt_pad,
		\u2_R5_reg[16]/NET0131 ,
		\u2_uk_K_r5_reg[31]/NET0131 ,
		\u2_uk_K_r5_reg[7]/NET0131 ,
		_w11050_
	);
	LUT4 #(
		.INIT('hc963)
	) name5224 (
		decrypt_pad,
		\u2_R5_reg[21]/NET0131 ,
		\u2_uk_K_r5_reg[15]/NET0131 ,
		\u2_uk_K_r5_reg[50]/NET0131 ,
		_w11051_
	);
	LUT3 #(
		.INIT('h04)
	) name5225 (
		_w11049_,
		_w11050_,
		_w11051_,
		_w11052_
	);
	LUT4 #(
		.INIT('h0010)
	) name5226 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11053_
	);
	LUT4 #(
		.INIT('h4000)
	) name5227 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11054_
	);
	LUT4 #(
		.INIT('hbc67)
	) name5228 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11055_
	);
	LUT4 #(
		.INIT('h5bf8)
	) name5229 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11056_
	);
	LUT4 #(
		.INIT('h2004)
	) name5230 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11057_
	);
	LUT4 #(
		.INIT('h00d8)
	) name5231 (
		_w11047_,
		_w11056_,
		_w11055_,
		_w11057_,
		_w11058_
	);
	LUT4 #(
		.INIT('hc963)
	) name5232 (
		decrypt_pad,
		\u2_R5_reg[20]/NET0131 ,
		\u2_uk_K_r5_reg[14]/NET0131 ,
		\u2_uk_K_r5_reg[49]/NET0131 ,
		_w11059_
	);
	LUT2 #(
		.INIT('h1)
	) name5233 (
		_w11058_,
		_w11059_,
		_w11060_
	);
	LUT4 #(
		.INIT('ha43f)
	) name5234 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11061_
	);
	LUT2 #(
		.INIT('h2)
	) name5235 (
		_w11047_,
		_w11061_,
		_w11062_
	);
	LUT3 #(
		.INIT('hde)
	) name5236 (
		_w11049_,
		_w11050_,
		_w11051_,
		_w11063_
	);
	LUT2 #(
		.INIT('h1)
	) name5237 (
		_w11047_,
		_w11048_,
		_w11064_
	);
	LUT2 #(
		.INIT('h4)
	) name5238 (
		_w11063_,
		_w11064_,
		_w11065_
	);
	LUT2 #(
		.INIT('h9)
	) name5239 (
		_w11048_,
		_w11049_,
		_w11066_
	);
	LUT4 #(
		.INIT('h0060)
	) name5240 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11067_
	);
	LUT4 #(
		.INIT('h7000)
	) name5241 (
		_w11047_,
		_w11048_,
		_w11050_,
		_w11051_,
		_w11068_
	);
	LUT3 #(
		.INIT('h13)
	) name5242 (
		_w11066_,
		_w11067_,
		_w11068_,
		_w11069_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5243 (
		_w11059_,
		_w11062_,
		_w11065_,
		_w11069_,
		_w11070_
	);
	LUT4 #(
		.INIT('h0040)
	) name5244 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11071_
	);
	LUT4 #(
		.INIT('hffbd)
	) name5245 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11072_
	);
	LUT4 #(
		.INIT('h0200)
	) name5246 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11073_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name5247 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11074_
	);
	LUT3 #(
		.INIT('hd8)
	) name5248 (
		_w11047_,
		_w11072_,
		_w11074_,
		_w11075_
	);
	LUT4 #(
		.INIT('h5655)
	) name5249 (
		\u2_L5_reg[14]/NET0131 ,
		_w11060_,
		_w11070_,
		_w11075_,
		_w11076_
	);
	LUT4 #(
		.INIT('h5f4f)
	) name5250 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11077_
	);
	LUT4 #(
		.INIT('h5a4f)
	) name5251 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11078_
	);
	LUT4 #(
		.INIT('h0002)
	) name5252 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11079_
	);
	LUT4 #(
		.INIT('h3302)
	) name5253 (
		_w10996_,
		_w10990_,
		_w11078_,
		_w11079_,
		_w11080_
	);
	LUT4 #(
		.INIT('h0800)
	) name5254 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11081_
	);
	LUT3 #(
		.INIT('h20)
	) name5255 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w11082_
	);
	LUT4 #(
		.INIT('h0400)
	) name5256 (
		_w10996_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11083_
	);
	LUT4 #(
		.INIT('h0002)
	) name5257 (
		_w10996_,
		_w10991_,
		_w10993_,
		_w10994_,
		_w11084_
	);
	LUT4 #(
		.INIT('h0040)
	) name5258 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11085_
	);
	LUT4 #(
		.INIT('h0001)
	) name5259 (
		_w11082_,
		_w11083_,
		_w11084_,
		_w11085_,
		_w11086_
	);
	LUT3 #(
		.INIT('h8a)
	) name5260 (
		_w10990_,
		_w11081_,
		_w11086_,
		_w11087_
	);
	LUT4 #(
		.INIT('h1040)
	) name5261 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11088_
	);
	LUT4 #(
		.INIT('h080a)
	) name5262 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10990_,
		_w11089_
	);
	LUT4 #(
		.INIT('h0001)
	) name5263 (
		_w10996_,
		_w11008_,
		_w11088_,
		_w11089_,
		_w11090_
	);
	LUT4 #(
		.INIT('h0100)
	) name5264 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11091_
	);
	LUT3 #(
		.INIT('h02)
	) name5265 (
		_w10996_,
		_w11000_,
		_w11091_,
		_w11092_
	);
	LUT2 #(
		.INIT('h1)
	) name5266 (
		_w11090_,
		_w11092_,
		_w11093_
	);
	LUT4 #(
		.INIT('h5556)
	) name5267 (
		\u2_L5_reg[15]/NET0131 ,
		_w11080_,
		_w11087_,
		_w11093_,
		_w11094_
	);
	LUT4 #(
		.INIT('hcff8)
	) name5268 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11095_
	);
	LUT3 #(
		.INIT('h8a)
	) name5269 (
		_w10894_,
		_w10895_,
		_w10896_,
		_w11096_
	);
	LUT4 #(
		.INIT('h8200)
	) name5270 (
		_w10894_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11097_
	);
	LUT4 #(
		.INIT('hf7df)
	) name5271 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11098_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5272 (
		_w10894_,
		_w11095_,
		_w11097_,
		_w11098_,
		_w11099_
	);
	LUT4 #(
		.INIT('h1000)
	) name5273 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11100_
	);
	LUT4 #(
		.INIT('hef11)
	) name5274 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11101_
	);
	LUT4 #(
		.INIT('h4401)
	) name5275 (
		_w10894_,
		_w10897_,
		_w10895_,
		_w10898_,
		_w11102_
	);
	LUT4 #(
		.INIT('h0400)
	) name5276 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11103_
	);
	LUT4 #(
		.INIT('h7b7f)
	) name5277 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11104_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5278 (
		_w10894_,
		_w11101_,
		_w11102_,
		_w11104_,
		_w11105_
	);
	LUT3 #(
		.INIT('hf9)
	) name5279 (
		_w10897_,
		_w10896_,
		_w10898_,
		_w11106_
	);
	LUT2 #(
		.INIT('h8)
	) name5280 (
		_w10894_,
		_w10895_,
		_w11107_
	);
	LUT2 #(
		.INIT('h4)
	) name5281 (
		_w11106_,
		_w11107_,
		_w11108_
	);
	LUT4 #(
		.INIT('h00e4)
	) name5282 (
		_w10893_,
		_w11099_,
		_w11105_,
		_w11108_,
		_w11109_
	);
	LUT2 #(
		.INIT('h9)
	) name5283 (
		\u2_L5_reg[17]/NET0131 ,
		_w11109_,
		_w11110_
	);
	LUT4 #(
		.INIT('haafb)
	) name5284 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11111_
	);
	LUT2 #(
		.INIT('h2)
	) name5285 (
		_w10967_,
		_w11111_,
		_w11112_
	);
	LUT3 #(
		.INIT('h20)
	) name5286 (
		_w10960_,
		_w10973_,
		_w11015_,
		_w11113_
	);
	LUT4 #(
		.INIT('h0080)
	) name5287 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11114_
	);
	LUT3 #(
		.INIT('h01)
	) name5288 (
		_w10960_,
		_w10977_,
		_w11114_,
		_w11115_
	);
	LUT3 #(
		.INIT('h0b)
	) name5289 (
		_w11112_,
		_w11113_,
		_w11115_,
		_w11116_
	);
	LUT3 #(
		.INIT('hac)
	) name5290 (
		_w10961_,
		_w10956_,
		_w10958_,
		_w11117_
	);
	LUT3 #(
		.INIT('h8c)
	) name5291 (
		_w10961_,
		_w10957_,
		_w10960_,
		_w11118_
	);
	LUT2 #(
		.INIT('h4)
	) name5292 (
		_w11117_,
		_w11118_,
		_w11119_
	);
	LUT2 #(
		.INIT('h9)
	) name5293 (
		_w10957_,
		_w10956_,
		_w11120_
	);
	LUT4 #(
		.INIT('h0700)
	) name5294 (
		_w10961_,
		_w10957_,
		_w10958_,
		_w10960_,
		_w11121_
	);
	LUT3 #(
		.INIT('h15)
	) name5295 (
		_w10967_,
		_w11120_,
		_w11121_,
		_w11122_
	);
	LUT4 #(
		.INIT('hd5fd)
	) name5296 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11123_
	);
	LUT4 #(
		.INIT('hef00)
	) name5297 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10967_,
		_w11124_
	);
	LUT4 #(
		.INIT('h3200)
	) name5298 (
		_w10960_,
		_w11114_,
		_w11123_,
		_w11124_,
		_w11125_
	);
	LUT4 #(
		.INIT('h00df)
	) name5299 (
		_w10982_,
		_w11119_,
		_w11122_,
		_w11125_,
		_w11126_
	);
	LUT3 #(
		.INIT('h56)
	) name5300 (
		\u2_L5_reg[1]/NET0131 ,
		_w11116_,
		_w11126_,
		_w11127_
	);
	LUT4 #(
		.INIT('h2c7f)
	) name5301 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11128_
	);
	LUT2 #(
		.INIT('h2)
	) name5302 (
		_w10996_,
		_w11128_,
		_w11129_
	);
	LUT4 #(
		.INIT('hf7dd)
	) name5303 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11130_
	);
	LUT2 #(
		.INIT('h1)
	) name5304 (
		_w10996_,
		_w11130_,
		_w11131_
	);
	LUT4 #(
		.INIT('h0084)
	) name5305 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11132_
	);
	LUT3 #(
		.INIT('h02)
	) name5306 (
		_w10990_,
		_w11091_,
		_w11132_,
		_w11133_
	);
	LUT3 #(
		.INIT('h10)
	) name5307 (
		_w11131_,
		_w11129_,
		_w11133_,
		_w11134_
	);
	LUT2 #(
		.INIT('h8)
	) name5308 (
		_w10991_,
		_w10994_,
		_w11135_
	);
	LUT3 #(
		.INIT('h31)
	) name5309 (
		_w10996_,
		_w10992_,
		_w10993_,
		_w11136_
	);
	LUT2 #(
		.INIT('h8)
	) name5310 (
		_w11135_,
		_w11136_,
		_w11137_
	);
	LUT4 #(
		.INIT('h00bf)
	) name5311 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10990_,
		_w11138_
	);
	LUT2 #(
		.INIT('h4)
	) name5312 (
		_w10996_,
		_w10994_,
		_w11139_
	);
	LUT4 #(
		.INIT('h1000)
	) name5313 (
		_w10996_,
		_w10991_,
		_w10992_,
		_w10994_,
		_w11140_
	);
	LUT4 #(
		.INIT('h0010)
	) name5314 (
		_w10996_,
		_w10991_,
		_w10993_,
		_w10994_,
		_w11141_
	);
	LUT3 #(
		.INIT('h10)
	) name5315 (
		_w11140_,
		_w11141_,
		_w11138_,
		_w11142_
	);
	LUT4 #(
		.INIT('hf757)
	) name5316 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11143_
	);
	LUT4 #(
		.INIT('h0009)
	) name5317 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11144_
	);
	LUT3 #(
		.INIT('h0d)
	) name5318 (
		_w10996_,
		_w11143_,
		_w11144_,
		_w11145_
	);
	LUT3 #(
		.INIT('h40)
	) name5319 (
		_w11137_,
		_w11142_,
		_w11145_,
		_w11146_
	);
	LUT4 #(
		.INIT('h0002)
	) name5320 (
		_w10996_,
		_w10991_,
		_w10992_,
		_w10993_,
		_w11147_
	);
	LUT3 #(
		.INIT('h07)
	) name5321 (
		_w11082_,
		_w11139_,
		_w11147_,
		_w11148_
	);
	LUT4 #(
		.INIT('ha955)
	) name5322 (
		\u2_L5_reg[21]/NET0131 ,
		_w11134_,
		_w11146_,
		_w11148_,
		_w11149_
	);
	LUT4 #(
		.INIT('h3ce4)
	) name5323 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11150_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name5324 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11151_
	);
	LUT4 #(
		.INIT('hbb7f)
	) name5325 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11152_
	);
	LUT4 #(
		.INIT('hd800)
	) name5326 (
		_w11047_,
		_w11150_,
		_w11151_,
		_w11152_,
		_w11153_
	);
	LUT2 #(
		.INIT('h2)
	) name5327 (
		_w11059_,
		_w11153_,
		_w11154_
	);
	LUT4 #(
		.INIT('hfe7d)
	) name5328 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11155_
	);
	LUT2 #(
		.INIT('h2)
	) name5329 (
		_w11047_,
		_w11155_,
		_w11156_
	);
	LUT3 #(
		.INIT('ha2)
	) name5330 (
		_w11047_,
		_w11049_,
		_w11051_,
		_w11157_
	);
	LUT4 #(
		.INIT('h2223)
	) name5331 (
		_w11047_,
		_w11048_,
		_w11049_,
		_w11050_,
		_w11158_
	);
	LUT2 #(
		.INIT('h4)
	) name5332 (
		_w11157_,
		_w11158_,
		_w11159_
	);
	LUT4 #(
		.INIT('h0010)
	) name5333 (
		_w11047_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11160_
	);
	LUT2 #(
		.INIT('h2)
	) name5334 (
		_w11047_,
		_w11051_,
		_w11161_
	);
	LUT3 #(
		.INIT('h08)
	) name5335 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11162_
	);
	LUT3 #(
		.INIT('h45)
	) name5336 (
		_w11160_,
		_w11161_,
		_w11162_,
		_w11163_
	);
	LUT4 #(
		.INIT('h0400)
	) name5337 (
		_w11047_,
		_w11048_,
		_w11049_,
		_w11050_,
		_w11164_
	);
	LUT2 #(
		.INIT('h1)
	) name5338 (
		_w11054_,
		_w11164_,
		_w11165_
	);
	LUT4 #(
		.INIT('hba00)
	) name5339 (
		_w11059_,
		_w11159_,
		_w11163_,
		_w11165_,
		_w11166_
	);
	LUT4 #(
		.INIT('h5655)
	) name5340 (
		\u2_L5_reg[25]/NET0131 ,
		_w11154_,
		_w11156_,
		_w11166_,
		_w11167_
	);
	LUT4 #(
		.INIT('hcfdf)
	) name5341 (
		_w10961_,
		_w10957_,
		_w10958_,
		_w10960_,
		_w11168_
	);
	LUT2 #(
		.INIT('h2)
	) name5342 (
		_w10956_,
		_w11168_,
		_w11169_
	);
	LUT4 #(
		.INIT('hff7d)
	) name5343 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11170_
	);
	LUT4 #(
		.INIT('h0100)
	) name5344 (
		_w10961_,
		_w10957_,
		_w10958_,
		_w10960_,
		_w11171_
	);
	LUT4 #(
		.INIT('h00d0)
	) name5345 (
		_w10961_,
		_w10957_,
		_w10958_,
		_w10960_,
		_w11172_
	);
	LUT4 #(
		.INIT('h1300)
	) name5346 (
		_w11120_,
		_w11171_,
		_w11172_,
		_w11170_,
		_w11173_
	);
	LUT3 #(
		.INIT('h8a)
	) name5347 (
		_w10967_,
		_w11169_,
		_w11173_,
		_w11174_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5348 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11175_
	);
	LUT4 #(
		.INIT('h0806)
	) name5349 (
		_w10961_,
		_w10957_,
		_w10956_,
		_w10958_,
		_w11176_
	);
	LUT4 #(
		.INIT('h5501)
	) name5350 (
		_w10960_,
		_w10967_,
		_w11175_,
		_w11176_,
		_w11177_
	);
	LUT2 #(
		.INIT('h4)
	) name5351 (
		_w10976_,
		_w11019_,
		_w11178_
	);
	LUT2 #(
		.INIT('h2)
	) name5352 (
		_w10971_,
		_w10980_,
		_w11179_
	);
	LUT3 #(
		.INIT('h01)
	) name5353 (
		_w10965_,
		_w10981_,
		_w10984_,
		_w11180_
	);
	LUT4 #(
		.INIT('h2322)
	) name5354 (
		_w10967_,
		_w11178_,
		_w11179_,
		_w11180_,
		_w11181_
	);
	LUT4 #(
		.INIT('h5655)
	) name5355 (
		\u2_L5_reg[26]/NET0131 ,
		_w11177_,
		_w11174_,
		_w11181_,
		_w11182_
	);
	LUT4 #(
		.INIT('hc693)
	) name5356 (
		decrypt_pad,
		\u2_R5_reg[8]/NET0131 ,
		\u2_uk_K_r5_reg[12]/NET0131 ,
		\u2_uk_K_r5_reg[34]/NET0131 ,
		_w11183_
	);
	LUT4 #(
		.INIT('hc693)
	) name5357 (
		decrypt_pad,
		\u2_R5_reg[4]/NET0131 ,
		\u2_uk_K_r5_reg[25]/NET0131 ,
		\u2_uk_K_r5_reg[47]/NET0131 ,
		_w11184_
	);
	LUT4 #(
		.INIT('hc693)
	) name5358 (
		decrypt_pad,
		\u2_R5_reg[9]/NET0131 ,
		\u2_uk_K_r5_reg[17]/NET0131 ,
		\u2_uk_K_r5_reg[39]/NET0131 ,
		_w11185_
	);
	LUT2 #(
		.INIT('h8)
	) name5359 (
		_w11184_,
		_w11185_,
		_w11186_
	);
	LUT4 #(
		.INIT('hc963)
	) name5360 (
		decrypt_pad,
		\u2_R5_reg[5]/NET0131 ,
		\u2_uk_K_r5_reg[26]/NET0131 ,
		\u2_uk_K_r5_reg[4]/NET0131 ,
		_w11187_
	);
	LUT4 #(
		.INIT('hc963)
	) name5361 (
		decrypt_pad,
		\u2_R5_reg[6]/NET0131 ,
		\u2_uk_K_r5_reg[17]/NET0131 ,
		\u2_uk_K_r5_reg[27]/NET0131 ,
		_w11188_
	);
	LUT4 #(
		.INIT('h0034)
	) name5362 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11189_
	);
	LUT4 #(
		.INIT('hc963)
	) name5363 (
		decrypt_pad,
		\u2_R5_reg[7]/NET0131 ,
		\u2_uk_K_r5_reg[11]/NET0131 ,
		\u2_uk_K_r5_reg[46]/NET0131 ,
		_w11190_
	);
	LUT2 #(
		.INIT('h8)
	) name5364 (
		_w11184_,
		_w11188_,
		_w11191_
	);
	LUT4 #(
		.INIT('h0800)
	) name5365 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11192_
	);
	LUT3 #(
		.INIT('h15)
	) name5366 (
		_w11189_,
		_w11190_,
		_w11192_,
		_w11193_
	);
	LUT2 #(
		.INIT('h2)
	) name5367 (
		_w11187_,
		_w11188_,
		_w11194_
	);
	LUT3 #(
		.INIT('h02)
	) name5368 (
		_w11185_,
		_w11188_,
		_w11190_,
		_w11195_
	);
	LUT3 #(
		.INIT('h40)
	) name5369 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11196_
	);
	LUT3 #(
		.INIT('h54)
	) name5370 (
		_w11194_,
		_w11195_,
		_w11196_,
		_w11197_
	);
	LUT3 #(
		.INIT('h09)
	) name5371 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11198_
	);
	LUT2 #(
		.INIT('h2)
	) name5372 (
		_w11184_,
		_w11188_,
		_w11199_
	);
	LUT2 #(
		.INIT('h1)
	) name5373 (
		_w11187_,
		_w11190_,
		_w11200_
	);
	LUT2 #(
		.INIT('h2)
	) name5374 (
		_w11184_,
		_w11190_,
		_w11201_
	);
	LUT4 #(
		.INIT('h00b1)
	) name5375 (
		_w11184_,
		_w11187_,
		_w11188_,
		_w11190_,
		_w11202_
	);
	LUT2 #(
		.INIT('h4)
	) name5376 (
		_w11198_,
		_w11202_,
		_w11203_
	);
	LUT4 #(
		.INIT('h5455)
	) name5377 (
		_w11183_,
		_w11197_,
		_w11203_,
		_w11193_,
		_w11204_
	);
	LUT4 #(
		.INIT('he6ee)
	) name5378 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11205_
	);
	LUT4 #(
		.INIT('h4044)
	) name5379 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11206_
	);
	LUT3 #(
		.INIT('h0d)
	) name5380 (
		_w11187_,
		_w11188_,
		_w11190_,
		_w11207_
	);
	LUT4 #(
		.INIT('hf200)
	) name5381 (
		_w11183_,
		_w11205_,
		_w11206_,
		_w11207_,
		_w11208_
	);
	LUT4 #(
		.INIT('h0100)
	) name5382 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11209_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name5383 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11210_
	);
	LUT2 #(
		.INIT('h2)
	) name5384 (
		_w11190_,
		_w11210_,
		_w11211_
	);
	LUT4 #(
		.INIT('h0080)
	) name5385 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11212_
	);
	LUT4 #(
		.INIT('h0002)
	) name5386 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11213_
	);
	LUT4 #(
		.INIT('h8c00)
	) name5387 (
		_w11184_,
		_w11187_,
		_w11188_,
		_w11190_,
		_w11214_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5388 (
		_w11183_,
		_w11213_,
		_w11214_,
		_w11212_,
		_w11215_
	);
	LUT3 #(
		.INIT('h01)
	) name5389 (
		_w11211_,
		_w11215_,
		_w11208_,
		_w11216_
	);
	LUT3 #(
		.INIT('h65)
	) name5390 (
		\u2_L5_reg[2]/NET0131 ,
		_w11204_,
		_w11216_,
		_w11217_
	);
	LUT4 #(
		.INIT('h67dc)
	) name5391 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11218_
	);
	LUT4 #(
		.INIT('hd2f7)
	) name5392 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11219_
	);
	LUT4 #(
		.INIT('h0040)
	) name5393 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11220_
	);
	LUT4 #(
		.INIT('h00d8)
	) name5394 (
		_w10929_,
		_w11218_,
		_w11219_,
		_w11220_,
		_w11221_
	);
	LUT4 #(
		.INIT('h9aff)
	) name5395 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11222_
	);
	LUT4 #(
		.INIT('haa02)
	) name5396 (
		_w10929_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11223_
	);
	LUT4 #(
		.INIT('h9297)
	) name5397 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11224_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name5398 (
		_w10929_,
		_w11222_,
		_w11223_,
		_w11224_,
		_w11225_
	);
	LUT4 #(
		.INIT('h0800)
	) name5399 (
		_w10929_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11226_
	);
	LUT2 #(
		.INIT('h1)
	) name5400 (
		_w10941_,
		_w11226_,
		_w11227_
	);
	LUT4 #(
		.INIT('hd800)
	) name5401 (
		_w10925_,
		_w11225_,
		_w11221_,
		_w11227_,
		_w11228_
	);
	LUT2 #(
		.INIT('h6)
	) name5402 (
		\u2_L5_reg[29]/NET0131 ,
		_w11228_,
		_w11229_
	);
	LUT4 #(
		.INIT('h2000)
	) name5403 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11230_
	);
	LUT4 #(
		.INIT('hdaff)
	) name5404 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11231_
	);
	LUT2 #(
		.INIT('h1)
	) name5405 (
		_w11190_,
		_w11231_,
		_w11232_
	);
	LUT4 #(
		.INIT('h2900)
	) name5406 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11233_
	);
	LUT3 #(
		.INIT('h51)
	) name5407 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11234_
	);
	LUT4 #(
		.INIT('h0b08)
	) name5408 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11235_
	);
	LUT3 #(
		.INIT('h01)
	) name5409 (
		_w11190_,
		_w11234_,
		_w11235_,
		_w11236_
	);
	LUT4 #(
		.INIT('h4051)
	) name5410 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11237_
	);
	LUT3 #(
		.INIT('h15)
	) name5411 (
		_w11183_,
		_w11190_,
		_w11237_,
		_w11238_
	);
	LUT3 #(
		.INIT('h10)
	) name5412 (
		_w11236_,
		_w11233_,
		_w11238_,
		_w11239_
	);
	LUT3 #(
		.INIT('h0d)
	) name5413 (
		_w11185_,
		_w11187_,
		_w11190_,
		_w11240_
	);
	LUT4 #(
		.INIT('h0400)
	) name5414 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11241_
	);
	LUT4 #(
		.INIT('h0a02)
	) name5415 (
		_w11183_,
		_w11199_,
		_w11241_,
		_w11240_,
		_w11242_
	);
	LUT4 #(
		.INIT('h283c)
	) name5416 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11243_
	);
	LUT3 #(
		.INIT('h45)
	) name5417 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11244_
	);
	LUT4 #(
		.INIT('hbbb1)
	) name5418 (
		_w11190_,
		_w11237_,
		_w11244_,
		_w11243_,
		_w11245_
	);
	LUT2 #(
		.INIT('h8)
	) name5419 (
		_w11242_,
		_w11245_,
		_w11246_
	);
	LUT4 #(
		.INIT('h6665)
	) name5420 (
		\u2_L5_reg[28]/NET0131 ,
		_w11232_,
		_w11239_,
		_w11246_,
		_w11247_
	);
	LUT4 #(
		.INIT('hd97b)
	) name5421 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11248_
	);
	LUT2 #(
		.INIT('h2)
	) name5422 (
		_w10929_,
		_w11248_,
		_w11249_
	);
	LUT4 #(
		.INIT('heebf)
	) name5423 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11250_
	);
	LUT4 #(
		.INIT('h0040)
	) name5424 (
		_w10929_,
		_w10926_,
		_w10931_,
		_w10927_,
		_w11251_
	);
	LUT4 #(
		.INIT('h0032)
	) name5425 (
		_w10929_,
		_w10941_,
		_w11250_,
		_w11251_,
		_w11252_
	);
	LUT3 #(
		.INIT('h45)
	) name5426 (
		_w10925_,
		_w11249_,
		_w11252_,
		_w11253_
	);
	LUT4 #(
		.INIT('h7c7f)
	) name5427 (
		_w10929_,
		_w10926_,
		_w10931_,
		_w10928_,
		_w11254_
	);
	LUT2 #(
		.INIT('h1)
	) name5428 (
		_w10927_,
		_w11254_,
		_w11255_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name5429 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11256_
	);
	LUT3 #(
		.INIT('h80)
	) name5430 (
		_w10931_,
		_w10927_,
		_w10928_,
		_w11257_
	);
	LUT3 #(
		.INIT('h0e)
	) name5431 (
		_w10929_,
		_w11256_,
		_w11257_,
		_w11258_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5432 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11259_
	);
	LUT4 #(
		.INIT('h5501)
	) name5433 (
		_w10929_,
		_w10926_,
		_w10931_,
		_w10927_,
		_w11260_
	);
	LUT3 #(
		.INIT('h9e)
	) name5434 (
		_w10926_,
		_w10931_,
		_w10928_,
		_w11261_
	);
	LUT2 #(
		.INIT('h8)
	) name5435 (
		_w10929_,
		_w10927_,
		_w11262_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5436 (
		_w11259_,
		_w11260_,
		_w11261_,
		_w11262_,
		_w11263_
	);
	LUT4 #(
		.INIT('h7500)
	) name5437 (
		_w10925_,
		_w11255_,
		_w11258_,
		_w11263_,
		_w11264_
	);
	LUT3 #(
		.INIT('h65)
	) name5438 (
		\u2_L5_reg[4]/NET0131 ,
		_w11253_,
		_w11264_,
		_w11265_
	);
	LUT3 #(
		.INIT('h40)
	) name5439 (
		_w11184_,
		_w11185_,
		_w11188_,
		_w11266_
	);
	LUT3 #(
		.INIT('h01)
	) name5440 (
		_w11185_,
		_w11187_,
		_w11188_,
		_w11267_
	);
	LUT4 #(
		.INIT('heee4)
	) name5441 (
		_w11190_,
		_w11235_,
		_w11267_,
		_w11266_,
		_w11268_
	);
	LUT4 #(
		.INIT('hdf6f)
	) name5442 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11269_
	);
	LUT4 #(
		.INIT('hab00)
	) name5443 (
		_w11194_,
		_w11195_,
		_w11196_,
		_w11269_,
		_w11270_
	);
	LUT3 #(
		.INIT('h8a)
	) name5444 (
		_w11183_,
		_w11268_,
		_w11270_,
		_w11271_
	);
	LUT4 #(
		.INIT('hf6d6)
	) name5445 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11272_
	);
	LUT2 #(
		.INIT('h2)
	) name5446 (
		_w11190_,
		_w11272_,
		_w11273_
	);
	LUT3 #(
		.INIT('hb0)
	) name5447 (
		_w11185_,
		_w11187_,
		_w11190_,
		_w11274_
	);
	LUT3 #(
		.INIT('h04)
	) name5448 (
		_w11184_,
		_w11185_,
		_w11188_,
		_w11275_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name5449 (
		_w11191_,
		_w11200_,
		_w11274_,
		_w11275_,
		_w11276_
	);
	LUT4 #(
		.INIT('hebed)
	) name5450 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11277_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name5451 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11278_
	);
	LUT4 #(
		.INIT('h0133)
	) name5452 (
		_w11183_,
		_w11190_,
		_w11277_,
		_w11278_,
		_w11279_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5453 (
		_w11183_,
		_w11273_,
		_w11276_,
		_w11279_,
		_w11280_
	);
	LUT3 #(
		.INIT('h9a)
	) name5454 (
		\u2_L5_reg[13]/NET0131 ,
		_w11271_,
		_w11280_,
		_w11281_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name5455 (
		_w10929_,
		_w10926_,
		_w10931_,
		_w10927_,
		_w11282_
	);
	LUT4 #(
		.INIT('hef00)
	) name5456 (
		_w10931_,
		_w10927_,
		_w10928_,
		_w10925_,
		_w11283_
	);
	LUT3 #(
		.INIT('he0)
	) name5457 (
		_w10928_,
		_w11282_,
		_w11283_,
		_w11284_
	);
	LUT4 #(
		.INIT('h4010)
	) name5458 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11285_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name5459 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11286_
	);
	LUT3 #(
		.INIT('h31)
	) name5460 (
		_w10929_,
		_w11285_,
		_w11286_,
		_w11287_
	);
	LUT4 #(
		.INIT('h4e55)
	) name5461 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11288_
	);
	LUT2 #(
		.INIT('h2)
	) name5462 (
		_w10929_,
		_w11288_,
		_w11289_
	);
	LUT4 #(
		.INIT('h1001)
	) name5463 (
		_w10929_,
		_w10926_,
		_w10931_,
		_w10928_,
		_w11290_
	);
	LUT4 #(
		.INIT('h8000)
	) name5464 (
		_w10926_,
		_w10931_,
		_w10927_,
		_w10928_,
		_w11291_
	);
	LUT3 #(
		.INIT('h01)
	) name5465 (
		_w10925_,
		_w11291_,
		_w11290_,
		_w11292_
	);
	LUT4 #(
		.INIT('h7077)
	) name5466 (
		_w11284_,
		_w11287_,
		_w11289_,
		_w11292_,
		_w11293_
	);
	LUT2 #(
		.INIT('h4)
	) name5467 (
		_w10928_,
		_w11251_,
		_w11294_
	);
	LUT2 #(
		.INIT('h1)
	) name5468 (
		_w10949_,
		_w11294_,
		_w11295_
	);
	LUT3 #(
		.INIT('h65)
	) name5469 (
		\u2_L5_reg[19]/NET0131 ,
		_w11293_,
		_w11295_,
		_w11296_
	);
	LUT4 #(
		.INIT('hfdc3)
	) name5470 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11297_
	);
	LUT4 #(
		.INIT('h7bff)
	) name5471 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11298_
	);
	LUT4 #(
		.INIT('h0233)
	) name5472 (
		_w10893_,
		_w10894_,
		_w11297_,
		_w11298_,
		_w11299_
	);
	LUT3 #(
		.INIT('h8a)
	) name5473 (
		_w10894_,
		_w10897_,
		_w10898_,
		_w11300_
	);
	LUT2 #(
		.INIT('h8)
	) name5474 (
		_w10912_,
		_w11300_,
		_w11301_
	);
	LUT3 #(
		.INIT('h07)
	) name5475 (
		_w10913_,
		_w10921_,
		_w11100_,
		_w11302_
	);
	LUT3 #(
		.INIT('h8a)
	) name5476 (
		_w10893_,
		_w11301_,
		_w11302_,
		_w11303_
	);
	LUT4 #(
		.INIT('h88a2)
	) name5477 (
		_w10894_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11304_
	);
	LUT4 #(
		.INIT('h5545)
	) name5478 (
		_w10894_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11305_
	);
	LUT3 #(
		.INIT('h01)
	) name5479 (
		_w10897_,
		_w11305_,
		_w11304_,
		_w11306_
	);
	LUT4 #(
		.INIT('h5400)
	) name5480 (
		_w10894_,
		_w10897_,
		_w10895_,
		_w10898_,
		_w11307_
	);
	LUT3 #(
		.INIT('h32)
	) name5481 (
		_w10921_,
		_w10905_,
		_w11307_,
		_w11308_
	);
	LUT3 #(
		.INIT('h01)
	) name5482 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w11309_
	);
	LUT4 #(
		.INIT('h0080)
	) name5483 (
		_w10894_,
		_w10897_,
		_w10896_,
		_w10898_,
		_w11310_
	);
	LUT3 #(
		.INIT('h01)
	) name5484 (
		_w10917_,
		_w11310_,
		_w11309_,
		_w11311_
	);
	LUT4 #(
		.INIT('h2322)
	) name5485 (
		_w10893_,
		_w11306_,
		_w11308_,
		_w11311_,
		_w11312_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5486 (
		\u2_L5_reg[23]/NET0131 ,
		_w11303_,
		_w11299_,
		_w11312_,
		_w11313_
	);
	LUT4 #(
		.INIT('h0e5e)
	) name5487 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11314_
	);
	LUT3 #(
		.INIT('h15)
	) name5488 (
		_w10996_,
		_w10991_,
		_w10994_,
		_w11315_
	);
	LUT2 #(
		.INIT('h4)
	) name5489 (
		_w11314_,
		_w11315_,
		_w11316_
	);
	LUT3 #(
		.INIT('ha2)
	) name5490 (
		_w10996_,
		_w10991_,
		_w10994_,
		_w11317_
	);
	LUT4 #(
		.INIT('hbcf7)
	) name5491 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11318_
	);
	LUT3 #(
		.INIT('hb0)
	) name5492 (
		_w11077_,
		_w11317_,
		_w11318_,
		_w11319_
	);
	LUT3 #(
		.INIT('h8a)
	) name5493 (
		_w10990_,
		_w11316_,
		_w11319_,
		_w11320_
	);
	LUT4 #(
		.INIT('hcf40)
	) name5494 (
		_w10991_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11321_
	);
	LUT4 #(
		.INIT('haa8a)
	) name5495 (
		_w10996_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11322_
	);
	LUT2 #(
		.INIT('h4)
	) name5496 (
		_w11321_,
		_w11322_,
		_w11323_
	);
	LUT4 #(
		.INIT('h4000)
	) name5497 (
		_w10996_,
		_w10991_,
		_w10992_,
		_w10994_,
		_w11324_
	);
	LUT3 #(
		.INIT('h01)
	) name5498 (
		_w11009_,
		_w11141_,
		_w11324_,
		_w11325_
	);
	LUT4 #(
		.INIT('h0008)
	) name5499 (
		_w10996_,
		_w10992_,
		_w10993_,
		_w10994_,
		_w11326_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5500 (
		_w10996_,
		_w10997_,
		_w11007_,
		_w11326_,
		_w11327_
	);
	LUT4 #(
		.INIT('hba00)
	) name5501 (
		_w10990_,
		_w11323_,
		_w11325_,
		_w11327_,
		_w11328_
	);
	LUT3 #(
		.INIT('h65)
	) name5502 (
		\u2_L5_reg[27]/NET0131 ,
		_w11320_,
		_w11328_,
		_w11329_
	);
	LUT3 #(
		.INIT('h20)
	) name5503 (
		_w10868_,
		_w10870_,
		_w10869_,
		_w11330_
	);
	LUT4 #(
		.INIT('h2000)
	) name5504 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11331_
	);
	LUT4 #(
		.INIT('hdeb9)
	) name5505 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11332_
	);
	LUT2 #(
		.INIT('h1)
	) name5506 (
		_w10866_,
		_w11332_,
		_w11333_
	);
	LUT3 #(
		.INIT('h08)
	) name5507 (
		_w10868_,
		_w10867_,
		_w10869_,
		_w11334_
	);
	LUT4 #(
		.INIT('hf3ee)
	) name5508 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11335_
	);
	LUT4 #(
		.INIT('h1f13)
	) name5509 (
		_w10870_,
		_w10866_,
		_w11334_,
		_w11335_,
		_w11336_
	);
	LUT3 #(
		.INIT('h8a)
	) name5510 (
		_w10865_,
		_w11333_,
		_w11336_,
		_w11337_
	);
	LUT4 #(
		.INIT('h6fb7)
	) name5511 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11338_
	);
	LUT4 #(
		.INIT('h4547)
	) name5512 (
		_w10866_,
		_w10876_,
		_w11043_,
		_w11330_,
		_w11339_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name5513 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11340_
	);
	LUT3 #(
		.INIT('h72)
	) name5514 (
		_w10866_,
		_w10882_,
		_w11340_,
		_w11341_
	);
	LUT4 #(
		.INIT('hea00)
	) name5515 (
		_w10865_,
		_w11338_,
		_w11339_,
		_w11341_,
		_w11342_
	);
	LUT3 #(
		.INIT('h65)
	) name5516 (
		\u2_L5_reg[32]/NET0131 ,
		_w11337_,
		_w11342_,
		_w11343_
	);
	LUT4 #(
		.INIT('hc963)
	) name5517 (
		decrypt_pad,
		\u2_R5_reg[12]/NET0131 ,
		\u2_uk_K_r5_reg[12]/NET0131 ,
		\u2_uk_K_r5_reg[47]/NET0131 ,
		_w11344_
	);
	LUT4 #(
		.INIT('hc963)
	) name5518 (
		decrypt_pad,
		\u2_R5_reg[13]/NET0131 ,
		\u2_uk_K_r5_reg[25]/NET0131 ,
		\u2_uk_K_r5_reg[3]/NET0131 ,
		_w11345_
	);
	LUT4 #(
		.INIT('hc693)
	) name5519 (
		decrypt_pad,
		\u2_R5_reg[8]/NET0131 ,
		\u2_uk_K_r5_reg[26]/NET0131 ,
		\u2_uk_K_r5_reg[48]/NET0131 ,
		_w11346_
	);
	LUT2 #(
		.INIT('h6)
	) name5520 (
		_w11345_,
		_w11346_,
		_w11347_
	);
	LUT4 #(
		.INIT('hc963)
	) name5521 (
		decrypt_pad,
		\u2_R5_reg[9]/NET0131 ,
		\u2_uk_K_r5_reg[20]/NET0131 ,
		\u2_uk_K_r5_reg[55]/NET0131 ,
		_w11348_
	);
	LUT4 #(
		.INIT('hc963)
	) name5522 (
		decrypt_pad,
		\u2_R5_reg[10]/NET0131 ,
		\u2_uk_K_r5_reg[53]/NET0131 ,
		\u2_uk_K_r5_reg[6]/NET0131 ,
		_w11349_
	);
	LUT4 #(
		.INIT('h2100)
	) name5523 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11350_
	);
	LUT3 #(
		.INIT('h08)
	) name5524 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11351_
	);
	LUT4 #(
		.INIT('hc693)
	) name5525 (
		decrypt_pad,
		\u2_R5_reg[11]/NET0131 ,
		\u2_uk_K_r5_reg[32]/NET0131 ,
		\u2_uk_K_r5_reg[54]/NET0131 ,
		_w11352_
	);
	LUT2 #(
		.INIT('h2)
	) name5526 (
		_w11349_,
		_w11352_,
		_w11353_
	);
	LUT3 #(
		.INIT('h40)
	) name5527 (
		_w11345_,
		_w11348_,
		_w11349_,
		_w11354_
	);
	LUT4 #(
		.INIT('h4000)
	) name5528 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11355_
	);
	LUT4 #(
		.INIT('h0007)
	) name5529 (
		_w11351_,
		_w11353_,
		_w11355_,
		_w11350_,
		_w11356_
	);
	LUT2 #(
		.INIT('h8)
	) name5530 (
		_w11345_,
		_w11352_,
		_w11357_
	);
	LUT3 #(
		.INIT('h46)
	) name5531 (
		_w11345_,
		_w11346_,
		_w11352_,
		_w11358_
	);
	LUT2 #(
		.INIT('h1)
	) name5532 (
		_w11348_,
		_w11349_,
		_w11359_
	);
	LUT2 #(
		.INIT('h8)
	) name5533 (
		_w11359_,
		_w11358_,
		_w11360_
	);
	LUT3 #(
		.INIT('hed)
	) name5534 (
		_w11348_,
		_w11349_,
		_w11358_,
		_w11361_
	);
	LUT3 #(
		.INIT('h15)
	) name5535 (
		_w11344_,
		_w11356_,
		_w11361_,
		_w11362_
	);
	LUT4 #(
		.INIT('h959d)
	) name5536 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11363_
	);
	LUT4 #(
		.INIT('h0001)
	) name5537 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11364_
	);
	LUT4 #(
		.INIT('hddfe)
	) name5538 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11365_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5539 (
		_w11363_,
		_w11344_,
		_w11365_,
		_w11352_,
		_w11366_
	);
	LUT2 #(
		.INIT('h8)
	) name5540 (
		_w11349_,
		_w11344_,
		_w11367_
	);
	LUT3 #(
		.INIT('h04)
	) name5541 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11368_
	);
	LUT2 #(
		.INIT('h2)
	) name5542 (
		_w11344_,
		_w11352_,
		_w11369_
	);
	LUT3 #(
		.INIT('h80)
	) name5543 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11370_
	);
	LUT4 #(
		.INIT('h6f67)
	) name5544 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11371_
	);
	LUT4 #(
		.INIT('h7707)
	) name5545 (
		_w11367_,
		_w11368_,
		_w11369_,
		_w11371_,
		_w11372_
	);
	LUT2 #(
		.INIT('h4)
	) name5546 (
		_w11366_,
		_w11372_,
		_w11373_
	);
	LUT3 #(
		.INIT('h65)
	) name5547 (
		\u2_L5_reg[6]/NET0131 ,
		_w11362_,
		_w11373_,
		_w11374_
	);
	LUT4 #(
		.INIT('h0a04)
	) name5548 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11375_
	);
	LUT3 #(
		.INIT('h48)
	) name5549 (
		_w10868_,
		_w10870_,
		_w10869_,
		_w11376_
	);
	LUT4 #(
		.INIT('h4080)
	) name5550 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11377_
	);
	LUT4 #(
		.INIT('h0010)
	) name5551 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11378_
	);
	LUT2 #(
		.INIT('h4)
	) name5552 (
		_w10865_,
		_w10866_,
		_w11379_
	);
	LUT2 #(
		.INIT('h2)
	) name5553 (
		_w10865_,
		_w10866_,
		_w11380_
	);
	LUT2 #(
		.INIT('h9)
	) name5554 (
		_w10865_,
		_w10866_,
		_w11381_
	);
	LUT4 #(
		.INIT('h0100)
	) name5555 (
		_w11378_,
		_w11377_,
		_w11375_,
		_w11381_,
		_w11382_
	);
	LUT3 #(
		.INIT('h41)
	) name5556 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w11383_
	);
	LUT4 #(
		.INIT('h0004)
	) name5557 (
		_w11334_,
		_w11380_,
		_w11376_,
		_w11383_,
		_w11384_
	);
	LUT4 #(
		.INIT('h957a)
	) name5558 (
		_w10868_,
		_w10870_,
		_w10867_,
		_w10869_,
		_w11385_
	);
	LUT3 #(
		.INIT('h04)
	) name5559 (
		_w11378_,
		_w11379_,
		_w11385_,
		_w11386_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5560 (
		_w11331_,
		_w11382_,
		_w11384_,
		_w11386_,
		_w11387_
	);
	LUT2 #(
		.INIT('h6)
	) name5561 (
		\u2_L5_reg[7]/NET0131 ,
		_w11387_,
		_w11388_
	);
	LUT4 #(
		.INIT('h3fef)
	) name5562 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11389_
	);
	LUT4 #(
		.INIT('hc2ff)
	) name5563 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11390_
	);
	LUT4 #(
		.INIT('hfb79)
	) name5564 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11391_
	);
	LUT4 #(
		.INIT('hd800)
	) name5565 (
		_w11047_,
		_w11389_,
		_w11390_,
		_w11391_,
		_w11392_
	);
	LUT4 #(
		.INIT('h0001)
	) name5566 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11393_
	);
	LUT4 #(
		.INIT('hcffe)
	) name5567 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11394_
	);
	LUT3 #(
		.INIT('h10)
	) name5568 (
		_w11047_,
		_w11048_,
		_w11050_,
		_w11395_
	);
	LUT4 #(
		.INIT('h00c4)
	) name5569 (
		_w11047_,
		_w11074_,
		_w11394_,
		_w11395_,
		_w11396_
	);
	LUT4 #(
		.INIT('hf977)
	) name5570 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11397_
	);
	LUT4 #(
		.INIT('hbf15)
	) name5571 (
		_w11047_,
		_w11048_,
		_w11052_,
		_w11397_,
		_w11398_
	);
	LUT4 #(
		.INIT('hd800)
	) name5572 (
		_w11059_,
		_w11396_,
		_w11392_,
		_w11398_,
		_w11399_
	);
	LUT2 #(
		.INIT('h9)
	) name5573 (
		\u2_L5_reg[8]/NET0131 ,
		_w11399_,
		_w11400_
	);
	LUT4 #(
		.INIT('hf700)
	) name5574 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11401_
	);
	LUT4 #(
		.INIT('h0400)
	) name5575 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11352_,
		_w11402_
	);
	LUT4 #(
		.INIT('h006d)
	) name5576 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11403_
	);
	LUT3 #(
		.INIT('h45)
	) name5577 (
		_w11401_,
		_w11402_,
		_w11403_,
		_w11404_
	);
	LUT4 #(
		.INIT('h0100)
	) name5578 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11405_
	);
	LUT3 #(
		.INIT('h14)
	) name5579 (
		_w11345_,
		_w11346_,
		_w11349_,
		_w11406_
	);
	LUT4 #(
		.INIT('hfd00)
	) name5580 (
		_w11352_,
		_w11355_,
		_w11405_,
		_w11406_,
		_w11407_
	);
	LUT3 #(
		.INIT('ha8)
	) name5581 (
		_w11344_,
		_w11404_,
		_w11407_,
		_w11408_
	);
	LUT3 #(
		.INIT('h40)
	) name5582 (
		_w11348_,
		_w11346_,
		_w11349_,
		_w11409_
	);
	LUT4 #(
		.INIT('h00bf)
	) name5583 (
		_w11348_,
		_w11346_,
		_w11349_,
		_w11352_,
		_w11410_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5584 (
		_w11352_,
		_w11355_,
		_w11405_,
		_w11410_,
		_w11411_
	);
	LUT4 #(
		.INIT('h7d78)
	) name5585 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11412_
	);
	LUT3 #(
		.INIT('he0)
	) name5586 (
		_w11345_,
		_w11346_,
		_w11352_,
		_w11413_
	);
	LUT4 #(
		.INIT('h6800)
	) name5587 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11352_,
		_w11414_
	);
	LUT4 #(
		.INIT('h0504)
	) name5588 (
		_w11364_,
		_w11352_,
		_w11414_,
		_w11412_,
		_w11415_
	);
	LUT3 #(
		.INIT('h32)
	) name5589 (
		_w11344_,
		_w11411_,
		_w11415_,
		_w11416_
	);
	LUT3 #(
		.INIT('h65)
	) name5590 (
		\u2_L5_reg[16]/NET0131 ,
		_w11408_,
		_w11416_,
		_w11417_
	);
	LUT2 #(
		.INIT('h4)
	) name5591 (
		_w11349_,
		_w11352_,
		_w11418_
	);
	LUT3 #(
		.INIT('h31)
	) name5592 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11419_
	);
	LUT2 #(
		.INIT('h8)
	) name5593 (
		_w11418_,
		_w11419_,
		_w11420_
	);
	LUT3 #(
		.INIT('h0e)
	) name5594 (
		_w11348_,
		_w11349_,
		_w11352_,
		_w11421_
	);
	LUT3 #(
		.INIT('hb0)
	) name5595 (
		_w11348_,
		_w11346_,
		_w11349_,
		_w11422_
	);
	LUT4 #(
		.INIT('h23af)
	) name5596 (
		_w11347_,
		_w11413_,
		_w11421_,
		_w11422_,
		_w11423_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5597 (
		_w11344_,
		_w11360_,
		_w11420_,
		_w11423_,
		_w11424_
	);
	LUT4 #(
		.INIT('hcaf1)
	) name5598 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11425_
	);
	LUT4 #(
		.INIT('h1000)
	) name5599 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11426_
	);
	LUT4 #(
		.INIT('h5504)
	) name5600 (
		_w11344_,
		_w11352_,
		_w11425_,
		_w11426_,
		_w11427_
	);
	LUT4 #(
		.INIT('h0021)
	) name5601 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11428_
	);
	LUT4 #(
		.INIT('hb59e)
	) name5602 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11429_
	);
	LUT2 #(
		.INIT('h1)
	) name5603 (
		_w11344_,
		_w11352_,
		_w11430_
	);
	LUT2 #(
		.INIT('h4)
	) name5604 (
		_w11429_,
		_w11430_,
		_w11431_
	);
	LUT3 #(
		.INIT('he7)
	) name5605 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11432_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name5606 (
		_w11349_,
		_w11352_,
		_w11370_,
		_w11432_,
		_w11433_
	);
	LUT3 #(
		.INIT('h10)
	) name5607 (
		_w11427_,
		_w11431_,
		_w11433_,
		_w11434_
	);
	LUT3 #(
		.INIT('h65)
	) name5608 (
		\u2_L5_reg[24]/NET0131 ,
		_w11424_,
		_w11434_,
		_w11435_
	);
	LUT4 #(
		.INIT('hfae5)
	) name5609 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11436_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name5610 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11437_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name5611 (
		_w11344_,
		_w11354_,
		_w11436_,
		_w11437_,
		_w11438_
	);
	LUT2 #(
		.INIT('h2)
	) name5612 (
		_w11352_,
		_w11438_,
		_w11439_
	);
	LUT4 #(
		.INIT('h0200)
	) name5613 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11440_
	);
	LUT3 #(
		.INIT('h0e)
	) name5614 (
		_w11348_,
		_w11346_,
		_w11352_,
		_w11441_
	);
	LUT4 #(
		.INIT('h0015)
	) name5615 (
		_w11428_,
		_w11437_,
		_w11441_,
		_w11440_,
		_w11442_
	);
	LUT2 #(
		.INIT('h1)
	) name5616 (
		_w11344_,
		_w11442_,
		_w11443_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name5617 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11349_,
		_w11444_
	);
	LUT2 #(
		.INIT('h2)
	) name5618 (
		_w11369_,
		_w11444_,
		_w11445_
	);
	LUT3 #(
		.INIT('h4c)
	) name5619 (
		_w11345_,
		_w11348_,
		_w11346_,
		_w11446_
	);
	LUT2 #(
		.INIT('h8)
	) name5620 (
		_w11367_,
		_w11446_,
		_w11447_
	);
	LUT4 #(
		.INIT('h0040)
	) name5621 (
		_w11345_,
		_w11348_,
		_w11349_,
		_w11352_,
		_w11448_
	);
	LUT3 #(
		.INIT('h07)
	) name5622 (
		_w11357_,
		_w11409_,
		_w11448_,
		_w11449_
	);
	LUT3 #(
		.INIT('h10)
	) name5623 (
		_w11445_,
		_w11447_,
		_w11449_,
		_w11450_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5624 (
		\u2_L5_reg[30]/NET0131 ,
		_w11439_,
		_w11443_,
		_w11450_,
		_w11451_
	);
	LUT4 #(
		.INIT('hfa3f)
	) name5625 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11452_
	);
	LUT2 #(
		.INIT('h2)
	) name5626 (
		_w11047_,
		_w11452_,
		_w11453_
	);
	LUT3 #(
		.INIT('ha2)
	) name5627 (
		_w11047_,
		_w11048_,
		_w11049_,
		_w11454_
	);
	LUT4 #(
		.INIT('h45f0)
	) name5628 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11455_
	);
	LUT3 #(
		.INIT('h54)
	) name5629 (
		_w11059_,
		_w11454_,
		_w11455_,
		_w11456_
	);
	LUT3 #(
		.INIT('h8c)
	) name5630 (
		_w11048_,
		_w11050_,
		_w11051_,
		_w11457_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5631 (
		_w11047_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11458_
	);
	LUT2 #(
		.INIT('h4)
	) name5632 (
		_w11457_,
		_w11458_,
		_w11459_
	);
	LUT4 #(
		.INIT('h0400)
	) name5633 (
		_w11047_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11460_
	);
	LUT4 #(
		.INIT('h0020)
	) name5634 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11461_
	);
	LUT4 #(
		.INIT('h0004)
	) name5635 (
		_w11054_,
		_w11059_,
		_w11461_,
		_w11460_,
		_w11462_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5636 (
		_w11453_,
		_w11456_,
		_w11459_,
		_w11462_,
		_w11463_
	);
	LUT4 #(
		.INIT('h2000)
	) name5637 (
		_w11048_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11464_
	);
	LUT4 #(
		.INIT('h0001)
	) name5638 (
		_w11047_,
		_w11071_,
		_w11393_,
		_w11464_,
		_w11465_
	);
	LUT3 #(
		.INIT('h02)
	) name5639 (
		_w11047_,
		_w11053_,
		_w11073_,
		_w11466_
	);
	LUT2 #(
		.INIT('h1)
	) name5640 (
		_w11465_,
		_w11466_,
		_w11467_
	);
	LUT3 #(
		.INIT('h56)
	) name5641 (
		\u2_L5_reg[3]/NET0131 ,
		_w11463_,
		_w11467_,
		_w11468_
	);
	LUT3 #(
		.INIT('he6)
	) name5642 (
		_w10895_,
		_w10896_,
		_w10898_,
		_w11469_
	);
	LUT4 #(
		.INIT('h5414)
	) name5643 (
		_w10894_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11470_
	);
	LUT4 #(
		.INIT('h080c)
	) name5644 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11471_
	);
	LUT4 #(
		.INIT('h9ffd)
	) name5645 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11472_
	);
	LUT4 #(
		.INIT('hce00)
	) name5646 (
		_w11096_,
		_w11470_,
		_w11471_,
		_w11472_,
		_w11473_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name5647 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11474_
	);
	LUT2 #(
		.INIT('h1)
	) name5648 (
		_w10894_,
		_w11474_,
		_w11475_
	);
	LUT4 #(
		.INIT('h8228)
	) name5649 (
		_w10897_,
		_w10895_,
		_w10896_,
		_w10898_,
		_w11476_
	);
	LUT4 #(
		.INIT('h0031)
	) name5650 (
		_w10902_,
		_w11103_,
		_w11469_,
		_w11476_,
		_w11477_
	);
	LUT4 #(
		.INIT('h3120)
	) name5651 (
		_w10893_,
		_w11475_,
		_w11477_,
		_w11473_,
		_w11478_
	);
	LUT2 #(
		.INIT('h9)
	) name5652 (
		\u2_L5_reg[9]/NET0131 ,
		_w11478_,
		_w11479_
	);
	LUT4 #(
		.INIT('h0a20)
	) name5653 (
		_w11183_,
		_w11184_,
		_w11185_,
		_w11187_,
		_w11480_
	);
	LUT4 #(
		.INIT('h8810)
	) name5654 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11481_
	);
	LUT3 #(
		.INIT('ha8)
	) name5655 (
		_w11190_,
		_w11480_,
		_w11481_,
		_w11482_
	);
	LUT4 #(
		.INIT('h0040)
	) name5656 (
		_w11184_,
		_w11185_,
		_w11187_,
		_w11190_,
		_w11483_
	);
	LUT4 #(
		.INIT('h5554)
	) name5657 (
		_w11183_,
		_w11185_,
		_w11187_,
		_w11188_,
		_w11484_
	);
	LUT2 #(
		.INIT('h4)
	) name5658 (
		_w11230_,
		_w11484_,
		_w11485_
	);
	LUT3 #(
		.INIT('h1b)
	) name5659 (
		_w11187_,
		_w11188_,
		_w11190_,
		_w11486_
	);
	LUT4 #(
		.INIT('h0141)
	) name5660 (
		_w11184_,
		_w11187_,
		_w11188_,
		_w11190_,
		_w11487_
	);
	LUT3 #(
		.INIT('h0d)
	) name5661 (
		_w11186_,
		_w11486_,
		_w11487_,
		_w11488_
	);
	LUT3 #(
		.INIT('he4)
	) name5662 (
		_w11185_,
		_w11187_,
		_w11188_,
		_w11489_
	);
	LUT4 #(
		.INIT('h0a02)
	) name5663 (
		_w11183_,
		_w11201_,
		_w11209_,
		_w11489_,
		_w11490_
	);
	LUT4 #(
		.INIT('h5540)
	) name5664 (
		_w11483_,
		_w11485_,
		_w11488_,
		_w11490_,
		_w11491_
	);
	LUT3 #(
		.INIT('h65)
	) name5665 (
		\u2_L5_reg[18]/NET0131 ,
		_w11482_,
		_w11491_,
		_w11492_
	);
	LUT4 #(
		.INIT('hc963)
	) name5666 (
		decrypt_pad,
		\u2_R4_reg[5]/NET0131 ,
		\u2_uk_K_r4_reg[47]/NET0131 ,
		\u2_uk_K_r4_reg[53]/NET0131 ,
		_w11493_
	);
	LUT4 #(
		.INIT('hc693)
	) name5667 (
		decrypt_pad,
		\u2_R4_reg[32]/NET0131 ,
		\u2_uk_K_r4_reg[34]/NET0131 ,
		\u2_uk_K_r4_reg[53]/NET0131 ,
		_w11494_
	);
	LUT2 #(
		.INIT('h1)
	) name5668 (
		_w11493_,
		_w11494_,
		_w11495_
	);
	LUT4 #(
		.INIT('hc963)
	) name5669 (
		decrypt_pad,
		\u2_R4_reg[1]/NET0131 ,
		\u2_uk_K_r4_reg[17]/NET0131 ,
		\u2_uk_K_r4_reg[55]/NET0131 ,
		_w11496_
	);
	LUT4 #(
		.INIT('hc963)
	) name5670 (
		decrypt_pad,
		\u2_R4_reg[3]/NET0131 ,
		\u2_uk_K_r4_reg[41]/NET0131 ,
		\u2_uk_K_r4_reg[47]/NET0131 ,
		_w11497_
	);
	LUT4 #(
		.INIT('hc693)
	) name5671 (
		decrypt_pad,
		\u2_R4_reg[2]/NET0131 ,
		\u2_uk_K_r4_reg[13]/NET0131 ,
		\u2_uk_K_r4_reg[32]/NET0131 ,
		_w11498_
	);
	LUT2 #(
		.INIT('h2)
	) name5672 (
		_w11497_,
		_w11498_,
		_w11499_
	);
	LUT4 #(
		.INIT('h003b)
	) name5673 (
		_w11497_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11500_
	);
	LUT3 #(
		.INIT('h01)
	) name5674 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11501_
	);
	LUT3 #(
		.INIT('h54)
	) name5675 (
		_w11495_,
		_w11500_,
		_w11501_,
		_w11502_
	);
	LUT4 #(
		.INIT('hdd8d)
	) name5676 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11503_
	);
	LUT3 #(
		.INIT('h04)
	) name5677 (
		_w11496_,
		_w11498_,
		_w11494_,
		_w11504_
	);
	LUT4 #(
		.INIT('hc963)
	) name5678 (
		decrypt_pad,
		\u2_R4_reg[4]/NET0131 ,
		\u2_uk_K_r4_reg[19]/NET0131 ,
		\u2_uk_K_r4_reg[25]/NET0131 ,
		_w11505_
	);
	LUT4 #(
		.INIT('hbf00)
	) name5679 (
		_w11497_,
		_w11496_,
		_w11494_,
		_w11505_,
		_w11506_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5680 (
		_w11497_,
		_w11503_,
		_w11504_,
		_w11506_,
		_w11507_
	);
	LUT2 #(
		.INIT('h4)
	) name5681 (
		_w11502_,
		_w11507_,
		_w11508_
	);
	LUT3 #(
		.INIT('h08)
	) name5682 (
		_w11497_,
		_w11498_,
		_w11494_,
		_w11509_
	);
	LUT4 #(
		.INIT('hff7c)
	) name5683 (
		_w11497_,
		_w11493_,
		_w11498_,
		_w11494_,
		_w11510_
	);
	LUT2 #(
		.INIT('h2)
	) name5684 (
		_w11496_,
		_w11510_,
		_w11511_
	);
	LUT2 #(
		.INIT('h8)
	) name5685 (
		_w11493_,
		_w11494_,
		_w11512_
	);
	LUT3 #(
		.INIT('hf4)
	) name5686 (
		_w11497_,
		_w11496_,
		_w11498_,
		_w11513_
	);
	LUT2 #(
		.INIT('h2)
	) name5687 (
		_w11512_,
		_w11513_,
		_w11514_
	);
	LUT2 #(
		.INIT('h8)
	) name5688 (
		_w11497_,
		_w11494_,
		_w11515_
	);
	LUT3 #(
		.INIT('h40)
	) name5689 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11516_
	);
	LUT3 #(
		.INIT('h15)
	) name5690 (
		_w11505_,
		_w11515_,
		_w11516_,
		_w11517_
	);
	LUT3 #(
		.INIT('h10)
	) name5691 (
		_w11511_,
		_w11514_,
		_w11517_,
		_w11518_
	);
	LUT2 #(
		.INIT('h1)
	) name5692 (
		_w11493_,
		_w11496_,
		_w11519_
	);
	LUT4 #(
		.INIT('heff2)
	) name5693 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11520_
	);
	LUT4 #(
		.INIT('h8000)
	) name5694 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11521_
	);
	LUT4 #(
		.INIT('h7bdb)
	) name5695 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11522_
	);
	LUT4 #(
		.INIT('h0155)
	) name5696 (
		_w11497_,
		_w11520_,
		_w11505_,
		_w11522_,
		_w11523_
	);
	LUT4 #(
		.INIT('h0200)
	) name5697 (
		_w11497_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11524_
	);
	LUT3 #(
		.INIT('h13)
	) name5698 (
		_w11519_,
		_w11524_,
		_w11509_,
		_w11525_
	);
	LUT2 #(
		.INIT('h4)
	) name5699 (
		_w11523_,
		_w11525_,
		_w11526_
	);
	LUT4 #(
		.INIT('ha955)
	) name5700 (
		\u2_L4_reg[31]/NET0131 ,
		_w11508_,
		_w11518_,
		_w11526_,
		_w11527_
	);
	LUT4 #(
		.INIT('hc963)
	) name5701 (
		decrypt_pad,
		\u2_R4_reg[24]/NET0131 ,
		\u2_uk_K_r4_reg[43]/NET0131 ,
		\u2_uk_K_r4_reg[51]/NET0131 ,
		_w11528_
	);
	LUT4 #(
		.INIT('hc963)
	) name5702 (
		decrypt_pad,
		\u2_R4_reg[20]/NET0131 ,
		\u2_uk_K_r4_reg[22]/NET0131 ,
		\u2_uk_K_r4_reg[30]/NET0131 ,
		_w11529_
	);
	LUT4 #(
		.INIT('hc963)
	) name5703 (
		decrypt_pad,
		\u2_R4_reg[22]/NET0131 ,
		\u2_uk_K_r4_reg[28]/NET0131 ,
		\u2_uk_K_r4_reg[36]/NET0131 ,
		_w11530_
	);
	LUT4 #(
		.INIT('hc693)
	) name5704 (
		decrypt_pad,
		\u2_R4_reg[21]/NET0131 ,
		\u2_uk_K_r4_reg[14]/NET0131 ,
		\u2_uk_K_r4_reg[37]/NET0131 ,
		_w11531_
	);
	LUT4 #(
		.INIT('hc963)
	) name5705 (
		decrypt_pad,
		\u2_R4_reg[23]/NET0131 ,
		\u2_uk_K_r4_reg[45]/NET0131 ,
		\u2_uk_K_r4_reg[49]/NET0131 ,
		_w11532_
	);
	LUT4 #(
		.INIT('h4155)
	) name5706 (
		_w11532_,
		_w11529_,
		_w11530_,
		_w11531_,
		_w11533_
	);
	LUT4 #(
		.INIT('hc693)
	) name5707 (
		decrypt_pad,
		\u2_R4_reg[25]/NET0131 ,
		\u2_uk_K_r4_reg[15]/NET0131 ,
		\u2_uk_K_r4_reg[7]/NET0131 ,
		_w11534_
	);
	LUT4 #(
		.INIT('haa8a)
	) name5708 (
		_w11532_,
		_w11529_,
		_w11534_,
		_w11531_,
		_w11535_
	);
	LUT3 #(
		.INIT('he6)
	) name5709 (
		_w11529_,
		_w11530_,
		_w11531_,
		_w11536_
	);
	LUT3 #(
		.INIT('h13)
	) name5710 (
		_w11535_,
		_w11533_,
		_w11536_,
		_w11537_
	);
	LUT4 #(
		.INIT('h0080)
	) name5711 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11538_
	);
	LUT2 #(
		.INIT('h2)
	) name5712 (
		_w11529_,
		_w11534_,
		_w11539_
	);
	LUT2 #(
		.INIT('h1)
	) name5713 (
		_w11532_,
		_w11530_,
		_w11540_
	);
	LUT3 #(
		.INIT('hce)
	) name5714 (
		_w11532_,
		_w11530_,
		_w11531_,
		_w11541_
	);
	LUT3 #(
		.INIT('h31)
	) name5715 (
		_w11539_,
		_w11538_,
		_w11541_,
		_w11542_
	);
	LUT3 #(
		.INIT('h45)
	) name5716 (
		_w11528_,
		_w11537_,
		_w11542_,
		_w11543_
	);
	LUT4 #(
		.INIT('h0002)
	) name5717 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11544_
	);
	LUT4 #(
		.INIT('h27fd)
	) name5718 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11545_
	);
	LUT2 #(
		.INIT('h2)
	) name5719 (
		_w11532_,
		_w11545_,
		_w11546_
	);
	LUT4 #(
		.INIT('h0415)
	) name5720 (
		_w11532_,
		_w11529_,
		_w11534_,
		_w11531_,
		_w11547_
	);
	LUT4 #(
		.INIT('h0b07)
	) name5721 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11548_
	);
	LUT3 #(
		.INIT('h0e)
	) name5722 (
		_w11540_,
		_w11547_,
		_w11548_,
		_w11549_
	);
	LUT3 #(
		.INIT('he0)
	) name5723 (
		_w11546_,
		_w11549_,
		_w11528_,
		_w11550_
	);
	LUT4 #(
		.INIT('h5155)
	) name5724 (
		_w11532_,
		_w11529_,
		_w11534_,
		_w11531_,
		_w11551_
	);
	LUT3 #(
		.INIT('h01)
	) name5725 (
		_w11530_,
		_w11551_,
		_w11535_,
		_w11552_
	);
	LUT4 #(
		.INIT('h7077)
	) name5726 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11553_
	);
	LUT4 #(
		.INIT('haa02)
	) name5727 (
		_w11532_,
		_w11529_,
		_w11534_,
		_w11530_,
		_w11554_
	);
	LUT3 #(
		.INIT('h01)
	) name5728 (
		_w11529_,
		_w11534_,
		_w11531_,
		_w11555_
	);
	LUT4 #(
		.INIT('h45cf)
	) name5729 (
		_w11540_,
		_w11553_,
		_w11554_,
		_w11555_,
		_w11556_
	);
	LUT2 #(
		.INIT('h4)
	) name5730 (
		_w11552_,
		_w11556_,
		_w11557_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5731 (
		\u2_L4_reg[11]/NET0131 ,
		_w11550_,
		_w11543_,
		_w11557_,
		_w11558_
	);
	LUT4 #(
		.INIT('hc693)
	) name5732 (
		decrypt_pad,
		\u2_R4_reg[28]/NET0131 ,
		\u2_uk_K_r4_reg[31]/P0001 ,
		\u2_uk_K_r4_reg[50]/NET0131 ,
		_w11559_
	);
	LUT4 #(
		.INIT('hc693)
	) name5733 (
		decrypt_pad,
		\u2_R4_reg[27]/NET0131 ,
		\u2_uk_K_r4_reg[16]/NET0131 ,
		\u2_uk_K_r4_reg[8]/NET0131 ,
		_w11560_
	);
	LUT4 #(
		.INIT('hc963)
	) name5734 (
		decrypt_pad,
		\u2_R4_reg[25]/NET0131 ,
		\u2_uk_K_r4_reg[14]/NET0131 ,
		\u2_uk_K_r4_reg[22]/NET0131 ,
		_w11561_
	);
	LUT4 #(
		.INIT('hc963)
	) name5735 (
		decrypt_pad,
		\u2_R4_reg[26]/NET0131 ,
		\u2_uk_K_r4_reg[30]/NET0131 ,
		\u2_uk_K_r4_reg[7]/NET0131 ,
		_w11562_
	);
	LUT4 #(
		.INIT('hc963)
	) name5736 (
		decrypt_pad,
		\u2_R4_reg[24]/NET0131 ,
		\u2_uk_K_r4_reg[38]/NET0131 ,
		\u2_uk_K_r4_reg[42]/NET0131 ,
		_w11563_
	);
	LUT4 #(
		.INIT('hc963)
	) name5737 (
		decrypt_pad,
		\u2_R4_reg[29]/NET0131 ,
		\u2_uk_K_r4_reg[42]/NET0131 ,
		\u2_uk_K_r4_reg[50]/NET0131 ,
		_w11564_
	);
	LUT4 #(
		.INIT('h1000)
	) name5738 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11565_
	);
	LUT2 #(
		.INIT('h4)
	) name5739 (
		_w11563_,
		_w11564_,
		_w11566_
	);
	LUT4 #(
		.INIT('he5ff)
	) name5740 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11567_
	);
	LUT2 #(
		.INIT('h1)
	) name5741 (
		_w11560_,
		_w11567_,
		_w11568_
	);
	LUT2 #(
		.INIT('h6)
	) name5742 (
		_w11561_,
		_w11562_,
		_w11569_
	);
	LUT4 #(
		.INIT('ha080)
	) name5743 (
		_w11560_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11570_
	);
	LUT4 #(
		.INIT('h0400)
	) name5744 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11571_
	);
	LUT4 #(
		.INIT('h0001)
	) name5745 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11572_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name5746 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11573_
	);
	LUT3 #(
		.INIT('h70)
	) name5747 (
		_w11569_,
		_w11570_,
		_w11573_,
		_w11574_
	);
	LUT3 #(
		.INIT('h8a)
	) name5748 (
		_w11559_,
		_w11568_,
		_w11574_,
		_w11575_
	);
	LUT4 #(
		.INIT('h0008)
	) name5749 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11576_
	);
	LUT4 #(
		.INIT('hfba6)
	) name5750 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11577_
	);
	LUT2 #(
		.INIT('h2)
	) name5751 (
		_w11560_,
		_w11577_,
		_w11578_
	);
	LUT4 #(
		.INIT('h80b0)
	) name5752 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11579_
	);
	LUT4 #(
		.INIT('h0004)
	) name5753 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11580_
	);
	LUT3 #(
		.INIT('h01)
	) name5754 (
		_w11560_,
		_w11579_,
		_w11580_,
		_w11581_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5755 (
		_w11560_,
		_w11561_,
		_w11562_,
		_w11563_,
		_w11582_
	);
	LUT2 #(
		.INIT('h1)
	) name5756 (
		_w11559_,
		_w11582_,
		_w11583_
	);
	LUT2 #(
		.INIT('h4)
	) name5757 (
		_w11559_,
		_w11564_,
		_w11584_
	);
	LUT4 #(
		.INIT('h8acf)
	) name5758 (
		_w11559_,
		_w11560_,
		_w11561_,
		_w11564_,
		_w11585_
	);
	LUT4 #(
		.INIT('hd00d)
	) name5759 (
		_w11560_,
		_w11561_,
		_w11562_,
		_w11563_,
		_w11586_
	);
	LUT2 #(
		.INIT('h4)
	) name5760 (
		_w11585_,
		_w11586_,
		_w11587_
	);
	LUT4 #(
		.INIT('h000b)
	) name5761 (
		_w11581_,
		_w11583_,
		_w11578_,
		_w11587_,
		_w11588_
	);
	LUT3 #(
		.INIT('h65)
	) name5762 (
		\u2_L4_reg[22]/NET0131 ,
		_w11575_,
		_w11588_,
		_w11589_
	);
	LUT4 #(
		.INIT('h0048)
	) name5763 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11590_
	);
	LUT4 #(
		.INIT('h28aa)
	) name5764 (
		_w11497_,
		_w11493_,
		_w11496_,
		_w11494_,
		_w11591_
	);
	LUT3 #(
		.INIT('h21)
	) name5765 (
		_w11493_,
		_w11496_,
		_w11494_,
		_w11592_
	);
	LUT4 #(
		.INIT('h5554)
	) name5766 (
		_w11497_,
		_w11493_,
		_w11498_,
		_w11494_,
		_w11593_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5767 (
		_w11590_,
		_w11591_,
		_w11592_,
		_w11593_,
		_w11594_
	);
	LUT4 #(
		.INIT('h4020)
	) name5768 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11595_
	);
	LUT2 #(
		.INIT('h1)
	) name5769 (
		_w11505_,
		_w11595_,
		_w11596_
	);
	LUT2 #(
		.INIT('h4)
	) name5770 (
		_w11594_,
		_w11596_,
		_w11597_
	);
	LUT4 #(
		.INIT('h0200)
	) name5771 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11598_
	);
	LUT4 #(
		.INIT('hfd03)
	) name5772 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11599_
	);
	LUT2 #(
		.INIT('h2)
	) name5773 (
		_w11497_,
		_w11599_,
		_w11600_
	);
	LUT4 #(
		.INIT('h0400)
	) name5774 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11601_
	);
	LUT4 #(
		.INIT('h0001)
	) name5775 (
		_w11497_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11602_
	);
	LUT3 #(
		.INIT('h80)
	) name5776 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11603_
	);
	LUT3 #(
		.INIT('h40)
	) name5777 (
		_w11497_,
		_w11498_,
		_w11494_,
		_w11604_
	);
	LUT4 #(
		.INIT('h0002)
	) name5778 (
		_w11505_,
		_w11602_,
		_w11603_,
		_w11604_,
		_w11605_
	);
	LUT3 #(
		.INIT('h10)
	) name5779 (
		_w11600_,
		_w11601_,
		_w11605_,
		_w11606_
	);
	LUT3 #(
		.INIT('ha9)
	) name5780 (
		\u2_L4_reg[17]/NET0131 ,
		_w11597_,
		_w11606_,
		_w11607_
	);
	LUT4 #(
		.INIT('hc693)
	) name5781 (
		decrypt_pad,
		\u2_R4_reg[13]/NET0131 ,
		\u2_uk_K_r4_reg[10]/NET0131 ,
		\u2_uk_K_r4_reg[4]/NET0131 ,
		_w11608_
	);
	LUT4 #(
		.INIT('hc963)
	) name5782 (
		decrypt_pad,
		\u2_R4_reg[12]/NET0131 ,
		\u2_uk_K_r4_reg[10]/NET0131 ,
		\u2_uk_K_r4_reg[48]/NET0131 ,
		_w11609_
	);
	LUT4 #(
		.INIT('hc963)
	) name5783 (
		decrypt_pad,
		\u2_R4_reg[17]/NET0131 ,
		\u2_uk_K_r4_reg[26]/NET0131 ,
		\u2_uk_K_r4_reg[32]/NET0131 ,
		_w11610_
	);
	LUT4 #(
		.INIT('hc963)
	) name5784 (
		decrypt_pad,
		\u2_R4_reg[15]/NET0131 ,
		\u2_uk_K_r4_reg[13]/NET0131 ,
		\u2_uk_K_r4_reg[19]/NET0131 ,
		_w11611_
	);
	LUT4 #(
		.INIT('h1000)
	) name5785 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11611_,
		_w11612_
	);
	LUT4 #(
		.INIT('hc693)
	) name5786 (
		decrypt_pad,
		\u2_R4_reg[16]/NET0131 ,
		\u2_uk_K_r4_reg[27]/P0001 ,
		\u2_uk_K_r4_reg[46]/NET0131 ,
		_w11613_
	);
	LUT4 #(
		.INIT('h0800)
	) name5787 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11611_,
		_w11614_
	);
	LUT2 #(
		.INIT('h4)
	) name5788 (
		_w11608_,
		_w11609_,
		_w11615_
	);
	LUT4 #(
		.INIT('hc693)
	) name5789 (
		decrypt_pad,
		\u2_R4_reg[14]/NET0131 ,
		\u2_uk_K_r4_reg[11]/NET0131 ,
		\u2_uk_K_r4_reg[5]/NET0131 ,
		_w11616_
	);
	LUT4 #(
		.INIT('h0006)
	) name5790 (
		_w11608_,
		_w11609_,
		_w11611_,
		_w11616_,
		_w11617_
	);
	LUT4 #(
		.INIT('h0004)
	) name5791 (
		_w11612_,
		_w11613_,
		_w11614_,
		_w11617_,
		_w11618_
	);
	LUT4 #(
		.INIT('h0020)
	) name5792 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11619_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name5793 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11620_
	);
	LUT4 #(
		.INIT('h0100)
	) name5794 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11621_
	);
	LUT3 #(
		.INIT('h8c)
	) name5795 (
		_w11611_,
		_w11620_,
		_w11621_,
		_w11622_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5796 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11611_,
		_w11623_
	);
	LUT4 #(
		.INIT('h7e00)
	) name5797 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11611_,
		_w11624_
	);
	LUT3 #(
		.INIT('h20)
	) name5798 (
		_w11609_,
		_w11610_,
		_w11616_,
		_w11625_
	);
	LUT3 #(
		.INIT('h0b)
	) name5799 (
		_w11608_,
		_w11610_,
		_w11611_,
		_w11626_
	);
	LUT3 #(
		.INIT('h45)
	) name5800 (
		_w11624_,
		_w11625_,
		_w11626_,
		_w11627_
	);
	LUT2 #(
		.INIT('h8)
	) name5801 (
		_w11611_,
		_w11616_,
		_w11628_
	);
	LUT4 #(
		.INIT('h2000)
	) name5802 (
		_w11608_,
		_w11609_,
		_w11611_,
		_w11616_,
		_w11629_
	);
	LUT4 #(
		.INIT('h0001)
	) name5803 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11630_
	);
	LUT4 #(
		.INIT('h0200)
	) name5804 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11631_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name5805 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11632_
	);
	LUT4 #(
		.INIT('h0100)
	) name5806 (
		_w11613_,
		_w11630_,
		_w11629_,
		_w11632_,
		_w11633_
	);
	LUT4 #(
		.INIT('h7077)
	) name5807 (
		_w11618_,
		_w11622_,
		_w11627_,
		_w11633_,
		_w11634_
	);
	LUT4 #(
		.INIT('h0400)
	) name5808 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11635_
	);
	LUT4 #(
		.INIT('hfff6)
	) name5809 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11636_
	);
	LUT4 #(
		.INIT('he4ee)
	) name5810 (
		_w11611_,
		_w11619_,
		_w11635_,
		_w11636_,
		_w11637_
	);
	LUT3 #(
		.INIT('h56)
	) name5811 (
		\u2_L4_reg[20]/NET0131 ,
		_w11634_,
		_w11637_,
		_w11638_
	);
	LUT4 #(
		.INIT('h67dc)
	) name5812 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11639_
	);
	LUT4 #(
		.INIT('hd2f7)
	) name5813 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11640_
	);
	LUT4 #(
		.INIT('h0040)
	) name5814 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11641_
	);
	LUT4 #(
		.INIT('h00d8)
	) name5815 (
		_w11532_,
		_w11639_,
		_w11640_,
		_w11641_,
		_w11642_
	);
	LUT4 #(
		.INIT('h9aff)
	) name5816 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11643_
	);
	LUT4 #(
		.INIT('haa02)
	) name5817 (
		_w11532_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11644_
	);
	LUT4 #(
		.INIT('h9297)
	) name5818 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11645_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name5819 (
		_w11532_,
		_w11643_,
		_w11644_,
		_w11645_,
		_w11646_
	);
	LUT4 #(
		.INIT('h0800)
	) name5820 (
		_w11532_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11647_
	);
	LUT2 #(
		.INIT('h1)
	) name5821 (
		_w11544_,
		_w11647_,
		_w11648_
	);
	LUT4 #(
		.INIT('hd800)
	) name5822 (
		_w11528_,
		_w11646_,
		_w11642_,
		_w11648_,
		_w11649_
	);
	LUT2 #(
		.INIT('h6)
	) name5823 (
		\u2_L4_reg[29]/NET0131 ,
		_w11649_,
		_w11650_
	);
	LUT4 #(
		.INIT('hc963)
	) name5824 (
		decrypt_pad,
		\u2_R4_reg[8]/NET0131 ,
		\u2_uk_K_r4_reg[20]/NET0131 ,
		\u2_uk_K_r4_reg[26]/NET0131 ,
		_w11651_
	);
	LUT4 #(
		.INIT('hc963)
	) name5825 (
		decrypt_pad,
		\u2_R4_reg[5]/NET0131 ,
		\u2_uk_K_r4_reg[12]/NET0131 ,
		\u2_uk_K_r4_reg[18]/NET0131 ,
		_w11652_
	);
	LUT4 #(
		.INIT('hc963)
	) name5826 (
		decrypt_pad,
		\u2_R4_reg[9]/NET0131 ,
		\u2_uk_K_r4_reg[25]/NET0131 ,
		\u2_uk_K_r4_reg[6]/NET0131 ,
		_w11653_
	);
	LUT4 #(
		.INIT('hc963)
	) name5827 (
		decrypt_pad,
		\u2_R4_reg[4]/NET0131 ,
		\u2_uk_K_r4_reg[33]/NET0131 ,
		\u2_uk_K_r4_reg[39]/NET0131 ,
		_w11654_
	);
	LUT3 #(
		.INIT('h04)
	) name5828 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11655_
	);
	LUT3 #(
		.INIT('hd9)
	) name5829 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11656_
	);
	LUT4 #(
		.INIT('hc963)
	) name5830 (
		decrypt_pad,
		\u2_R4_reg[6]/NET0131 ,
		\u2_uk_K_r4_reg[3]/NET0131 ,
		\u2_uk_K_r4_reg[41]/NET0131 ,
		_w11657_
	);
	LUT4 #(
		.INIT('h0026)
	) name5831 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11658_
	);
	LUT4 #(
		.INIT('hc693)
	) name5832 (
		decrypt_pad,
		\u2_R4_reg[7]/NET0131 ,
		\u2_uk_K_r4_reg[3]/NET0131 ,
		\u2_uk_K_r4_reg[54]/NET0131 ,
		_w11659_
	);
	LUT4 #(
		.INIT('h4000)
	) name5833 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11660_
	);
	LUT3 #(
		.INIT('h15)
	) name5834 (
		_w11658_,
		_w11659_,
		_w11660_,
		_w11661_
	);
	LUT2 #(
		.INIT('h8)
	) name5835 (
		_w11654_,
		_w11657_,
		_w11662_
	);
	LUT4 #(
		.INIT('h4bfb)
	) name5836 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11663_
	);
	LUT3 #(
		.INIT('hcd)
	) name5837 (
		_w11652_,
		_w11657_,
		_w11659_,
		_w11664_
	);
	LUT2 #(
		.INIT('h2)
	) name5838 (
		_w11653_,
		_w11654_,
		_w11665_
	);
	LUT4 #(
		.INIT('h084c)
	) name5839 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11666_
	);
	LUT4 #(
		.INIT('h0eee)
	) name5840 (
		_w11659_,
		_w11663_,
		_w11664_,
		_w11666_,
		_w11667_
	);
	LUT3 #(
		.INIT('h15)
	) name5841 (
		_w11651_,
		_w11661_,
		_w11667_,
		_w11668_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name5842 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11669_
	);
	LUT4 #(
		.INIT('h080c)
	) name5843 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11670_
	);
	LUT3 #(
		.INIT('h0d)
	) name5844 (
		_w11652_,
		_w11657_,
		_w11659_,
		_w11671_
	);
	LUT4 #(
		.INIT('hf200)
	) name5845 (
		_w11651_,
		_w11669_,
		_w11670_,
		_w11671_,
		_w11672_
	);
	LUT4 #(
		.INIT('h0080)
	) name5846 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11673_
	);
	LUT4 #(
		.INIT('h0010)
	) name5847 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11674_
	);
	LUT4 #(
		.INIT('h8a00)
	) name5848 (
		_w11652_,
		_w11654_,
		_w11657_,
		_w11659_,
		_w11675_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5849 (
		_w11651_,
		_w11674_,
		_w11675_,
		_w11673_,
		_w11676_
	);
	LUT4 #(
		.INIT('hfc54)
	) name5850 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11677_
	);
	LUT4 #(
		.INIT('hdc00)
	) name5851 (
		_w11652_,
		_w11654_,
		_w11657_,
		_w11659_,
		_w11678_
	);
	LUT2 #(
		.INIT('h4)
	) name5852 (
		_w11677_,
		_w11678_,
		_w11679_
	);
	LUT3 #(
		.INIT('h01)
	) name5853 (
		_w11676_,
		_w11679_,
		_w11672_,
		_w11680_
	);
	LUT3 #(
		.INIT('h65)
	) name5854 (
		\u2_L4_reg[2]/NET0131 ,
		_w11668_,
		_w11680_,
		_w11681_
	);
	LUT4 #(
		.INIT('hd97b)
	) name5855 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11682_
	);
	LUT2 #(
		.INIT('h2)
	) name5856 (
		_w11532_,
		_w11682_,
		_w11683_
	);
	LUT4 #(
		.INIT('heebf)
	) name5857 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11684_
	);
	LUT4 #(
		.INIT('h0040)
	) name5858 (
		_w11532_,
		_w11529_,
		_w11534_,
		_w11530_,
		_w11685_
	);
	LUT4 #(
		.INIT('h0032)
	) name5859 (
		_w11532_,
		_w11544_,
		_w11684_,
		_w11685_,
		_w11686_
	);
	LUT3 #(
		.INIT('h45)
	) name5860 (
		_w11528_,
		_w11683_,
		_w11686_,
		_w11687_
	);
	LUT4 #(
		.INIT('h7c7f)
	) name5861 (
		_w11532_,
		_w11529_,
		_w11534_,
		_w11531_,
		_w11688_
	);
	LUT2 #(
		.INIT('h1)
	) name5862 (
		_w11530_,
		_w11688_,
		_w11689_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name5863 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11690_
	);
	LUT3 #(
		.INIT('h80)
	) name5864 (
		_w11534_,
		_w11530_,
		_w11531_,
		_w11691_
	);
	LUT3 #(
		.INIT('h0e)
	) name5865 (
		_w11532_,
		_w11690_,
		_w11691_,
		_w11692_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5866 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11693_
	);
	LUT4 #(
		.INIT('h5501)
	) name5867 (
		_w11532_,
		_w11529_,
		_w11534_,
		_w11530_,
		_w11694_
	);
	LUT3 #(
		.INIT('h9e)
	) name5868 (
		_w11529_,
		_w11534_,
		_w11531_,
		_w11695_
	);
	LUT2 #(
		.INIT('h8)
	) name5869 (
		_w11532_,
		_w11530_,
		_w11696_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name5870 (
		_w11693_,
		_w11694_,
		_w11695_,
		_w11696_,
		_w11697_
	);
	LUT4 #(
		.INIT('h7500)
	) name5871 (
		_w11528_,
		_w11689_,
		_w11692_,
		_w11697_,
		_w11698_
	);
	LUT3 #(
		.INIT('h65)
	) name5872 (
		\u2_L4_reg[4]/NET0131 ,
		_w11687_,
		_w11698_,
		_w11699_
	);
	LUT4 #(
		.INIT('hc963)
	) name5873 (
		decrypt_pad,
		\u2_R4_reg[32]/NET0131 ,
		\u2_uk_K_r4_reg[15]/NET0131 ,
		\u2_uk_K_r4_reg[23]/NET0131 ,
		_w11700_
	);
	LUT4 #(
		.INIT('hc693)
	) name5874 (
		decrypt_pad,
		\u2_R4_reg[31]/P0001 ,
		\u2_uk_K_r4_reg[45]/NET0131 ,
		\u2_uk_K_r4_reg[9]/NET0131 ,
		_w11701_
	);
	LUT4 #(
		.INIT('hc693)
	) name5875 (
		decrypt_pad,
		\u2_R4_reg[28]/NET0131 ,
		\u2_uk_K_r4_reg[1]/NET0131 ,
		\u2_uk_K_r4_reg[52]/NET0131 ,
		_w11702_
	);
	LUT4 #(
		.INIT('hc693)
	) name5876 (
		decrypt_pad,
		\u2_R4_reg[29]/NET0131 ,
		\u2_uk_K_r4_reg[28]/NET0131 ,
		\u2_uk_K_r4_reg[51]/NET0131 ,
		_w11703_
	);
	LUT4 #(
		.INIT('hc963)
	) name5877 (
		decrypt_pad,
		\u2_R4_reg[1]/NET0131 ,
		\u2_uk_K_r4_reg[36]/NET0131 ,
		\u2_uk_K_r4_reg[44]/NET0131 ,
		_w11704_
	);
	LUT4 #(
		.INIT('hc963)
	) name5878 (
		decrypt_pad,
		\u2_R4_reg[30]/NET0131 ,
		\u2_uk_K_r4_reg[21]/NET0131 ,
		\u2_uk_K_r4_reg[29]/NET0131 ,
		_w11705_
	);
	LUT4 #(
		.INIT('h1000)
	) name5879 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11706_
	);
	LUT4 #(
		.INIT('hebfb)
	) name5880 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11707_
	);
	LUT2 #(
		.INIT('h2)
	) name5881 (
		_w11702_,
		_w11705_,
		_w11708_
	);
	LUT2 #(
		.INIT('h4)
	) name5882 (
		_w11702_,
		_w11705_,
		_w11709_
	);
	LUT4 #(
		.INIT('h7407)
	) name5883 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11710_
	);
	LUT3 #(
		.INIT('h08)
	) name5884 (
		_w11703_,
		_w11702_,
		_w11705_,
		_w11711_
	);
	LUT4 #(
		.INIT('h0020)
	) name5885 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11712_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name5886 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11713_
	);
	LUT4 #(
		.INIT('he400)
	) name5887 (
		_w11701_,
		_w11710_,
		_w11707_,
		_w11713_,
		_w11714_
	);
	LUT2 #(
		.INIT('h1)
	) name5888 (
		_w11700_,
		_w11714_,
		_w11715_
	);
	LUT4 #(
		.INIT('hcf45)
	) name5889 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11716_
	);
	LUT4 #(
		.INIT('h22d2)
	) name5890 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11717_
	);
	LUT4 #(
		.INIT('h0001)
	) name5891 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11718_
	);
	LUT4 #(
		.INIT('h0400)
	) name5892 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11719_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name5893 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11720_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5894 (
		_w11700_,
		_w11716_,
		_w11717_,
		_w11720_,
		_w11721_
	);
	LUT4 #(
		.INIT('h0800)
	) name5895 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11722_
	);
	LUT2 #(
		.INIT('h8)
	) name5896 (
		_w11700_,
		_w11722_,
		_w11723_
	);
	LUT4 #(
		.INIT('h2002)
	) name5897 (
		_w11700_,
		_w11703_,
		_w11702_,
		_w11705_,
		_w11724_
	);
	LUT2 #(
		.INIT('h1)
	) name5898 (
		_w11724_,
		_w11712_,
		_w11725_
	);
	LUT4 #(
		.INIT('h5404)
	) name5899 (
		_w11723_,
		_w11725_,
		_w11701_,
		_w11721_,
		_w11726_
	);
	LUT3 #(
		.INIT('h9a)
	) name5900 (
		\u2_L4_reg[5]/NET0131 ,
		_w11715_,
		_w11726_,
		_w11727_
	);
	LUT4 #(
		.INIT('hfdbd)
	) name5901 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11728_
	);
	LUT2 #(
		.INIT('h2)
	) name5902 (
		_w11611_,
		_w11728_,
		_w11729_
	);
	LUT4 #(
		.INIT('h6fff)
	) name5903 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11730_
	);
	LUT4 #(
		.INIT('hf353)
	) name5904 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11731_
	);
	LUT3 #(
		.INIT('h08)
	) name5905 (
		_w11608_,
		_w11609_,
		_w11616_,
		_w11732_
	);
	LUT4 #(
		.INIT('h0f07)
	) name5906 (
		_w11608_,
		_w11609_,
		_w11611_,
		_w11616_,
		_w11733_
	);
	LUT3 #(
		.INIT('h8a)
	) name5907 (
		_w11730_,
		_w11731_,
		_w11733_,
		_w11734_
	);
	LUT3 #(
		.INIT('h8a)
	) name5908 (
		_w11613_,
		_w11729_,
		_w11734_,
		_w11735_
	);
	LUT4 #(
		.INIT('hcefe)
	) name5909 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11611_,
		_w11736_
	);
	LUT2 #(
		.INIT('h1)
	) name5910 (
		_w11628_,
		_w11736_,
		_w11737_
	);
	LUT3 #(
		.INIT('hc4)
	) name5911 (
		_w11610_,
		_w11611_,
		_w11616_,
		_w11738_
	);
	LUT2 #(
		.INIT('h8)
	) name5912 (
		_w11615_,
		_w11738_,
		_w11739_
	);
	LUT4 #(
		.INIT('h0008)
	) name5913 (
		_w11609_,
		_w11610_,
		_w11611_,
		_w11616_,
		_w11740_
	);
	LUT3 #(
		.INIT('h01)
	) name5914 (
		_w11631_,
		_w11740_,
		_w11732_,
		_w11741_
	);
	LUT4 #(
		.INIT('h5455)
	) name5915 (
		_w11613_,
		_w11737_,
		_w11739_,
		_w11741_,
		_w11742_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name5916 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11743_
	);
	LUT2 #(
		.INIT('h1)
	) name5917 (
		_w11611_,
		_w11743_,
		_w11744_
	);
	LUT3 #(
		.INIT('h0b)
	) name5918 (
		_w11616_,
		_w11614_,
		_w11629_,
		_w11745_
	);
	LUT2 #(
		.INIT('h4)
	) name5919 (
		_w11744_,
		_w11745_,
		_w11746_
	);
	LUT4 #(
		.INIT('h5655)
	) name5920 (
		\u2_L4_reg[10]/NET0131 ,
		_w11742_,
		_w11735_,
		_w11746_,
		_w11747_
	);
	LUT4 #(
		.INIT('h0006)
	) name5921 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11748_
	);
	LUT3 #(
		.INIT('h1d)
	) name5922 (
		_w11560_,
		_w11561_,
		_w11562_,
		_w11749_
	);
	LUT4 #(
		.INIT('h4000)
	) name5923 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11750_
	);
	LUT4 #(
		.INIT('h000d)
	) name5924 (
		_w11566_,
		_w11749_,
		_w11748_,
		_w11750_,
		_w11751_
	);
	LUT4 #(
		.INIT('h5455)
	) name5925 (
		_w11559_,
		_w11561_,
		_w11562_,
		_w11563_,
		_w11752_
	);
	LUT2 #(
		.INIT('h6)
	) name5926 (
		_w11561_,
		_w11564_,
		_w11753_
	);
	LUT4 #(
		.INIT('h152a)
	) name5927 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11754_
	);
	LUT4 #(
		.INIT('hfca8)
	) name5928 (
		_w11560_,
		_w11584_,
		_w11752_,
		_w11754_,
		_w11755_
	);
	LUT3 #(
		.INIT('h2a)
	) name5929 (
		_w11560_,
		_w11561_,
		_w11563_,
		_w11756_
	);
	LUT4 #(
		.INIT('he0ee)
	) name5930 (
		_w11560_,
		_w11571_,
		_w11572_,
		_w11756_,
		_w11757_
	);
	LUT4 #(
		.INIT('h0240)
	) name5931 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11758_
	);
	LUT4 #(
		.INIT('h0002)
	) name5932 (
		_w11559_,
		_w11576_,
		_w11565_,
		_w11758_,
		_w11759_
	);
	LUT4 #(
		.INIT('h7077)
	) name5933 (
		_w11751_,
		_w11755_,
		_w11757_,
		_w11759_,
		_w11760_
	);
	LUT2 #(
		.INIT('h6)
	) name5934 (
		\u2_L4_reg[12]/NET0131 ,
		_w11760_,
		_w11761_
	);
	LUT4 #(
		.INIT('h2000)
	) name5935 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11762_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name5936 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11763_
	);
	LUT4 #(
		.INIT('h0400)
	) name5937 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11764_
	);
	LUT4 #(
		.INIT('hf9ed)
	) name5938 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11765_
	);
	LUT4 #(
		.INIT('h0313)
	) name5939 (
		_w11651_,
		_w11659_,
		_w11763_,
		_w11765_,
		_w11766_
	);
	LUT3 #(
		.INIT('h8e)
	) name5940 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11767_
	);
	LUT4 #(
		.INIT('h3010)
	) name5941 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11768_
	);
	LUT3 #(
		.INIT('h02)
	) name5942 (
		_w11659_,
		_w11767_,
		_w11768_,
		_w11769_
	);
	LUT3 #(
		.INIT('hd0)
	) name5943 (
		_w11652_,
		_w11653_,
		_w11659_,
		_w11770_
	);
	LUT2 #(
		.INIT('h8)
	) name5944 (
		_w11662_,
		_w11770_,
		_w11771_
	);
	LUT3 #(
		.INIT('h51)
	) name5945 (
		_w11651_,
		_w11665_,
		_w11664_,
		_w11772_
	);
	LUT3 #(
		.INIT('h10)
	) name5946 (
		_w11771_,
		_w11769_,
		_w11772_,
		_w11773_
	);
	LUT4 #(
		.INIT('h0002)
	) name5947 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11774_
	);
	LUT4 #(
		.INIT('h002a)
	) name5948 (
		_w11651_,
		_w11664_,
		_w11666_,
		_w11774_,
		_w11775_
	);
	LUT4 #(
		.INIT('h5140)
	) name5949 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11776_
	);
	LUT3 #(
		.INIT('h01)
	) name5950 (
		_w11652_,
		_w11653_,
		_w11657_,
		_w11777_
	);
	LUT4 #(
		.INIT('hf3ee)
	) name5951 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11778_
	);
	LUT4 #(
		.INIT('h80c4)
	) name5952 (
		_w11659_,
		_w11763_,
		_w11778_,
		_w11776_,
		_w11779_
	);
	LUT2 #(
		.INIT('h8)
	) name5953 (
		_w11775_,
		_w11779_,
		_w11780_
	);
	LUT4 #(
		.INIT('h999a)
	) name5954 (
		\u2_L4_reg[13]/NET0131 ,
		_w11766_,
		_w11773_,
		_w11780_,
		_w11781_
	);
	LUT4 #(
		.INIT('h02a0)
	) name5955 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11782_
	);
	LUT4 #(
		.INIT('h0100)
	) name5956 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11701_,
		_w11783_
	);
	LUT4 #(
		.INIT('h4000)
	) name5957 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11784_
	);
	LUT4 #(
		.INIT('h0040)
	) name5958 (
		_w11703_,
		_w11704_,
		_w11705_,
		_w11701_,
		_w11785_
	);
	LUT4 #(
		.INIT('h0002)
	) name5959 (
		_w11700_,
		_w11784_,
		_w11783_,
		_w11785_,
		_w11786_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name5960 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11787_
	);
	LUT4 #(
		.INIT('h5b59)
	) name5961 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11788_
	);
	LUT4 #(
		.INIT('h0010)
	) name5962 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11789_
	);
	LUT4 #(
		.INIT('h0501)
	) name5963 (
		_w11700_,
		_w11701_,
		_w11789_,
		_w11788_,
		_w11790_
	);
	LUT3 #(
		.INIT('h0b)
	) name5964 (
		_w11782_,
		_w11786_,
		_w11790_,
		_w11791_
	);
	LUT4 #(
		.INIT('h0009)
	) name5965 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11792_
	);
	LUT4 #(
		.INIT('h3010)
	) name5966 (
		_w11700_,
		_w11703_,
		_w11702_,
		_w11705_,
		_w11793_
	);
	LUT4 #(
		.INIT('h0200)
	) name5967 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11794_
	);
	LUT4 #(
		.INIT('h0001)
	) name5968 (
		_w11701_,
		_w11794_,
		_w11792_,
		_w11793_,
		_w11795_
	);
	LUT4 #(
		.INIT('h0004)
	) name5969 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11796_
	);
	LUT3 #(
		.INIT('h04)
	) name5970 (
		_w11722_,
		_w11701_,
		_w11796_,
		_w11797_
	);
	LUT2 #(
		.INIT('h1)
	) name5971 (
		_w11795_,
		_w11797_,
		_w11798_
	);
	LUT3 #(
		.INIT('h56)
	) name5972 (
		\u2_L4_reg[15]/NET0131 ,
		_w11791_,
		_w11798_,
		_w11799_
	);
	LUT4 #(
		.INIT('hc963)
	) name5973 (
		decrypt_pad,
		\u2_R4_reg[20]/NET0131 ,
		\u2_uk_K_r4_reg[0]/P0001 ,
		\u2_uk_K_r4_reg[8]/NET0131 ,
		_w11800_
	);
	LUT4 #(
		.INIT('hc963)
	) name5974 (
		decrypt_pad,
		\u2_R4_reg[19]/NET0131 ,
		\u2_uk_K_r4_reg[16]/NET0131 ,
		\u2_uk_K_r4_reg[52]/NET0131 ,
		_w11801_
	);
	LUT4 #(
		.INIT('hc963)
	) name5975 (
		decrypt_pad,
		\u2_R4_reg[18]/NET0131 ,
		\u2_uk_K_r4_reg[29]/NET0131 ,
		\u2_uk_K_r4_reg[37]/NET0131 ,
		_w11802_
	);
	LUT4 #(
		.INIT('hc963)
	) name5976 (
		decrypt_pad,
		\u2_R4_reg[21]/NET0131 ,
		\u2_uk_K_r4_reg[1]/NET0131 ,
		\u2_uk_K_r4_reg[9]/NET0131 ,
		_w11803_
	);
	LUT4 #(
		.INIT('hc693)
	) name5977 (
		decrypt_pad,
		\u2_R4_reg[16]/NET0131 ,
		\u2_uk_K_r4_reg[21]/NET0131 ,
		\u2_uk_K_r4_reg[44]/NET0131 ,
		_w11804_
	);
	LUT4 #(
		.INIT('hc963)
	) name5978 (
		decrypt_pad,
		\u2_R4_reg[17]/NET0131 ,
		\u2_uk_K_r4_reg[35]/NET0131 ,
		\u2_uk_K_r4_reg[43]/NET0131 ,
		_w11805_
	);
	LUT4 #(
		.INIT('h0004)
	) name5979 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11806_
	);
	LUT4 #(
		.INIT('h0080)
	) name5980 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11807_
	);
	LUT4 #(
		.INIT('had79)
	) name5981 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11808_
	);
	LUT2 #(
		.INIT('h1)
	) name5982 (
		_w11801_,
		_w11808_,
		_w11809_
	);
	LUT4 #(
		.INIT('h0810)
	) name5983 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11810_
	);
	LUT4 #(
		.INIT('h46ce)
	) name5984 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11811_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5985 (
		_w11801_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11812_
	);
	LUT3 #(
		.INIT('h45)
	) name5986 (
		_w11810_,
		_w11811_,
		_w11812_,
		_w11813_
	);
	LUT3 #(
		.INIT('h45)
	) name5987 (
		_w11800_,
		_w11809_,
		_w11813_,
		_w11814_
	);
	LUT3 #(
		.INIT('h04)
	) name5988 (
		_w11804_,
		_w11805_,
		_w11802_,
		_w11815_
	);
	LUT4 #(
		.INIT('h9d35)
	) name5989 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11816_
	);
	LUT2 #(
		.INIT('h2)
	) name5990 (
		_w11801_,
		_w11816_,
		_w11817_
	);
	LUT2 #(
		.INIT('h1)
	) name5991 (
		_w11801_,
		_w11802_,
		_w11818_
	);
	LUT3 #(
		.INIT('hde)
	) name5992 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11819_
	);
	LUT2 #(
		.INIT('h2)
	) name5993 (
		_w11818_,
		_w11819_,
		_w11820_
	);
	LUT4 #(
		.INIT('h0400)
	) name5994 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11821_
	);
	LUT4 #(
		.INIT('hfbf7)
	) name5995 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11822_
	);
	LUT2 #(
		.INIT('h4)
	) name5996 (
		_w11801_,
		_w11802_,
		_w11823_
	);
	LUT3 #(
		.INIT('h80)
	) name5997 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11824_
	);
	LUT4 #(
		.INIT('h0040)
	) name5998 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11825_
	);
	LUT4 #(
		.INIT('h0700)
	) name5999 (
		_w11823_,
		_w11824_,
		_w11825_,
		_w11822_,
		_w11826_
	);
	LUT4 #(
		.INIT('hef00)
	) name6000 (
		_w11817_,
		_w11820_,
		_w11826_,
		_w11800_,
		_w11827_
	);
	LUT4 #(
		.INIT('h0200)
	) name6001 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11828_
	);
	LUT4 #(
		.INIT('h1200)
	) name6002 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11829_
	);
	LUT4 #(
		.INIT('hfebf)
	) name6003 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11830_
	);
	LUT3 #(
		.INIT('hb1)
	) name6004 (
		_w11801_,
		_w11829_,
		_w11830_,
		_w11831_
	);
	LUT4 #(
		.INIT('h5655)
	) name6005 (
		\u2_L4_reg[14]/NET0131 ,
		_w11827_,
		_w11814_,
		_w11831_,
		_w11832_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name6006 (
		_w11532_,
		_w11529_,
		_w11534_,
		_w11530_,
		_w11833_
	);
	LUT4 #(
		.INIT('hef00)
	) name6007 (
		_w11534_,
		_w11530_,
		_w11531_,
		_w11528_,
		_w11834_
	);
	LUT3 #(
		.INIT('he0)
	) name6008 (
		_w11531_,
		_w11833_,
		_w11834_,
		_w11835_
	);
	LUT4 #(
		.INIT('h4010)
	) name6009 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11836_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name6010 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11837_
	);
	LUT3 #(
		.INIT('h31)
	) name6011 (
		_w11532_,
		_w11836_,
		_w11837_,
		_w11838_
	);
	LUT4 #(
		.INIT('h4e55)
	) name6012 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11839_
	);
	LUT2 #(
		.INIT('h2)
	) name6013 (
		_w11532_,
		_w11839_,
		_w11840_
	);
	LUT4 #(
		.INIT('h1001)
	) name6014 (
		_w11532_,
		_w11529_,
		_w11534_,
		_w11531_,
		_w11841_
	);
	LUT4 #(
		.INIT('h8000)
	) name6015 (
		_w11529_,
		_w11534_,
		_w11530_,
		_w11531_,
		_w11842_
	);
	LUT3 #(
		.INIT('h01)
	) name6016 (
		_w11528_,
		_w11842_,
		_w11841_,
		_w11843_
	);
	LUT4 #(
		.INIT('h7077)
	) name6017 (
		_w11835_,
		_w11838_,
		_w11840_,
		_w11843_,
		_w11844_
	);
	LUT2 #(
		.INIT('h4)
	) name6018 (
		_w11531_,
		_w11685_,
		_w11845_
	);
	LUT2 #(
		.INIT('h1)
	) name6019 (
		_w11552_,
		_w11845_,
		_w11846_
	);
	LUT3 #(
		.INIT('h65)
	) name6020 (
		\u2_L4_reg[19]/NET0131 ,
		_w11844_,
		_w11846_,
		_w11847_
	);
	LUT4 #(
		.INIT('hafab)
	) name6021 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11848_
	);
	LUT4 #(
		.INIT('h6dff)
	) name6022 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11849_
	);
	LUT4 #(
		.INIT('h08aa)
	) name6023 (
		_w11611_,
		_w11613_,
		_w11848_,
		_w11849_,
		_w11850_
	);
	LUT4 #(
		.INIT('h404c)
	) name6024 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11851_
	);
	LUT3 #(
		.INIT('h01)
	) name6025 (
		_w11609_,
		_w11610_,
		_w11616_,
		_w11852_
	);
	LUT4 #(
		.INIT('hfad8)
	) name6026 (
		_w11611_,
		_w11635_,
		_w11851_,
		_w11852_,
		_w11853_
	);
	LUT4 #(
		.INIT('h7fd7)
	) name6027 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11854_
	);
	LUT3 #(
		.INIT('h45)
	) name6028 (
		_w11613_,
		_w11853_,
		_w11854_,
		_w11855_
	);
	LUT4 #(
		.INIT('hdf5d)
	) name6029 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11856_
	);
	LUT4 #(
		.INIT('he6ff)
	) name6030 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11857_
	);
	LUT4 #(
		.INIT('h04cc)
	) name6031 (
		_w11611_,
		_w11613_,
		_w11856_,
		_w11857_,
		_w11858_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name6032 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11859_
	);
	LUT2 #(
		.INIT('h1)
	) name6033 (
		_w11611_,
		_w11859_,
		_w11860_
	);
	LUT2 #(
		.INIT('h1)
	) name6034 (
		_w11858_,
		_w11860_,
		_w11861_
	);
	LUT4 #(
		.INIT('h5655)
	) name6035 (
		\u2_L4_reg[1]/NET0131 ,
		_w11855_,
		_w11850_,
		_w11861_,
		_w11862_
	);
	LUT4 #(
		.INIT('h00fb)
	) name6036 (
		_w11704_,
		_w11702_,
		_w11705_,
		_w11701_,
		_w11863_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6037 (
		_w11703_,
		_w11702_,
		_w11705_,
		_w11701_,
		_w11864_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name6038 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11865_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name6039 (
		_w11784_,
		_w11863_,
		_w11864_,
		_w11865_,
		_w11866_
	);
	LUT4 #(
		.INIT('h2100)
	) name6040 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11867_
	);
	LUT3 #(
		.INIT('h02)
	) name6041 (
		_w11700_,
		_w11796_,
		_w11867_,
		_w11868_
	);
	LUT2 #(
		.INIT('h4)
	) name6042 (
		_w11866_,
		_w11868_,
		_w11869_
	);
	LUT2 #(
		.INIT('h2)
	) name6043 (
		_w11704_,
		_w11701_,
		_w11870_
	);
	LUT3 #(
		.INIT('h73)
	) name6044 (
		_w11703_,
		_w11704_,
		_w11701_,
		_w11871_
	);
	LUT2 #(
		.INIT('h2)
	) name6045 (
		_w11708_,
		_w11871_,
		_w11872_
	);
	LUT3 #(
		.INIT('h51)
	) name6046 (
		_w11703_,
		_w11704_,
		_w11701_,
		_w11873_
	);
	LUT3 #(
		.INIT('h31)
	) name6047 (
		_w11709_,
		_w11706_,
		_w11873_,
		_w11874_
	);
	LUT4 #(
		.INIT('h8fdf)
	) name6048 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11875_
	);
	LUT2 #(
		.INIT('h2)
	) name6049 (
		_w11701_,
		_w11875_,
		_w11876_
	);
	LUT4 #(
		.INIT('h0002)
	) name6050 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11701_,
		_w11877_
	);
	LUT3 #(
		.INIT('h01)
	) name6051 (
		_w11700_,
		_w11718_,
		_w11877_,
		_w11878_
	);
	LUT4 #(
		.INIT('h1000)
	) name6052 (
		_w11876_,
		_w11872_,
		_w11878_,
		_w11874_,
		_w11879_
	);
	LUT4 #(
		.INIT('h0100)
	) name6053 (
		_w11703_,
		_w11702_,
		_w11705_,
		_w11701_,
		_w11880_
	);
	LUT3 #(
		.INIT('h13)
	) name6054 (
		_w11711_,
		_w11880_,
		_w11870_,
		_w11881_
	);
	LUT4 #(
		.INIT('ha955)
	) name6055 (
		\u2_L4_reg[21]/NET0131 ,
		_w11869_,
		_w11879_,
		_w11881_,
		_w11882_
	);
	LUT4 #(
		.INIT('h004c)
	) name6056 (
		_w11519_,
		_w11505_,
		_w11509_,
		_w11598_,
		_w11883_
	);
	LUT4 #(
		.INIT('h0080)
	) name6057 (
		_w11497_,
		_w11493_,
		_w11496_,
		_w11494_,
		_w11884_
	);
	LUT3 #(
		.INIT('h07)
	) name6058 (
		_w11515_,
		_w11516_,
		_w11884_,
		_w11885_
	);
	LUT4 #(
		.INIT('h4080)
	) name6059 (
		_w11497_,
		_w11493_,
		_w11498_,
		_w11494_,
		_w11886_
	);
	LUT3 #(
		.INIT('h04)
	) name6060 (
		_w11493_,
		_w11496_,
		_w11494_,
		_w11887_
	);
	LUT4 #(
		.INIT('h0020)
	) name6061 (
		_w11497_,
		_w11493_,
		_w11496_,
		_w11494_,
		_w11888_
	);
	LUT4 #(
		.INIT('h00bf)
	) name6062 (
		_w11497_,
		_w11496_,
		_w11494_,
		_w11505_,
		_w11889_
	);
	LUT3 #(
		.INIT('h7e)
	) name6063 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11890_
	);
	LUT4 #(
		.INIT('h1000)
	) name6064 (
		_w11886_,
		_w11888_,
		_w11889_,
		_w11890_,
		_w11891_
	);
	LUT3 #(
		.INIT('h07)
	) name6065 (
		_w11883_,
		_w11885_,
		_w11891_,
		_w11892_
	);
	LUT4 #(
		.INIT('hef99)
	) name6066 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11893_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name6067 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w11894_
	);
	LUT4 #(
		.INIT('h0455)
	) name6068 (
		_w11497_,
		_w11505_,
		_w11893_,
		_w11894_,
		_w11895_
	);
	LUT2 #(
		.INIT('h4)
	) name6069 (
		_w11497_,
		_w11521_,
		_w11896_
	);
	LUT3 #(
		.INIT('h15)
	) name6070 (
		_w11524_,
		_w11499_,
		_w11887_,
		_w11897_
	);
	LUT3 #(
		.INIT('h10)
	) name6071 (
		_w11895_,
		_w11896_,
		_w11897_,
		_w11898_
	);
	LUT3 #(
		.INIT('h9a)
	) name6072 (
		\u2_L4_reg[23]/NET0131 ,
		_w11892_,
		_w11898_,
		_w11899_
	);
	LUT4 #(
		.INIT('h0010)
	) name6073 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11900_
	);
	LUT4 #(
		.INIT('h070f)
	) name6074 (
		_w11609_,
		_w11610_,
		_w11611_,
		_w11616_,
		_w11901_
	);
	LUT3 #(
		.INIT('h45)
	) name6075 (
		_w11623_,
		_w11900_,
		_w11901_,
		_w11902_
	);
	LUT4 #(
		.INIT('h0002)
	) name6076 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11903_
	);
	LUT4 #(
		.INIT('hc7d7)
	) name6077 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11611_,
		_w11904_
	);
	LUT3 #(
		.INIT('h31)
	) name6078 (
		_w11616_,
		_w11903_,
		_w11904_,
		_w11905_
	);
	LUT3 #(
		.INIT('h8a)
	) name6079 (
		_w11613_,
		_w11902_,
		_w11905_,
		_w11906_
	);
	LUT4 #(
		.INIT('h0086)
	) name6080 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11611_,
		_w11907_
	);
	LUT3 #(
		.INIT('h9b)
	) name6081 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11908_
	);
	LUT3 #(
		.INIT('h70)
	) name6082 (
		_w11610_,
		_w11611_,
		_w11613_,
		_w11909_
	);
	LUT4 #(
		.INIT('h4445)
	) name6083 (
		_w11616_,
		_w11907_,
		_w11908_,
		_w11909_,
		_w11910_
	);
	LUT4 #(
		.INIT('heafa)
	) name6084 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11616_,
		_w11911_
	);
	LUT2 #(
		.INIT('h1)
	) name6085 (
		_w11611_,
		_w11911_,
		_w11912_
	);
	LUT3 #(
		.INIT('h8a)
	) name6086 (
		_w11608_,
		_w11609_,
		_w11610_,
		_w11913_
	);
	LUT3 #(
		.INIT('h15)
	) name6087 (
		_w11614_,
		_w11628_,
		_w11913_,
		_w11914_
	);
	LUT4 #(
		.INIT('h2322)
	) name6088 (
		_w11613_,
		_w11910_,
		_w11912_,
		_w11914_,
		_w11915_
	);
	LUT3 #(
		.INIT('h65)
	) name6089 (
		\u2_L4_reg[26]/NET0131 ,
		_w11906_,
		_w11915_,
		_w11916_
	);
	LUT4 #(
		.INIT('h5515)
	) name6090 (
		_w11801_,
		_w11803_,
		_w11804_,
		_w11805_,
		_w11917_
	);
	LUT4 #(
		.INIT('h1105)
	) name6091 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11918_
	);
	LUT4 #(
		.INIT('h2aa0)
	) name6092 (
		_w11801_,
		_w11803_,
		_w11804_,
		_w11805_,
		_w11919_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6093 (
		_w11815_,
		_w11917_,
		_w11918_,
		_w11919_,
		_w11920_
	);
	LUT4 #(
		.INIT('h4000)
	) name6094 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11921_
	);
	LUT4 #(
		.INIT('hf700)
	) name6095 (
		_w11803_,
		_w11805_,
		_w11802_,
		_w11800_,
		_w11922_
	);
	LUT2 #(
		.INIT('h4)
	) name6096 (
		_w11921_,
		_w11922_,
		_w11923_
	);
	LUT3 #(
		.INIT('h8a)
	) name6097 (
		_w11801_,
		_w11803_,
		_w11805_,
		_w11924_
	);
	LUT4 #(
		.INIT('h00ab)
	) name6098 (
		_w11801_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11925_
	);
	LUT2 #(
		.INIT('h4)
	) name6099 (
		_w11924_,
		_w11925_,
		_w11926_
	);
	LUT2 #(
		.INIT('h2)
	) name6100 (
		_w11801_,
		_w11803_,
		_w11927_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name6101 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11928_
	);
	LUT3 #(
		.INIT('h54)
	) name6102 (
		_w11800_,
		_w11927_,
		_w11928_,
		_w11929_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6103 (
		_w11920_,
		_w11923_,
		_w11926_,
		_w11929_,
		_w11930_
	);
	LUT4 #(
		.INIT('hbefd)
	) name6104 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11931_
	);
	LUT4 #(
		.INIT('h0400)
	) name6105 (
		_w11801_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11932_
	);
	LUT4 #(
		.INIT('h0031)
	) name6106 (
		_w11801_,
		_w11807_,
		_w11931_,
		_w11932_,
		_w11933_
	);
	LUT3 #(
		.INIT('h65)
	) name6107 (
		\u2_L4_reg[25]/NET0131 ,
		_w11930_,
		_w11933_,
		_w11934_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name6108 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11935_
	);
	LUT2 #(
		.INIT('h8)
	) name6109 (
		_w11659_,
		_w11935_,
		_w11936_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name6110 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11937_
	);
	LUT3 #(
		.INIT('h10)
	) name6111 (
		_w11652_,
		_w11654_,
		_w11657_,
		_w11938_
	);
	LUT4 #(
		.INIT('h0001)
	) name6112 (
		_w11655_,
		_w11659_,
		_w11762_,
		_w11938_,
		_w11939_
	);
	LUT4 #(
		.INIT('h6100)
	) name6113 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11940_
	);
	LUT2 #(
		.INIT('h1)
	) name6114 (
		_w11651_,
		_w11940_,
		_w11941_
	);
	LUT4 #(
		.INIT('hba00)
	) name6115 (
		_w11936_,
		_w11937_,
		_w11939_,
		_w11941_,
		_w11942_
	);
	LUT4 #(
		.INIT('h0010)
	) name6116 (
		_w11659_,
		_w11762_,
		_w11935_,
		_w11938_,
		_w11943_
	);
	LUT4 #(
		.INIT('h8280)
	) name6117 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w11944_
	);
	LUT4 #(
		.INIT('hef00)
	) name6118 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11659_,
		_w11945_
	);
	LUT2 #(
		.INIT('h4)
	) name6119 (
		_w11944_,
		_w11945_,
		_w11946_
	);
	LUT3 #(
		.INIT('h0b)
	) name6120 (
		_w11652_,
		_w11653_,
		_w11659_,
		_w11947_
	);
	LUT2 #(
		.INIT('h2)
	) name6121 (
		_w11654_,
		_w11657_,
		_w11948_
	);
	LUT4 #(
		.INIT('h2022)
	) name6122 (
		_w11651_,
		_w11764_,
		_w11947_,
		_w11948_,
		_w11949_
	);
	LUT3 #(
		.INIT('he0)
	) name6123 (
		_w11943_,
		_w11946_,
		_w11949_,
		_w11950_
	);
	LUT3 #(
		.INIT('ha9)
	) name6124 (
		\u2_L4_reg[28]/NET0131 ,
		_w11942_,
		_w11950_,
		_w11951_
	);
	LUT3 #(
		.INIT('h02)
	) name6125 (
		_w11801_,
		_w11824_,
		_w11806_,
		_w11952_
	);
	LUT4 #(
		.INIT('h2022)
	) name6126 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11953_
	);
	LUT2 #(
		.INIT('h2)
	) name6127 (
		_w11917_,
		_w11953_,
		_w11954_
	);
	LUT4 #(
		.INIT('hbecf)
	) name6128 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11955_
	);
	LUT4 #(
		.INIT('h0155)
	) name6129 (
		_w11800_,
		_w11952_,
		_w11954_,
		_w11955_,
		_w11956_
	);
	LUT4 #(
		.INIT('hf7f6)
	) name6130 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11957_
	);
	LUT3 #(
		.INIT('h04)
	) name6131 (
		_w11801_,
		_w11804_,
		_w11802_,
		_w11958_
	);
	LUT4 #(
		.INIT('h0031)
	) name6132 (
		_w11801_,
		_w11829_,
		_w11957_,
		_w11958_,
		_w11959_
	);
	LUT4 #(
		.INIT('haddf)
	) name6133 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11960_
	);
	LUT3 #(
		.INIT('hb1)
	) name6134 (
		_w11801_,
		_w11821_,
		_w11960_,
		_w11961_
	);
	LUT3 #(
		.INIT('hd0)
	) name6135 (
		_w11800_,
		_w11959_,
		_w11961_,
		_w11962_
	);
	LUT3 #(
		.INIT('h65)
	) name6136 (
		\u2_L4_reg[8]/NET0131 ,
		_w11956_,
		_w11962_,
		_w11963_
	);
	LUT4 #(
		.INIT('hd7d2)
	) name6137 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11964_
	);
	LUT2 #(
		.INIT('h1)
	) name6138 (
		_w11701_,
		_w11964_,
		_w11965_
	);
	LUT3 #(
		.INIT('hb0)
	) name6139 (
		_w11704_,
		_w11702_,
		_w11701_,
		_w11966_
	);
	LUT4 #(
		.INIT('he7bb)
	) name6140 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11967_
	);
	LUT3 #(
		.INIT('hb0)
	) name6141 (
		_w11787_,
		_w11966_,
		_w11967_,
		_w11968_
	);
	LUT3 #(
		.INIT('h8a)
	) name6142 (
		_w11700_,
		_w11965_,
		_w11968_,
		_w11969_
	);
	LUT4 #(
		.INIT('hce44)
	) name6143 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11970_
	);
	LUT4 #(
		.INIT('hfd00)
	) name6144 (
		_w11703_,
		_w11704_,
		_w11705_,
		_w11701_,
		_w11971_
	);
	LUT2 #(
		.INIT('h4)
	) name6145 (
		_w11970_,
		_w11971_,
		_w11972_
	);
	LUT4 #(
		.INIT('h0080)
	) name6146 (
		_w11704_,
		_w11702_,
		_w11705_,
		_w11701_,
		_w11973_
	);
	LUT3 #(
		.INIT('h01)
	) name6147 (
		_w11719_,
		_w11877_,
		_w11973_,
		_w11974_
	);
	LUT4 #(
		.INIT('h1000)
	) name6148 (
		_w11703_,
		_w11704_,
		_w11705_,
		_w11701_,
		_w11975_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name6149 (
		_w11703_,
		_w11704_,
		_w11702_,
		_w11705_,
		_w11976_
	);
	LUT3 #(
		.INIT('h32)
	) name6150 (
		_w11701_,
		_w11975_,
		_w11976_,
		_w11977_
	);
	LUT4 #(
		.INIT('hba00)
	) name6151 (
		_w11700_,
		_w11972_,
		_w11974_,
		_w11977_,
		_w11978_
	);
	LUT3 #(
		.INIT('h65)
	) name6152 (
		\u2_L4_reg[27]/NET0131 ,
		_w11969_,
		_w11978_,
		_w11979_
	);
	LUT4 #(
		.INIT('hb005)
	) name6153 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11980_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name6154 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11981_
	);
	LUT3 #(
		.INIT('h01)
	) name6155 (
		_w11560_,
		_w11981_,
		_w11980_,
		_w11982_
	);
	LUT4 #(
		.INIT('hddfa)
	) name6156 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11983_
	);
	LUT3 #(
		.INIT('h08)
	) name6157 (
		_w11562_,
		_w11563_,
		_w11564_,
		_w11984_
	);
	LUT4 #(
		.INIT('h11f5)
	) name6158 (
		_w11560_,
		_w11561_,
		_w11983_,
		_w11984_,
		_w11985_
	);
	LUT3 #(
		.INIT('h8a)
	) name6159 (
		_w11559_,
		_w11982_,
		_w11985_,
		_w11986_
	);
	LUT3 #(
		.INIT('h4c)
	) name6160 (
		_w11561_,
		_w11563_,
		_w11564_,
		_w11987_
	);
	LUT4 #(
		.INIT('h2808)
	) name6161 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11988_
	);
	LUT4 #(
		.INIT('h5504)
	) name6162 (
		_w11560_,
		_w11752_,
		_w11753_,
		_w11988_,
		_w11989_
	);
	LUT2 #(
		.INIT('h2)
	) name6163 (
		_w11559_,
		_w11560_,
		_w11990_
	);
	LUT2 #(
		.INIT('h2)
	) name6164 (
		_w11571_,
		_w11990_,
		_w11991_
	);
	LUT4 #(
		.INIT('h8008)
	) name6165 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w11992_
	);
	LUT4 #(
		.INIT('hee0e)
	) name6166 (
		_w11560_,
		_w11561_,
		_w11562_,
		_w11564_,
		_w11993_
	);
	LUT4 #(
		.INIT('h5450)
	) name6167 (
		_w11559_,
		_w11987_,
		_w11992_,
		_w11993_,
		_w11994_
	);
	LUT3 #(
		.INIT('h01)
	) name6168 (
		_w11991_,
		_w11989_,
		_w11994_,
		_w11995_
	);
	LUT3 #(
		.INIT('h65)
	) name6169 (
		\u2_L4_reg[32]/NET0131 ,
		_w11986_,
		_w11995_,
		_w11996_
	);
	LUT3 #(
		.INIT('h04)
	) name6170 (
		_w11821_,
		_w11800_,
		_w11807_,
		_w11997_
	);
	LUT4 #(
		.INIT('h0400)
	) name6171 (
		_w11801_,
		_w11803_,
		_w11804_,
		_w11805_,
		_w11998_
	);
	LUT4 #(
		.INIT('hcf45)
	) name6172 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w11999_
	);
	LUT3 #(
		.INIT('ha2)
	) name6173 (
		_w11801_,
		_w11803_,
		_w11804_,
		_w12000_
	);
	LUT3 #(
		.INIT('h45)
	) name6174 (
		_w11998_,
		_w11999_,
		_w12000_,
		_w12001_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name6175 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w12002_
	);
	LUT2 #(
		.INIT('h2)
	) name6176 (
		_w11801_,
		_w12002_,
		_w12003_
	);
	LUT3 #(
		.INIT('h8a)
	) name6177 (
		_w11801_,
		_w11805_,
		_w11802_,
		_w12004_
	);
	LUT4 #(
		.INIT('h44e6)
	) name6178 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w12005_
	);
	LUT3 #(
		.INIT('h54)
	) name6179 (
		_w11800_,
		_w12004_,
		_w12005_,
		_w12006_
	);
	LUT4 #(
		.INIT('h7077)
	) name6180 (
		_w11997_,
		_w12001_,
		_w12003_,
		_w12006_,
		_w12007_
	);
	LUT3 #(
		.INIT('h02)
	) name6181 (
		_w11801_,
		_w11806_,
		_w11828_,
		_w12008_
	);
	LUT4 #(
		.INIT('hffbe)
	) name6182 (
		_w11803_,
		_w11804_,
		_w11805_,
		_w11802_,
		_w12009_
	);
	LUT3 #(
		.INIT('he0)
	) name6183 (
		_w11818_,
		_w11917_,
		_w12009_,
		_w12010_
	);
	LUT2 #(
		.INIT('h1)
	) name6184 (
		_w12008_,
		_w12010_,
		_w12011_
	);
	LUT3 #(
		.INIT('h56)
	) name6185 (
		\u2_L4_reg[3]/NET0131 ,
		_w12007_,
		_w12011_,
		_w12012_
	);
	LUT4 #(
		.INIT('hc963)
	) name6186 (
		decrypt_pad,
		\u2_R4_reg[11]/NET0131 ,
		\u2_uk_K_r4_reg[40]/NET0131 ,
		\u2_uk_K_r4_reg[46]/NET0131 ,
		_w12013_
	);
	LUT4 #(
		.INIT('hc693)
	) name6187 (
		decrypt_pad,
		\u2_R4_reg[12]/NET0131 ,
		\u2_uk_K_r4_reg[4]/NET0131 ,
		\u2_uk_K_r4_reg[55]/NET0131 ,
		_w12014_
	);
	LUT4 #(
		.INIT('hc963)
	) name6188 (
		decrypt_pad,
		\u2_R4_reg[13]/NET0131 ,
		\u2_uk_K_r4_reg[11]/NET0131 ,
		\u2_uk_K_r4_reg[17]/NET0131 ,
		_w12015_
	);
	LUT4 #(
		.INIT('hc693)
	) name6189 (
		decrypt_pad,
		\u2_R4_reg[9]/NET0131 ,
		\u2_uk_K_r4_reg[12]/NET0131 ,
		\u2_uk_K_r4_reg[6]/NET0131 ,
		_w12016_
	);
	LUT4 #(
		.INIT('hc963)
	) name6190 (
		decrypt_pad,
		\u2_R4_reg[8]/NET0131 ,
		\u2_uk_K_r4_reg[34]/NET0131 ,
		\u2_uk_K_r4_reg[40]/NET0131 ,
		_w12017_
	);
	LUT2 #(
		.INIT('h2)
	) name6191 (
		_w12015_,
		_w12017_,
		_w12018_
	);
	LUT4 #(
		.INIT('hc693)
	) name6192 (
		decrypt_pad,
		\u2_R4_reg[10]/NET0131 ,
		\u2_uk_K_r4_reg[20]/NET0131 ,
		\u2_uk_K_r4_reg[39]/NET0131 ,
		_w12019_
	);
	LUT4 #(
		.INIT('h95b5)
	) name6193 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12020_
	);
	LUT4 #(
		.INIT('h0001)
	) name6194 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12021_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name6195 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12022_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6196 (
		_w12014_,
		_w12013_,
		_w12020_,
		_w12022_,
		_w12023_
	);
	LUT4 #(
		.INIT('h0900)
	) name6197 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12024_
	);
	LUT3 #(
		.INIT('h20)
	) name6198 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12025_
	);
	LUT2 #(
		.INIT('h4)
	) name6199 (
		_w12013_,
		_w12019_,
		_w12026_
	);
	LUT4 #(
		.INIT('h4000)
	) name6200 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12027_
	);
	LUT4 #(
		.INIT('h0007)
	) name6201 (
		_w12025_,
		_w12026_,
		_w12024_,
		_w12027_,
		_w12028_
	);
	LUT2 #(
		.INIT('h1)
	) name6202 (
		_w12016_,
		_w12019_,
		_w12029_
	);
	LUT2 #(
		.INIT('h8)
	) name6203 (
		_w12015_,
		_w12013_,
		_w12030_
	);
	LUT3 #(
		.INIT('h46)
	) name6204 (
		_w12015_,
		_w12017_,
		_w12013_,
		_w12031_
	);
	LUT2 #(
		.INIT('h8)
	) name6205 (
		_w12029_,
		_w12031_,
		_w12032_
	);
	LUT3 #(
		.INIT('hed)
	) name6206 (
		_w12016_,
		_w12019_,
		_w12031_,
		_w12033_
	);
	LUT2 #(
		.INIT('h8)
	) name6207 (
		_w12014_,
		_w12019_,
		_w12034_
	);
	LUT3 #(
		.INIT('h10)
	) name6208 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12035_
	);
	LUT3 #(
		.INIT('h51)
	) name6209 (
		_w12017_,
		_w12016_,
		_w12019_,
		_w12036_
	);
	LUT2 #(
		.INIT('h2)
	) name6210 (
		_w12014_,
		_w12013_,
		_w12037_
	);
	LUT4 #(
		.INIT('h0082)
	) name6211 (
		_w12014_,
		_w12015_,
		_w12016_,
		_w12013_,
		_w12038_
	);
	LUT4 #(
		.INIT('h7077)
	) name6212 (
		_w12034_,
		_w12035_,
		_w12036_,
		_w12038_,
		_w12039_
	);
	LUT4 #(
		.INIT('hea00)
	) name6213 (
		_w12014_,
		_w12028_,
		_w12033_,
		_w12039_,
		_w12040_
	);
	LUT3 #(
		.INIT('h65)
	) name6214 (
		\u2_L4_reg[6]/NET0131 ,
		_w12023_,
		_w12040_,
		_w12041_
	);
	LUT4 #(
		.INIT('h0770)
	) name6215 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w12042_
	);
	LUT4 #(
		.INIT('h3882)
	) name6216 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w12043_
	);
	LUT2 #(
		.INIT('h4)
	) name6217 (
		_w11559_,
		_w11560_,
		_w12044_
	);
	LUT2 #(
		.INIT('h9)
	) name6218 (
		_w11559_,
		_w11560_,
		_w12045_
	);
	LUT3 #(
		.INIT('h10)
	) name6219 (
		_w11750_,
		_w12043_,
		_w12045_,
		_w12046_
	);
	LUT4 #(
		.INIT('h800c)
	) name6220 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w12047_
	);
	LUT3 #(
		.INIT('h02)
	) name6221 (
		_w12044_,
		_w12042_,
		_w12047_,
		_w12048_
	);
	LUT4 #(
		.INIT('h0ae0)
	) name6222 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w11564_,
		_w12049_
	);
	LUT3 #(
		.INIT('h09)
	) name6223 (
		_w11561_,
		_w11562_,
		_w11563_,
		_w12050_
	);
	LUT4 #(
		.INIT('h0004)
	) name6224 (
		_w11750_,
		_w11990_,
		_w12050_,
		_w12049_,
		_w12051_
	);
	LUT4 #(
		.INIT('h00ab)
	) name6225 (
		_w11580_,
		_w12046_,
		_w12048_,
		_w12051_,
		_w12052_
	);
	LUT2 #(
		.INIT('h6)
	) name6226 (
		\u2_L4_reg[7]/NET0131 ,
		_w12052_,
		_w12053_
	);
	LUT4 #(
		.INIT('h9060)
	) name6227 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w12054_
	);
	LUT3 #(
		.INIT('he6)
	) name6228 (
		_w11493_,
		_w11496_,
		_w11494_,
		_w12055_
	);
	LUT4 #(
		.INIT('h0031)
	) name6229 (
		_w11499_,
		_w11601_,
		_w12055_,
		_w12054_,
		_w12056_
	);
	LUT4 #(
		.INIT('hf77f)
	) name6230 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w12057_
	);
	LUT2 #(
		.INIT('h1)
	) name6231 (
		_w11497_,
		_w12057_,
		_w12058_
	);
	LUT4 #(
		.INIT('h5414)
	) name6232 (
		_w11497_,
		_w11493_,
		_w11496_,
		_w11494_,
		_w12059_
	);
	LUT4 #(
		.INIT('h82a2)
	) name6233 (
		_w11497_,
		_w11493_,
		_w11496_,
		_w11498_,
		_w12060_
	);
	LUT4 #(
		.INIT('hd7ef)
	) name6234 (
		_w11493_,
		_w11496_,
		_w11498_,
		_w11494_,
		_w12061_
	);
	LUT4 #(
		.INIT('hdc00)
	) name6235 (
		_w11887_,
		_w12059_,
		_w12060_,
		_w12061_,
		_w12062_
	);
	LUT4 #(
		.INIT('h3210)
	) name6236 (
		_w11505_,
		_w12058_,
		_w12062_,
		_w12056_,
		_w12063_
	);
	LUT2 #(
		.INIT('h9)
	) name6237 (
		\u2_L4_reg[9]/NET0131 ,
		_w12063_,
		_w12064_
	);
	LUT3 #(
		.INIT('h80)
	) name6238 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12065_
	);
	LUT3 #(
		.INIT('h68)
	) name6239 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12066_
	);
	LUT4 #(
		.INIT('h0111)
	) name6240 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12013_,
		_w12067_
	);
	LUT3 #(
		.INIT('h01)
	) name6241 (
		_w12019_,
		_w12067_,
		_w12066_,
		_w12068_
	);
	LUT4 #(
		.INIT('h0104)
	) name6242 (
		_w12015_,
		_w12017_,
		_w12013_,
		_w12019_,
		_w12069_
	);
	LUT4 #(
		.INIT('h2000)
	) name6243 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12070_
	);
	LUT3 #(
		.INIT('h02)
	) name6244 (
		_w12014_,
		_w12070_,
		_w12069_,
		_w12071_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name6245 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12072_
	);
	LUT2 #(
		.INIT('h1)
	) name6246 (
		_w12013_,
		_w12072_,
		_w12073_
	);
	LUT4 #(
		.INIT('h6800)
	) name6247 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12013_,
		_w12074_
	);
	LUT3 #(
		.INIT('h01)
	) name6248 (
		_w12014_,
		_w12021_,
		_w12074_,
		_w12075_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6249 (
		_w12068_,
		_w12071_,
		_w12073_,
		_w12075_,
		_w12076_
	);
	LUT3 #(
		.INIT('h20)
	) name6250 (
		_w12017_,
		_w12016_,
		_w12019_,
		_w12077_
	);
	LUT4 #(
		.INIT('h0200)
	) name6251 (
		_w12017_,
		_w12016_,
		_w12013_,
		_w12019_,
		_w12078_
	);
	LUT4 #(
		.INIT('hbeff)
	) name6252 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12079_
	);
	LUT3 #(
		.INIT('h31)
	) name6253 (
		_w12013_,
		_w12078_,
		_w12079_,
		_w12080_
	);
	LUT3 #(
		.INIT('h65)
	) name6254 (
		\u2_L4_reg[16]/NET0131 ,
		_w12076_,
		_w12080_,
		_w12081_
	);
	LUT4 #(
		.INIT('hef2f)
	) name6255 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w12082_
	);
	LUT4 #(
		.INIT('h0100)
	) name6256 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w12083_
	);
	LUT4 #(
		.INIT('h0b08)
	) name6257 (
		_w11656_,
		_w11659_,
		_w12083_,
		_w12082_,
		_w12084_
	);
	LUT4 #(
		.INIT('h0121)
	) name6258 (
		_w11652_,
		_w11654_,
		_w11657_,
		_w11659_,
		_w12085_
	);
	LUT4 #(
		.INIT('h9fff)
	) name6259 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w12086_
	);
	LUT4 #(
		.INIT('h8000)
	) name6260 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11659_,
		_w12087_
	);
	LUT4 #(
		.INIT('h0100)
	) name6261 (
		_w11777_,
		_w12087_,
		_w12085_,
		_w12086_,
		_w12088_
	);
	LUT4 #(
		.INIT('h0008)
	) name6262 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11659_,
		_w12089_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name6263 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11657_,
		_w12090_
	);
	LUT3 #(
		.INIT('h31)
	) name6264 (
		_w11659_,
		_w12089_,
		_w12090_,
		_w12091_
	);
	LUT4 #(
		.INIT('hd800)
	) name6265 (
		_w11651_,
		_w12084_,
		_w12088_,
		_w12091_,
		_w12092_
	);
	LUT2 #(
		.INIT('h9)
	) name6266 (
		\u2_L4_reg[18]/P0001 ,
		_w12092_,
		_w12093_
	);
	LUT4 #(
		.INIT('he2cd)
	) name6267 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12094_
	);
	LUT4 #(
		.INIT('h0400)
	) name6268 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12095_
	);
	LUT4 #(
		.INIT('h5504)
	) name6269 (
		_w12014_,
		_w12013_,
		_w12094_,
		_w12095_,
		_w12096_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name6270 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12097_
	);
	LUT3 #(
		.INIT('hc8)
	) name6271 (
		_w12016_,
		_w12013_,
		_w12019_,
		_w12098_
	);
	LUT4 #(
		.INIT('h0054)
	) name6272 (
		_w12018_,
		_w12013_,
		_w12097_,
		_w12098_,
		_w12099_
	);
	LUT3 #(
		.INIT('ha8)
	) name6273 (
		_w12014_,
		_w12032_,
		_w12099_,
		_w12100_
	);
	LUT4 #(
		.INIT('h1dff)
	) name6274 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12101_
	);
	LUT4 #(
		.INIT('hffdb)
	) name6275 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12102_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6276 (
		_w12014_,
		_w12013_,
		_w12101_,
		_w12102_,
		_w12103_
	);
	LUT4 #(
		.INIT('h9db6)
	) name6277 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12104_
	);
	LUT2 #(
		.INIT('h1)
	) name6278 (
		_w12014_,
		_w12013_,
		_w12105_
	);
	LUT4 #(
		.INIT('h7077)
	) name6279 (
		_w12026_,
		_w12065_,
		_w12104_,
		_w12105_,
		_w12106_
	);
	LUT2 #(
		.INIT('h4)
	) name6280 (
		_w12103_,
		_w12106_,
		_w12107_
	);
	LUT4 #(
		.INIT('h5655)
	) name6281 (
		\u2_L4_reg[24]/NET0131 ,
		_w12096_,
		_w12100_,
		_w12107_,
		_w12108_
	);
	LUT4 #(
		.INIT('h73af)
	) name6282 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12109_
	);
	LUT3 #(
		.INIT('h0b)
	) name6283 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12110_
	);
	LUT4 #(
		.INIT('h22ad)
	) name6284 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12111_
	);
	LUT4 #(
		.INIT('h08dd)
	) name6285 (
		_w12013_,
		_w12109_,
		_w12110_,
		_w12111_,
		_w12112_
	);
	LUT2 #(
		.INIT('h1)
	) name6286 (
		_w12014_,
		_w12112_,
		_w12113_
	);
	LUT4 #(
		.INIT('heed9)
	) name6287 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12114_
	);
	LUT2 #(
		.INIT('h8)
	) name6288 (
		_w12014_,
		_w12013_,
		_w12115_
	);
	LUT2 #(
		.INIT('h4)
	) name6289 (
		_w12114_,
		_w12115_,
		_w12116_
	);
	LUT4 #(
		.INIT('h23ef)
	) name6290 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12019_,
		_w12117_
	);
	LUT2 #(
		.INIT('h2)
	) name6291 (
		_w12037_,
		_w12117_,
		_w12118_
	);
	LUT3 #(
		.INIT('h70)
	) name6292 (
		_w12015_,
		_w12017_,
		_w12016_,
		_w12119_
	);
	LUT2 #(
		.INIT('h8)
	) name6293 (
		_w12034_,
		_w12119_,
		_w12120_
	);
	LUT4 #(
		.INIT('h0400)
	) name6294 (
		_w12015_,
		_w12016_,
		_w12013_,
		_w12019_,
		_w12121_
	);
	LUT3 #(
		.INIT('h07)
	) name6295 (
		_w12030_,
		_w12077_,
		_w12121_,
		_w12122_
	);
	LUT4 #(
		.INIT('h0100)
	) name6296 (
		_w12118_,
		_w12120_,
		_w12116_,
		_w12122_,
		_w12123_
	);
	LUT3 #(
		.INIT('h9a)
	) name6297 (
		\u2_L4_reg[30]/NET0131 ,
		_w12113_,
		_w12123_,
		_w12124_
	);
	LUT4 #(
		.INIT('hc693)
	) name6298 (
		decrypt_pad,
		\u2_R3_reg[27]/NET0131 ,
		\u2_uk_K_r3_reg[30]/NET0131 ,
		\u2_uk_K_r3_reg[49]/NET0131 ,
		_w12125_
	);
	LUT4 #(
		.INIT('hc963)
	) name6299 (
		decrypt_pad,
		\u2_R3_reg[25]/NET0131 ,
		\u2_uk_K_r3_reg[0]/NET0131 ,
		\u2_uk_K_r3_reg[36]/NET0131 ,
		_w12126_
	);
	LUT4 #(
		.INIT('hc963)
	) name6300 (
		decrypt_pad,
		\u2_R3_reg[26]/NET0131 ,
		\u2_uk_K_r3_reg[16]/NET0131 ,
		\u2_uk_K_r3_reg[21]/NET0131 ,
		_w12127_
	);
	LUT4 #(
		.INIT('hc693)
	) name6301 (
		decrypt_pad,
		\u2_R3_reg[24]/NET0131 ,
		\u2_uk_K_r3_reg[1]/NET0131 ,
		\u2_uk_K_r3_reg[51]/NET0131 ,
		_w12128_
	);
	LUT4 #(
		.INIT('hc963)
	) name6302 (
		decrypt_pad,
		\u2_R3_reg[29]/NET0131 ,
		\u2_uk_K_r3_reg[28]/NET0131 ,
		\u2_uk_K_r3_reg[9]/NET0131 ,
		_w12129_
	);
	LUT3 #(
		.INIT('h02)
	) name6303 (
		_w12127_,
		_w12128_,
		_w12129_,
		_w12130_
	);
	LUT4 #(
		.INIT('h0002)
	) name6304 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12131_
	);
	LUT2 #(
		.INIT('h6)
	) name6305 (
		_w12127_,
		_w12128_,
		_w12132_
	);
	LUT4 #(
		.INIT('h5a2d)
	) name6306 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12133_
	);
	LUT4 #(
		.INIT('h0200)
	) name6307 (
		_w12125_,
		_w12127_,
		_w12126_,
		_w12128_,
		_w12134_
	);
	LUT4 #(
		.INIT('h8400)
	) name6308 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12135_
	);
	LUT4 #(
		.INIT('h000e)
	) name6309 (
		_w12125_,
		_w12133_,
		_w12134_,
		_w12135_,
		_w12136_
	);
	LUT4 #(
		.INIT('hc963)
	) name6310 (
		decrypt_pad,
		\u2_R3_reg[28]/NET0131 ,
		\u2_uk_K_r3_reg[36]/NET0131 ,
		\u2_uk_K_r3_reg[45]/P0001 ,
		_w12137_
	);
	LUT2 #(
		.INIT('h1)
	) name6311 (
		_w12136_,
		_w12137_,
		_w12138_
	);
	LUT4 #(
		.INIT('h1000)
	) name6312 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12139_
	);
	LUT2 #(
		.INIT('h4)
	) name6313 (
		_w12128_,
		_w12129_,
		_w12140_
	);
	LUT4 #(
		.INIT('he3ff)
	) name6314 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12141_
	);
	LUT2 #(
		.INIT('h1)
	) name6315 (
		_w12125_,
		_w12141_,
		_w12142_
	);
	LUT2 #(
		.INIT('h6)
	) name6316 (
		_w12127_,
		_w12126_,
		_w12143_
	);
	LUT4 #(
		.INIT('ha080)
	) name6317 (
		_w12125_,
		_w12127_,
		_w12128_,
		_w12129_,
		_w12144_
	);
	LUT4 #(
		.INIT('h0200)
	) name6318 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12145_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name6319 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12146_
	);
	LUT3 #(
		.INIT('h70)
	) name6320 (
		_w12143_,
		_w12144_,
		_w12146_,
		_w12147_
	);
	LUT4 #(
		.INIT('h0008)
	) name6321 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12148_
	);
	LUT4 #(
		.INIT('hfdc7)
	) name6322 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12149_
	);
	LUT4 #(
		.INIT('h4010)
	) name6323 (
		_w12125_,
		_w12127_,
		_w12126_,
		_w12128_,
		_w12150_
	);
	LUT4 #(
		.INIT('h0002)
	) name6324 (
		_w12125_,
		_w12127_,
		_w12126_,
		_w12129_,
		_w12151_
	);
	LUT4 #(
		.INIT('h0031)
	) name6325 (
		_w12125_,
		_w12150_,
		_w12149_,
		_w12151_,
		_w12152_
	);
	LUT4 #(
		.INIT('h7500)
	) name6326 (
		_w12137_,
		_w12142_,
		_w12147_,
		_w12152_,
		_w12153_
	);
	LUT3 #(
		.INIT('h65)
	) name6327 (
		\u2_L3_reg[22]/NET0131 ,
		_w12138_,
		_w12153_,
		_w12154_
	);
	LUT4 #(
		.INIT('hc693)
	) name6328 (
		decrypt_pad,
		\u2_R3_reg[4]/NET0131 ,
		\u2_uk_K_r3_reg[39]/NET0131 ,
		\u2_uk_K_r3_reg[5]/NET0131 ,
		_w12155_
	);
	LUT4 #(
		.INIT('hc963)
	) name6329 (
		decrypt_pad,
		\u2_R3_reg[3]/NET0131 ,
		\u2_uk_K_r3_reg[27]/NET0131 ,
		\u2_uk_K_r3_reg[4]/NET0131 ,
		_w12156_
	);
	LUT4 #(
		.INIT('hc963)
	) name6330 (
		decrypt_pad,
		\u2_R3_reg[2]/NET0131 ,
		\u2_uk_K_r3_reg[18]/NET0131 ,
		\u2_uk_K_r3_reg[27]/NET0131 ,
		_w12157_
	);
	LUT4 #(
		.INIT('hc963)
	) name6331 (
		decrypt_pad,
		\u2_R3_reg[32]/NET0131 ,
		\u2_uk_K_r3_reg[39]/NET0131 ,
		\u2_uk_K_r3_reg[48]/NET0131 ,
		_w12158_
	);
	LUT4 #(
		.INIT('hc693)
	) name6332 (
		decrypt_pad,
		\u2_R3_reg[1]/NET0131 ,
		\u2_uk_K_r3_reg[12]/NET0131 ,
		\u2_uk_K_r3_reg[3]/NET0131 ,
		_w12159_
	);
	LUT4 #(
		.INIT('hc693)
	) name6333 (
		decrypt_pad,
		\u2_R3_reg[5]/NET0131 ,
		\u2_uk_K_r3_reg[10]/NET0131 ,
		\u2_uk_K_r3_reg[33]/NET0131 ,
		_w12160_
	);
	LUT4 #(
		.INIT('hfdba)
	) name6334 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12161_
	);
	LUT2 #(
		.INIT('h1)
	) name6335 (
		_w12156_,
		_w12161_,
		_w12162_
	);
	LUT2 #(
		.INIT('h2)
	) name6336 (
		_w12160_,
		_w12158_,
		_w12163_
	);
	LUT4 #(
		.INIT('h0800)
	) name6337 (
		_w12157_,
		_w12160_,
		_w12158_,
		_w12156_,
		_w12164_
	);
	LUT4 #(
		.INIT('hf6fe)
	) name6338 (
		_w12157_,
		_w12160_,
		_w12158_,
		_w12156_,
		_w12165_
	);
	LUT2 #(
		.INIT('h2)
	) name6339 (
		_w12159_,
		_w12165_,
		_w12166_
	);
	LUT4 #(
		.INIT('h0800)
	) name6340 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12167_
	);
	LUT2 #(
		.INIT('h8)
	) name6341 (
		_w12160_,
		_w12158_,
		_w12168_
	);
	LUT2 #(
		.INIT('h4)
	) name6342 (
		_w12157_,
		_w12156_,
		_w12169_
	);
	LUT3 #(
		.INIT('hae)
	) name6343 (
		_w12157_,
		_w12159_,
		_w12156_,
		_w12170_
	);
	LUT4 #(
		.INIT('h7707)
	) name6344 (
		_w12167_,
		_w12156_,
		_w12168_,
		_w12170_,
		_w12171_
	);
	LUT4 #(
		.INIT('h5455)
	) name6345 (
		_w12155_,
		_w12162_,
		_w12166_,
		_w12171_,
		_w12172_
	);
	LUT3 #(
		.INIT('h02)
	) name6346 (
		_w12157_,
		_w12160_,
		_w12158_,
		_w12173_
	);
	LUT4 #(
		.INIT('hcfc5)
	) name6347 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12174_
	);
	LUT2 #(
		.INIT('h2)
	) name6348 (
		_w12156_,
		_w12174_,
		_w12175_
	);
	LUT3 #(
		.INIT('h8c)
	) name6349 (
		_w12157_,
		_w12159_,
		_w12156_,
		_w12176_
	);
	LUT4 #(
		.INIT('h0100)
	) name6350 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12177_
	);
	LUT2 #(
		.INIT('h2)
	) name6351 (
		_w12158_,
		_w12156_,
		_w12178_
	);
	LUT4 #(
		.INIT('h02c2)
	) name6352 (
		_w12157_,
		_w12159_,
		_w12158_,
		_w12156_,
		_w12179_
	);
	LUT4 #(
		.INIT('h0301)
	) name6353 (
		_w12163_,
		_w12177_,
		_w12179_,
		_w12176_,
		_w12180_
	);
	LUT2 #(
		.INIT('h4)
	) name6354 (
		_w12159_,
		_w12156_,
		_w12181_
	);
	LUT3 #(
		.INIT('had)
	) name6355 (
		_w12157_,
		_w12160_,
		_w12158_,
		_w12182_
	);
	LUT3 #(
		.INIT('h80)
	) name6356 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12183_
	);
	LUT4 #(
		.INIT('h7bdb)
	) name6357 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12184_
	);
	LUT4 #(
		.INIT('hfbc8)
	) name6358 (
		_w12159_,
		_w12156_,
		_w12182_,
		_w12184_,
		_w12185_
	);
	LUT4 #(
		.INIT('h7500)
	) name6359 (
		_w12155_,
		_w12175_,
		_w12180_,
		_w12185_,
		_w12186_
	);
	LUT3 #(
		.INIT('h65)
	) name6360 (
		\u2_L3_reg[31]/NET0131 ,
		_w12172_,
		_w12186_,
		_w12187_
	);
	LUT4 #(
		.INIT('hc963)
	) name6361 (
		decrypt_pad,
		\u2_R3_reg[24]/NET0131 ,
		\u2_uk_K_r3_reg[29]/NET0131 ,
		\u2_uk_K_r3_reg[38]/NET0131 ,
		_w12188_
	);
	LUT4 #(
		.INIT('hc693)
	) name6362 (
		decrypt_pad,
		\u2_R3_reg[20]/NET0131 ,
		\u2_uk_K_r3_reg[44]/NET0131 ,
		\u2_uk_K_r3_reg[8]/NET0131 ,
		_w12189_
	);
	LUT4 #(
		.INIT('hc963)
	) name6363 (
		decrypt_pad,
		\u2_R3_reg[22]/NET0131 ,
		\u2_uk_K_r3_reg[14]/NET0131 ,
		\u2_uk_K_r3_reg[50]/NET0131 ,
		_w12190_
	);
	LUT4 #(
		.INIT('hc963)
	) name6364 (
		decrypt_pad,
		\u2_R3_reg[21]/NET0131 ,
		\u2_uk_K_r3_reg[23]/NET0131 ,
		\u2_uk_K_r3_reg[28]/NET0131 ,
		_w12191_
	);
	LUT4 #(
		.INIT('hc963)
	) name6365 (
		decrypt_pad,
		\u2_R3_reg[23]/NET0131 ,
		\u2_uk_K_r3_reg[31]/NET0131 ,
		\u2_uk_K_r3_reg[8]/NET0131 ,
		_w12192_
	);
	LUT4 #(
		.INIT('h4155)
	) name6366 (
		_w12192_,
		_w12189_,
		_w12190_,
		_w12191_,
		_w12193_
	);
	LUT4 #(
		.INIT('hc693)
	) name6367 (
		decrypt_pad,
		\u2_R3_reg[25]/NET0131 ,
		\u2_uk_K_r3_reg[29]/NET0131 ,
		\u2_uk_K_r3_reg[52]/NET0131 ,
		_w12194_
	);
	LUT4 #(
		.INIT('haa8a)
	) name6368 (
		_w12192_,
		_w12189_,
		_w12194_,
		_w12191_,
		_w12195_
	);
	LUT3 #(
		.INIT('he6)
	) name6369 (
		_w12189_,
		_w12190_,
		_w12191_,
		_w12196_
	);
	LUT3 #(
		.INIT('h13)
	) name6370 (
		_w12195_,
		_w12193_,
		_w12196_,
		_w12197_
	);
	LUT4 #(
		.INIT('h0080)
	) name6371 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12198_
	);
	LUT2 #(
		.INIT('h2)
	) name6372 (
		_w12189_,
		_w12194_,
		_w12199_
	);
	LUT2 #(
		.INIT('h1)
	) name6373 (
		_w12192_,
		_w12190_,
		_w12200_
	);
	LUT3 #(
		.INIT('hce)
	) name6374 (
		_w12192_,
		_w12190_,
		_w12191_,
		_w12201_
	);
	LUT3 #(
		.INIT('h31)
	) name6375 (
		_w12199_,
		_w12198_,
		_w12201_,
		_w12202_
	);
	LUT3 #(
		.INIT('h45)
	) name6376 (
		_w12188_,
		_w12197_,
		_w12202_,
		_w12203_
	);
	LUT4 #(
		.INIT('h0002)
	) name6377 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12204_
	);
	LUT4 #(
		.INIT('h27fd)
	) name6378 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12205_
	);
	LUT2 #(
		.INIT('h2)
	) name6379 (
		_w12192_,
		_w12205_,
		_w12206_
	);
	LUT4 #(
		.INIT('h0415)
	) name6380 (
		_w12192_,
		_w12189_,
		_w12194_,
		_w12191_,
		_w12207_
	);
	LUT4 #(
		.INIT('h0b07)
	) name6381 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12208_
	);
	LUT3 #(
		.INIT('h0e)
	) name6382 (
		_w12200_,
		_w12207_,
		_w12208_,
		_w12209_
	);
	LUT3 #(
		.INIT('he0)
	) name6383 (
		_w12206_,
		_w12209_,
		_w12188_,
		_w12210_
	);
	LUT4 #(
		.INIT('h5155)
	) name6384 (
		_w12192_,
		_w12189_,
		_w12194_,
		_w12191_,
		_w12211_
	);
	LUT3 #(
		.INIT('h01)
	) name6385 (
		_w12190_,
		_w12211_,
		_w12195_,
		_w12212_
	);
	LUT4 #(
		.INIT('h7077)
	) name6386 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12213_
	);
	LUT4 #(
		.INIT('haa02)
	) name6387 (
		_w12192_,
		_w12189_,
		_w12194_,
		_w12190_,
		_w12214_
	);
	LUT3 #(
		.INIT('h01)
	) name6388 (
		_w12189_,
		_w12194_,
		_w12191_,
		_w12215_
	);
	LUT4 #(
		.INIT('h45cf)
	) name6389 (
		_w12200_,
		_w12213_,
		_w12214_,
		_w12215_,
		_w12216_
	);
	LUT2 #(
		.INIT('h4)
	) name6390 (
		_w12212_,
		_w12216_,
		_w12217_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6391 (
		\u2_L3_reg[11]/NET0131 ,
		_w12210_,
		_w12203_,
		_w12217_,
		_w12218_
	);
	LUT4 #(
		.INIT('hc963)
	) name6392 (
		decrypt_pad,
		\u2_R3_reg[12]/NET0131 ,
		\u2_uk_K_r3_reg[53]/NET0131 ,
		\u2_uk_K_r3_reg[5]/NET0131 ,
		_w12219_
	);
	LUT4 #(
		.INIT('hc693)
	) name6393 (
		decrypt_pad,
		\u2_R3_reg[13]/NET0131 ,
		\u2_uk_K_r3_reg[24]/NET0131 ,
		\u2_uk_K_r3_reg[47]/NET0131 ,
		_w12220_
	);
	LUT2 #(
		.INIT('h4)
	) name6394 (
		_w12219_,
		_w12220_,
		_w12221_
	);
	LUT2 #(
		.INIT('h2)
	) name6395 (
		_w12219_,
		_w12220_,
		_w12222_
	);
	LUT2 #(
		.INIT('h9)
	) name6396 (
		_w12219_,
		_w12220_,
		_w12223_
	);
	LUT4 #(
		.INIT('hc963)
	) name6397 (
		decrypt_pad,
		\u2_R3_reg[15]/NET0131 ,
		\u2_uk_K_r3_reg[24]/NET0131 ,
		\u2_uk_K_r3_reg[33]/NET0131 ,
		_w12224_
	);
	LUT4 #(
		.INIT('hc693)
	) name6398 (
		decrypt_pad,
		\u2_R3_reg[14]/NET0131 ,
		\u2_uk_K_r3_reg[25]/NET0131 ,
		\u2_uk_K_r3_reg[48]/NET0131 ,
		_w12225_
	);
	LUT4 #(
		.INIT('h0012)
	) name6399 (
		_w12219_,
		_w12224_,
		_w12220_,
		_w12225_,
		_w12226_
	);
	LUT4 #(
		.INIT('hc963)
	) name6400 (
		decrypt_pad,
		\u2_R3_reg[17]/NET0131 ,
		\u2_uk_K_r3_reg[12]/NET0131 ,
		\u2_uk_K_r3_reg[46]/NET0131 ,
		_w12227_
	);
	LUT2 #(
		.INIT('h4)
	) name6401 (
		_w12219_,
		_w12227_,
		_w12228_
	);
	LUT4 #(
		.INIT('h0040)
	) name6402 (
		_w12219_,
		_w12227_,
		_w12224_,
		_w12220_,
		_w12229_
	);
	LUT4 #(
		.INIT('h2000)
	) name6403 (
		_w12219_,
		_w12227_,
		_w12224_,
		_w12220_,
		_w12230_
	);
	LUT4 #(
		.INIT('hc963)
	) name6404 (
		decrypt_pad,
		\u2_R3_reg[16]/NET0131 ,
		\u2_uk_K_r3_reg[32]/NET0131 ,
		\u2_uk_K_r3_reg[41]/NET0131 ,
		_w12231_
	);
	LUT4 #(
		.INIT('h0010)
	) name6405 (
		_w12229_,
		_w12230_,
		_w12231_,
		_w12226_,
		_w12232_
	);
	LUT4 #(
		.INIT('h0001)
	) name6406 (
		_w12219_,
		_w12227_,
		_w12224_,
		_w12220_,
		_w12233_
	);
	LUT4 #(
		.INIT('h0040)
	) name6407 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12234_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name6408 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12235_
	);
	LUT3 #(
		.INIT('h70)
	) name6409 (
		_w12233_,
		_w12225_,
		_w12235_,
		_w12236_
	);
	LUT2 #(
		.INIT('h8)
	) name6410 (
		_w12232_,
		_w12236_,
		_w12237_
	);
	LUT3 #(
		.INIT('h02)
	) name6411 (
		_w12219_,
		_w12220_,
		_w12225_,
		_w12238_
	);
	LUT4 #(
		.INIT('h0008)
	) name6412 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12239_
	);
	LUT4 #(
		.INIT('h8000)
	) name6413 (
		_w12219_,
		_w12227_,
		_w12224_,
		_w12220_,
		_w12240_
	);
	LUT3 #(
		.INIT('h01)
	) name6414 (
		_w12231_,
		_w12239_,
		_w12240_,
		_w12241_
	);
	LUT4 #(
		.INIT('h0010)
	) name6415 (
		_w12219_,
		_w12227_,
		_w12224_,
		_w12220_,
		_w12242_
	);
	LUT3 #(
		.INIT('h80)
	) name6416 (
		_w12224_,
		_w12220_,
		_w12225_,
		_w12243_
	);
	LUT4 #(
		.INIT('h4000)
	) name6417 (
		_w12219_,
		_w12224_,
		_w12220_,
		_w12225_,
		_w12244_
	);
	LUT2 #(
		.INIT('h1)
	) name6418 (
		_w12242_,
		_w12244_,
		_w12245_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name6419 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12246_
	);
	LUT4 #(
		.INIT('heffe)
	) name6420 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12247_
	);
	LUT3 #(
		.INIT('he0)
	) name6421 (
		_w12224_,
		_w12246_,
		_w12247_,
		_w12248_
	);
	LUT3 #(
		.INIT('h80)
	) name6422 (
		_w12241_,
		_w12245_,
		_w12248_,
		_w12249_
	);
	LUT4 #(
		.INIT('h0200)
	) name6423 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12250_
	);
	LUT4 #(
		.INIT('h0020)
	) name6424 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12251_
	);
	LUT4 #(
		.INIT('hfdde)
	) name6425 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12252_
	);
	LUT3 #(
		.INIT('h02)
	) name6426 (
		_w12227_,
		_w12224_,
		_w12225_,
		_w12253_
	);
	LUT4 #(
		.INIT('h31f5)
	) name6427 (
		_w12224_,
		_w12221_,
		_w12252_,
		_w12253_,
		_w12254_
	);
	LUT4 #(
		.INIT('ha955)
	) name6428 (
		\u2_L3_reg[20]/NET0131 ,
		_w12237_,
		_w12249_,
		_w12254_,
		_w12255_
	);
	LUT4 #(
		.INIT('hc963)
	) name6429 (
		decrypt_pad,
		\u2_R3_reg[32]/NET0131 ,
		\u2_uk_K_r3_reg[1]/NET0131 ,
		\u2_uk_K_r3_reg[37]/NET0131 ,
		_w12256_
	);
	LUT4 #(
		.INIT('hc963)
	) name6430 (
		decrypt_pad,
		\u2_R3_reg[1]/NET0131 ,
		\u2_uk_K_r3_reg[22]/NET0131 ,
		\u2_uk_K_r3_reg[31]/NET0131 ,
		_w12257_
	);
	LUT4 #(
		.INIT('hc693)
	) name6431 (
		decrypt_pad,
		\u2_R3_reg[28]/NET0131 ,
		\u2_uk_K_r3_reg[15]/NET0131 ,
		\u2_uk_K_r3_reg[38]/NET0131 ,
		_w12258_
	);
	LUT4 #(
		.INIT('hc693)
	) name6432 (
		decrypt_pad,
		\u2_R3_reg[30]/NET0131 ,
		\u2_uk_K_r3_reg[43]/NET0131 ,
		\u2_uk_K_r3_reg[7]/NET0131 ,
		_w12259_
	);
	LUT4 #(
		.INIT('hc963)
	) name6433 (
		decrypt_pad,
		\u2_R3_reg[29]/NET0131 ,
		\u2_uk_K_r3_reg[37]/NET0131 ,
		\u2_uk_K_r3_reg[42]/NET0131 ,
		_w12260_
	);
	LUT3 #(
		.INIT('h08)
	) name6434 (
		_w12259_,
		_w12258_,
		_w12260_,
		_w12261_
	);
	LUT4 #(
		.INIT('h0020)
	) name6435 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12262_
	);
	LUT4 #(
		.INIT('hc693)
	) name6436 (
		decrypt_pad,
		\u2_R3_reg[31]/P0001 ,
		\u2_uk_K_r3_reg[0]/NET0131 ,
		\u2_uk_K_r3_reg[50]/NET0131 ,
		_w12263_
	);
	LUT4 #(
		.INIT('hfd00)
	) name6437 (
		_w12257_,
		_w12258_,
		_w12260_,
		_w12263_,
		_w12264_
	);
	LUT3 #(
		.INIT('h02)
	) name6438 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12265_
	);
	LUT3 #(
		.INIT('h07)
	) name6439 (
		_w12257_,
		_w12260_,
		_w12263_,
		_w12266_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6440 (
		_w12262_,
		_w12264_,
		_w12265_,
		_w12266_,
		_w12267_
	);
	LUT2 #(
		.INIT('h4)
	) name6441 (
		_w12257_,
		_w12260_,
		_w12268_
	);
	LUT2 #(
		.INIT('h1)
	) name6442 (
		_w12259_,
		_w12263_,
		_w12269_
	);
	LUT4 #(
		.INIT('h6f2a)
	) name6443 (
		_w12259_,
		_w12257_,
		_w12260_,
		_w12263_,
		_w12270_
	);
	LUT2 #(
		.INIT('h2)
	) name6444 (
		_w12258_,
		_w12270_,
		_w12271_
	);
	LUT3 #(
		.INIT('h54)
	) name6445 (
		_w12256_,
		_w12267_,
		_w12271_,
		_w12272_
	);
	LUT4 #(
		.INIT('h0800)
	) name6446 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12273_
	);
	LUT4 #(
		.INIT('h00fe)
	) name6447 (
		_w12259_,
		_w12258_,
		_w12260_,
		_w12263_,
		_w12274_
	);
	LUT2 #(
		.INIT('h4)
	) name6448 (
		_w12259_,
		_w12258_,
		_w12275_
	);
	LUT4 #(
		.INIT('h1331)
	) name6449 (
		_w12263_,
		_w12274_,
		_w12268_,
		_w12275_,
		_w12276_
	);
	LUT3 #(
		.INIT('he0)
	) name6450 (
		_w12273_,
		_w12276_,
		_w12256_,
		_w12277_
	);
	LUT3 #(
		.INIT('h20)
	) name6451 (
		_w12259_,
		_w12258_,
		_w12260_,
		_w12278_
	);
	LUT2 #(
		.INIT('h8)
	) name6452 (
		_w12257_,
		_w12258_,
		_w12279_
	);
	LUT4 #(
		.INIT('h0008)
	) name6453 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12280_
	);
	LUT4 #(
		.INIT('hfdb6)
	) name6454 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12281_
	);
	LUT2 #(
		.INIT('h2)
	) name6455 (
		_w12263_,
		_w12281_,
		_w12282_
	);
	LUT2 #(
		.INIT('h4)
	) name6456 (
		_w12263_,
		_w12256_,
		_w12283_
	);
	LUT3 #(
		.INIT('h40)
	) name6457 (
		_w12257_,
		_w12258_,
		_w12260_,
		_w12284_
	);
	LUT4 #(
		.INIT('h135f)
	) name6458 (
		_w12261_,
		_w12269_,
		_w12283_,
		_w12284_,
		_w12285_
	);
	LUT2 #(
		.INIT('h4)
	) name6459 (
		_w12282_,
		_w12285_,
		_w12286_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6460 (
		\u2_L3_reg[5]/NET0131 ,
		_w12277_,
		_w12272_,
		_w12286_,
		_w12287_
	);
	LUT3 #(
		.INIT('hc4)
	) name6461 (
		_w12227_,
		_w12224_,
		_w12225_,
		_w12288_
	);
	LUT4 #(
		.INIT('h0040)
	) name6462 (
		_w12219_,
		_w12227_,
		_w12224_,
		_w12225_,
		_w12289_
	);
	LUT4 #(
		.INIT('h0105)
	) name6463 (
		_w12233_,
		_w12222_,
		_w12289_,
		_w12288_,
		_w12290_
	);
	LUT4 #(
		.INIT('hff0d)
	) name6464 (
		_w12227_,
		_w12224_,
		_w12220_,
		_w12225_,
		_w12291_
	);
	LUT3 #(
		.INIT('hc4)
	) name6465 (
		_w12219_,
		_w12247_,
		_w12291_,
		_w12292_
	);
	LUT3 #(
		.INIT('h15)
	) name6466 (
		_w12231_,
		_w12290_,
		_w12292_,
		_w12293_
	);
	LUT4 #(
		.INIT('hefe7)
	) name6467 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12294_
	);
	LUT4 #(
		.INIT('h7bff)
	) name6468 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12295_
	);
	LUT4 #(
		.INIT('hddbd)
	) name6469 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12296_
	);
	LUT4 #(
		.INIT('hc840)
	) name6470 (
		_w12224_,
		_w12295_,
		_w12296_,
		_w12294_,
		_w12297_
	);
	LUT4 #(
		.INIT('h7bfe)
	) name6471 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12298_
	);
	LUT4 #(
		.INIT('h1302)
	) name6472 (
		_w12224_,
		_w12244_,
		_w12251_,
		_w12298_,
		_w12299_
	);
	LUT3 #(
		.INIT('hd0)
	) name6473 (
		_w12231_,
		_w12297_,
		_w12299_,
		_w12300_
	);
	LUT3 #(
		.INIT('h65)
	) name6474 (
		\u2_L3_reg[10]/NET0131 ,
		_w12293_,
		_w12300_,
		_w12301_
	);
	LUT4 #(
		.INIT('h2000)
	) name6475 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12302_
	);
	LUT4 #(
		.INIT('h00bf)
	) name6476 (
		_w12125_,
		_w12127_,
		_w12128_,
		_w12137_,
		_w12303_
	);
	LUT2 #(
		.INIT('h4)
	) name6477 (
		_w12302_,
		_w12303_,
		_w12304_
	);
	LUT3 #(
		.INIT('h35)
	) name6478 (
		_w12125_,
		_w12127_,
		_w12126_,
		_w12305_
	);
	LUT3 #(
		.INIT('h41)
	) name6479 (
		_w12125_,
		_w12126_,
		_w12129_,
		_w12306_
	);
	LUT3 #(
		.INIT('h02)
	) name6480 (
		_w12126_,
		_w12128_,
		_w12129_,
		_w12307_
	);
	LUT4 #(
		.INIT('hffe9)
	) name6481 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12308_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6482 (
		_w12140_,
		_w12305_,
		_w12306_,
		_w12308_,
		_w12309_
	);
	LUT2 #(
		.INIT('h8)
	) name6483 (
		_w12304_,
		_w12309_,
		_w12310_
	);
	LUT4 #(
		.INIT('h0020)
	) name6484 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12311_
	);
	LUT4 #(
		.INIT('h000b)
	) name6485 (
		_w12125_,
		_w12145_,
		_w12148_,
		_w12311_,
		_w12312_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name6486 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12313_
	);
	LUT2 #(
		.INIT('h2)
	) name6487 (
		_w12125_,
		_w12313_,
		_w12314_
	);
	LUT4 #(
		.INIT('h0400)
	) name6488 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12315_
	);
	LUT3 #(
		.INIT('h02)
	) name6489 (
		_w12137_,
		_w12139_,
		_w12315_,
		_w12316_
	);
	LUT3 #(
		.INIT('h40)
	) name6490 (
		_w12314_,
		_w12316_,
		_w12312_,
		_w12317_
	);
	LUT3 #(
		.INIT('ha9)
	) name6491 (
		\u2_L3_reg[12]/NET0131 ,
		_w12310_,
		_w12317_,
		_w12318_
	);
	LUT4 #(
		.INIT('hc963)
	) name6492 (
		decrypt_pad,
		\u2_R3_reg[19]/NET0131 ,
		\u2_uk_K_r3_reg[2]/NET0131 ,
		\u2_uk_K_r3_reg[7]/NET0131 ,
		_w12319_
	);
	LUT4 #(
		.INIT('hc963)
	) name6493 (
		decrypt_pad,
		\u2_R3_reg[18]/NET0131 ,
		\u2_uk_K_r3_reg[15]/NET0131 ,
		\u2_uk_K_r3_reg[51]/NET0131 ,
		_w12320_
	);
	LUT4 #(
		.INIT('hc963)
	) name6494 (
		decrypt_pad,
		\u2_R3_reg[17]/NET0131 ,
		\u2_uk_K_r3_reg[21]/NET0131 ,
		\u2_uk_K_r3_reg[2]/NET0131 ,
		_w12321_
	);
	LUT4 #(
		.INIT('hc963)
	) name6495 (
		decrypt_pad,
		\u2_R3_reg[16]/NET0131 ,
		\u2_uk_K_r3_reg[30]/NET0131 ,
		\u2_uk_K_r3_reg[35]/NET0131 ,
		_w12322_
	);
	LUT4 #(
		.INIT('hc693)
	) name6496 (
		decrypt_pad,
		\u2_R3_reg[21]/NET0131 ,
		\u2_uk_K_r3_reg[23]/NET0131 ,
		\u2_uk_K_r3_reg[42]/NET0131 ,
		_w12323_
	);
	LUT3 #(
		.INIT('h04)
	) name6497 (
		_w12321_,
		_w12322_,
		_w12323_,
		_w12324_
	);
	LUT4 #(
		.INIT('h0010)
	) name6498 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12325_
	);
	LUT4 #(
		.INIT('h4000)
	) name6499 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12326_
	);
	LUT4 #(
		.INIT('hbc67)
	) name6500 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12327_
	);
	LUT4 #(
		.INIT('h5bf8)
	) name6501 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12328_
	);
	LUT4 #(
		.INIT('h2004)
	) name6502 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12329_
	);
	LUT4 #(
		.INIT('h00d8)
	) name6503 (
		_w12319_,
		_w12328_,
		_w12327_,
		_w12329_,
		_w12330_
	);
	LUT4 #(
		.INIT('hc693)
	) name6504 (
		decrypt_pad,
		\u2_R3_reg[20]/NET0131 ,
		\u2_uk_K_r3_reg[22]/NET0131 ,
		\u2_uk_K_r3_reg[45]/P0001 ,
		_w12331_
	);
	LUT2 #(
		.INIT('h1)
	) name6505 (
		_w12330_,
		_w12331_,
		_w12332_
	);
	LUT4 #(
		.INIT('ha43f)
	) name6506 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12333_
	);
	LUT2 #(
		.INIT('h2)
	) name6507 (
		_w12319_,
		_w12333_,
		_w12334_
	);
	LUT3 #(
		.INIT('hde)
	) name6508 (
		_w12321_,
		_w12322_,
		_w12323_,
		_w12335_
	);
	LUT2 #(
		.INIT('h1)
	) name6509 (
		_w12319_,
		_w12320_,
		_w12336_
	);
	LUT2 #(
		.INIT('h4)
	) name6510 (
		_w12335_,
		_w12336_,
		_w12337_
	);
	LUT2 #(
		.INIT('h9)
	) name6511 (
		_w12320_,
		_w12321_,
		_w12338_
	);
	LUT4 #(
		.INIT('h0060)
	) name6512 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12339_
	);
	LUT4 #(
		.INIT('h7000)
	) name6513 (
		_w12319_,
		_w12320_,
		_w12322_,
		_w12323_,
		_w12340_
	);
	LUT3 #(
		.INIT('h13)
	) name6514 (
		_w12338_,
		_w12339_,
		_w12340_,
		_w12341_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6515 (
		_w12331_,
		_w12334_,
		_w12337_,
		_w12341_,
		_w12342_
	);
	LUT4 #(
		.INIT('h0040)
	) name6516 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12343_
	);
	LUT4 #(
		.INIT('hffbd)
	) name6517 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12344_
	);
	LUT4 #(
		.INIT('h0200)
	) name6518 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12345_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name6519 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12346_
	);
	LUT3 #(
		.INIT('hd8)
	) name6520 (
		_w12319_,
		_w12344_,
		_w12346_,
		_w12347_
	);
	LUT4 #(
		.INIT('h5655)
	) name6521 (
		\u2_L3_reg[14]/NET0131 ,
		_w12332_,
		_w12342_,
		_w12347_,
		_w12348_
	);
	LUT4 #(
		.INIT('h1000)
	) name6522 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12349_
	);
	LUT4 #(
		.INIT('hef11)
	) name6523 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12350_
	);
	LUT4 #(
		.INIT('h00a1)
	) name6524 (
		_w12157_,
		_w12159_,
		_w12158_,
		_w12156_,
		_w12351_
	);
	LUT4 #(
		.INIT('h0400)
	) name6525 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12352_
	);
	LUT4 #(
		.INIT('h7b7f)
	) name6526 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12353_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6527 (
		_w12156_,
		_w12350_,
		_w12351_,
		_w12353_,
		_w12354_
	);
	LUT4 #(
		.INIT('h0048)
	) name6528 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12355_
	);
	LUT4 #(
		.INIT('h4100)
	) name6529 (
		_w12155_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12356_
	);
	LUT3 #(
		.INIT('ha8)
	) name6530 (
		_w12156_,
		_w12355_,
		_w12356_,
		_w12357_
	);
	LUT4 #(
		.INIT('hccc8)
	) name6531 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12358_
	);
	LUT3 #(
		.INIT('h09)
	) name6532 (
		_w12160_,
		_w12158_,
		_w12156_,
		_w12359_
	);
	LUT4 #(
		.INIT('hf7df)
	) name6533 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12360_
	);
	LUT3 #(
		.INIT('hb0)
	) name6534 (
		_w12358_,
		_w12359_,
		_w12360_,
		_w12361_
	);
	LUT4 #(
		.INIT('h3210)
	) name6535 (
		_w12155_,
		_w12357_,
		_w12361_,
		_w12354_,
		_w12362_
	);
	LUT2 #(
		.INIT('h9)
	) name6536 (
		\u2_L3_reg[17]/NET0131 ,
		_w12362_,
		_w12363_
	);
	LUT4 #(
		.INIT('h0010)
	) name6537 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12364_
	);
	LUT4 #(
		.INIT('h0ef3)
	) name6538 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12365_
	);
	LUT4 #(
		.INIT('h3032)
	) name6539 (
		_w12263_,
		_w12256_,
		_w12364_,
		_w12365_,
		_w12366_
	);
	LUT4 #(
		.INIT('hf95e)
	) name6540 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12367_
	);
	LUT2 #(
		.INIT('h1)
	) name6541 (
		_w12263_,
		_w12367_,
		_w12368_
	);
	LUT4 #(
		.INIT('hadff)
	) name6542 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12369_
	);
	LUT4 #(
		.INIT('h0100)
	) name6543 (
		_w12257_,
		_w12258_,
		_w12260_,
		_w12263_,
		_w12370_
	);
	LUT3 #(
		.INIT('h08)
	) name6544 (
		_w12259_,
		_w12257_,
		_w12260_,
		_w12371_
	);
	LUT2 #(
		.INIT('h4)
	) name6545 (
		_w12258_,
		_w12263_,
		_w12372_
	);
	LUT4 #(
		.INIT('h5100)
	) name6546 (
		_w12370_,
		_w12371_,
		_w12372_,
		_w12369_,
		_w12373_
	);
	LUT4 #(
		.INIT('hf7fb)
	) name6547 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12374_
	);
	LUT4 #(
		.INIT('h0002)
	) name6548 (
		_w12258_,
		_w12260_,
		_w12263_,
		_w12256_,
		_w12375_
	);
	LUT3 #(
		.INIT('h0d)
	) name6549 (
		_w12263_,
		_w12374_,
		_w12375_,
		_w12376_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6550 (
		_w12256_,
		_w12373_,
		_w12368_,
		_w12376_,
		_w12377_
	);
	LUT3 #(
		.INIT('h65)
	) name6551 (
		\u2_L3_reg[15]/NET0131 ,
		_w12366_,
		_w12377_,
		_w12378_
	);
	LUT4 #(
		.INIT('h082a)
	) name6552 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12379_
	);
	LUT3 #(
		.INIT('h01)
	) name6553 (
		_w12219_,
		_w12227_,
		_w12225_,
		_w12380_
	);
	LUT4 #(
		.INIT('hfad8)
	) name6554 (
		_w12224_,
		_w12250_,
		_w12379_,
		_w12380_,
		_w12381_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name6555 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12382_
	);
	LUT3 #(
		.INIT('h45)
	) name6556 (
		_w12231_,
		_w12381_,
		_w12382_,
		_w12383_
	);
	LUT4 #(
		.INIT('hbf2f)
	) name6557 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12384_
	);
	LUT4 #(
		.INIT('h2000)
	) name6558 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12385_
	);
	LUT4 #(
		.INIT('hdaff)
	) name6559 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12386_
	);
	LUT4 #(
		.INIT('h04cc)
	) name6560 (
		_w12224_,
		_w12231_,
		_w12384_,
		_w12386_,
		_w12387_
	);
	LUT4 #(
		.INIT('h6bff)
	) name6561 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12388_
	);
	LUT2 #(
		.INIT('h2)
	) name6562 (
		_w12224_,
		_w12388_,
		_w12389_
	);
	LUT2 #(
		.INIT('h4)
	) name6563 (
		_w12224_,
		_w12385_,
		_w12390_
	);
	LUT4 #(
		.INIT('hf3f1)
	) name6564 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12391_
	);
	LUT2 #(
		.INIT('h8)
	) name6565 (
		_w12224_,
		_w12231_,
		_w12392_
	);
	LUT4 #(
		.INIT('h7077)
	) name6566 (
		_w12233_,
		_w12225_,
		_w12391_,
		_w12392_,
		_w12393_
	);
	LUT4 #(
		.INIT('h0100)
	) name6567 (
		_w12389_,
		_w12390_,
		_w12387_,
		_w12393_,
		_w12394_
	);
	LUT3 #(
		.INIT('h65)
	) name6568 (
		\u2_L3_reg[1]/NET0131 ,
		_w12383_,
		_w12394_,
		_w12395_
	);
	LUT4 #(
		.INIT('h53bb)
	) name6569 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12396_
	);
	LUT4 #(
		.INIT('hef6f)
	) name6570 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12397_
	);
	LUT4 #(
		.INIT('hdff9)
	) name6571 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12398_
	);
	LUT4 #(
		.INIT('he400)
	) name6572 (
		_w12263_,
		_w12397_,
		_w12396_,
		_w12398_,
		_w12399_
	);
	LUT2 #(
		.INIT('h2)
	) name6573 (
		_w12256_,
		_w12399_,
		_w12400_
	);
	LUT3 #(
		.INIT('hba)
	) name6574 (
		_w12259_,
		_w12260_,
		_w12263_,
		_w12401_
	);
	LUT4 #(
		.INIT('hffde)
	) name6575 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12402_
	);
	LUT3 #(
		.INIT('hd0)
	) name6576 (
		_w12279_,
		_w12401_,
		_w12402_,
		_w12403_
	);
	LUT4 #(
		.INIT('hcf5f)
	) name6577 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12404_
	);
	LUT2 #(
		.INIT('h2)
	) name6578 (
		_w12263_,
		_w12404_,
		_w12405_
	);
	LUT4 #(
		.INIT('h0010)
	) name6579 (
		_w12257_,
		_w12258_,
		_w12260_,
		_w12263_,
		_w12406_
	);
	LUT4 #(
		.INIT('h0008)
	) name6580 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12263_,
		_w12407_
	);
	LUT3 #(
		.INIT('h01)
	) name6581 (
		_w12278_,
		_w12407_,
		_w12406_,
		_w12408_
	);
	LUT4 #(
		.INIT('h4555)
	) name6582 (
		_w12256_,
		_w12405_,
		_w12408_,
		_w12403_,
		_w12409_
	);
	LUT3 #(
		.INIT('h80)
	) name6583 (
		_w12257_,
		_w12258_,
		_w12260_,
		_w12410_
	);
	LUT4 #(
		.INIT('h0100)
	) name6584 (
		_w12259_,
		_w12258_,
		_w12260_,
		_w12263_,
		_w12411_
	);
	LUT3 #(
		.INIT('h07)
	) name6585 (
		_w12269_,
		_w12410_,
		_w12411_,
		_w12412_
	);
	LUT4 #(
		.INIT('h5655)
	) name6586 (
		\u2_L3_reg[21]/NET0131 ,
		_w12409_,
		_w12400_,
		_w12412_,
		_w12413_
	);
	LUT4 #(
		.INIT('hf8fc)
	) name6587 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12414_
	);
	LUT4 #(
		.INIT('h0092)
	) name6588 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12415_
	);
	LUT4 #(
		.INIT('h5501)
	) name6589 (
		_w12224_,
		_w12231_,
		_w12414_,
		_w12415_,
		_w12416_
	);
	LUT4 #(
		.INIT('h0010)
	) name6590 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12417_
	);
	LUT4 #(
		.INIT('h0002)
	) name6591 (
		_w12231_,
		_w12242_,
		_w12385_,
		_w12417_,
		_w12418_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name6592 (
		_w12219_,
		_w12227_,
		_w12224_,
		_w12220_,
		_w12419_
	);
	LUT4 #(
		.INIT('h77fb)
	) name6593 (
		_w12219_,
		_w12227_,
		_w12220_,
		_w12225_,
		_w12420_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name6594 (
		_w12224_,
		_w12225_,
		_w12419_,
		_w12420_,
		_w12421_
	);
	LUT2 #(
		.INIT('h4)
	) name6595 (
		_w12228_,
		_w12243_,
		_w12422_
	);
	LUT4 #(
		.INIT('h0001)
	) name6596 (
		_w12234_,
		_w12230_,
		_w12231_,
		_w12238_,
		_w12423_
	);
	LUT4 #(
		.INIT('h7077)
	) name6597 (
		_w12418_,
		_w12421_,
		_w12422_,
		_w12423_,
		_w12424_
	);
	LUT3 #(
		.INIT('h08)
	) name6598 (
		_w12227_,
		_w12224_,
		_w12225_,
		_w12425_
	);
	LUT2 #(
		.INIT('h4)
	) name6599 (
		_w12223_,
		_w12425_,
		_w12426_
	);
	LUT4 #(
		.INIT('h5556)
	) name6600 (
		\u2_L3_reg[26]/NET0131 ,
		_w12424_,
		_w12416_,
		_w12426_,
		_w12427_
	);
	LUT4 #(
		.INIT('h67dc)
	) name6601 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12428_
	);
	LUT4 #(
		.INIT('hd2f7)
	) name6602 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12429_
	);
	LUT4 #(
		.INIT('h0040)
	) name6603 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12430_
	);
	LUT4 #(
		.INIT('h00d8)
	) name6604 (
		_w12192_,
		_w12428_,
		_w12429_,
		_w12430_,
		_w12431_
	);
	LUT4 #(
		.INIT('h9aff)
	) name6605 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12432_
	);
	LUT4 #(
		.INIT('haa02)
	) name6606 (
		_w12192_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12433_
	);
	LUT4 #(
		.INIT('h9297)
	) name6607 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12434_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name6608 (
		_w12192_,
		_w12432_,
		_w12433_,
		_w12434_,
		_w12435_
	);
	LUT4 #(
		.INIT('h0800)
	) name6609 (
		_w12192_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12436_
	);
	LUT2 #(
		.INIT('h1)
	) name6610 (
		_w12204_,
		_w12436_,
		_w12437_
	);
	LUT4 #(
		.INIT('hd800)
	) name6611 (
		_w12188_,
		_w12435_,
		_w12431_,
		_w12437_,
		_w12438_
	);
	LUT2 #(
		.INIT('h6)
	) name6612 (
		\u2_L3_reg[29]/NET0131 ,
		_w12438_,
		_w12439_
	);
	LUT4 #(
		.INIT('h3ce4)
	) name6613 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12440_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name6614 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12441_
	);
	LUT4 #(
		.INIT('hbb7f)
	) name6615 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12442_
	);
	LUT4 #(
		.INIT('hd800)
	) name6616 (
		_w12319_,
		_w12440_,
		_w12441_,
		_w12442_,
		_w12443_
	);
	LUT2 #(
		.INIT('h2)
	) name6617 (
		_w12331_,
		_w12443_,
		_w12444_
	);
	LUT4 #(
		.INIT('hfe7d)
	) name6618 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12445_
	);
	LUT2 #(
		.INIT('h2)
	) name6619 (
		_w12319_,
		_w12445_,
		_w12446_
	);
	LUT3 #(
		.INIT('ha2)
	) name6620 (
		_w12319_,
		_w12321_,
		_w12323_,
		_w12447_
	);
	LUT4 #(
		.INIT('h2223)
	) name6621 (
		_w12319_,
		_w12320_,
		_w12321_,
		_w12322_,
		_w12448_
	);
	LUT2 #(
		.INIT('h4)
	) name6622 (
		_w12447_,
		_w12448_,
		_w12449_
	);
	LUT4 #(
		.INIT('h0010)
	) name6623 (
		_w12319_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12450_
	);
	LUT2 #(
		.INIT('h2)
	) name6624 (
		_w12319_,
		_w12323_,
		_w12451_
	);
	LUT3 #(
		.INIT('h08)
	) name6625 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12452_
	);
	LUT3 #(
		.INIT('h45)
	) name6626 (
		_w12450_,
		_w12451_,
		_w12452_,
		_w12453_
	);
	LUT4 #(
		.INIT('h0400)
	) name6627 (
		_w12319_,
		_w12320_,
		_w12321_,
		_w12322_,
		_w12454_
	);
	LUT2 #(
		.INIT('h1)
	) name6628 (
		_w12326_,
		_w12454_,
		_w12455_
	);
	LUT4 #(
		.INIT('hba00)
	) name6629 (
		_w12331_,
		_w12449_,
		_w12453_,
		_w12455_,
		_w12456_
	);
	LUT4 #(
		.INIT('h5655)
	) name6630 (
		\u2_L3_reg[25]/NET0131 ,
		_w12444_,
		_w12446_,
		_w12456_,
		_w12457_
	);
	LUT4 #(
		.INIT('hc693)
	) name6631 (
		decrypt_pad,
		\u2_R3_reg[8]/NET0131 ,
		\u2_uk_K_r3_reg[40]/NET0131 ,
		\u2_uk_K_r3_reg[6]/NET0131 ,
		_w12458_
	);
	LUT4 #(
		.INIT('hc693)
	) name6632 (
		decrypt_pad,
		\u2_R3_reg[5]/NET0131 ,
		\u2_uk_K_r3_reg[32]/NET0131 ,
		\u2_uk_K_r3_reg[55]/NET0131 ,
		_w12459_
	);
	LUT4 #(
		.INIT('hc963)
	) name6633 (
		decrypt_pad,
		\u2_R3_reg[9]/NET0131 ,
		\u2_uk_K_r3_reg[11]/NET0131 ,
		\u2_uk_K_r3_reg[20]/NET0131 ,
		_w12460_
	);
	LUT4 #(
		.INIT('hc963)
	) name6634 (
		decrypt_pad,
		\u2_R3_reg[4]/NET0131 ,
		\u2_uk_K_r3_reg[19]/NET0131 ,
		\u2_uk_K_r3_reg[53]/NET0131 ,
		_w12461_
	);
	LUT3 #(
		.INIT('h04)
	) name6635 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12462_
	);
	LUT3 #(
		.INIT('hd9)
	) name6636 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12463_
	);
	LUT4 #(
		.INIT('hc963)
	) name6637 (
		decrypt_pad,
		\u2_R3_reg[6]/NET0131 ,
		\u2_uk_K_r3_reg[46]/NET0131 ,
		\u2_uk_K_r3_reg[55]/NET0131 ,
		_w12464_
	);
	LUT4 #(
		.INIT('h0026)
	) name6638 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12465_
	);
	LUT4 #(
		.INIT('hc693)
	) name6639 (
		decrypt_pad,
		\u2_R3_reg[7]/NET0131 ,
		\u2_uk_K_r3_reg[17]/NET0131 ,
		\u2_uk_K_r3_reg[40]/NET0131 ,
		_w12466_
	);
	LUT4 #(
		.INIT('h4000)
	) name6640 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12467_
	);
	LUT3 #(
		.INIT('h15)
	) name6641 (
		_w12465_,
		_w12466_,
		_w12467_,
		_w12468_
	);
	LUT2 #(
		.INIT('h8)
	) name6642 (
		_w12461_,
		_w12464_,
		_w12469_
	);
	LUT4 #(
		.INIT('h4bfb)
	) name6643 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12470_
	);
	LUT3 #(
		.INIT('hcd)
	) name6644 (
		_w12459_,
		_w12464_,
		_w12466_,
		_w12471_
	);
	LUT2 #(
		.INIT('h2)
	) name6645 (
		_w12460_,
		_w12461_,
		_w12472_
	);
	LUT4 #(
		.INIT('h084c)
	) name6646 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12473_
	);
	LUT4 #(
		.INIT('h0eee)
	) name6647 (
		_w12466_,
		_w12470_,
		_w12471_,
		_w12473_,
		_w12474_
	);
	LUT3 #(
		.INIT('h15)
	) name6648 (
		_w12458_,
		_w12468_,
		_w12474_,
		_w12475_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name6649 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12476_
	);
	LUT4 #(
		.INIT('h080c)
	) name6650 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12477_
	);
	LUT3 #(
		.INIT('h0d)
	) name6651 (
		_w12459_,
		_w12464_,
		_w12466_,
		_w12478_
	);
	LUT4 #(
		.INIT('hf200)
	) name6652 (
		_w12458_,
		_w12476_,
		_w12477_,
		_w12478_,
		_w12479_
	);
	LUT4 #(
		.INIT('h0080)
	) name6653 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12480_
	);
	LUT4 #(
		.INIT('h0010)
	) name6654 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12481_
	);
	LUT4 #(
		.INIT('h8a00)
	) name6655 (
		_w12459_,
		_w12461_,
		_w12464_,
		_w12466_,
		_w12482_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6656 (
		_w12458_,
		_w12481_,
		_w12482_,
		_w12480_,
		_w12483_
	);
	LUT4 #(
		.INIT('hfc54)
	) name6657 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12484_
	);
	LUT4 #(
		.INIT('hdc00)
	) name6658 (
		_w12459_,
		_w12461_,
		_w12464_,
		_w12466_,
		_w12485_
	);
	LUT2 #(
		.INIT('h4)
	) name6659 (
		_w12484_,
		_w12485_,
		_w12486_
	);
	LUT3 #(
		.INIT('h01)
	) name6660 (
		_w12483_,
		_w12486_,
		_w12479_,
		_w12487_
	);
	LUT3 #(
		.INIT('h65)
	) name6661 (
		\u2_L3_reg[2]/NET0131 ,
		_w12475_,
		_w12487_,
		_w12488_
	);
	LUT4 #(
		.INIT('hd97b)
	) name6662 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12489_
	);
	LUT2 #(
		.INIT('h2)
	) name6663 (
		_w12192_,
		_w12489_,
		_w12490_
	);
	LUT4 #(
		.INIT('heebf)
	) name6664 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12491_
	);
	LUT4 #(
		.INIT('h0040)
	) name6665 (
		_w12192_,
		_w12189_,
		_w12194_,
		_w12190_,
		_w12492_
	);
	LUT4 #(
		.INIT('h0032)
	) name6666 (
		_w12192_,
		_w12204_,
		_w12491_,
		_w12492_,
		_w12493_
	);
	LUT3 #(
		.INIT('h45)
	) name6667 (
		_w12188_,
		_w12490_,
		_w12493_,
		_w12494_
	);
	LUT4 #(
		.INIT('h7c7f)
	) name6668 (
		_w12192_,
		_w12189_,
		_w12194_,
		_w12191_,
		_w12495_
	);
	LUT2 #(
		.INIT('h1)
	) name6669 (
		_w12190_,
		_w12495_,
		_w12496_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name6670 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12497_
	);
	LUT3 #(
		.INIT('h80)
	) name6671 (
		_w12194_,
		_w12190_,
		_w12191_,
		_w12498_
	);
	LUT3 #(
		.INIT('h0e)
	) name6672 (
		_w12192_,
		_w12497_,
		_w12498_,
		_w12499_
	);
	LUT4 #(
		.INIT('h70d0)
	) name6673 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12500_
	);
	LUT4 #(
		.INIT('h5501)
	) name6674 (
		_w12192_,
		_w12189_,
		_w12194_,
		_w12190_,
		_w12501_
	);
	LUT3 #(
		.INIT('h9e)
	) name6675 (
		_w12189_,
		_w12194_,
		_w12191_,
		_w12502_
	);
	LUT2 #(
		.INIT('h8)
	) name6676 (
		_w12192_,
		_w12190_,
		_w12503_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6677 (
		_w12500_,
		_w12501_,
		_w12502_,
		_w12503_,
		_w12504_
	);
	LUT4 #(
		.INIT('h7500)
	) name6678 (
		_w12188_,
		_w12496_,
		_w12499_,
		_w12504_,
		_w12505_
	);
	LUT3 #(
		.INIT('h65)
	) name6679 (
		\u2_L3_reg[4]/NET0131 ,
		_w12494_,
		_w12505_,
		_w12506_
	);
	LUT4 #(
		.INIT('h2000)
	) name6680 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12507_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name6681 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12508_
	);
	LUT4 #(
		.INIT('h0400)
	) name6682 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12509_
	);
	LUT4 #(
		.INIT('hf9ed)
	) name6683 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12510_
	);
	LUT4 #(
		.INIT('h0313)
	) name6684 (
		_w12458_,
		_w12466_,
		_w12508_,
		_w12510_,
		_w12511_
	);
	LUT3 #(
		.INIT('h8e)
	) name6685 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12512_
	);
	LUT4 #(
		.INIT('h3010)
	) name6686 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12513_
	);
	LUT3 #(
		.INIT('h02)
	) name6687 (
		_w12466_,
		_w12512_,
		_w12513_,
		_w12514_
	);
	LUT3 #(
		.INIT('hd0)
	) name6688 (
		_w12459_,
		_w12460_,
		_w12466_,
		_w12515_
	);
	LUT2 #(
		.INIT('h8)
	) name6689 (
		_w12469_,
		_w12515_,
		_w12516_
	);
	LUT3 #(
		.INIT('h51)
	) name6690 (
		_w12458_,
		_w12472_,
		_w12471_,
		_w12517_
	);
	LUT3 #(
		.INIT('h10)
	) name6691 (
		_w12516_,
		_w12514_,
		_w12517_,
		_w12518_
	);
	LUT4 #(
		.INIT('h0002)
	) name6692 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12519_
	);
	LUT4 #(
		.INIT('h002a)
	) name6693 (
		_w12458_,
		_w12471_,
		_w12473_,
		_w12519_,
		_w12520_
	);
	LUT4 #(
		.INIT('h5140)
	) name6694 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12521_
	);
	LUT3 #(
		.INIT('h01)
	) name6695 (
		_w12459_,
		_w12460_,
		_w12464_,
		_w12522_
	);
	LUT4 #(
		.INIT('hf3ee)
	) name6696 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12523_
	);
	LUT4 #(
		.INIT('h80c4)
	) name6697 (
		_w12466_,
		_w12508_,
		_w12523_,
		_w12521_,
		_w12524_
	);
	LUT2 #(
		.INIT('h8)
	) name6698 (
		_w12520_,
		_w12524_,
		_w12525_
	);
	LUT4 #(
		.INIT('h999a)
	) name6699 (
		\u2_L3_reg[13]/NET0131 ,
		_w12511_,
		_w12518_,
		_w12525_,
		_w12526_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name6700 (
		_w12192_,
		_w12189_,
		_w12194_,
		_w12190_,
		_w12527_
	);
	LUT4 #(
		.INIT('hef00)
	) name6701 (
		_w12194_,
		_w12190_,
		_w12191_,
		_w12188_,
		_w12528_
	);
	LUT3 #(
		.INIT('he0)
	) name6702 (
		_w12191_,
		_w12527_,
		_w12528_,
		_w12529_
	);
	LUT4 #(
		.INIT('h4010)
	) name6703 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12530_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name6704 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12531_
	);
	LUT3 #(
		.INIT('h31)
	) name6705 (
		_w12192_,
		_w12530_,
		_w12531_,
		_w12532_
	);
	LUT4 #(
		.INIT('h4e55)
	) name6706 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12533_
	);
	LUT2 #(
		.INIT('h2)
	) name6707 (
		_w12192_,
		_w12533_,
		_w12534_
	);
	LUT4 #(
		.INIT('h1001)
	) name6708 (
		_w12192_,
		_w12189_,
		_w12194_,
		_w12191_,
		_w12535_
	);
	LUT4 #(
		.INIT('h8000)
	) name6709 (
		_w12189_,
		_w12194_,
		_w12190_,
		_w12191_,
		_w12536_
	);
	LUT3 #(
		.INIT('h01)
	) name6710 (
		_w12188_,
		_w12536_,
		_w12535_,
		_w12537_
	);
	LUT4 #(
		.INIT('h7077)
	) name6711 (
		_w12529_,
		_w12532_,
		_w12534_,
		_w12537_,
		_w12538_
	);
	LUT2 #(
		.INIT('h4)
	) name6712 (
		_w12191_,
		_w12492_,
		_w12539_
	);
	LUT2 #(
		.INIT('h1)
	) name6713 (
		_w12212_,
		_w12539_,
		_w12540_
	);
	LUT3 #(
		.INIT('h65)
	) name6714 (
		\u2_L3_reg[19]/NET0131 ,
		_w12538_,
		_w12540_,
		_w12541_
	);
	LUT4 #(
		.INIT('hf73f)
	) name6715 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12542_
	);
	LUT2 #(
		.INIT('h2)
	) name6716 (
		_w12156_,
		_w12542_,
		_w12543_
	);
	LUT3 #(
		.INIT('h07)
	) name6717 (
		_w12173_,
		_w12181_,
		_w12349_,
		_w12544_
	);
	LUT3 #(
		.INIT('h8a)
	) name6718 (
		_w12155_,
		_w12543_,
		_w12544_,
		_w12545_
	);
	LUT4 #(
		.INIT('h7bef)
	) name6719 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12546_
	);
	LUT2 #(
		.INIT('h1)
	) name6720 (
		_w12156_,
		_w12546_,
		_w12547_
	);
	LUT3 #(
		.INIT('h01)
	) name6721 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12548_
	);
	LUT3 #(
		.INIT('h01)
	) name6722 (
		_w12164_,
		_w12183_,
		_w12548_,
		_w12549_
	);
	LUT3 #(
		.INIT('h02)
	) name6723 (
		_w12159_,
		_w12160_,
		_w12158_,
		_w12550_
	);
	LUT4 #(
		.INIT('h0200)
	) name6724 (
		_w12159_,
		_w12160_,
		_w12158_,
		_w12156_,
		_w12551_
	);
	LUT3 #(
		.INIT('hec)
	) name6725 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12552_
	);
	LUT3 #(
		.INIT('h13)
	) name6726 (
		_w12178_,
		_w12551_,
		_w12552_,
		_w12553_
	);
	LUT3 #(
		.INIT('had)
	) name6727 (
		_w12159_,
		_w12160_,
		_w12158_,
		_w12554_
	);
	LUT4 #(
		.INIT('hfdc3)
	) name6728 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12555_
	);
	LUT2 #(
		.INIT('h2)
	) name6729 (
		_w12155_,
		_w12156_,
		_w12556_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name6730 (
		_w12169_,
		_w12554_,
		_w12555_,
		_w12556_,
		_w12557_
	);
	LUT4 #(
		.INIT('hea00)
	) name6731 (
		_w12155_,
		_w12549_,
		_w12553_,
		_w12557_,
		_w12558_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6732 (
		\u2_L3_reg[23]/NET0131 ,
		_w12547_,
		_w12545_,
		_w12558_,
		_w12559_
	);
	LUT3 #(
		.INIT('h9f)
	) name6733 (
		_w12257_,
		_w12258_,
		_w12260_,
		_w12560_
	);
	LUT4 #(
		.INIT('h0100)
	) name6734 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12561_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6735 (
		_w12257_,
		_w12258_,
		_w12260_,
		_w12263_,
		_w12562_
	);
	LUT4 #(
		.INIT('h7077)
	) name6736 (
		_w12274_,
		_w12560_,
		_w12561_,
		_w12562_,
		_w12563_
	);
	LUT4 #(
		.INIT('hf79b)
	) name6737 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12564_
	);
	LUT3 #(
		.INIT('h8a)
	) name6738 (
		_w12256_,
		_w12563_,
		_w12564_,
		_w12565_
	);
	LUT4 #(
		.INIT('hef00)
	) name6739 (
		_w12259_,
		_w12257_,
		_w12260_,
		_w12263_,
		_w12566_
	);
	LUT4 #(
		.INIT('h7533)
	) name6740 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12567_
	);
	LUT2 #(
		.INIT('h8)
	) name6741 (
		_w12566_,
		_w12567_,
		_w12568_
	);
	LUT4 #(
		.INIT('h0080)
	) name6742 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12263_,
		_w12569_
	);
	LUT3 #(
		.INIT('h01)
	) name6743 (
		_w12280_,
		_w12406_,
		_w12569_,
		_w12570_
	);
	LUT3 #(
		.INIT('h45)
	) name6744 (
		_w12256_,
		_w12568_,
		_w12570_,
		_w12571_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name6745 (
		_w12259_,
		_w12257_,
		_w12258_,
		_w12260_,
		_w12572_
	);
	LUT2 #(
		.INIT('h1)
	) name6746 (
		_w12263_,
		_w12572_,
		_w12573_
	);
	LUT4 #(
		.INIT('h0200)
	) name6747 (
		_w12259_,
		_w12257_,
		_w12260_,
		_w12263_,
		_w12574_
	);
	LUT3 #(
		.INIT('h07)
	) name6748 (
		_w12269_,
		_w12284_,
		_w12574_,
		_w12575_
	);
	LUT2 #(
		.INIT('h4)
	) name6749 (
		_w12573_,
		_w12575_,
		_w12576_
	);
	LUT4 #(
		.INIT('h5655)
	) name6750 (
		\u2_L3_reg[27]/NET0131 ,
		_w12571_,
		_w12565_,
		_w12576_,
		_w12577_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name6751 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12578_
	);
	LUT2 #(
		.INIT('h8)
	) name6752 (
		_w12466_,
		_w12578_,
		_w12579_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name6753 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12580_
	);
	LUT3 #(
		.INIT('h10)
	) name6754 (
		_w12459_,
		_w12461_,
		_w12464_,
		_w12581_
	);
	LUT4 #(
		.INIT('h0001)
	) name6755 (
		_w12462_,
		_w12466_,
		_w12507_,
		_w12581_,
		_w12582_
	);
	LUT4 #(
		.INIT('h6100)
	) name6756 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12583_
	);
	LUT2 #(
		.INIT('h1)
	) name6757 (
		_w12458_,
		_w12583_,
		_w12584_
	);
	LUT4 #(
		.INIT('hba00)
	) name6758 (
		_w12579_,
		_w12580_,
		_w12582_,
		_w12584_,
		_w12585_
	);
	LUT4 #(
		.INIT('h0010)
	) name6759 (
		_w12466_,
		_w12507_,
		_w12578_,
		_w12581_,
		_w12586_
	);
	LUT4 #(
		.INIT('h8280)
	) name6760 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12587_
	);
	LUT4 #(
		.INIT('hef00)
	) name6761 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12466_,
		_w12588_
	);
	LUT2 #(
		.INIT('h4)
	) name6762 (
		_w12587_,
		_w12588_,
		_w12589_
	);
	LUT3 #(
		.INIT('h0b)
	) name6763 (
		_w12459_,
		_w12460_,
		_w12466_,
		_w12590_
	);
	LUT2 #(
		.INIT('h2)
	) name6764 (
		_w12461_,
		_w12464_,
		_w12591_
	);
	LUT4 #(
		.INIT('h2022)
	) name6765 (
		_w12458_,
		_w12509_,
		_w12590_,
		_w12591_,
		_w12592_
	);
	LUT3 #(
		.INIT('he0)
	) name6766 (
		_w12586_,
		_w12589_,
		_w12592_,
		_w12593_
	);
	LUT3 #(
		.INIT('ha9)
	) name6767 (
		\u2_L3_reg[28]/NET0131 ,
		_w12585_,
		_w12593_,
		_w12594_
	);
	LUT4 #(
		.INIT('h0080)
	) name6768 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12595_
	);
	LUT4 #(
		.INIT('h00a3)
	) name6769 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12596_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name6770 (
		_w12125_,
		_w12127_,
		_w12126_,
		_w12129_,
		_w12597_
	);
	LUT2 #(
		.INIT('h4)
	) name6771 (
		_w12596_,
		_w12597_,
		_w12598_
	);
	LUT4 #(
		.INIT('h0110)
	) name6772 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12599_
	);
	LUT4 #(
		.INIT('h0001)
	) name6773 (
		_w12125_,
		_w12302_,
		_w12307_,
		_w12599_,
		_w12600_
	);
	LUT4 #(
		.INIT('h888a)
	) name6774 (
		_w12137_,
		_w12595_,
		_w12598_,
		_w12600_,
		_w12601_
	);
	LUT4 #(
		.INIT('h8000)
	) name6775 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12602_
	);
	LUT4 #(
		.INIT('h7db7)
	) name6776 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12603_
	);
	LUT3 #(
		.INIT('h40)
	) name6777 (
		_w12126_,
		_w12128_,
		_w12129_,
		_w12604_
	);
	LUT3 #(
		.INIT('h04)
	) name6778 (
		_w12127_,
		_w12128_,
		_w12129_,
		_w12605_
	);
	LUT4 #(
		.INIT('h5513)
	) name6779 (
		_w12125_,
		_w12306_,
		_w12604_,
		_w12605_,
		_w12606_
	);
	LUT4 #(
		.INIT('h4404)
	) name6780 (
		_w12125_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12607_
	);
	LUT4 #(
		.INIT('h135f)
	) name6781 (
		_w12125_,
		_w12132_,
		_w12145_,
		_w12607_,
		_w12608_
	);
	LUT4 #(
		.INIT('hea00)
	) name6782 (
		_w12137_,
		_w12603_,
		_w12606_,
		_w12608_,
		_w12609_
	);
	LUT3 #(
		.INIT('h65)
	) name6783 (
		\u2_L3_reg[32]/NET0131 ,
		_w12601_,
		_w12609_,
		_w12610_
	);
	LUT4 #(
		.INIT('hc693)
	) name6784 (
		decrypt_pad,
		\u2_R3_reg[12]/NET0131 ,
		\u2_uk_K_r3_reg[18]/NET0131 ,
		\u2_uk_K_r3_reg[41]/NET0131 ,
		_w12611_
	);
	LUT4 #(
		.INIT('hc963)
	) name6785 (
		decrypt_pad,
		\u2_R3_reg[13]/NET0131 ,
		\u2_uk_K_r3_reg[54]/NET0131 ,
		\u2_uk_K_r3_reg[6]/NET0131 ,
		_w12612_
	);
	LUT4 #(
		.INIT('hc963)
	) name6786 (
		decrypt_pad,
		\u2_R3_reg[8]/NET0131 ,
		\u2_uk_K_r3_reg[20]/NET0131 ,
		\u2_uk_K_r3_reg[54]/NET0131 ,
		_w12613_
	);
	LUT2 #(
		.INIT('h6)
	) name6787 (
		_w12612_,
		_w12613_,
		_w12614_
	);
	LUT4 #(
		.INIT('hc963)
	) name6788 (
		decrypt_pad,
		\u2_R3_reg[9]/NET0131 ,
		\u2_uk_K_r3_reg[17]/NET0131 ,
		\u2_uk_K_r3_reg[26]/NET0131 ,
		_w12615_
	);
	LUT4 #(
		.INIT('hc963)
	) name6789 (
		decrypt_pad,
		\u2_R3_reg[10]/NET0131 ,
		\u2_uk_K_r3_reg[25]/NET0131 ,
		\u2_uk_K_r3_reg[34]/NET0131 ,
		_w12616_
	);
	LUT4 #(
		.INIT('h2100)
	) name6790 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12617_
	);
	LUT3 #(
		.INIT('h08)
	) name6791 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12618_
	);
	LUT4 #(
		.INIT('hc963)
	) name6792 (
		decrypt_pad,
		\u2_R3_reg[11]/P0001 ,
		\u2_uk_K_r3_reg[26]/NET0131 ,
		\u2_uk_K_r3_reg[3]/NET0131 ,
		_w12619_
	);
	LUT2 #(
		.INIT('h2)
	) name6793 (
		_w12616_,
		_w12619_,
		_w12620_
	);
	LUT3 #(
		.INIT('h40)
	) name6794 (
		_w12612_,
		_w12615_,
		_w12616_,
		_w12621_
	);
	LUT4 #(
		.INIT('h4000)
	) name6795 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12622_
	);
	LUT4 #(
		.INIT('h0007)
	) name6796 (
		_w12618_,
		_w12620_,
		_w12622_,
		_w12617_,
		_w12623_
	);
	LUT2 #(
		.INIT('h8)
	) name6797 (
		_w12612_,
		_w12619_,
		_w12624_
	);
	LUT3 #(
		.INIT('h46)
	) name6798 (
		_w12612_,
		_w12613_,
		_w12619_,
		_w12625_
	);
	LUT2 #(
		.INIT('h1)
	) name6799 (
		_w12615_,
		_w12616_,
		_w12626_
	);
	LUT2 #(
		.INIT('h8)
	) name6800 (
		_w12626_,
		_w12625_,
		_w12627_
	);
	LUT3 #(
		.INIT('hed)
	) name6801 (
		_w12615_,
		_w12616_,
		_w12625_,
		_w12628_
	);
	LUT3 #(
		.INIT('h15)
	) name6802 (
		_w12611_,
		_w12623_,
		_w12628_,
		_w12629_
	);
	LUT4 #(
		.INIT('h959d)
	) name6803 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12630_
	);
	LUT4 #(
		.INIT('h0001)
	) name6804 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12631_
	);
	LUT4 #(
		.INIT('hddfe)
	) name6805 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12632_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6806 (
		_w12630_,
		_w12611_,
		_w12632_,
		_w12619_,
		_w12633_
	);
	LUT2 #(
		.INIT('h8)
	) name6807 (
		_w12616_,
		_w12611_,
		_w12634_
	);
	LUT3 #(
		.INIT('h04)
	) name6808 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12635_
	);
	LUT2 #(
		.INIT('h2)
	) name6809 (
		_w12611_,
		_w12619_,
		_w12636_
	);
	LUT3 #(
		.INIT('h80)
	) name6810 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12637_
	);
	LUT4 #(
		.INIT('h6f67)
	) name6811 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12638_
	);
	LUT4 #(
		.INIT('h7707)
	) name6812 (
		_w12634_,
		_w12635_,
		_w12636_,
		_w12638_,
		_w12639_
	);
	LUT2 #(
		.INIT('h4)
	) name6813 (
		_w12633_,
		_w12639_,
		_w12640_
	);
	LUT3 #(
		.INIT('h65)
	) name6814 (
		\u2_L3_reg[6]/NET0131 ,
		_w12629_,
		_w12640_,
		_w12641_
	);
	LUT4 #(
		.INIT('h0770)
	) name6815 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12642_
	);
	LUT2 #(
		.INIT('h2)
	) name6816 (
		_w12125_,
		_w12137_,
		_w12643_
	);
	LUT4 #(
		.INIT('h0010)
	) name6817 (
		_w12130_,
		_w12602_,
		_w12643_,
		_w12642_,
		_w12644_
	);
	LUT4 #(
		.INIT('h5884)
	) name6818 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12645_
	);
	LUT2 #(
		.INIT('h4)
	) name6819 (
		_w12125_,
		_w12137_,
		_w12646_
	);
	LUT2 #(
		.INIT('h9)
	) name6820 (
		_w12125_,
		_w12137_,
		_w12647_
	);
	LUT3 #(
		.INIT('h10)
	) name6821 (
		_w12302_,
		_w12645_,
		_w12647_,
		_w12648_
	);
	LUT3 #(
		.INIT('h28)
	) name6822 (
		_w12126_,
		_w12128_,
		_w12129_,
		_w12649_
	);
	LUT3 #(
		.INIT('h09)
	) name6823 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12650_
	);
	LUT4 #(
		.INIT('h20a0)
	) name6824 (
		_w12127_,
		_w12126_,
		_w12128_,
		_w12129_,
		_w12651_
	);
	LUT4 #(
		.INIT('h0002)
	) name6825 (
		_w12646_,
		_w12651_,
		_w12650_,
		_w12649_,
		_w12652_
	);
	LUT4 #(
		.INIT('h00ab)
	) name6826 (
		_w12131_,
		_w12644_,
		_w12648_,
		_w12652_,
		_w12653_
	);
	LUT2 #(
		.INIT('h6)
	) name6827 (
		\u2_L3_reg[7]/NET0131 ,
		_w12653_,
		_w12654_
	);
	LUT4 #(
		.INIT('h3fef)
	) name6828 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12655_
	);
	LUT4 #(
		.INIT('hc2ff)
	) name6829 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12656_
	);
	LUT4 #(
		.INIT('hfb79)
	) name6830 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12657_
	);
	LUT4 #(
		.INIT('hd800)
	) name6831 (
		_w12319_,
		_w12655_,
		_w12656_,
		_w12657_,
		_w12658_
	);
	LUT4 #(
		.INIT('h0001)
	) name6832 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12659_
	);
	LUT4 #(
		.INIT('hcffe)
	) name6833 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12660_
	);
	LUT3 #(
		.INIT('h10)
	) name6834 (
		_w12319_,
		_w12320_,
		_w12322_,
		_w12661_
	);
	LUT4 #(
		.INIT('h00c4)
	) name6835 (
		_w12319_,
		_w12346_,
		_w12660_,
		_w12661_,
		_w12662_
	);
	LUT4 #(
		.INIT('hf977)
	) name6836 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12663_
	);
	LUT4 #(
		.INIT('hbf15)
	) name6837 (
		_w12319_,
		_w12320_,
		_w12324_,
		_w12663_,
		_w12664_
	);
	LUT4 #(
		.INIT('hd800)
	) name6838 (
		_w12331_,
		_w12662_,
		_w12658_,
		_w12664_,
		_w12665_
	);
	LUT2 #(
		.INIT('h9)
	) name6839 (
		\u2_L3_reg[8]/NET0131 ,
		_w12665_,
		_w12666_
	);
	LUT4 #(
		.INIT('hf700)
	) name6840 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12667_
	);
	LUT4 #(
		.INIT('h0400)
	) name6841 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12619_,
		_w12668_
	);
	LUT4 #(
		.INIT('h006d)
	) name6842 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12669_
	);
	LUT3 #(
		.INIT('h45)
	) name6843 (
		_w12667_,
		_w12668_,
		_w12669_,
		_w12670_
	);
	LUT4 #(
		.INIT('h0100)
	) name6844 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12671_
	);
	LUT3 #(
		.INIT('h14)
	) name6845 (
		_w12612_,
		_w12613_,
		_w12616_,
		_w12672_
	);
	LUT4 #(
		.INIT('hfd00)
	) name6846 (
		_w12619_,
		_w12622_,
		_w12671_,
		_w12672_,
		_w12673_
	);
	LUT3 #(
		.INIT('ha8)
	) name6847 (
		_w12611_,
		_w12670_,
		_w12673_,
		_w12674_
	);
	LUT3 #(
		.INIT('h40)
	) name6848 (
		_w12615_,
		_w12613_,
		_w12616_,
		_w12675_
	);
	LUT4 #(
		.INIT('h00bf)
	) name6849 (
		_w12615_,
		_w12613_,
		_w12616_,
		_w12619_,
		_w12676_
	);
	LUT4 #(
		.INIT('h00fd)
	) name6850 (
		_w12619_,
		_w12622_,
		_w12671_,
		_w12676_,
		_w12677_
	);
	LUT4 #(
		.INIT('h7d78)
	) name6851 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12678_
	);
	LUT3 #(
		.INIT('he0)
	) name6852 (
		_w12612_,
		_w12613_,
		_w12619_,
		_w12679_
	);
	LUT4 #(
		.INIT('h6800)
	) name6853 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12619_,
		_w12680_
	);
	LUT4 #(
		.INIT('h0504)
	) name6854 (
		_w12631_,
		_w12619_,
		_w12680_,
		_w12678_,
		_w12681_
	);
	LUT3 #(
		.INIT('h32)
	) name6855 (
		_w12611_,
		_w12677_,
		_w12681_,
		_w12682_
	);
	LUT3 #(
		.INIT('h65)
	) name6856 (
		\u2_L3_reg[16]/NET0131 ,
		_w12674_,
		_w12682_,
		_w12683_
	);
	LUT2 #(
		.INIT('h4)
	) name6857 (
		_w12616_,
		_w12619_,
		_w12684_
	);
	LUT3 #(
		.INIT('h31)
	) name6858 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12685_
	);
	LUT2 #(
		.INIT('h8)
	) name6859 (
		_w12684_,
		_w12685_,
		_w12686_
	);
	LUT3 #(
		.INIT('h0e)
	) name6860 (
		_w12615_,
		_w12616_,
		_w12619_,
		_w12687_
	);
	LUT3 #(
		.INIT('hb0)
	) name6861 (
		_w12615_,
		_w12613_,
		_w12616_,
		_w12688_
	);
	LUT4 #(
		.INIT('h23af)
	) name6862 (
		_w12614_,
		_w12679_,
		_w12687_,
		_w12688_,
		_w12689_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6863 (
		_w12611_,
		_w12627_,
		_w12686_,
		_w12689_,
		_w12690_
	);
	LUT4 #(
		.INIT('hcaf1)
	) name6864 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12691_
	);
	LUT4 #(
		.INIT('h1000)
	) name6865 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12692_
	);
	LUT4 #(
		.INIT('h5504)
	) name6866 (
		_w12611_,
		_w12619_,
		_w12691_,
		_w12692_,
		_w12693_
	);
	LUT4 #(
		.INIT('h0021)
	) name6867 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12694_
	);
	LUT4 #(
		.INIT('hb59e)
	) name6868 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12695_
	);
	LUT2 #(
		.INIT('h1)
	) name6869 (
		_w12611_,
		_w12619_,
		_w12696_
	);
	LUT2 #(
		.INIT('h4)
	) name6870 (
		_w12695_,
		_w12696_,
		_w12697_
	);
	LUT3 #(
		.INIT('he7)
	) name6871 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12698_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name6872 (
		_w12616_,
		_w12619_,
		_w12637_,
		_w12698_,
		_w12699_
	);
	LUT3 #(
		.INIT('h10)
	) name6873 (
		_w12693_,
		_w12697_,
		_w12699_,
		_w12700_
	);
	LUT3 #(
		.INIT('h65)
	) name6874 (
		\u2_L3_reg[24]/NET0131 ,
		_w12690_,
		_w12700_,
		_w12701_
	);
	LUT4 #(
		.INIT('hfae5)
	) name6875 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12702_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name6876 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12703_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name6877 (
		_w12611_,
		_w12621_,
		_w12702_,
		_w12703_,
		_w12704_
	);
	LUT2 #(
		.INIT('h2)
	) name6878 (
		_w12619_,
		_w12704_,
		_w12705_
	);
	LUT4 #(
		.INIT('h0200)
	) name6879 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12706_
	);
	LUT3 #(
		.INIT('h0e)
	) name6880 (
		_w12615_,
		_w12613_,
		_w12619_,
		_w12707_
	);
	LUT4 #(
		.INIT('h0015)
	) name6881 (
		_w12694_,
		_w12703_,
		_w12707_,
		_w12706_,
		_w12708_
	);
	LUT2 #(
		.INIT('h1)
	) name6882 (
		_w12611_,
		_w12708_,
		_w12709_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name6883 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12616_,
		_w12710_
	);
	LUT2 #(
		.INIT('h2)
	) name6884 (
		_w12636_,
		_w12710_,
		_w12711_
	);
	LUT3 #(
		.INIT('h4c)
	) name6885 (
		_w12612_,
		_w12615_,
		_w12613_,
		_w12712_
	);
	LUT2 #(
		.INIT('h8)
	) name6886 (
		_w12634_,
		_w12712_,
		_w12713_
	);
	LUT4 #(
		.INIT('h0040)
	) name6887 (
		_w12612_,
		_w12615_,
		_w12616_,
		_w12619_,
		_w12714_
	);
	LUT3 #(
		.INIT('h07)
	) name6888 (
		_w12624_,
		_w12675_,
		_w12714_,
		_w12715_
	);
	LUT3 #(
		.INIT('h10)
	) name6889 (
		_w12711_,
		_w12713_,
		_w12715_,
		_w12716_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6890 (
		\u2_L3_reg[30]/NET0131 ,
		_w12705_,
		_w12709_,
		_w12716_,
		_w12717_
	);
	LUT4 #(
		.INIT('hfa3f)
	) name6891 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12718_
	);
	LUT2 #(
		.INIT('h2)
	) name6892 (
		_w12319_,
		_w12718_,
		_w12719_
	);
	LUT3 #(
		.INIT('ha2)
	) name6893 (
		_w12319_,
		_w12320_,
		_w12321_,
		_w12720_
	);
	LUT4 #(
		.INIT('h45f0)
	) name6894 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12721_
	);
	LUT3 #(
		.INIT('h54)
	) name6895 (
		_w12331_,
		_w12720_,
		_w12721_,
		_w12722_
	);
	LUT3 #(
		.INIT('h8c)
	) name6896 (
		_w12320_,
		_w12322_,
		_w12323_,
		_w12723_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6897 (
		_w12319_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12724_
	);
	LUT2 #(
		.INIT('h4)
	) name6898 (
		_w12723_,
		_w12724_,
		_w12725_
	);
	LUT4 #(
		.INIT('h0400)
	) name6899 (
		_w12319_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12726_
	);
	LUT4 #(
		.INIT('h0020)
	) name6900 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12727_
	);
	LUT4 #(
		.INIT('h0004)
	) name6901 (
		_w12326_,
		_w12331_,
		_w12727_,
		_w12726_,
		_w12728_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6902 (
		_w12719_,
		_w12722_,
		_w12725_,
		_w12728_,
		_w12729_
	);
	LUT4 #(
		.INIT('h2000)
	) name6903 (
		_w12320_,
		_w12321_,
		_w12322_,
		_w12323_,
		_w12730_
	);
	LUT4 #(
		.INIT('h0001)
	) name6904 (
		_w12319_,
		_w12343_,
		_w12659_,
		_w12730_,
		_w12731_
	);
	LUT3 #(
		.INIT('h02)
	) name6905 (
		_w12319_,
		_w12325_,
		_w12345_,
		_w12732_
	);
	LUT2 #(
		.INIT('h1)
	) name6906 (
		_w12731_,
		_w12732_,
		_w12733_
	);
	LUT3 #(
		.INIT('h56)
	) name6907 (
		\u2_L3_reg[3]/NET0131 ,
		_w12729_,
		_w12733_,
		_w12734_
	);
	LUT4 #(
		.INIT('h8228)
	) name6908 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12735_
	);
	LUT3 #(
		.INIT('he6)
	) name6909 (
		_w12159_,
		_w12160_,
		_w12158_,
		_w12736_
	);
	LUT4 #(
		.INIT('h0031)
	) name6910 (
		_w12169_,
		_w12352_,
		_w12736_,
		_w12735_,
		_w12737_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name6911 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12738_
	);
	LUT2 #(
		.INIT('h1)
	) name6912 (
		_w12156_,
		_w12738_,
		_w12739_
	);
	LUT4 #(
		.INIT('h00e6)
	) name6913 (
		_w12159_,
		_w12160_,
		_w12158_,
		_w12156_,
		_w12740_
	);
	LUT4 #(
		.INIT('hc700)
	) name6914 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12156_,
		_w12741_
	);
	LUT4 #(
		.INIT('h9ffd)
	) name6915 (
		_w12157_,
		_w12159_,
		_w12160_,
		_w12158_,
		_w12742_
	);
	LUT4 #(
		.INIT('hdc00)
	) name6916 (
		_w12550_,
		_w12740_,
		_w12741_,
		_w12742_,
		_w12743_
	);
	LUT4 #(
		.INIT('h3210)
	) name6917 (
		_w12155_,
		_w12739_,
		_w12743_,
		_w12737_,
		_w12744_
	);
	LUT2 #(
		.INIT('h9)
	) name6918 (
		\u2_L3_reg[9]/NET0131 ,
		_w12744_,
		_w12745_
	);
	LUT4 #(
		.INIT('hef2f)
	) name6919 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12746_
	);
	LUT4 #(
		.INIT('h0100)
	) name6920 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12747_
	);
	LUT4 #(
		.INIT('h0b08)
	) name6921 (
		_w12463_,
		_w12466_,
		_w12747_,
		_w12746_,
		_w12748_
	);
	LUT4 #(
		.INIT('h0121)
	) name6922 (
		_w12459_,
		_w12461_,
		_w12464_,
		_w12466_,
		_w12749_
	);
	LUT4 #(
		.INIT('h9fff)
	) name6923 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12750_
	);
	LUT4 #(
		.INIT('h8000)
	) name6924 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12466_,
		_w12751_
	);
	LUT4 #(
		.INIT('h0100)
	) name6925 (
		_w12522_,
		_w12751_,
		_w12749_,
		_w12750_,
		_w12752_
	);
	LUT4 #(
		.INIT('h0008)
	) name6926 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12466_,
		_w12753_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name6927 (
		_w12459_,
		_w12460_,
		_w12461_,
		_w12464_,
		_w12754_
	);
	LUT3 #(
		.INIT('h31)
	) name6928 (
		_w12466_,
		_w12753_,
		_w12754_,
		_w12755_
	);
	LUT4 #(
		.INIT('hd800)
	) name6929 (
		_w12458_,
		_w12748_,
		_w12752_,
		_w12755_,
		_w12756_
	);
	LUT2 #(
		.INIT('h9)
	) name6930 (
		\u2_L3_reg[18]/P0001 ,
		_w12756_,
		_w12757_
	);
	LUT4 #(
		.INIT('hc693)
	) name6931 (
		decrypt_pad,
		\u2_R2_reg[1]/NET0131 ,
		\u2_uk_K_r2_reg[26]/NET0131 ,
		\u2_uk_K_r2_reg[46]/NET0131 ,
		_w12758_
	);
	LUT4 #(
		.INIT('hc963)
	) name6932 (
		decrypt_pad,
		\u2_R2_reg[5]/NET0131 ,
		\u2_uk_K_r2_reg[19]/NET0131 ,
		\u2_uk_K_r2_reg[24]/NET0131 ,
		_w12759_
	);
	LUT4 #(
		.INIT('hc693)
	) name6933 (
		decrypt_pad,
		\u2_R2_reg[2]/NET0131 ,
		\u2_uk_K_r2_reg[41]/NET0131 ,
		\u2_uk_K_r2_reg[4]/NET0131 ,
		_w12760_
	);
	LUT4 #(
		.INIT('hc963)
	) name6934 (
		decrypt_pad,
		\u2_R2_reg[32]/NET0131 ,
		\u2_uk_K_r2_reg[25]/NET0131 ,
		\u2_uk_K_r2_reg[5]/NET0131 ,
		_w12761_
	);
	LUT4 #(
		.INIT('hbb83)
	) name6935 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12762_
	);
	LUT4 #(
		.INIT('hc963)
	) name6936 (
		decrypt_pad,
		\u2_R2_reg[3]/NET0131 ,
		\u2_uk_K_r2_reg[13]/NET0131 ,
		\u2_uk_K_r2_reg[18]/NET0131 ,
		_w12763_
	);
	LUT2 #(
		.INIT('h4)
	) name6937 (
		_w12762_,
		_w12763_,
		_w12764_
	);
	LUT4 #(
		.INIT('h04a4)
	) name6938 (
		_w12758_,
		_w12760_,
		_w12761_,
		_w12763_,
		_w12765_
	);
	LUT2 #(
		.INIT('h8)
	) name6939 (
		_w12759_,
		_w12761_,
		_w12766_
	);
	LUT2 #(
		.INIT('h6)
	) name6940 (
		_w12759_,
		_w12761_,
		_w12767_
	);
	LUT4 #(
		.INIT('h0144)
	) name6941 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12768_
	);
	LUT4 #(
		.INIT('hc963)
	) name6942 (
		decrypt_pad,
		\u2_R2_reg[4]/NET0131 ,
		\u2_uk_K_r2_reg[48]/NET0131 ,
		\u2_uk_K_r2_reg[53]/P0001 ,
		_w12769_
	);
	LUT3 #(
		.INIT('h10)
	) name6943 (
		_w12768_,
		_w12765_,
		_w12769_,
		_w12770_
	);
	LUT2 #(
		.INIT('h8)
	) name6944 (
		_w12760_,
		_w12763_,
		_w12771_
	);
	LUT3 #(
		.INIT('h20)
	) name6945 (
		_w12760_,
		_w12761_,
		_w12763_,
		_w12772_
	);
	LUT4 #(
		.INIT('h0800)
	) name6946 (
		_w12759_,
		_w12760_,
		_w12761_,
		_w12763_,
		_w12773_
	);
	LUT4 #(
		.INIT('hb6fe)
	) name6947 (
		_w12759_,
		_w12760_,
		_w12761_,
		_w12763_,
		_w12774_
	);
	LUT2 #(
		.INIT('h2)
	) name6948 (
		_w12758_,
		_w12774_,
		_w12775_
	);
	LUT2 #(
		.INIT('h4)
	) name6949 (
		_w12760_,
		_w12763_,
		_w12776_
	);
	LUT3 #(
		.INIT('hce)
	) name6950 (
		_w12758_,
		_w12760_,
		_w12763_,
		_w12777_
	);
	LUT3 #(
		.INIT('h31)
	) name6951 (
		_w12766_,
		_w12769_,
		_w12777_,
		_w12778_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6952 (
		_w12764_,
		_w12770_,
		_w12775_,
		_w12778_,
		_w12779_
	);
	LUT4 #(
		.INIT('heff4)
	) name6953 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12780_
	);
	LUT4 #(
		.INIT('h7dbd)
	) name6954 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12781_
	);
	LUT4 #(
		.INIT('h0155)
	) name6955 (
		_w12763_,
		_w12769_,
		_w12780_,
		_w12781_,
		_w12782_
	);
	LUT2 #(
		.INIT('h1)
	) name6956 (
		_w12758_,
		_w12759_,
		_w12783_
	);
	LUT4 #(
		.INIT('h1000)
	) name6957 (
		_w12758_,
		_w12760_,
		_w12761_,
		_w12763_,
		_w12784_
	);
	LUT3 #(
		.INIT('h07)
	) name6958 (
		_w12772_,
		_w12783_,
		_w12784_,
		_w12785_
	);
	LUT2 #(
		.INIT('h4)
	) name6959 (
		_w12782_,
		_w12785_,
		_w12786_
	);
	LUT3 #(
		.INIT('h65)
	) name6960 (
		\u2_L2_reg[31]/NET0131 ,
		_w12779_,
		_w12786_,
		_w12787_
	);
	LUT4 #(
		.INIT('hc963)
	) name6961 (
		decrypt_pad,
		\u2_R2_reg[24]/NET0131 ,
		\u2_uk_K_r2_reg[15]/NET0131 ,
		\u2_uk_K_r2_reg[52]/NET0131 ,
		_w12788_
	);
	LUT4 #(
		.INIT('hc693)
	) name6962 (
		decrypt_pad,
		\u2_R2_reg[20]/NET0131 ,
		\u2_uk_K_r2_reg[31]/NET0131 ,
		\u2_uk_K_r2_reg[49]/NET0131 ,
		_w12789_
	);
	LUT4 #(
		.INIT('hc963)
	) name6963 (
		decrypt_pad,
		\u2_R2_reg[22]/NET0131 ,
		\u2_uk_K_r2_reg[0]/NET0131 ,
		\u2_uk_K_r2_reg[9]/NET0131 ,
		_w12790_
	);
	LUT4 #(
		.INIT('hc693)
	) name6964 (
		decrypt_pad,
		\u2_R2_reg[21]/NET0131 ,
		\u2_uk_K_r2_reg[42]/NET0131 ,
		\u2_uk_K_r2_reg[9]/NET0131 ,
		_w12791_
	);
	LUT4 #(
		.INIT('hc693)
	) name6965 (
		decrypt_pad,
		\u2_R2_reg[23]/NET0131 ,
		\u2_uk_K_r2_reg[22]/NET0131 ,
		\u2_uk_K_r2_reg[44]/NET0131 ,
		_w12792_
	);
	LUT4 #(
		.INIT('h4155)
	) name6966 (
		_w12792_,
		_w12789_,
		_w12790_,
		_w12791_,
		_w12793_
	);
	LUT4 #(
		.INIT('hc963)
	) name6967 (
		decrypt_pad,
		\u2_R2_reg[25]/NET0131 ,
		\u2_uk_K_r2_reg[38]/NET0131 ,
		\u2_uk_K_r2_reg[43]/NET0131 ,
		_w12794_
	);
	LUT4 #(
		.INIT('haa8a)
	) name6968 (
		_w12792_,
		_w12789_,
		_w12794_,
		_w12791_,
		_w12795_
	);
	LUT3 #(
		.INIT('he6)
	) name6969 (
		_w12789_,
		_w12790_,
		_w12791_,
		_w12796_
	);
	LUT3 #(
		.INIT('h13)
	) name6970 (
		_w12795_,
		_w12793_,
		_w12796_,
		_w12797_
	);
	LUT4 #(
		.INIT('h0080)
	) name6971 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12798_
	);
	LUT2 #(
		.INIT('h2)
	) name6972 (
		_w12789_,
		_w12794_,
		_w12799_
	);
	LUT2 #(
		.INIT('h1)
	) name6973 (
		_w12792_,
		_w12790_,
		_w12800_
	);
	LUT3 #(
		.INIT('hce)
	) name6974 (
		_w12792_,
		_w12790_,
		_w12791_,
		_w12801_
	);
	LUT3 #(
		.INIT('h31)
	) name6975 (
		_w12799_,
		_w12798_,
		_w12801_,
		_w12802_
	);
	LUT3 #(
		.INIT('h45)
	) name6976 (
		_w12788_,
		_w12797_,
		_w12802_,
		_w12803_
	);
	LUT4 #(
		.INIT('h0002)
	) name6977 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12804_
	);
	LUT4 #(
		.INIT('h27fd)
	) name6978 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12805_
	);
	LUT2 #(
		.INIT('h2)
	) name6979 (
		_w12792_,
		_w12805_,
		_w12806_
	);
	LUT4 #(
		.INIT('h0415)
	) name6980 (
		_w12792_,
		_w12789_,
		_w12794_,
		_w12791_,
		_w12807_
	);
	LUT4 #(
		.INIT('h0b07)
	) name6981 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12808_
	);
	LUT3 #(
		.INIT('h0e)
	) name6982 (
		_w12800_,
		_w12807_,
		_w12808_,
		_w12809_
	);
	LUT3 #(
		.INIT('he0)
	) name6983 (
		_w12806_,
		_w12809_,
		_w12788_,
		_w12810_
	);
	LUT4 #(
		.INIT('h5155)
	) name6984 (
		_w12792_,
		_w12789_,
		_w12794_,
		_w12791_,
		_w12811_
	);
	LUT3 #(
		.INIT('h01)
	) name6985 (
		_w12790_,
		_w12811_,
		_w12795_,
		_w12812_
	);
	LUT4 #(
		.INIT('h7077)
	) name6986 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12813_
	);
	LUT4 #(
		.INIT('haa02)
	) name6987 (
		_w12792_,
		_w12789_,
		_w12794_,
		_w12790_,
		_w12814_
	);
	LUT3 #(
		.INIT('h01)
	) name6988 (
		_w12789_,
		_w12794_,
		_w12791_,
		_w12815_
	);
	LUT4 #(
		.INIT('h45cf)
	) name6989 (
		_w12800_,
		_w12813_,
		_w12814_,
		_w12815_,
		_w12816_
	);
	LUT2 #(
		.INIT('h4)
	) name6990 (
		_w12812_,
		_w12816_,
		_w12817_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6991 (
		\u2_L2_reg[11]/NET0131 ,
		_w12810_,
		_w12803_,
		_w12817_,
		_w12818_
	);
	LUT4 #(
		.INIT('hc693)
	) name6992 (
		decrypt_pad,
		\u2_R2_reg[28]/NET0131 ,
		\u2_uk_K_r2_reg[0]/NET0131 ,
		\u2_uk_K_r2_reg[22]/NET0131 ,
		_w12819_
	);
	LUT4 #(
		.INIT('hc963)
	) name6993 (
		decrypt_pad,
		\u2_R2_reg[25]/NET0131 ,
		\u2_uk_K_r2_reg[45]/NET0131 ,
		\u2_uk_K_r2_reg[50]/NET0131 ,
		_w12820_
	);
	LUT4 #(
		.INIT('hc693)
	) name6994 (
		decrypt_pad,
		\u2_R2_reg[24]/NET0131 ,
		\u2_uk_K_r2_reg[15]/NET0131 ,
		\u2_uk_K_r2_reg[37]/NET0131 ,
		_w12821_
	);
	LUT4 #(
		.INIT('hc963)
	) name6995 (
		decrypt_pad,
		\u2_R2_reg[29]/NET0131 ,
		\u2_uk_K_r2_reg[14]/NET0131 ,
		\u2_uk_K_r2_reg[23]/NET0131 ,
		_w12822_
	);
	LUT2 #(
		.INIT('h4)
	) name6996 (
		_w12821_,
		_w12822_,
		_w12823_
	);
	LUT3 #(
		.INIT('h40)
	) name6997 (
		_w12820_,
		_w12821_,
		_w12822_,
		_w12824_
	);
	LUT3 #(
		.INIT('h9f)
	) name6998 (
		_w12820_,
		_w12821_,
		_w12822_,
		_w12825_
	);
	LUT4 #(
		.INIT('hc963)
	) name6999 (
		decrypt_pad,
		\u2_R2_reg[27]/NET0131 ,
		\u2_uk_K_r2_reg[35]/NET0131 ,
		\u2_uk_K_r2_reg[44]/NET0131 ,
		_w12826_
	);
	LUT4 #(
		.INIT('hc963)
	) name7000 (
		decrypt_pad,
		\u2_R2_reg[26]/NET0131 ,
		\u2_uk_K_r2_reg[2]/NET0131 ,
		\u2_uk_K_r2_reg[35]/NET0131 ,
		_w12827_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name7001 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12828_
	);
	LUT3 #(
		.INIT('h01)
	) name7002 (
		_w12826_,
		_w12828_,
		_w12825_,
		_w12829_
	);
	LUT3 #(
		.INIT('h9b)
	) name7003 (
		_w12820_,
		_w12827_,
		_w12822_,
		_w12830_
	);
	LUT2 #(
		.INIT('h8)
	) name7004 (
		_w12826_,
		_w12821_,
		_w12831_
	);
	LUT4 #(
		.INIT('h1000)
	) name7005 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12832_
	);
	LUT4 #(
		.INIT('heffe)
	) name7006 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12833_
	);
	LUT3 #(
		.INIT('hb0)
	) name7007 (
		_w12830_,
		_w12831_,
		_w12833_,
		_w12834_
	);
	LUT3 #(
		.INIT('h8a)
	) name7008 (
		_w12819_,
		_w12829_,
		_w12834_,
		_w12835_
	);
	LUT3 #(
		.INIT('hd8)
	) name7009 (
		_w12820_,
		_w12826_,
		_w12827_,
		_w12836_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name7010 (
		_w12826_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12837_
	);
	LUT2 #(
		.INIT('h4)
	) name7011 (
		_w12836_,
		_w12837_,
		_w12838_
	);
	LUT4 #(
		.INIT('h0010)
	) name7012 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12839_
	);
	LUT2 #(
		.INIT('h9)
	) name7013 (
		_w12821_,
		_w12827_,
		_w12840_
	);
	LUT3 #(
		.INIT('hb0)
	) name7014 (
		_w12820_,
		_w12826_,
		_w12822_,
		_w12841_
	);
	LUT4 #(
		.INIT('h23af)
	) name7015 (
		_w12826_,
		_w12840_,
		_w12839_,
		_w12841_,
		_w12842_
	);
	LUT4 #(
		.INIT('h2002)
	) name7016 (
		_w12820_,
		_w12826_,
		_w12821_,
		_w12827_,
		_w12843_
	);
	LUT4 #(
		.INIT('h0020)
	) name7017 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12844_
	);
	LUT4 #(
		.INIT('hefdf)
	) name7018 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12845_
	);
	LUT4 #(
		.INIT('hef9a)
	) name7019 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12846_
	);
	LUT3 #(
		.INIT('h31)
	) name7020 (
		_w12826_,
		_w12843_,
		_w12846_,
		_w12847_
	);
	LUT4 #(
		.INIT('hba00)
	) name7021 (
		_w12819_,
		_w12838_,
		_w12842_,
		_w12847_,
		_w12848_
	);
	LUT3 #(
		.INIT('h65)
	) name7022 (
		\u2_L2_reg[22]/NET0131 ,
		_w12835_,
		_w12848_,
		_w12849_
	);
	LUT4 #(
		.INIT('h0400)
	) name7023 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12850_
	);
	LUT4 #(
		.INIT('hfb05)
	) name7024 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12851_
	);
	LUT4 #(
		.INIT('h00c1)
	) name7025 (
		_w12758_,
		_w12760_,
		_w12761_,
		_w12763_,
		_w12852_
	);
	LUT3 #(
		.INIT('h10)
	) name7026 (
		_w12759_,
		_w12760_,
		_w12761_,
		_w12853_
	);
	LUT4 #(
		.INIT('h0200)
	) name7027 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12854_
	);
	LUT4 #(
		.INIT('h7d7f)
	) name7028 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12855_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7029 (
		_w12763_,
		_w12851_,
		_w12852_,
		_w12855_,
		_w12856_
	);
	LUT4 #(
		.INIT('h0028)
	) name7030 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12857_
	);
	LUT4 #(
		.INIT('h0090)
	) name7031 (
		_w12758_,
		_w12759_,
		_w12761_,
		_w12769_,
		_w12858_
	);
	LUT3 #(
		.INIT('ha8)
	) name7032 (
		_w12763_,
		_w12857_,
		_w12858_,
		_w12859_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7033 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12860_
	);
	LUT3 #(
		.INIT('h09)
	) name7034 (
		_w12759_,
		_w12761_,
		_w12763_,
		_w12861_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name7035 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w12862_
	);
	LUT3 #(
		.INIT('hb0)
	) name7036 (
		_w12860_,
		_w12861_,
		_w12862_,
		_w12863_
	);
	LUT4 #(
		.INIT('h3210)
	) name7037 (
		_w12769_,
		_w12859_,
		_w12863_,
		_w12856_,
		_w12864_
	);
	LUT2 #(
		.INIT('h9)
	) name7038 (
		\u2_L2_reg[17]/NET0131 ,
		_w12864_,
		_w12865_
	);
	LUT4 #(
		.INIT('hc963)
	) name7039 (
		decrypt_pad,
		\u2_R2_reg[15]/NET0131 ,
		\u2_uk_K_r2_reg[10]/NET0131 ,
		\u2_uk_K_r2_reg[47]/NET0131 ,
		_w12866_
	);
	LUT4 #(
		.INIT('hc693)
	) name7040 (
		decrypt_pad,
		\u2_R2_reg[13]/NET0131 ,
		\u2_uk_K_r2_reg[13]/NET0131 ,
		\u2_uk_K_r2_reg[33]/NET0131 ,
		_w12867_
	);
	LUT4 #(
		.INIT('hc693)
	) name7041 (
		decrypt_pad,
		\u2_R2_reg[17]/NET0131 ,
		\u2_uk_K_r2_reg[3]/NET0131 ,
		\u2_uk_K_r2_reg[55]/NET0131 ,
		_w12868_
	);
	LUT4 #(
		.INIT('hc693)
	) name7042 (
		decrypt_pad,
		\u2_R2_reg[12]/NET0131 ,
		\u2_uk_K_r2_reg[19]/NET0131 ,
		\u2_uk_K_r2_reg[39]/NET0131 ,
		_w12869_
	);
	LUT4 #(
		.INIT('h8000)
	) name7043 (
		_w12866_,
		_w12868_,
		_w12869_,
		_w12867_,
		_w12870_
	);
	LUT2 #(
		.INIT('h2)
	) name7044 (
		_w12866_,
		_w12868_,
		_w12871_
	);
	LUT4 #(
		.INIT('h0002)
	) name7045 (
		_w12866_,
		_w12868_,
		_w12869_,
		_w12867_,
		_w12872_
	);
	LUT4 #(
		.INIT('hc963)
	) name7046 (
		decrypt_pad,
		\u2_R2_reg[16]/NET0131 ,
		\u2_uk_K_r2_reg[18]/NET0131 ,
		\u2_uk_K_r2_reg[55]/NET0131 ,
		_w12873_
	);
	LUT4 #(
		.INIT('hc963)
	) name7047 (
		decrypt_pad,
		\u2_R2_reg[14]/NET0131 ,
		\u2_uk_K_r2_reg[34]/NET0131 ,
		\u2_uk_K_r2_reg[39]/NET0131 ,
		_w12874_
	);
	LUT4 #(
		.INIT('h2000)
	) name7048 (
		_w12866_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12875_
	);
	LUT4 #(
		.INIT('h0008)
	) name7049 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12876_
	);
	LUT4 #(
		.INIT('h0001)
	) name7050 (
		_w12872_,
		_w12875_,
		_w12876_,
		_w12873_,
		_w12877_
	);
	LUT4 #(
		.INIT('hb1f5)
	) name7051 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12878_
	);
	LUT3 #(
		.INIT('h10)
	) name7052 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12879_
	);
	LUT4 #(
		.INIT('h0001)
	) name7053 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12880_
	);
	LUT4 #(
		.INIT('heffe)
	) name7054 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12881_
	);
	LUT3 #(
		.INIT('he0)
	) name7055 (
		_w12866_,
		_w12878_,
		_w12881_,
		_w12882_
	);
	LUT3 #(
		.INIT('h40)
	) name7056 (
		_w12870_,
		_w12877_,
		_w12882_,
		_w12883_
	);
	LUT2 #(
		.INIT('h1)
	) name7057 (
		_w12866_,
		_w12868_,
		_w12884_
	);
	LUT4 #(
		.INIT('h0001)
	) name7058 (
		_w12866_,
		_w12868_,
		_w12869_,
		_w12867_,
		_w12885_
	);
	LUT4 #(
		.INIT('h3ffe)
	) name7059 (
		_w12866_,
		_w12868_,
		_w12869_,
		_w12867_,
		_w12886_
	);
	LUT2 #(
		.INIT('h2)
	) name7060 (
		_w12874_,
		_w12886_,
		_w12887_
	);
	LUT2 #(
		.INIT('h2)
	) name7061 (
		_w12868_,
		_w12869_,
		_w12888_
	);
	LUT4 #(
		.INIT('h0008)
	) name7062 (
		_w12866_,
		_w12868_,
		_w12869_,
		_w12867_,
		_w12889_
	);
	LUT2 #(
		.INIT('h2)
	) name7063 (
		_w12873_,
		_w12889_,
		_w12890_
	);
	LUT4 #(
		.INIT('h2000)
	) name7064 (
		_w12866_,
		_w12868_,
		_w12869_,
		_w12867_,
		_w12891_
	);
	LUT4 #(
		.INIT('h0020)
	) name7065 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12892_
	);
	LUT4 #(
		.INIT('h0014)
	) name7066 (
		_w12866_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12893_
	);
	LUT3 #(
		.INIT('h01)
	) name7067 (
		_w12891_,
		_w12892_,
		_w12893_,
		_w12894_
	);
	LUT3 #(
		.INIT('h40)
	) name7068 (
		_w12887_,
		_w12890_,
		_w12894_,
		_w12895_
	);
	LUT4 #(
		.INIT('h0400)
	) name7069 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12896_
	);
	LUT4 #(
		.INIT('hfad8)
	) name7070 (
		_w12866_,
		_w12880_,
		_w12892_,
		_w12896_,
		_w12897_
	);
	LUT3 #(
		.INIT('h08)
	) name7071 (
		_w12869_,
		_w12867_,
		_w12874_,
		_w12898_
	);
	LUT2 #(
		.INIT('h8)
	) name7072 (
		_w12871_,
		_w12898_,
		_w12899_
	);
	LUT2 #(
		.INIT('h1)
	) name7073 (
		_w12897_,
		_w12899_,
		_w12900_
	);
	LUT4 #(
		.INIT('ha955)
	) name7074 (
		\u2_L2_reg[20]/NET0131 ,
		_w12883_,
		_w12895_,
		_w12900_,
		_w12901_
	);
	LUT4 #(
		.INIT('h67dc)
	) name7075 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12902_
	);
	LUT4 #(
		.INIT('hd2f7)
	) name7076 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12903_
	);
	LUT4 #(
		.INIT('h0040)
	) name7077 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12904_
	);
	LUT4 #(
		.INIT('h00d8)
	) name7078 (
		_w12792_,
		_w12902_,
		_w12903_,
		_w12904_,
		_w12905_
	);
	LUT4 #(
		.INIT('h9aff)
	) name7079 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12906_
	);
	LUT4 #(
		.INIT('haa02)
	) name7080 (
		_w12792_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12907_
	);
	LUT4 #(
		.INIT('h9297)
	) name7081 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12908_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name7082 (
		_w12792_,
		_w12906_,
		_w12907_,
		_w12908_,
		_w12909_
	);
	LUT4 #(
		.INIT('h0800)
	) name7083 (
		_w12792_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w12910_
	);
	LUT2 #(
		.INIT('h1)
	) name7084 (
		_w12804_,
		_w12910_,
		_w12911_
	);
	LUT4 #(
		.INIT('hd800)
	) name7085 (
		_w12788_,
		_w12909_,
		_w12905_,
		_w12911_,
		_w12912_
	);
	LUT2 #(
		.INIT('h6)
	) name7086 (
		\u2_L2_reg[29]/NET0131 ,
		_w12912_,
		_w12913_
	);
	LUT4 #(
		.INIT('hc963)
	) name7087 (
		decrypt_pad,
		\u2_R2_reg[8]/NET0131 ,
		\u2_uk_K_r2_reg[17]/NET0131 ,
		\u2_uk_K_r2_reg[54]/NET0131 ,
		_w12914_
	);
	LUT4 #(
		.INIT('hc963)
	) name7088 (
		decrypt_pad,
		\u2_R2_reg[5]/NET0131 ,
		\u2_uk_K_r2_reg[41]/NET0131 ,
		\u2_uk_K_r2_reg[46]/NET0131 ,
		_w12915_
	);
	LUT4 #(
		.INIT('hc693)
	) name7089 (
		decrypt_pad,
		\u2_R2_reg[9]/NET0131 ,
		\u2_uk_K_r2_reg[34]/NET0131 ,
		\u2_uk_K_r2_reg[54]/NET0131 ,
		_w12916_
	);
	LUT4 #(
		.INIT('hc693)
	) name7090 (
		decrypt_pad,
		\u2_R2_reg[4]/NET0131 ,
		\u2_uk_K_r2_reg[10]/NET0131 ,
		\u2_uk_K_r2_reg[5]/NET0131 ,
		_w12917_
	);
	LUT3 #(
		.INIT('h04)
	) name7091 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12918_
	);
	LUT3 #(
		.INIT('hd9)
	) name7092 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12919_
	);
	LUT4 #(
		.INIT('hc693)
	) name7093 (
		decrypt_pad,
		\u2_R2_reg[6]/NET0131 ,
		\u2_uk_K_r2_reg[12]/NET0131 ,
		\u2_uk_K_r2_reg[32]/NET0131 ,
		_w12920_
	);
	LUT4 #(
		.INIT('h0026)
	) name7094 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12921_
	);
	LUT4 #(
		.INIT('hc963)
	) name7095 (
		decrypt_pad,
		\u2_R2_reg[7]/NET0131 ,
		\u2_uk_K_r2_reg[26]/NET0131 ,
		\u2_uk_K_r2_reg[6]/NET0131 ,
		_w12922_
	);
	LUT4 #(
		.INIT('h4000)
	) name7096 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12923_
	);
	LUT3 #(
		.INIT('h15)
	) name7097 (
		_w12921_,
		_w12922_,
		_w12923_,
		_w12924_
	);
	LUT2 #(
		.INIT('h8)
	) name7098 (
		_w12917_,
		_w12920_,
		_w12925_
	);
	LUT4 #(
		.INIT('h4bfb)
	) name7099 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12926_
	);
	LUT3 #(
		.INIT('hcd)
	) name7100 (
		_w12915_,
		_w12920_,
		_w12922_,
		_w12927_
	);
	LUT2 #(
		.INIT('h2)
	) name7101 (
		_w12916_,
		_w12917_,
		_w12928_
	);
	LUT4 #(
		.INIT('h084c)
	) name7102 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12929_
	);
	LUT4 #(
		.INIT('h0eee)
	) name7103 (
		_w12922_,
		_w12926_,
		_w12927_,
		_w12929_,
		_w12930_
	);
	LUT3 #(
		.INIT('h15)
	) name7104 (
		_w12914_,
		_w12924_,
		_w12930_,
		_w12931_
	);
	LUT4 #(
		.INIT('hbcfc)
	) name7105 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12932_
	);
	LUT4 #(
		.INIT('h080c)
	) name7106 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12933_
	);
	LUT3 #(
		.INIT('h0d)
	) name7107 (
		_w12915_,
		_w12920_,
		_w12922_,
		_w12934_
	);
	LUT4 #(
		.INIT('hf200)
	) name7108 (
		_w12914_,
		_w12932_,
		_w12933_,
		_w12934_,
		_w12935_
	);
	LUT4 #(
		.INIT('h0080)
	) name7109 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12936_
	);
	LUT4 #(
		.INIT('h0010)
	) name7110 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12937_
	);
	LUT4 #(
		.INIT('h8a00)
	) name7111 (
		_w12915_,
		_w12917_,
		_w12920_,
		_w12922_,
		_w12938_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7112 (
		_w12914_,
		_w12937_,
		_w12938_,
		_w12936_,
		_w12939_
	);
	LUT4 #(
		.INIT('hfc54)
	) name7113 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12940_
	);
	LUT4 #(
		.INIT('hdc00)
	) name7114 (
		_w12915_,
		_w12917_,
		_w12920_,
		_w12922_,
		_w12941_
	);
	LUT2 #(
		.INIT('h4)
	) name7115 (
		_w12940_,
		_w12941_,
		_w12942_
	);
	LUT3 #(
		.INIT('h01)
	) name7116 (
		_w12939_,
		_w12942_,
		_w12935_,
		_w12943_
	);
	LUT3 #(
		.INIT('h65)
	) name7117 (
		\u2_L2_reg[2]/NET0131 ,
		_w12931_,
		_w12943_,
		_w12944_
	);
	LUT4 #(
		.INIT('h0040)
	) name7118 (
		_w12866_,
		_w12868_,
		_w12869_,
		_w12874_,
		_w12945_
	);
	LUT3 #(
		.INIT('h01)
	) name7119 (
		_w12885_,
		_w12898_,
		_w12945_,
		_w12946_
	);
	LUT3 #(
		.INIT('hce)
	) name7120 (
		_w12868_,
		_w12867_,
		_w12874_,
		_w12947_
	);
	LUT2 #(
		.INIT('h8)
	) name7121 (
		_w12866_,
		_w12869_,
		_w12948_
	);
	LUT4 #(
		.INIT('h0008)
	) name7122 (
		_w12866_,
		_w12868_,
		_w12869_,
		_w12874_,
		_w12949_
	);
	LUT3 #(
		.INIT('h0b)
	) name7123 (
		_w12947_,
		_w12948_,
		_w12949_,
		_w12950_
	);
	LUT4 #(
		.INIT('h1333)
	) name7124 (
		_w12881_,
		_w12873_,
		_w12946_,
		_w12950_,
		_w12951_
	);
	LUT3 #(
		.INIT('h02)
	) name7125 (
		_w12866_,
		_w12879_,
		_w12876_,
		_w12952_
	);
	LUT4 #(
		.INIT('h4404)
	) name7126 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12953_
	);
	LUT3 #(
		.INIT('h01)
	) name7127 (
		_w12866_,
		_w12892_,
		_w12953_,
		_w12954_
	);
	LUT3 #(
		.INIT('h90)
	) name7128 (
		_w12869_,
		_w12867_,
		_w12874_,
		_w12955_
	);
	LUT4 #(
		.INIT('h8200)
	) name7129 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12956_
	);
	LUT4 #(
		.INIT('haa02)
	) name7130 (
		_w12873_,
		_w12952_,
		_w12954_,
		_w12956_,
		_w12957_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name7131 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w12958_
	);
	LUT2 #(
		.INIT('h1)
	) name7132 (
		_w12866_,
		_w12958_,
		_w12959_
	);
	LUT3 #(
		.INIT('h13)
	) name7133 (
		_w12871_,
		_w12875_,
		_w12898_,
		_w12960_
	);
	LUT2 #(
		.INIT('h4)
	) name7134 (
		_w12959_,
		_w12960_,
		_w12961_
	);
	LUT4 #(
		.INIT('h5655)
	) name7135 (
		\u2_L2_reg[10]/NET0131 ,
		_w12957_,
		_w12951_,
		_w12961_,
		_w12962_
	);
	LUT3 #(
		.INIT('h02)
	) name7136 (
		_w12821_,
		_w12827_,
		_w12822_,
		_w12963_
	);
	LUT4 #(
		.INIT('h4004)
	) name7137 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12964_
	);
	LUT4 #(
		.INIT('h0012)
	) name7138 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12965_
	);
	LUT4 #(
		.INIT('h00bf)
	) name7139 (
		_w12826_,
		_w12821_,
		_w12827_,
		_w12819_,
		_w12966_
	);
	LUT2 #(
		.INIT('h4)
	) name7140 (
		_w12965_,
		_w12966_,
		_w12967_
	);
	LUT3 #(
		.INIT('h21)
	) name7141 (
		_w12820_,
		_w12826_,
		_w12822_,
		_w12968_
	);
	LUT3 #(
		.INIT('h1b)
	) name7142 (
		_w12820_,
		_w12826_,
		_w12827_,
		_w12969_
	);
	LUT3 #(
		.INIT('h31)
	) name7143 (
		_w12823_,
		_w12968_,
		_w12969_,
		_w12970_
	);
	LUT3 #(
		.INIT('h40)
	) name7144 (
		_w12964_,
		_w12967_,
		_w12970_,
		_w12971_
	);
	LUT4 #(
		.INIT('h3332)
	) name7145 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12972_
	);
	LUT3 #(
		.INIT('h8c)
	) name7146 (
		_w12820_,
		_w12826_,
		_w12821_,
		_w12973_
	);
	LUT2 #(
		.INIT('h4)
	) name7147 (
		_w12972_,
		_w12973_,
		_w12974_
	);
	LUT4 #(
		.INIT('h0600)
	) name7148 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w12975_
	);
	LUT2 #(
		.INIT('h9)
	) name7149 (
		_w12821_,
		_w12822_,
		_w12976_
	);
	LUT4 #(
		.INIT('h5100)
	) name7150 (
		_w12820_,
		_w12826_,
		_w12821_,
		_w12827_,
		_w12977_
	);
	LUT4 #(
		.INIT('h2022)
	) name7151 (
		_w12819_,
		_w12844_,
		_w12976_,
		_w12977_,
		_w12978_
	);
	LUT3 #(
		.INIT('h10)
	) name7152 (
		_w12975_,
		_w12974_,
		_w12978_,
		_w12979_
	);
	LUT3 #(
		.INIT('ha9)
	) name7153 (
		\u2_L2_reg[12]/NET0131 ,
		_w12971_,
		_w12979_,
		_w12980_
	);
	LUT4 #(
		.INIT('h2000)
	) name7154 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12981_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name7155 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12982_
	);
	LUT4 #(
		.INIT('h0400)
	) name7156 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12983_
	);
	LUT4 #(
		.INIT('hf9ed)
	) name7157 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12984_
	);
	LUT4 #(
		.INIT('h0313)
	) name7158 (
		_w12914_,
		_w12922_,
		_w12982_,
		_w12984_,
		_w12985_
	);
	LUT3 #(
		.INIT('h8e)
	) name7159 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12986_
	);
	LUT4 #(
		.INIT('h3010)
	) name7160 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12987_
	);
	LUT3 #(
		.INIT('h02)
	) name7161 (
		_w12922_,
		_w12986_,
		_w12987_,
		_w12988_
	);
	LUT3 #(
		.INIT('hd0)
	) name7162 (
		_w12915_,
		_w12916_,
		_w12922_,
		_w12989_
	);
	LUT2 #(
		.INIT('h8)
	) name7163 (
		_w12925_,
		_w12989_,
		_w12990_
	);
	LUT3 #(
		.INIT('h51)
	) name7164 (
		_w12914_,
		_w12928_,
		_w12927_,
		_w12991_
	);
	LUT3 #(
		.INIT('h10)
	) name7165 (
		_w12990_,
		_w12988_,
		_w12991_,
		_w12992_
	);
	LUT4 #(
		.INIT('h0002)
	) name7166 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12993_
	);
	LUT4 #(
		.INIT('h002a)
	) name7167 (
		_w12914_,
		_w12927_,
		_w12929_,
		_w12993_,
		_w12994_
	);
	LUT4 #(
		.INIT('h5140)
	) name7168 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12995_
	);
	LUT3 #(
		.INIT('h01)
	) name7169 (
		_w12915_,
		_w12916_,
		_w12920_,
		_w12996_
	);
	LUT4 #(
		.INIT('hf3ee)
	) name7170 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w12997_
	);
	LUT4 #(
		.INIT('h80c4)
	) name7171 (
		_w12922_,
		_w12982_,
		_w12997_,
		_w12995_,
		_w12998_
	);
	LUT2 #(
		.INIT('h8)
	) name7172 (
		_w12994_,
		_w12998_,
		_w12999_
	);
	LUT4 #(
		.INIT('h999a)
	) name7173 (
		\u2_L2_reg[13]/NET0131 ,
		_w12985_,
		_w12992_,
		_w12999_,
		_w13000_
	);
	LUT4 #(
		.INIT('hc963)
	) name7174 (
		decrypt_pad,
		\u2_R2_reg[20]/NET0131 ,
		\u2_uk_K_r2_reg[31]/NET0131 ,
		\u2_uk_K_r2_reg[36]/NET0131 ,
		_w13001_
	);
	LUT4 #(
		.INIT('hc693)
	) name7175 (
		decrypt_pad,
		\u2_R2_reg[19]/NET0131 ,
		\u2_uk_K_r2_reg[21]/NET0131 ,
		\u2_uk_K_r2_reg[43]/NET0131 ,
		_w13002_
	);
	LUT4 #(
		.INIT('hc963)
	) name7176 (
		decrypt_pad,
		\u2_R2_reg[16]/NET0131 ,
		\u2_uk_K_r2_reg[16]/NET0131 ,
		\u2_uk_K_r2_reg[49]/NET0131 ,
		_w13003_
	);
	LUT4 #(
		.INIT('hc693)
	) name7177 (
		decrypt_pad,
		\u2_R2_reg[17]/NET0131 ,
		\u2_uk_K_r2_reg[16]/NET0131 ,
		\u2_uk_K_r2_reg[7]/NET0131 ,
		_w13004_
	);
	LUT4 #(
		.INIT('hc963)
	) name7178 (
		decrypt_pad,
		\u2_R2_reg[18]/NET0131 ,
		\u2_uk_K_r2_reg[1]/NET0131 ,
		\u2_uk_K_r2_reg[38]/NET0131 ,
		_w13005_
	);
	LUT4 #(
		.INIT('hc963)
	) name7179 (
		decrypt_pad,
		\u2_R2_reg[21]/NET0131 ,
		\u2_uk_K_r2_reg[28]/NET0131 ,
		\u2_uk_K_r2_reg[37]/NET0131 ,
		_w13006_
	);
	LUT4 #(
		.INIT('h30d0)
	) name7180 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13007_
	);
	LUT4 #(
		.INIT('hc52f)
	) name7181 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13008_
	);
	LUT2 #(
		.INIT('h2)
	) name7182 (
		_w13002_,
		_w13008_,
		_w13009_
	);
	LUT2 #(
		.INIT('h1)
	) name7183 (
		_w13002_,
		_w13005_,
		_w13010_
	);
	LUT3 #(
		.INIT('hf6)
	) name7184 (
		_w13004_,
		_w13006_,
		_w13003_,
		_w13011_
	);
	LUT2 #(
		.INIT('h2)
	) name7185 (
		_w13010_,
		_w13011_,
		_w13012_
	);
	LUT2 #(
		.INIT('h9)
	) name7186 (
		_w13004_,
		_w13005_,
		_w13013_
	);
	LUT4 #(
		.INIT('h0600)
	) name7187 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13014_
	);
	LUT4 #(
		.INIT('h1000)
	) name7188 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13015_
	);
	LUT3 #(
		.INIT('h80)
	) name7189 (
		_w13004_,
		_w13006_,
		_w13003_,
		_w13016_
	);
	LUT2 #(
		.INIT('h4)
	) name7190 (
		_w13002_,
		_w13005_,
		_w13017_
	);
	LUT4 #(
		.INIT('h0013)
	) name7191 (
		_w13016_,
		_w13015_,
		_w13017_,
		_w13014_,
		_w13018_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7192 (
		_w13001_,
		_w13009_,
		_w13012_,
		_w13018_,
		_w13019_
	);
	LUT4 #(
		.INIT('h2000)
	) name7193 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13020_
	);
	LUT4 #(
		.INIT('h0100)
	) name7194 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13021_
	);
	LUT3 #(
		.INIT('h08)
	) name7195 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13022_
	);
	LUT4 #(
		.INIT('hd6a7)
	) name7196 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13023_
	);
	LUT2 #(
		.INIT('h1)
	) name7197 (
		_w13002_,
		_w13023_,
		_w13024_
	);
	LUT3 #(
		.INIT('h8a)
	) name7198 (
		_w13002_,
		_w13006_,
		_w13003_,
		_w13025_
	);
	LUT4 #(
		.INIT('h4000)
	) name7199 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13026_
	);
	LUT4 #(
		.INIT('hbffd)
	) name7200 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13027_
	);
	LUT4 #(
		.INIT('hef00)
	) name7201 (
		_w13022_,
		_w13007_,
		_w13025_,
		_w13027_,
		_w13028_
	);
	LUT4 #(
		.INIT('hfdfb)
	) name7202 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13029_
	);
	LUT4 #(
		.INIT('h0040)
	) name7203 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13030_
	);
	LUT4 #(
		.INIT('hffb7)
	) name7204 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13031_
	);
	LUT3 #(
		.INIT('hd8)
	) name7205 (
		_w13002_,
		_w13029_,
		_w13031_,
		_w13032_
	);
	LUT4 #(
		.INIT('hf400)
	) name7206 (
		_w13024_,
		_w13028_,
		_w13001_,
		_w13032_,
		_w13033_
	);
	LUT3 #(
		.INIT('h65)
	) name7207 (
		\u2_L2_reg[14]/NET0131 ,
		_w13019_,
		_w13033_,
		_w13034_
	);
	LUT4 #(
		.INIT('hc693)
	) name7208 (
		decrypt_pad,
		\u2_R2_reg[28]/NET0131 ,
		\u2_uk_K_r2_reg[29]/NET0131 ,
		\u2_uk_K_r2_reg[51]/NET0131 ,
		_w13035_
	);
	LUT4 #(
		.INIT('hc693)
	) name7209 (
		decrypt_pad,
		\u2_R2_reg[30]/NET0131 ,
		\u2_uk_K_r2_reg[2]/NET0131 ,
		\u2_uk_K_r2_reg[52]/NET0131 ,
		_w13036_
	);
	LUT4 #(
		.INIT('hc693)
	) name7210 (
		decrypt_pad,
		\u2_R2_reg[1]/NET0131 ,
		\u2_uk_K_r2_reg[45]/NET0131 ,
		\u2_uk_K_r2_reg[8]/NET0131 ,
		_w13037_
	);
	LUT4 #(
		.INIT('hc693)
	) name7211 (
		decrypt_pad,
		\u2_R2_reg[29]/NET0131 ,
		\u2_uk_K_r2_reg[1]/NET0131 ,
		\u2_uk_K_r2_reg[23]/NET0131 ,
		_w13038_
	);
	LUT4 #(
		.INIT('h2600)
	) name7212 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13039_
	);
	LUT4 #(
		.INIT('hc963)
	) name7213 (
		decrypt_pad,
		\u2_R2_reg[32]/NET0131 ,
		\u2_uk_K_r2_reg[42]/NET0131 ,
		\u2_uk_K_r2_reg[51]/NET0131 ,
		_w13040_
	);
	LUT2 #(
		.INIT('h4)
	) name7214 (
		_w13039_,
		_w13040_,
		_w13041_
	);
	LUT2 #(
		.INIT('h1)
	) name7215 (
		_w13037_,
		_w13038_,
		_w13042_
	);
	LUT4 #(
		.INIT('hc693)
	) name7216 (
		decrypt_pad,
		\u2_R2_reg[31]/P0001 ,
		\u2_uk_K_r2_reg[14]/NET0131 ,
		\u2_uk_K_r2_reg[36]/NET0131 ,
		_w13043_
	);
	LUT4 #(
		.INIT('h0100)
	) name7217 (
		_w13035_,
		_w13037_,
		_w13038_,
		_w13043_,
		_w13044_
	);
	LUT2 #(
		.INIT('h2)
	) name7218 (
		_w13037_,
		_w13038_,
		_w13045_
	);
	LUT3 #(
		.INIT('h73)
	) name7219 (
		_w13035_,
		_w13036_,
		_w13043_,
		_w13046_
	);
	LUT3 #(
		.INIT('h51)
	) name7220 (
		_w13044_,
		_w13045_,
		_w13046_,
		_w13047_
	);
	LUT4 #(
		.INIT('hfef0)
	) name7221 (
		_w13036_,
		_w13037_,
		_w13038_,
		_w13043_,
		_w13048_
	);
	LUT2 #(
		.INIT('h2)
	) name7222 (
		_w13035_,
		_w13048_,
		_w13049_
	);
	LUT3 #(
		.INIT('h4b)
	) name7223 (
		_w13035_,
		_w13037_,
		_w13038_,
		_w13050_
	);
	LUT4 #(
		.INIT('hbf00)
	) name7224 (
		_w13035_,
		_w13036_,
		_w13038_,
		_w13043_,
		_w13051_
	);
	LUT3 #(
		.INIT('h45)
	) name7225 (
		_w13040_,
		_w13050_,
		_w13051_,
		_w13052_
	);
	LUT4 #(
		.INIT('h7077)
	) name7226 (
		_w13041_,
		_w13047_,
		_w13049_,
		_w13052_,
		_w13053_
	);
	LUT4 #(
		.INIT('h1089)
	) name7227 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13054_
	);
	LUT4 #(
		.INIT('h0400)
	) name7228 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13055_
	);
	LUT3 #(
		.INIT('h01)
	) name7229 (
		_w13043_,
		_w13055_,
		_w13054_,
		_w13056_
	);
	LUT4 #(
		.INIT('h0010)
	) name7230 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13057_
	);
	LUT4 #(
		.INIT('h4000)
	) name7231 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13058_
	);
	LUT3 #(
		.INIT('h02)
	) name7232 (
		_w13043_,
		_w13058_,
		_w13057_,
		_w13059_
	);
	LUT2 #(
		.INIT('h1)
	) name7233 (
		_w13056_,
		_w13059_,
		_w13060_
	);
	LUT3 #(
		.INIT('h56)
	) name7234 (
		\u2_L2_reg[15]/NET0131 ,
		_w13053_,
		_w13060_,
		_w13061_
	);
	LUT3 #(
		.INIT('h01)
	) name7235 (
		_w12868_,
		_w12869_,
		_w12874_,
		_w13062_
	);
	LUT4 #(
		.INIT('h084c)
	) name7236 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13063_
	);
	LUT4 #(
		.INIT('hfda8)
	) name7237 (
		_w12866_,
		_w12896_,
		_w13062_,
		_w13063_,
		_w13064_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name7238 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13065_
	);
	LUT3 #(
		.INIT('h45)
	) name7239 (
		_w12873_,
		_w13064_,
		_w13065_,
		_w13066_
	);
	LUT4 #(
		.INIT('hf5f1)
	) name7240 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13067_
	);
	LUT4 #(
		.INIT('h6dff)
	) name7241 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13068_
	);
	LUT4 #(
		.INIT('h08aa)
	) name7242 (
		_w12866_,
		_w12873_,
		_w13067_,
		_w13068_,
		_w13069_
	);
	LUT2 #(
		.INIT('h8)
	) name7243 (
		_w12884_,
		_w12955_,
		_w13070_
	);
	LUT4 #(
		.INIT('hdf4f)
	) name7244 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13071_
	);
	LUT4 #(
		.INIT('h4000)
	) name7245 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13072_
	);
	LUT4 #(
		.INIT('hbcff)
	) name7246 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13073_
	);
	LUT4 #(
		.INIT('h04cc)
	) name7247 (
		_w12866_,
		_w12873_,
		_w13071_,
		_w13073_,
		_w13074_
	);
	LUT3 #(
		.INIT('h01)
	) name7248 (
		_w13070_,
		_w13069_,
		_w13074_,
		_w13075_
	);
	LUT3 #(
		.INIT('h65)
	) name7249 (
		\u2_L2_reg[1]/NET0131 ,
		_w13066_,
		_w13075_,
		_w13076_
	);
	LUT3 #(
		.INIT('h06)
	) name7250 (
		_w13035_,
		_w13036_,
		_w13043_,
		_w13077_
	);
	LUT3 #(
		.INIT('h06)
	) name7251 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13078_
	);
	LUT3 #(
		.INIT('h0e)
	) name7252 (
		_w13042_,
		_w13077_,
		_w13078_,
		_w13079_
	);
	LUT2 #(
		.INIT('h1)
	) name7253 (
		_w13036_,
		_w13038_,
		_w13080_
	);
	LUT2 #(
		.INIT('h8)
	) name7254 (
		_w13037_,
		_w13038_,
		_w13081_
	);
	LUT4 #(
		.INIT('h2a00)
	) name7255 (
		_w13035_,
		_w13037_,
		_w13038_,
		_w13043_,
		_w13082_
	);
	LUT2 #(
		.INIT('h4)
	) name7256 (
		_w13080_,
		_w13082_,
		_w13083_
	);
	LUT4 #(
		.INIT('h00bf)
	) name7257 (
		_w13035_,
		_w13036_,
		_w13038_,
		_w13040_,
		_w13084_
	);
	LUT4 #(
		.INIT('h0010)
	) name7258 (
		_w13035_,
		_w13037_,
		_w13038_,
		_w13043_,
		_w13085_
	);
	LUT4 #(
		.INIT('h2000)
	) name7259 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13086_
	);
	LUT3 #(
		.INIT('h10)
	) name7260 (
		_w13085_,
		_w13086_,
		_w13084_,
		_w13087_
	);
	LUT3 #(
		.INIT('h10)
	) name7261 (
		_w13079_,
		_w13083_,
		_w13087_,
		_w13088_
	);
	LUT3 #(
		.INIT('h02)
	) name7262 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13089_
	);
	LUT4 #(
		.INIT('h0080)
	) name7263 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13090_
	);
	LUT3 #(
		.INIT('h01)
	) name7264 (
		_w13043_,
		_w13090_,
		_w13089_,
		_w13091_
	);
	LUT4 #(
		.INIT('hd800)
	) name7265 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13092_
	);
	LUT4 #(
		.INIT('hfb00)
	) name7266 (
		_w13036_,
		_w13037_,
		_w13038_,
		_w13043_,
		_w13093_
	);
	LUT2 #(
		.INIT('h4)
	) name7267 (
		_w13092_,
		_w13093_,
		_w13094_
	);
	LUT4 #(
		.INIT('h0804)
	) name7268 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13095_
	);
	LUT3 #(
		.INIT('h02)
	) name7269 (
		_w13040_,
		_w13057_,
		_w13095_,
		_w13096_
	);
	LUT3 #(
		.INIT('he0)
	) name7270 (
		_w13091_,
		_w13094_,
		_w13096_,
		_w13097_
	);
	LUT4 #(
		.INIT('h0100)
	) name7271 (
		_w13035_,
		_w13036_,
		_w13038_,
		_w13043_,
		_w13098_
	);
	LUT3 #(
		.INIT('h0b)
	) name7272 (
		_w13043_,
		_w13086_,
		_w13098_,
		_w13099_
	);
	LUT4 #(
		.INIT('ha955)
	) name7273 (
		\u2_L2_reg[21]/NET0131 ,
		_w13088_,
		_w13097_,
		_w13099_,
		_w13100_
	);
	LUT4 #(
		.INIT('hef99)
	) name7274 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w13101_
	);
	LUT4 #(
		.INIT('hfdfb)
	) name7275 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w13102_
	);
	LUT4 #(
		.INIT('h0455)
	) name7276 (
		_w12763_,
		_w12769_,
		_w13101_,
		_w13102_,
		_w13103_
	);
	LUT4 #(
		.INIT('h8000)
	) name7277 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w13104_
	);
	LUT4 #(
		.INIT('h5200)
	) name7278 (
		_w12758_,
		_w12759_,
		_w12761_,
		_w12763_,
		_w13105_
	);
	LUT2 #(
		.INIT('h1)
	) name7279 (
		_w13104_,
		_w13105_,
		_w13106_
	);
	LUT3 #(
		.INIT('h45)
	) name7280 (
		_w12771_,
		_w13103_,
		_w13106_,
		_w13107_
	);
	LUT4 #(
		.INIT('h8a00)
	) name7281 (
		_w12758_,
		_w12760_,
		_w12761_,
		_w12763_,
		_w13108_
	);
	LUT2 #(
		.INIT('h8)
	) name7282 (
		_w12767_,
		_w13108_,
		_w13109_
	);
	LUT4 #(
		.INIT('h002a)
	) name7283 (
		_w12769_,
		_w12772_,
		_w12783_,
		_w12850_,
		_w13110_
	);
	LUT4 #(
		.INIT('h0200)
	) name7284 (
		_w12758_,
		_w12759_,
		_w12761_,
		_w12763_,
		_w13111_
	);
	LUT3 #(
		.INIT('h01)
	) name7285 (
		_w12769_,
		_w12773_,
		_w13111_,
		_w13112_
	);
	LUT4 #(
		.INIT('h00e0)
	) name7286 (
		_w12758_,
		_w12760_,
		_w12761_,
		_w12763_,
		_w13113_
	);
	LUT3 #(
		.INIT('h81)
	) name7287 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w13114_
	);
	LUT3 #(
		.INIT('h0b)
	) name7288 (
		_w12783_,
		_w13113_,
		_w13114_,
		_w13115_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7289 (
		_w13109_,
		_w13110_,
		_w13112_,
		_w13115_,
		_w13116_
	);
	LUT3 #(
		.INIT('ha9)
	) name7290 (
		\u2_L2_reg[23]/NET0131 ,
		_w13107_,
		_w13116_,
		_w13117_
	);
	LUT4 #(
		.INIT('h5ea2)
	) name7291 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13118_
	);
	LUT4 #(
		.INIT('hafdd)
	) name7292 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13119_
	);
	LUT4 #(
		.INIT('hd7df)
	) name7293 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13120_
	);
	LUT4 #(
		.INIT('hd800)
	) name7294 (
		_w13002_,
		_w13118_,
		_w13119_,
		_w13120_,
		_w13121_
	);
	LUT2 #(
		.INIT('h2)
	) name7295 (
		_w13001_,
		_w13121_,
		_w13122_
	);
	LUT4 #(
		.INIT('hf7eb)
	) name7296 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13123_
	);
	LUT2 #(
		.INIT('h2)
	) name7297 (
		_w13002_,
		_w13123_,
		_w13124_
	);
	LUT3 #(
		.INIT('ha2)
	) name7298 (
		_w13002_,
		_w13004_,
		_w13005_,
		_w13125_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name7299 (
		_w13002_,
		_w13004_,
		_w13006_,
		_w13003_,
		_w13126_
	);
	LUT3 #(
		.INIT('h2a)
	) name7300 (
		_w13002_,
		_w13004_,
		_w13006_,
		_w13127_
	);
	LUT3 #(
		.INIT('h09)
	) name7301 (
		_w13004_,
		_w13005_,
		_w13003_,
		_w13128_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name7302 (
		_w13125_,
		_w13126_,
		_w13127_,
		_w13128_,
		_w13129_
	);
	LUT4 #(
		.INIT('h1000)
	) name7303 (
		_w13002_,
		_w13004_,
		_w13005_,
		_w13003_,
		_w13130_
	);
	LUT2 #(
		.INIT('h1)
	) name7304 (
		_w13020_,
		_w13130_,
		_w13131_
	);
	LUT4 #(
		.INIT('h0e00)
	) name7305 (
		_w13001_,
		_w13129_,
		_w13124_,
		_w13131_,
		_w13132_
	);
	LUT3 #(
		.INIT('h65)
	) name7306 (
		\u2_L2_reg[25]/NET0131 ,
		_w13122_,
		_w13132_,
		_w13133_
	);
	LUT3 #(
		.INIT('h02)
	) name7307 (
		_w12866_,
		_w12876_,
		_w12892_,
		_w13134_
	);
	LUT4 #(
		.INIT('h0094)
	) name7308 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13135_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name7309 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13136_
	);
	LUT4 #(
		.INIT('h0504)
	) name7310 (
		_w12866_,
		_w12873_,
		_w13135_,
		_w13136_,
		_w13137_
	);
	LUT2 #(
		.INIT('h1)
	) name7311 (
		_w13134_,
		_w13137_,
		_w13138_
	);
	LUT4 #(
		.INIT('h0010)
	) name7312 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13139_
	);
	LUT4 #(
		.INIT('h0004)
	) name7313 (
		_w12872_,
		_w12873_,
		_w13072_,
		_w13139_,
		_w13140_
	);
	LUT4 #(
		.INIT('hf3f7)
	) name7314 (
		_w12866_,
		_w12868_,
		_w12869_,
		_w12867_,
		_w13141_
	);
	LUT4 #(
		.INIT('h7775)
	) name7315 (
		_w12868_,
		_w12869_,
		_w12867_,
		_w12874_,
		_w13142_
	);
	LUT3 #(
		.INIT('h51)
	) name7316 (
		_w12866_,
		_w12869_,
		_w12874_,
		_w13143_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name7317 (
		_w12874_,
		_w13141_,
		_w13142_,
		_w13143_,
		_w13144_
	);
	LUT3 #(
		.INIT('h80)
	) name7318 (
		_w12866_,
		_w12867_,
		_w12874_,
		_w13145_
	);
	LUT2 #(
		.INIT('h4)
	) name7319 (
		_w12888_,
		_w13145_,
		_w13146_
	);
	LUT4 #(
		.INIT('h00fd)
	) name7320 (
		_w12869_,
		_w12867_,
		_w12874_,
		_w12873_,
		_w13147_
	);
	LUT3 #(
		.INIT('h10)
	) name7321 (
		_w12891_,
		_w12892_,
		_w13147_,
		_w13148_
	);
	LUT4 #(
		.INIT('h7077)
	) name7322 (
		_w13140_,
		_w13144_,
		_w13146_,
		_w13148_,
		_w13149_
	);
	LUT3 #(
		.INIT('h56)
	) name7323 (
		\u2_L2_reg[26]/NET0131 ,
		_w13138_,
		_w13149_,
		_w13150_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name7324 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w13151_
	);
	LUT2 #(
		.INIT('h8)
	) name7325 (
		_w12922_,
		_w13151_,
		_w13152_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name7326 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w13153_
	);
	LUT3 #(
		.INIT('h10)
	) name7327 (
		_w12915_,
		_w12917_,
		_w12920_,
		_w13154_
	);
	LUT4 #(
		.INIT('h0001)
	) name7328 (
		_w12918_,
		_w12922_,
		_w12981_,
		_w13154_,
		_w13155_
	);
	LUT4 #(
		.INIT('h6100)
	) name7329 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w13156_
	);
	LUT2 #(
		.INIT('h1)
	) name7330 (
		_w12914_,
		_w13156_,
		_w13157_
	);
	LUT4 #(
		.INIT('hba00)
	) name7331 (
		_w13152_,
		_w13153_,
		_w13155_,
		_w13157_,
		_w13158_
	);
	LUT4 #(
		.INIT('h0010)
	) name7332 (
		_w12922_,
		_w12981_,
		_w13151_,
		_w13154_,
		_w13159_
	);
	LUT4 #(
		.INIT('h8280)
	) name7333 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w13160_
	);
	LUT4 #(
		.INIT('hef00)
	) name7334 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12922_,
		_w13161_
	);
	LUT2 #(
		.INIT('h4)
	) name7335 (
		_w13160_,
		_w13161_,
		_w13162_
	);
	LUT3 #(
		.INIT('h0b)
	) name7336 (
		_w12915_,
		_w12916_,
		_w12922_,
		_w13163_
	);
	LUT2 #(
		.INIT('h2)
	) name7337 (
		_w12917_,
		_w12920_,
		_w13164_
	);
	LUT4 #(
		.INIT('h2022)
	) name7338 (
		_w12914_,
		_w12983_,
		_w13163_,
		_w13164_,
		_w13165_
	);
	LUT3 #(
		.INIT('he0)
	) name7339 (
		_w13159_,
		_w13162_,
		_w13165_,
		_w13166_
	);
	LUT3 #(
		.INIT('ha9)
	) name7340 (
		\u2_L2_reg[28]/NET0131 ,
		_w13158_,
		_w13166_,
		_w13167_
	);
	LUT4 #(
		.INIT('hd97b)
	) name7341 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w13168_
	);
	LUT2 #(
		.INIT('h2)
	) name7342 (
		_w12792_,
		_w13168_,
		_w13169_
	);
	LUT4 #(
		.INIT('heebf)
	) name7343 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w13170_
	);
	LUT4 #(
		.INIT('h0040)
	) name7344 (
		_w12792_,
		_w12789_,
		_w12794_,
		_w12790_,
		_w13171_
	);
	LUT4 #(
		.INIT('h0032)
	) name7345 (
		_w12792_,
		_w12804_,
		_w13170_,
		_w13171_,
		_w13172_
	);
	LUT3 #(
		.INIT('h45)
	) name7346 (
		_w12788_,
		_w13169_,
		_w13172_,
		_w13173_
	);
	LUT4 #(
		.INIT('h7c7f)
	) name7347 (
		_w12792_,
		_w12789_,
		_w12794_,
		_w12791_,
		_w13174_
	);
	LUT2 #(
		.INIT('h1)
	) name7348 (
		_w12790_,
		_w13174_,
		_w13175_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name7349 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w13176_
	);
	LUT3 #(
		.INIT('h80)
	) name7350 (
		_w12794_,
		_w12790_,
		_w12791_,
		_w13177_
	);
	LUT3 #(
		.INIT('h0e)
	) name7351 (
		_w12792_,
		_w13176_,
		_w13177_,
		_w13178_
	);
	LUT4 #(
		.INIT('h70d0)
	) name7352 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w13179_
	);
	LUT4 #(
		.INIT('h5501)
	) name7353 (
		_w12792_,
		_w12789_,
		_w12794_,
		_w12790_,
		_w13180_
	);
	LUT3 #(
		.INIT('h9e)
	) name7354 (
		_w12789_,
		_w12794_,
		_w12791_,
		_w13181_
	);
	LUT2 #(
		.INIT('h8)
	) name7355 (
		_w12792_,
		_w12790_,
		_w13182_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name7356 (
		_w13179_,
		_w13180_,
		_w13181_,
		_w13182_,
		_w13183_
	);
	LUT4 #(
		.INIT('h7500)
	) name7357 (
		_w12788_,
		_w13175_,
		_w13178_,
		_w13183_,
		_w13184_
	);
	LUT3 #(
		.INIT('h65)
	) name7358 (
		\u2_L2_reg[4]/NET0131 ,
		_w13173_,
		_w13184_,
		_w13185_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name7359 (
		_w12792_,
		_w12789_,
		_w12794_,
		_w12790_,
		_w13186_
	);
	LUT4 #(
		.INIT('hef00)
	) name7360 (
		_w12794_,
		_w12790_,
		_w12791_,
		_w12788_,
		_w13187_
	);
	LUT3 #(
		.INIT('he0)
	) name7361 (
		_w12791_,
		_w13186_,
		_w13187_,
		_w13188_
	);
	LUT4 #(
		.INIT('h4010)
	) name7362 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w13189_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name7363 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w13190_
	);
	LUT3 #(
		.INIT('h31)
	) name7364 (
		_w12792_,
		_w13189_,
		_w13190_,
		_w13191_
	);
	LUT4 #(
		.INIT('h4e55)
	) name7365 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w13192_
	);
	LUT2 #(
		.INIT('h2)
	) name7366 (
		_w12792_,
		_w13192_,
		_w13193_
	);
	LUT4 #(
		.INIT('h1001)
	) name7367 (
		_w12792_,
		_w12789_,
		_w12794_,
		_w12791_,
		_w13194_
	);
	LUT4 #(
		.INIT('h8000)
	) name7368 (
		_w12789_,
		_w12794_,
		_w12790_,
		_w12791_,
		_w13195_
	);
	LUT3 #(
		.INIT('h01)
	) name7369 (
		_w12788_,
		_w13195_,
		_w13194_,
		_w13196_
	);
	LUT4 #(
		.INIT('h7077)
	) name7370 (
		_w13188_,
		_w13191_,
		_w13193_,
		_w13196_,
		_w13197_
	);
	LUT2 #(
		.INIT('h4)
	) name7371 (
		_w12791_,
		_w13171_,
		_w13198_
	);
	LUT2 #(
		.INIT('h1)
	) name7372 (
		_w12812_,
		_w13198_,
		_w13199_
	);
	LUT3 #(
		.INIT('h65)
	) name7373 (
		\u2_L2_reg[19]/NET0131 ,
		_w13197_,
		_w13199_,
		_w13200_
	);
	LUT2 #(
		.INIT('h9)
	) name7374 (
		_w13035_,
		_w13037_,
		_w13201_
	);
	LUT4 #(
		.INIT('ha5ee)
	) name7375 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13202_
	);
	LUT2 #(
		.INIT('h1)
	) name7376 (
		_w13043_,
		_w13202_,
		_w13203_
	);
	LUT4 #(
		.INIT('hbfcf)
	) name7377 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13204_
	);
	LUT3 #(
		.INIT('h02)
	) name7378 (
		_w13036_,
		_w13037_,
		_w13038_,
		_w13205_
	);
	LUT4 #(
		.INIT('h0008)
	) name7379 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13206_
	);
	LUT4 #(
		.INIT('hb000)
	) name7380 (
		_w13035_,
		_w13036_,
		_w13038_,
		_w13043_,
		_w13207_
	);
	LUT4 #(
		.INIT('h1300)
	) name7381 (
		_w13201_,
		_w13206_,
		_w13207_,
		_w13204_,
		_w13208_
	);
	LUT3 #(
		.INIT('h8a)
	) name7382 (
		_w13040_,
		_w13203_,
		_w13208_,
		_w13209_
	);
	LUT4 #(
		.INIT('h0700)
	) name7383 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13210_
	);
	LUT4 #(
		.INIT('h7300)
	) name7384 (
		_w13036_,
		_w13037_,
		_w13038_,
		_w13043_,
		_w13211_
	);
	LUT2 #(
		.INIT('h4)
	) name7385 (
		_w13210_,
		_w13211_,
		_w13212_
	);
	LUT4 #(
		.INIT('h0040)
	) name7386 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13213_
	);
	LUT4 #(
		.INIT('h0080)
	) name7387 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13043_,
		_w13214_
	);
	LUT3 #(
		.INIT('h01)
	) name7388 (
		_w13085_,
		_w13214_,
		_w13213_,
		_w13215_
	);
	LUT4 #(
		.INIT('h0200)
	) name7389 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13216_
	);
	LUT2 #(
		.INIT('h4)
	) name7390 (
		_w13043_,
		_w13216_,
		_w13217_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name7391 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13218_
	);
	LUT4 #(
		.INIT('h0420)
	) name7392 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13219_
	);
	LUT4 #(
		.INIT('h2227)
	) name7393 (
		_w13043_,
		_w13205_,
		_w13219_,
		_w13216_,
		_w13220_
	);
	LUT4 #(
		.INIT('hba00)
	) name7394 (
		_w13040_,
		_w13212_,
		_w13215_,
		_w13220_,
		_w13221_
	);
	LUT3 #(
		.INIT('h65)
	) name7395 (
		\u2_L2_reg[27]/NET0131 ,
		_w13209_,
		_w13221_,
		_w13222_
	);
	LUT4 #(
		.INIT('h4022)
	) name7396 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13223_
	);
	LUT4 #(
		.INIT('h0104)
	) name7397 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13224_
	);
	LUT3 #(
		.INIT('h01)
	) name7398 (
		_w12826_,
		_w13224_,
		_w13223_,
		_w13225_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name7399 (
		_w12820_,
		_w12826_,
		_w12827_,
		_w12822_,
		_w13226_
	);
	LUT4 #(
		.INIT('hff2e)
	) name7400 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13227_
	);
	LUT2 #(
		.INIT('h8)
	) name7401 (
		_w13226_,
		_w13227_,
		_w13228_
	);
	LUT4 #(
		.INIT('h0080)
	) name7402 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13229_
	);
	LUT2 #(
		.INIT('h2)
	) name7403 (
		_w12819_,
		_w13229_,
		_w13230_
	);
	LUT3 #(
		.INIT('he0)
	) name7404 (
		_w13225_,
		_w13228_,
		_w13230_,
		_w13231_
	);
	LUT4 #(
		.INIT('h8008)
	) name7405 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13232_
	);
	LUT3 #(
		.INIT('h04)
	) name7406 (
		_w12819_,
		_w12845_,
		_w13232_,
		_w13233_
	);
	LUT4 #(
		.INIT('h5507)
	) name7407 (
		_w12826_,
		_w12824_,
		_w12968_,
		_w12963_,
		_w13234_
	);
	LUT2 #(
		.INIT('h8)
	) name7408 (
		_w13233_,
		_w13234_,
		_w13235_
	);
	LUT4 #(
		.INIT('h2202)
	) name7409 (
		_w12820_,
		_w12826_,
		_w12821_,
		_w12822_,
		_w13236_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name7410 (
		_w12826_,
		_w12840_,
		_w12832_,
		_w13236_,
		_w13237_
	);
	LUT4 #(
		.INIT('ha955)
	) name7411 (
		\u2_L2_reg[32]/NET0131 ,
		_w13231_,
		_w13235_,
		_w13237_,
		_w13238_
	);
	LUT4 #(
		.INIT('hc693)
	) name7412 (
		decrypt_pad,
		\u2_R2_reg[13]/NET0131 ,
		\u2_uk_K_r2_reg[20]/NET0131 ,
		\u2_uk_K_r2_reg[40]/NET0131 ,
		_w13239_
	);
	LUT4 #(
		.INIT('hc963)
	) name7413 (
		decrypt_pad,
		\u2_R2_reg[9]/NET0131 ,
		\u2_uk_K_r2_reg[3]/NET0131 ,
		\u2_uk_K_r2_reg[40]/NET0131 ,
		_w13240_
	);
	LUT4 #(
		.INIT('hc963)
	) name7414 (
		decrypt_pad,
		\u2_R2_reg[11]/NET0131 ,
		\u2_uk_K_r2_reg[12]/NET0131 ,
		\u2_uk_K_r2_reg[17]/NET0131 ,
		_w13241_
	);
	LUT3 #(
		.INIT('h0b)
	) name7415 (
		_w13239_,
		_w13240_,
		_w13241_,
		_w13242_
	);
	LUT4 #(
		.INIT('hc963)
	) name7416 (
		decrypt_pad,
		\u2_R2_reg[10]/NET0131 ,
		\u2_uk_K_r2_reg[11]/NET0131 ,
		\u2_uk_K_r2_reg[48]/NET0131 ,
		_w13243_
	);
	LUT4 #(
		.INIT('hc693)
	) name7417 (
		decrypt_pad,
		\u2_R2_reg[8]/NET0131 ,
		\u2_uk_K_r2_reg[11]/NET0131 ,
		\u2_uk_K_r2_reg[6]/NET0131 ,
		_w13244_
	);
	LUT4 #(
		.INIT('h3b0b)
	) name7418 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13245_
	);
	LUT4 #(
		.INIT('h1000)
	) name7419 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13246_
	);
	LUT4 #(
		.INIT('hc963)
	) name7420 (
		decrypt_pad,
		\u2_R2_reg[12]/NET0131 ,
		\u2_uk_K_r2_reg[27]/NET0131 ,
		\u2_uk_K_r2_reg[32]/NET0131 ,
		_w13247_
	);
	LUT4 #(
		.INIT('h5100)
	) name7421 (
		_w13246_,
		_w13242_,
		_w13245_,
		_w13247_,
		_w13248_
	);
	LUT2 #(
		.INIT('h6)
	) name7422 (
		_w13239_,
		_w13244_,
		_w13249_
	);
	LUT4 #(
		.INIT('h9990)
	) name7423 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13250_
	);
	LUT4 #(
		.INIT('h0990)
	) name7424 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13251_
	);
	LUT4 #(
		.INIT('h4000)
	) name7425 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13252_
	);
	LUT4 #(
		.INIT('h0400)
	) name7426 (
		_w13244_,
		_w13240_,
		_w13243_,
		_w13241_,
		_w13253_
	);
	LUT3 #(
		.INIT('h01)
	) name7427 (
		_w13247_,
		_w13253_,
		_w13252_,
		_w13254_
	);
	LUT4 #(
		.INIT('h2000)
	) name7428 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13255_
	);
	LUT4 #(
		.INIT('h0203)
	) name7429 (
		_w13244_,
		_w13240_,
		_w13243_,
		_w13241_,
		_w13256_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7430 (
		_w13241_,
		_w13255_,
		_w13249_,
		_w13256_,
		_w13257_
	);
	LUT4 #(
		.INIT('h4555)
	) name7431 (
		_w13248_,
		_w13251_,
		_w13254_,
		_w13257_,
		_w13258_
	);
	LUT4 #(
		.INIT('h95b5)
	) name7432 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13259_
	);
	LUT4 #(
		.INIT('h0001)
	) name7433 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13260_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name7434 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13261_
	);
	LUT4 #(
		.INIT('h08aa)
	) name7435 (
		_w13241_,
		_w13247_,
		_w13259_,
		_w13261_,
		_w13262_
	);
	LUT3 #(
		.INIT('h56)
	) name7436 (
		\u2_L2_reg[6]/NET0131 ,
		_w13258_,
		_w13262_,
		_w13263_
	);
	LUT3 #(
		.INIT('h02)
	) name7437 (
		_w13002_,
		_w13021_,
		_w13016_,
		_w13264_
	);
	LUT4 #(
		.INIT('h00b0)
	) name7438 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13265_
	);
	LUT4 #(
		.INIT('h4555)
	) name7439 (
		_w13002_,
		_w13004_,
		_w13006_,
		_w13003_,
		_w13266_
	);
	LUT2 #(
		.INIT('h4)
	) name7440 (
		_w13265_,
		_w13266_,
		_w13267_
	);
	LUT4 #(
		.INIT('hf7d9)
	) name7441 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13268_
	);
	LUT4 #(
		.INIT('h0155)
	) name7442 (
		_w13001_,
		_w13264_,
		_w13267_,
		_w13268_,
		_w13269_
	);
	LUT4 #(
		.INIT('h0400)
	) name7443 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13270_
	);
	LUT2 #(
		.INIT('h1)
	) name7444 (
		_w13002_,
		_w13270_,
		_w13271_
	);
	LUT3 #(
		.INIT('ha2)
	) name7445 (
		_w13002_,
		_w13006_,
		_w13003_,
		_w13272_
	);
	LUT3 #(
		.INIT('h54)
	) name7446 (
		_w13022_,
		_w13013_,
		_w13272_,
		_w13273_
	);
	LUT4 #(
		.INIT('haffe)
	) name7447 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13274_
	);
	LUT3 #(
		.INIT('h10)
	) name7448 (
		_w13002_,
		_w13005_,
		_w13003_,
		_w13275_
	);
	LUT4 #(
		.INIT('h00c4)
	) name7449 (
		_w13002_,
		_w13031_,
		_w13274_,
		_w13275_,
		_w13276_
	);
	LUT4 #(
		.INIT('hfc54)
	) name7450 (
		_w13001_,
		_w13271_,
		_w13273_,
		_w13276_,
		_w13277_
	);
	LUT3 #(
		.INIT('h65)
	) name7451 (
		\u2_L2_reg[8]/NET0131 ,
		_w13269_,
		_w13277_,
		_w13278_
	);
	LUT3 #(
		.INIT('h28)
	) name7452 (
		_w12820_,
		_w12821_,
		_w12822_,
		_w13279_
	);
	LUT4 #(
		.INIT('h6080)
	) name7453 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13280_
	);
	LUT4 #(
		.INIT('h0c02)
	) name7454 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13281_
	);
	LUT2 #(
		.INIT('h2)
	) name7455 (
		_w12826_,
		_w13281_,
		_w13282_
	);
	LUT3 #(
		.INIT('h21)
	) name7456 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w13283_
	);
	LUT4 #(
		.INIT('h5515)
	) name7457 (
		_w12826_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13284_
	);
	LUT3 #(
		.INIT('h10)
	) name7458 (
		_w13279_,
		_w13283_,
		_w13284_,
		_w13285_
	);
	LUT4 #(
		.INIT('h888a)
	) name7459 (
		_w12819_,
		_w13280_,
		_w13282_,
		_w13285_,
		_w13286_
	);
	LUT4 #(
		.INIT('h2080)
	) name7460 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13287_
	);
	LUT4 #(
		.INIT('h4c03)
	) name7461 (
		_w12820_,
		_w12821_,
		_w12827_,
		_w12822_,
		_w13288_
	);
	LUT4 #(
		.INIT('h3332)
	) name7462 (
		_w12819_,
		_w12839_,
		_w13288_,
		_w13287_,
		_w13289_
	);
	LUT4 #(
		.INIT('h3130)
	) name7463 (
		_w12826_,
		_w12819_,
		_w12839_,
		_w13281_,
		_w13290_
	);
	LUT4 #(
		.INIT('h00b1)
	) name7464 (
		_w12826_,
		_w13280_,
		_w13289_,
		_w13290_,
		_w13291_
	);
	LUT3 #(
		.INIT('h65)
	) name7465 (
		\u2_L2_reg[7]/NET0131 ,
		_w13286_,
		_w13291_,
		_w13292_
	);
	LUT4 #(
		.INIT('h9060)
	) name7466 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w13293_
	);
	LUT3 #(
		.INIT('h19)
	) name7467 (
		_w12758_,
		_w12759_,
		_w12761_,
		_w13294_
	);
	LUT4 #(
		.INIT('h0013)
	) name7468 (
		_w12776_,
		_w12854_,
		_w13294_,
		_w13293_,
		_w13295_
	);
	LUT4 #(
		.INIT('h0019)
	) name7469 (
		_w12758_,
		_w12759_,
		_w12761_,
		_w12763_,
		_w13296_
	);
	LUT3 #(
		.INIT('h60)
	) name7470 (
		_w12758_,
		_w12759_,
		_w12763_,
		_w13297_
	);
	LUT4 #(
		.INIT('hb7ef)
	) name7471 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w13298_
	);
	LUT4 #(
		.INIT('h0b00)
	) name7472 (
		_w12853_,
		_w13297_,
		_w13296_,
		_w13298_,
		_w13299_
	);
	LUT4 #(
		.INIT('hf77f)
	) name7473 (
		_w12758_,
		_w12759_,
		_w12760_,
		_w12761_,
		_w13300_
	);
	LUT2 #(
		.INIT('h1)
	) name7474 (
		_w12763_,
		_w13300_,
		_w13301_
	);
	LUT4 #(
		.INIT('h0e04)
	) name7475 (
		_w12769_,
		_w13299_,
		_w13301_,
		_w13295_,
		_w13302_
	);
	LUT2 #(
		.INIT('h9)
	) name7476 (
		\u2_L2_reg[9]/NET0131 ,
		_w13302_,
		_w13303_
	);
	LUT4 #(
		.INIT('h6979)
	) name7477 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13241_,
		_w13304_
	);
	LUT3 #(
		.INIT('h07)
	) name7478 (
		_w13244_,
		_w13243_,
		_w13241_,
		_w13305_
	);
	LUT4 #(
		.INIT('h0014)
	) name7479 (
		_w13239_,
		_w13244_,
		_w13243_,
		_w13241_,
		_w13306_
	);
	LUT4 #(
		.INIT('h0032)
	) name7480 (
		_w13243_,
		_w13255_,
		_w13304_,
		_w13306_,
		_w13307_
	);
	LUT3 #(
		.INIT('he0)
	) name7481 (
		_w13239_,
		_w13244_,
		_w13241_,
		_w13308_
	);
	LUT4 #(
		.INIT('h6800)
	) name7482 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13241_,
		_w13309_
	);
	LUT3 #(
		.INIT('h0d)
	) name7483 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13310_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name7484 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13311_
	);
	LUT4 #(
		.INIT('h0f02)
	) name7485 (
		_w13241_,
		_w13260_,
		_w13309_,
		_w13311_,
		_w13312_
	);
	LUT3 #(
		.INIT('h08)
	) name7486 (
		_w13244_,
		_w13243_,
		_w13241_,
		_w13313_
	);
	LUT4 #(
		.INIT('h0020)
	) name7487 (
		_w13244_,
		_w13240_,
		_w13243_,
		_w13241_,
		_w13314_
	);
	LUT4 #(
		.INIT('hbeff)
	) name7488 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13315_
	);
	LUT3 #(
		.INIT('h31)
	) name7489 (
		_w13241_,
		_w13314_,
		_w13315_,
		_w13316_
	);
	LUT4 #(
		.INIT('hd800)
	) name7490 (
		_w13247_,
		_w13307_,
		_w13312_,
		_w13316_,
		_w13317_
	);
	LUT2 #(
		.INIT('h9)
	) name7491 (
		\u2_L2_reg[16]/NET0131 ,
		_w13317_,
		_w13318_
	);
	LUT4 #(
		.INIT('hef2f)
	) name7492 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w13319_
	);
	LUT4 #(
		.INIT('h0100)
	) name7493 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w13320_
	);
	LUT4 #(
		.INIT('h0b08)
	) name7494 (
		_w12919_,
		_w12922_,
		_w13320_,
		_w13319_,
		_w13321_
	);
	LUT4 #(
		.INIT('h0121)
	) name7495 (
		_w12915_,
		_w12917_,
		_w12920_,
		_w12922_,
		_w13322_
	);
	LUT4 #(
		.INIT('h9fff)
	) name7496 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w13323_
	);
	LUT4 #(
		.INIT('h8000)
	) name7497 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12922_,
		_w13324_
	);
	LUT4 #(
		.INIT('h0100)
	) name7498 (
		_w12996_,
		_w13324_,
		_w13322_,
		_w13323_,
		_w13325_
	);
	LUT4 #(
		.INIT('h0008)
	) name7499 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12922_,
		_w13326_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name7500 (
		_w12915_,
		_w12916_,
		_w12917_,
		_w12920_,
		_w13327_
	);
	LUT3 #(
		.INIT('h31)
	) name7501 (
		_w12922_,
		_w13326_,
		_w13327_,
		_w13328_
	);
	LUT4 #(
		.INIT('hd800)
	) name7502 (
		_w12914_,
		_w13321_,
		_w13325_,
		_w13328_,
		_w13329_
	);
	LUT2 #(
		.INIT('h9)
	) name7503 (
		\u2_L2_reg[18]/P0001 ,
		_w13329_,
		_w13330_
	);
	LUT3 #(
		.INIT('hed)
	) name7504 (
		_w13239_,
		_w13244_,
		_w13243_,
		_w13331_
	);
	LUT3 #(
		.INIT('h20)
	) name7505 (
		_w13244_,
		_w13240_,
		_w13243_,
		_w13332_
	);
	LUT4 #(
		.INIT('hef00)
	) name7506 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13241_,
		_w13333_
	);
	LUT3 #(
		.INIT('h20)
	) name7507 (
		_w13331_,
		_w13332_,
		_w13333_,
		_w13334_
	);
	LUT4 #(
		.INIT('h0009)
	) name7508 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13335_
	);
	LUT4 #(
		.INIT('h6640)
	) name7509 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13336_
	);
	LUT3 #(
		.INIT('h01)
	) name7510 (
		_w13241_,
		_w13336_,
		_w13335_,
		_w13337_
	);
	LUT3 #(
		.INIT('h54)
	) name7511 (
		_w13247_,
		_w13334_,
		_w13337_,
		_w13338_
	);
	LUT2 #(
		.INIT('h4)
	) name7512 (
		_w13241_,
		_w13250_,
		_w13339_
	);
	LUT3 #(
		.INIT('h2a)
	) name7513 (
		_w13247_,
		_w13249_,
		_w13256_,
		_w13340_
	);
	LUT3 #(
		.INIT('hd0)
	) name7514 (
		_w13244_,
		_w13240_,
		_w13243_,
		_w13341_
	);
	LUT2 #(
		.INIT('h4)
	) name7515 (
		_w13243_,
		_w13241_,
		_w13342_
	);
	LUT4 #(
		.INIT('h153f)
	) name7516 (
		_w13308_,
		_w13310_,
		_w13342_,
		_w13341_,
		_w13343_
	);
	LUT3 #(
		.INIT('h40)
	) name7517 (
		_w13339_,
		_w13340_,
		_w13343_,
		_w13344_
	);
	LUT2 #(
		.INIT('h8)
	) name7518 (
		_w13239_,
		_w13240_,
		_w13345_
	);
	LUT3 #(
		.INIT('h53)
	) name7519 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13346_
	);
	LUT4 #(
		.INIT('h0700)
	) name7520 (
		_w13239_,
		_w13244_,
		_w13243_,
		_w13241_,
		_w13347_
	);
	LUT4 #(
		.INIT('h7077)
	) name7521 (
		_w13313_,
		_w13345_,
		_w13346_,
		_w13347_,
		_w13348_
	);
	LUT4 #(
		.INIT('ha955)
	) name7522 (
		\u2_L2_reg[24]/NET0131 ,
		_w13338_,
		_w13344_,
		_w13348_,
		_w13349_
	);
	LUT4 #(
		.INIT('h8c00)
	) name7523 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13350_
	);
	LUT4 #(
		.INIT('h00fb)
	) name7524 (
		_w13239_,
		_w13240_,
		_w13243_,
		_w13247_,
		_w13351_
	);
	LUT2 #(
		.INIT('h4)
	) name7525 (
		_w13350_,
		_w13351_,
		_w13352_
	);
	LUT4 #(
		.INIT('h0004)
	) name7526 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13353_
	);
	LUT4 #(
		.INIT('haa2a)
	) name7527 (
		_w13241_,
		_w13247_,
		_w13331_,
		_w13353_,
		_w13354_
	);
	LUT2 #(
		.INIT('h4)
	) name7528 (
		_w13352_,
		_w13354_,
		_w13355_
	);
	LUT4 #(
		.INIT('h23ef)
	) name7529 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13356_
	);
	LUT4 #(
		.INIT('h7000)
	) name7530 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13357_
	);
	LUT4 #(
		.INIT('h0c08)
	) name7531 (
		_w13241_,
		_w13247_,
		_w13357_,
		_w13356_,
		_w13358_
	);
	LUT2 #(
		.INIT('h1)
	) name7532 (
		_w13247_,
		_w13335_,
		_w13359_
	);
	LUT4 #(
		.INIT('h0200)
	) name7533 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13243_,
		_w13360_
	);
	LUT3 #(
		.INIT('h0d)
	) name7534 (
		_w13305_,
		_w13346_,
		_w13360_,
		_w13361_
	);
	LUT4 #(
		.INIT('hf700)
	) name7535 (
		_w13239_,
		_w13244_,
		_w13240_,
		_w13241_,
		_w13362_
	);
	LUT4 #(
		.INIT('hf040)
	) name7536 (
		_w13239_,
		_w13240_,
		_w13243_,
		_w13241_,
		_w13363_
	);
	LUT2 #(
		.INIT('h4)
	) name7537 (
		_w13362_,
		_w13363_,
		_w13364_
	);
	LUT4 #(
		.INIT('h00ea)
	) name7538 (
		_w13358_,
		_w13359_,
		_w13361_,
		_w13364_,
		_w13365_
	);
	LUT3 #(
		.INIT('h9a)
	) name7539 (
		\u2_L2_reg[30]/NET0131 ,
		_w13355_,
		_w13365_,
		_w13366_
	);
	LUT3 #(
		.INIT('h8a)
	) name7540 (
		_w13002_,
		_w13004_,
		_w13005_,
		_w13367_
	);
	LUT4 #(
		.INIT('h2f30)
	) name7541 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13368_
	);
	LUT2 #(
		.INIT('h1)
	) name7542 (
		_w13367_,
		_w13368_,
		_w13369_
	);
	LUT4 #(
		.INIT('hf5cf)
	) name7543 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13370_
	);
	LUT3 #(
		.INIT('h31)
	) name7544 (
		_w13002_,
		_w13001_,
		_w13370_,
		_w13371_
	);
	LUT3 #(
		.INIT('hb0)
	) name7545 (
		_w13005_,
		_w13006_,
		_w13003_,
		_w13372_
	);
	LUT4 #(
		.INIT('haa08)
	) name7546 (
		_w13002_,
		_w13004_,
		_w13006_,
		_w13003_,
		_w13373_
	);
	LUT2 #(
		.INIT('h4)
	) name7547 (
		_w13372_,
		_w13373_,
		_w13374_
	);
	LUT4 #(
		.INIT('h0040)
	) name7548 (
		_w13002_,
		_w13004_,
		_w13006_,
		_w13003_,
		_w13375_
	);
	LUT4 #(
		.INIT('h0004)
	) name7549 (
		_w13020_,
		_w13001_,
		_w13270_,
		_w13375_,
		_w13376_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name7550 (
		_w13369_,
		_w13371_,
		_w13374_,
		_w13376_,
		_w13377_
	);
	LUT3 #(
		.INIT('h02)
	) name7551 (
		_w13002_,
		_w13021_,
		_w13030_,
		_w13378_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name7552 (
		_w13004_,
		_w13005_,
		_w13006_,
		_w13003_,
		_w13379_
	);
	LUT3 #(
		.INIT('h10)
	) name7553 (
		_w13002_,
		_w13026_,
		_w13379_,
		_w13380_
	);
	LUT2 #(
		.INIT('h1)
	) name7554 (
		_w13378_,
		_w13380_,
		_w13381_
	);
	LUT3 #(
		.INIT('h56)
	) name7555 (
		\u2_L2_reg[3]/NET0131 ,
		_w13377_,
		_w13381_,
		_w13382_
	);
	LUT4 #(
		.INIT('hc963)
	) name7556 (
		decrypt_pad,
		\u2_R1_reg[26]/NET0131 ,
		\u2_uk_K_r1_reg[43]/NET0131 ,
		\u2_uk_K_r1_reg[49]/NET0131 ,
		_w13383_
	);
	LUT4 #(
		.INIT('hc963)
	) name7557 (
		decrypt_pad,
		\u2_R1_reg[25]/NET0131 ,
		\u2_uk_K_r1_reg[31]/NET0131 ,
		\u2_uk_K_r1_reg[9]/NET0131 ,
		_w13384_
	);
	LUT4 #(
		.INIT('hc963)
	) name7558 (
		decrypt_pad,
		\u2_R1_reg[24]/NET0131 ,
		\u2_uk_K_r1_reg[23]/NET0131 ,
		\u2_uk_K_r1_reg[29]/NET0131 ,
		_w13385_
	);
	LUT4 #(
		.INIT('hc963)
	) name7559 (
		decrypt_pad,
		\u2_R1_reg[29]/NET0131 ,
		\u2_uk_K_r1_reg[0]/NET0131 ,
		\u2_uk_K_r1_reg[37]/NET0131 ,
		_w13386_
	);
	LUT2 #(
		.INIT('h4)
	) name7560 (
		_w13385_,
		_w13386_,
		_w13387_
	);
	LUT4 #(
		.INIT('h0200)
	) name7561 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13388_
	);
	LUT4 #(
		.INIT('h0008)
	) name7562 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13389_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name7563 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13390_
	);
	LUT4 #(
		.INIT('hc693)
	) name7564 (
		decrypt_pad,
		\u2_R1_reg[28]/NET0131 ,
		\u2_uk_K_r1_reg[14]/NET0131 ,
		\u2_uk_K_r1_reg[8]/NET0131 ,
		_w13391_
	);
	LUT4 #(
		.INIT('h9cfc)
	) name7565 (
		_w13383_,
		_w13384_,
		_w13386_,
		_w13391_,
		_w13392_
	);
	LUT4 #(
		.INIT('hc963)
	) name7566 (
		decrypt_pad,
		\u2_R1_reg[27]/NET0131 ,
		\u2_uk_K_r1_reg[21]/NET0131 ,
		\u2_uk_K_r1_reg[31]/NET0131 ,
		_w13393_
	);
	LUT4 #(
		.INIT('h3b00)
	) name7567 (
		_w13385_,
		_w13390_,
		_w13392_,
		_w13393_,
		_w13394_
	);
	LUT2 #(
		.INIT('h4)
	) name7568 (
		_w13384_,
		_w13393_,
		_w13395_
	);
	LUT4 #(
		.INIT('heef2)
	) name7569 (
		_w13383_,
		_w13384_,
		_w13386_,
		_w13393_,
		_w13396_
	);
	LUT2 #(
		.INIT('h6)
	) name7570 (
		_w13383_,
		_w13385_,
		_w13397_
	);
	LUT4 #(
		.INIT('h0002)
	) name7571 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13398_
	);
	LUT4 #(
		.INIT('h5afd)
	) name7572 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13399_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name7573 (
		_w13385_,
		_w13395_,
		_w13396_,
		_w13399_,
		_w13400_
	);
	LUT4 #(
		.INIT('h1000)
	) name7574 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13401_
	);
	LUT4 #(
		.INIT('he3ff)
	) name7575 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13402_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name7576 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13403_
	);
	LUT3 #(
		.INIT('he0)
	) name7577 (
		_w13393_,
		_w13402_,
		_w13403_,
		_w13404_
	);
	LUT4 #(
		.INIT('h0100)
	) name7578 (
		_w13383_,
		_w13384_,
		_w13386_,
		_w13393_,
		_w13405_
	);
	LUT4 #(
		.INIT('h0084)
	) name7579 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13393_,
		_w13406_
	);
	LUT2 #(
		.INIT('h1)
	) name7580 (
		_w13405_,
		_w13406_,
		_w13407_
	);
	LUT4 #(
		.INIT('he400)
	) name7581 (
		_w13391_,
		_w13400_,
		_w13404_,
		_w13407_,
		_w13408_
	);
	LUT3 #(
		.INIT('h65)
	) name7582 (
		\u2_L1_reg[22]/NET0131 ,
		_w13394_,
		_w13408_,
		_w13409_
	);
	LUT4 #(
		.INIT('hc693)
	) name7583 (
		decrypt_pad,
		\u2_R1_reg[4]/NET0131 ,
		\u2_uk_K_r1_reg[10]/P0001 ,
		\u2_uk_K_r1_reg[34]/NET0131 ,
		_w13410_
	);
	LUT4 #(
		.INIT('hc963)
	) name7584 (
		decrypt_pad,
		\u2_R1_reg[3]/NET0131 ,
		\u2_uk_K_r1_reg[24]/NET0131 ,
		\u2_uk_K_r1_reg[32]/NET0131 ,
		_w13411_
	);
	LUT4 #(
		.INIT('hc963)
	) name7585 (
		decrypt_pad,
		\u2_R1_reg[2]/NET0131 ,
		\u2_uk_K_r1_reg[47]/NET0131 ,
		\u2_uk_K_r1_reg[55]/NET0131 ,
		_w13412_
	);
	LUT4 #(
		.INIT('hc963)
	) name7586 (
		decrypt_pad,
		\u2_R1_reg[32]/NET0131 ,
		\u2_uk_K_r1_reg[11]/NET0131 ,
		\u2_uk_K_r1_reg[19]/NET0131 ,
		_w13413_
	);
	LUT4 #(
		.INIT('hc963)
	) name7587 (
		decrypt_pad,
		\u2_R1_reg[1]/NET0131 ,
		\u2_uk_K_r1_reg[32]/NET0131 ,
		\u2_uk_K_r1_reg[40]/NET0131 ,
		_w13414_
	);
	LUT4 #(
		.INIT('hc693)
	) name7588 (
		decrypt_pad,
		\u2_R1_reg[5]/NET0131 ,
		\u2_uk_K_r1_reg[13]/NET0131 ,
		\u2_uk_K_r1_reg[5]/NET0131 ,
		_w13415_
	);
	LUT4 #(
		.INIT('hfdba)
	) name7589 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13416_
	);
	LUT2 #(
		.INIT('h1)
	) name7590 (
		_w13411_,
		_w13416_,
		_w13417_
	);
	LUT2 #(
		.INIT('h2)
	) name7591 (
		_w13415_,
		_w13413_,
		_w13418_
	);
	LUT4 #(
		.INIT('h0800)
	) name7592 (
		_w13412_,
		_w13415_,
		_w13413_,
		_w13411_,
		_w13419_
	);
	LUT4 #(
		.INIT('hf6fe)
	) name7593 (
		_w13412_,
		_w13415_,
		_w13413_,
		_w13411_,
		_w13420_
	);
	LUT2 #(
		.INIT('h2)
	) name7594 (
		_w13414_,
		_w13420_,
		_w13421_
	);
	LUT4 #(
		.INIT('h0800)
	) name7595 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13422_
	);
	LUT2 #(
		.INIT('h8)
	) name7596 (
		_w13415_,
		_w13413_,
		_w13423_
	);
	LUT2 #(
		.INIT('h4)
	) name7597 (
		_w13412_,
		_w13411_,
		_w13424_
	);
	LUT3 #(
		.INIT('hae)
	) name7598 (
		_w13412_,
		_w13414_,
		_w13411_,
		_w13425_
	);
	LUT4 #(
		.INIT('h7707)
	) name7599 (
		_w13422_,
		_w13411_,
		_w13423_,
		_w13425_,
		_w13426_
	);
	LUT4 #(
		.INIT('h5455)
	) name7600 (
		_w13410_,
		_w13417_,
		_w13421_,
		_w13426_,
		_w13427_
	);
	LUT3 #(
		.INIT('h02)
	) name7601 (
		_w13412_,
		_w13415_,
		_w13413_,
		_w13428_
	);
	LUT4 #(
		.INIT('hcfc5)
	) name7602 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13429_
	);
	LUT2 #(
		.INIT('h2)
	) name7603 (
		_w13411_,
		_w13429_,
		_w13430_
	);
	LUT4 #(
		.INIT('h0100)
	) name7604 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13431_
	);
	LUT2 #(
		.INIT('h6)
	) name7605 (
		_w13414_,
		_w13413_,
		_w13432_
	);
	LUT2 #(
		.INIT('h8)
	) name7606 (
		_w13414_,
		_w13411_,
		_w13433_
	);
	LUT4 #(
		.INIT('h02c2)
	) name7607 (
		_w13412_,
		_w13414_,
		_w13413_,
		_w13411_,
		_w13434_
	);
	LUT3 #(
		.INIT('h8c)
	) name7608 (
		_w13412_,
		_w13414_,
		_w13411_,
		_w13435_
	);
	LUT4 #(
		.INIT('h0031)
	) name7609 (
		_w13418_,
		_w13434_,
		_w13435_,
		_w13431_,
		_w13436_
	);
	LUT4 #(
		.INIT('h7bdb)
	) name7610 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13437_
	);
	LUT2 #(
		.INIT('h4)
	) name7611 (
		_w13414_,
		_w13411_,
		_w13438_
	);
	LUT3 #(
		.INIT('had)
	) name7612 (
		_w13412_,
		_w13415_,
		_w13413_,
		_w13439_
	);
	LUT4 #(
		.INIT('hfcb8)
	) name7613 (
		_w13414_,
		_w13411_,
		_w13437_,
		_w13439_,
		_w13440_
	);
	LUT4 #(
		.INIT('h7500)
	) name7614 (
		_w13410_,
		_w13430_,
		_w13436_,
		_w13440_,
		_w13441_
	);
	LUT3 #(
		.INIT('h65)
	) name7615 (
		\u2_L1_reg[31]/NET0131 ,
		_w13427_,
		_w13441_,
		_w13442_
	);
	LUT4 #(
		.INIT('hc963)
	) name7616 (
		decrypt_pad,
		\u2_R1_reg[24]/NET0131 ,
		\u2_uk_K_r1_reg[1]/NET0131 ,
		\u2_uk_K_r1_reg[7]/P0001 ,
		_w13443_
	);
	LUT4 #(
		.INIT('hc963)
	) name7617 (
		decrypt_pad,
		\u2_R1_reg[23]/NET0131 ,
		\u2_uk_K_r1_reg[30]/NET0131 ,
		\u2_uk_K_r1_reg[36]/NET0131 ,
		_w13444_
	);
	LUT4 #(
		.INIT('hc693)
	) name7618 (
		decrypt_pad,
		\u2_R1_reg[22]/NET0131 ,
		\u2_uk_K_r1_reg[23]/NET0131 ,
		\u2_uk_K_r1_reg[45]/NET0131 ,
		_w13445_
	);
	LUT4 #(
		.INIT('hc963)
	) name7619 (
		decrypt_pad,
		\u2_R1_reg[20]/NET0131 ,
		\u2_uk_K_r1_reg[35]/NET0131 ,
		\u2_uk_K_r1_reg[45]/NET0131 ,
		_w13446_
	);
	LUT4 #(
		.INIT('hc693)
	) name7620 (
		decrypt_pad,
		\u2_R1_reg[21]/NET0131 ,
		\u2_uk_K_r1_reg[1]/NET0131 ,
		\u2_uk_K_r1_reg[50]/NET0131 ,
		_w13447_
	);
	LUT4 #(
		.INIT('hc693)
	) name7621 (
		decrypt_pad,
		\u2_R1_reg[25]/NET0131 ,
		\u2_uk_K_r1_reg[2]/NET0131 ,
		\u2_uk_K_r1_reg[51]/NET0131 ,
		_w13448_
	);
	LUT4 #(
		.INIT('hf1aa)
	) name7622 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13449_
	);
	LUT2 #(
		.INIT('h2)
	) name7623 (
		_w13444_,
		_w13449_,
		_w13450_
	);
	LUT4 #(
		.INIT('h1040)
	) name7624 (
		_w13444_,
		_w13446_,
		_w13447_,
		_w13445_,
		_w13451_
	);
	LUT2 #(
		.INIT('h2)
	) name7625 (
		_w13446_,
		_w13448_,
		_w13452_
	);
	LUT2 #(
		.INIT('h1)
	) name7626 (
		_w13444_,
		_w13445_,
		_w13453_
	);
	LUT3 #(
		.INIT('hf2)
	) name7627 (
		_w13444_,
		_w13447_,
		_w13445_,
		_w13454_
	);
	LUT4 #(
		.INIT('h0800)
	) name7628 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13455_
	);
	LUT4 #(
		.INIT('h0031)
	) name7629 (
		_w13452_,
		_w13451_,
		_w13454_,
		_w13455_,
		_w13456_
	);
	LUT3 #(
		.INIT('h45)
	) name7630 (
		_w13443_,
		_w13450_,
		_w13456_,
		_w13457_
	);
	LUT4 #(
		.INIT('h0002)
	) name7631 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13458_
	);
	LUT4 #(
		.INIT('h2f7d)
	) name7632 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13459_
	);
	LUT2 #(
		.INIT('h2)
	) name7633 (
		_w13444_,
		_w13459_,
		_w13460_
	);
	LUT4 #(
		.INIT('h00b7)
	) name7634 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13461_
	);
	LUT3 #(
		.INIT('h80)
	) name7635 (
		_w13446_,
		_w13448_,
		_w13445_,
		_w13462_
	);
	LUT4 #(
		.INIT('h4555)
	) name7636 (
		_w13444_,
		_w13446_,
		_w13447_,
		_w13445_,
		_w13463_
	);
	LUT3 #(
		.INIT('h10)
	) name7637 (
		_w13462_,
		_w13461_,
		_w13463_,
		_w13464_
	);
	LUT3 #(
		.INIT('he0)
	) name7638 (
		_w13460_,
		_w13464_,
		_w13443_,
		_w13465_
	);
	LUT3 #(
		.INIT('hde)
	) name7639 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13466_
	);
	LUT2 #(
		.INIT('h2)
	) name7640 (
		_w13453_,
		_w13466_,
		_w13467_
	);
	LUT4 #(
		.INIT('h0004)
	) name7641 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13468_
	);
	LUT4 #(
		.INIT('h0010)
	) name7642 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13469_
	);
	LUT4 #(
		.INIT('h77ef)
	) name7643 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13470_
	);
	LUT3 #(
		.INIT('h75)
	) name7644 (
		_w13444_,
		_w13468_,
		_w13470_,
		_w13471_
	);
	LUT2 #(
		.INIT('h4)
	) name7645 (
		_w13467_,
		_w13471_,
		_w13472_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name7646 (
		\u2_L1_reg[11]/NET0131 ,
		_w13465_,
		_w13457_,
		_w13472_,
		_w13473_
	);
	LUT4 #(
		.INIT('hc963)
	) name7647 (
		decrypt_pad,
		\u2_R1_reg[32]/NET0131 ,
		\u2_uk_K_r1_reg[28]/NET0131 ,
		\u2_uk_K_r1_reg[38]/NET0131 ,
		_w13474_
	);
	LUT4 #(
		.INIT('hc963)
	) name7648 (
		decrypt_pad,
		\u2_R1_reg[31]/P0001 ,
		\u2_uk_K_r1_reg[22]/NET0131 ,
		\u2_uk_K_r1_reg[28]/NET0131 ,
		_w13475_
	);
	LUT4 #(
		.INIT('hc963)
	) name7649 (
		decrypt_pad,
		\u2_R1_reg[28]/NET0131 ,
		\u2_uk_K_r1_reg[37]/NET0131 ,
		\u2_uk_K_r1_reg[43]/NET0131 ,
		_w13476_
	);
	LUT4 #(
		.INIT('hc693)
	) name7650 (
		decrypt_pad,
		\u2_R1_reg[29]/NET0131 ,
		\u2_uk_K_r1_reg[15]/NET0131 ,
		\u2_uk_K_r1_reg[9]/NET0131 ,
		_w13477_
	);
	LUT4 #(
		.INIT('hc693)
	) name7651 (
		decrypt_pad,
		\u2_R1_reg[1]/NET0131 ,
		\u2_uk_K_r1_reg[0]/NET0131 ,
		\u2_uk_K_r1_reg[49]/NET0131 ,
		_w13478_
	);
	LUT4 #(
		.INIT('hc693)
	) name7652 (
		decrypt_pad,
		\u2_R1_reg[30]/NET0131 ,
		\u2_uk_K_r1_reg[16]/NET0131 ,
		\u2_uk_K_r1_reg[38]/NET0131 ,
		_w13479_
	);
	LUT4 #(
		.INIT('h1000)
	) name7653 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13480_
	);
	LUT4 #(
		.INIT('hebfb)
	) name7654 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13481_
	);
	LUT2 #(
		.INIT('h2)
	) name7655 (
		_w13476_,
		_w13479_,
		_w13482_
	);
	LUT2 #(
		.INIT('h4)
	) name7656 (
		_w13476_,
		_w13479_,
		_w13483_
	);
	LUT4 #(
		.INIT('h7407)
	) name7657 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13484_
	);
	LUT3 #(
		.INIT('h08)
	) name7658 (
		_w13477_,
		_w13476_,
		_w13479_,
		_w13485_
	);
	LUT4 #(
		.INIT('h0020)
	) name7659 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13486_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name7660 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13487_
	);
	LUT4 #(
		.INIT('he400)
	) name7661 (
		_w13475_,
		_w13484_,
		_w13481_,
		_w13487_,
		_w13488_
	);
	LUT2 #(
		.INIT('h1)
	) name7662 (
		_w13474_,
		_w13488_,
		_w13489_
	);
	LUT4 #(
		.INIT('hcf45)
	) name7663 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13490_
	);
	LUT4 #(
		.INIT('h22d2)
	) name7664 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13491_
	);
	LUT4 #(
		.INIT('h0001)
	) name7665 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13492_
	);
	LUT4 #(
		.INIT('h0400)
	) name7666 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13493_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name7667 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13494_
	);
	LUT4 #(
		.INIT('h1f00)
	) name7668 (
		_w13474_,
		_w13490_,
		_w13491_,
		_w13494_,
		_w13495_
	);
	LUT4 #(
		.INIT('h0800)
	) name7669 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13496_
	);
	LUT2 #(
		.INIT('h8)
	) name7670 (
		_w13474_,
		_w13496_,
		_w13497_
	);
	LUT4 #(
		.INIT('h2002)
	) name7671 (
		_w13474_,
		_w13477_,
		_w13476_,
		_w13479_,
		_w13498_
	);
	LUT2 #(
		.INIT('h1)
	) name7672 (
		_w13498_,
		_w13486_,
		_w13499_
	);
	LUT4 #(
		.INIT('h5404)
	) name7673 (
		_w13497_,
		_w13499_,
		_w13475_,
		_w13495_,
		_w13500_
	);
	LUT3 #(
		.INIT('h9a)
	) name7674 (
		\u2_L1_reg[5]/NET0131 ,
		_w13489_,
		_w13500_,
		_w13501_
	);
	LUT4 #(
		.INIT('h2006)
	) name7675 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13502_
	);
	LUT4 #(
		.INIT('h134c)
	) name7676 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13503_
	);
	LUT2 #(
		.INIT('h1)
	) name7677 (
		_w13393_,
		_w13503_,
		_w13504_
	);
	LUT3 #(
		.INIT('h47)
	) name7678 (
		_w13383_,
		_w13384_,
		_w13393_,
		_w13505_
	);
	LUT4 #(
		.INIT('h0010)
	) name7679 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13506_
	);
	LUT4 #(
		.INIT('h0301)
	) name7680 (
		_w13387_,
		_w13391_,
		_w13506_,
		_w13505_,
		_w13507_
	);
	LUT3 #(
		.INIT('h10)
	) name7681 (
		_w13504_,
		_w13502_,
		_w13507_,
		_w13508_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name7682 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13509_
	);
	LUT2 #(
		.INIT('h2)
	) name7683 (
		_w13393_,
		_w13509_,
		_w13510_
	);
	LUT3 #(
		.INIT('h04)
	) name7684 (
		_w13389_,
		_w13391_,
		_w13401_,
		_w13511_
	);
	LUT4 #(
		.INIT('h0420)
	) name7685 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13512_
	);
	LUT3 #(
		.INIT('h0d)
	) name7686 (
		_w13388_,
		_w13393_,
		_w13512_,
		_w13513_
	);
	LUT3 #(
		.INIT('h40)
	) name7687 (
		_w13510_,
		_w13511_,
		_w13513_,
		_w13514_
	);
	LUT3 #(
		.INIT('ha9)
	) name7688 (
		\u2_L1_reg[12]/NET0131 ,
		_w13508_,
		_w13514_,
		_w13515_
	);
	LUT4 #(
		.INIT('hcff8)
	) name7689 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13516_
	);
	LUT3 #(
		.INIT('h6f)
	) name7690 (
		_w13414_,
		_w13415_,
		_w13413_,
		_w13517_
	);
	LUT4 #(
		.INIT('hf7df)
	) name7691 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13518_
	);
	LUT4 #(
		.INIT('hd800)
	) name7692 (
		_w13411_,
		_w13517_,
		_w13516_,
		_w13518_,
		_w13519_
	);
	LUT3 #(
		.INIT('hf9)
	) name7693 (
		_w13412_,
		_w13415_,
		_w13413_,
		_w13520_
	);
	LUT2 #(
		.INIT('h2)
	) name7694 (
		_w13433_,
		_w13520_,
		_w13521_
	);
	LUT4 #(
		.INIT('h1000)
	) name7695 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13522_
	);
	LUT4 #(
		.INIT('hef11)
	) name7696 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13523_
	);
	LUT4 #(
		.INIT('h00a1)
	) name7697 (
		_w13412_,
		_w13414_,
		_w13413_,
		_w13411_,
		_w13524_
	);
	LUT4 #(
		.INIT('h0400)
	) name7698 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13525_
	);
	LUT4 #(
		.INIT('h7b7f)
	) name7699 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13526_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7700 (
		_w13411_,
		_w13523_,
		_w13524_,
		_w13526_,
		_w13527_
	);
	LUT4 #(
		.INIT('h3120)
	) name7701 (
		_w13410_,
		_w13521_,
		_w13527_,
		_w13519_,
		_w13528_
	);
	LUT2 #(
		.INIT('h9)
	) name7702 (
		\u2_L1_reg[17]/NET0131 ,
		_w13528_,
		_w13529_
	);
	LUT4 #(
		.INIT('hc693)
	) name7703 (
		decrypt_pad,
		\u2_R1_reg[17]/NET0131 ,
		\u2_uk_K_r1_reg[17]/NET0131 ,
		\u2_uk_K_r1_reg[41]/NET0131 ,
		_w13530_
	);
	LUT4 #(
		.INIT('hc963)
	) name7704 (
		decrypt_pad,
		\u2_R1_reg[12]/NET0131 ,
		\u2_uk_K_r1_reg[25]/NET0131 ,
		\u2_uk_K_r1_reg[33]/NET0131 ,
		_w13531_
	);
	LUT4 #(
		.INIT('hc963)
	) name7705 (
		decrypt_pad,
		\u2_R1_reg[13]/NET0131 ,
		\u2_uk_K_r1_reg[19]/NET0131 ,
		\u2_uk_K_r1_reg[27]/NET0131 ,
		_w13532_
	);
	LUT4 #(
		.INIT('hc693)
	) name7706 (
		decrypt_pad,
		\u2_R1_reg[15]/NET0131 ,
		\u2_uk_K_r1_reg[4]/NET0131 ,
		\u2_uk_K_r1_reg[53]/NET0131 ,
		_w13533_
	);
	LUT4 #(
		.INIT('h7e00)
	) name7707 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13533_,
		_w13534_
	);
	LUT4 #(
		.INIT('hc963)
	) name7708 (
		decrypt_pad,
		\u2_R1_reg[14]/NET0131 ,
		\u2_uk_K_r1_reg[20]/NET0131 ,
		\u2_uk_K_r1_reg[53]/NET0131 ,
		_w13535_
	);
	LUT3 #(
		.INIT('h40)
	) name7709 (
		_w13530_,
		_w13531_,
		_w13535_,
		_w13536_
	);
	LUT3 #(
		.INIT('h0d)
	) name7710 (
		_w13530_,
		_w13532_,
		_w13533_,
		_w13537_
	);
	LUT3 #(
		.INIT('h45)
	) name7711 (
		_w13534_,
		_w13536_,
		_w13537_,
		_w13538_
	);
	LUT3 #(
		.INIT('h01)
	) name7712 (
		_w13530_,
		_w13531_,
		_w13535_,
		_w13539_
	);
	LUT4 #(
		.INIT('heffe)
	) name7713 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13540_
	);
	LUT4 #(
		.INIT('h0008)
	) name7714 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13541_
	);
	LUT4 #(
		.INIT('hc693)
	) name7715 (
		decrypt_pad,
		\u2_R1_reg[16]/NET0131 ,
		\u2_uk_K_r1_reg[12]/NET0131 ,
		\u2_uk_K_r1_reg[4]/NET0131 ,
		_w13542_
	);
	LUT3 #(
		.INIT('h80)
	) name7716 (
		_w13532_,
		_w13535_,
		_w13533_,
		_w13543_
	);
	LUT4 #(
		.INIT('h4000)
	) name7717 (
		_w13531_,
		_w13532_,
		_w13535_,
		_w13533_,
		_w13544_
	);
	LUT4 #(
		.INIT('h0002)
	) name7718 (
		_w13540_,
		_w13542_,
		_w13544_,
		_w13541_,
		_w13545_
	);
	LUT2 #(
		.INIT('h4)
	) name7719 (
		_w13538_,
		_w13545_,
		_w13546_
	);
	LUT4 #(
		.INIT('h8000)
	) name7720 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13547_
	);
	LUT2 #(
		.INIT('h1)
	) name7721 (
		_w13532_,
		_w13533_,
		_w13548_
	);
	LUT4 #(
		.INIT('h0001)
	) name7722 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13533_,
		_w13549_
	);
	LUT2 #(
		.INIT('h4)
	) name7723 (
		_w13532_,
		_w13533_,
		_w13550_
	);
	LUT2 #(
		.INIT('h2)
	) name7724 (
		_w13530_,
		_w13531_,
		_w13551_
	);
	LUT4 #(
		.INIT('h0200)
	) name7725 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13533_,
		_w13552_
	);
	LUT4 #(
		.INIT('h040c)
	) name7726 (
		_w13535_,
		_w13542_,
		_w13552_,
		_w13549_,
		_w13553_
	);
	LUT4 #(
		.INIT('h4000)
	) name7727 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13533_,
		_w13554_
	);
	LUT4 #(
		.INIT('h0020)
	) name7728 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13555_
	);
	LUT2 #(
		.INIT('h1)
	) name7729 (
		_w13554_,
		_w13555_,
		_w13556_
	);
	LUT3 #(
		.INIT('hf9)
	) name7730 (
		_w13531_,
		_w13532_,
		_w13535_,
		_w13557_
	);
	LUT4 #(
		.INIT('h0006)
	) name7731 (
		_w13531_,
		_w13532_,
		_w13535_,
		_w13533_,
		_w13558_
	);
	LUT3 #(
		.INIT('h01)
	) name7732 (
		_w13554_,
		_w13555_,
		_w13558_,
		_w13559_
	);
	LUT3 #(
		.INIT('h40)
	) name7733 (
		_w13547_,
		_w13553_,
		_w13559_,
		_w13560_
	);
	LUT2 #(
		.INIT('h4)
	) name7734 (
		_w13533_,
		_w13555_,
		_w13561_
	);
	LUT3 #(
		.INIT('hbe)
	) name7735 (
		_w13530_,
		_w13531_,
		_w13535_,
		_w13562_
	);
	LUT4 #(
		.INIT('haf23)
	) name7736 (
		_w13535_,
		_w13550_,
		_w13554_,
		_w13562_,
		_w13563_
	);
	LUT2 #(
		.INIT('h4)
	) name7737 (
		_w13561_,
		_w13563_,
		_w13564_
	);
	LUT4 #(
		.INIT('ha955)
	) name7738 (
		\u2_L1_reg[20]/NET0131 ,
		_w13546_,
		_w13560_,
		_w13564_,
		_w13565_
	);
	LUT4 #(
		.INIT('hc693)
	) name7739 (
		decrypt_pad,
		\u2_R1_reg[8]/NET0131 ,
		\u2_uk_K_r1_reg[11]/NET0131 ,
		\u2_uk_K_r1_reg[3]/NET0131 ,
		_w13566_
	);
	LUT4 #(
		.INIT('hc963)
	) name7740 (
		decrypt_pad,
		\u2_R1_reg[7]/NET0131 ,
		\u2_uk_K_r1_reg[12]/NET0131 ,
		\u2_uk_K_r1_reg[20]/NET0131 ,
		_w13567_
	);
	LUT4 #(
		.INIT('hc963)
	) name7741 (
		decrypt_pad,
		\u2_R1_reg[5]/NET0131 ,
		\u2_uk_K_r1_reg[27]/NET0131 ,
		\u2_uk_K_r1_reg[3]/NET0131 ,
		_w13568_
	);
	LUT4 #(
		.INIT('hc963)
	) name7742 (
		decrypt_pad,
		\u2_R1_reg[6]/NET0131 ,
		\u2_uk_K_r1_reg[18]/NET0131 ,
		\u2_uk_K_r1_reg[26]/NET0131 ,
		_w13569_
	);
	LUT4 #(
		.INIT('hc693)
	) name7743 (
		decrypt_pad,
		\u2_R1_reg[4]/NET0131 ,
		\u2_uk_K_r1_reg[24]/NET0131 ,
		\u2_uk_K_r1_reg[48]/NET0131 ,
		_w13570_
	);
	LUT4 #(
		.INIT('hc963)
	) name7744 (
		decrypt_pad,
		\u2_R1_reg[9]/NET0131 ,
		\u2_uk_K_r1_reg[40]/NET0131 ,
		\u2_uk_K_r1_reg[48]/NET0131 ,
		_w13571_
	);
	LUT4 #(
		.INIT('h5fa7)
	) name7745 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13572_
	);
	LUT2 #(
		.INIT('h2)
	) name7746 (
		_w13567_,
		_w13572_,
		_w13573_
	);
	LUT4 #(
		.INIT('hf5fc)
	) name7747 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13574_
	);
	LUT2 #(
		.INIT('h1)
	) name7748 (
		_w13567_,
		_w13574_,
		_w13575_
	);
	LUT2 #(
		.INIT('h4)
	) name7749 (
		_w13569_,
		_w13570_,
		_w13576_
	);
	LUT4 #(
		.INIT('h00bf)
	) name7750 (
		_w13568_,
		_w13570_,
		_w13571_,
		_w13567_,
		_w13577_
	);
	LUT3 #(
		.INIT('h10)
	) name7751 (
		_w13568_,
		_w13570_,
		_w13571_,
		_w13578_
	);
	LUT4 #(
		.INIT('h0400)
	) name7752 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13579_
	);
	LUT3 #(
		.INIT('h0d)
	) name7753 (
		_w13576_,
		_w13577_,
		_w13579_,
		_w13580_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7754 (
		_w13566_,
		_w13575_,
		_w13573_,
		_w13580_,
		_w13581_
	);
	LUT4 #(
		.INIT('hfb7b)
	) name7755 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13582_
	);
	LUT2 #(
		.INIT('h1)
	) name7756 (
		_w13582_,
		_w13567_,
		_w13583_
	);
	LUT2 #(
		.INIT('h8)
	) name7757 (
		_w13567_,
		_w13574_,
		_w13584_
	);
	LUT3 #(
		.INIT('h04)
	) name7758 (
		_w13569_,
		_w13570_,
		_w13571_,
		_w13585_
	);
	LUT3 #(
		.INIT('h07)
	) name7759 (
		_w13568_,
		_w13570_,
		_w13567_,
		_w13586_
	);
	LUT3 #(
		.INIT('h10)
	) name7760 (
		_w13585_,
		_w13578_,
		_w13586_,
		_w13587_
	);
	LUT4 #(
		.INIT('hbf7b)
	) name7761 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13588_
	);
	LUT4 #(
		.INIT('h0155)
	) name7762 (
		_w13566_,
		_w13584_,
		_w13587_,
		_w13588_,
		_w13589_
	);
	LUT4 #(
		.INIT('h5556)
	) name7763 (
		\u2_L1_reg[28]/NET0131 ,
		_w13583_,
		_w13589_,
		_w13581_,
		_w13590_
	);
	LUT4 #(
		.INIT('h6d7c)
	) name7764 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13591_
	);
	LUT4 #(
		.INIT('h00d8)
	) name7765 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13592_
	);
	LUT4 #(
		.INIT('hdf27)
	) name7766 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13593_
	);
	LUT4 #(
		.INIT('h0400)
	) name7767 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13594_
	);
	LUT4 #(
		.INIT('h00e4)
	) name7768 (
		_w13444_,
		_w13593_,
		_w13591_,
		_w13594_,
		_w13595_
	);
	LUT2 #(
		.INIT('h1)
	) name7769 (
		_w13443_,
		_w13595_,
		_w13596_
	);
	LUT4 #(
		.INIT('h9faf)
	) name7770 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13597_
	);
	LUT2 #(
		.INIT('h2)
	) name7771 (
		_w13444_,
		_w13597_,
		_w13598_
	);
	LUT3 #(
		.INIT('h60)
	) name7772 (
		_w13446_,
		_w13448_,
		_w13445_,
		_w13599_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name7773 (
		_w13444_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13600_
	);
	LUT3 #(
		.INIT('h01)
	) name7774 (
		_w13592_,
		_w13600_,
		_w13599_,
		_w13601_
	);
	LUT4 #(
		.INIT('h0080)
	) name7775 (
		_w13444_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13602_
	);
	LUT2 #(
		.INIT('h1)
	) name7776 (
		_w13458_,
		_w13602_,
		_w13603_
	);
	LUT4 #(
		.INIT('h5700)
	) name7777 (
		_w13443_,
		_w13598_,
		_w13601_,
		_w13603_,
		_w13604_
	);
	LUT3 #(
		.INIT('h9a)
	) name7778 (
		\u2_L1_reg[29]/NET0131 ,
		_w13596_,
		_w13604_,
		_w13605_
	);
	LUT4 #(
		.INIT('h7a3f)
	) name7779 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13606_
	);
	LUT2 #(
		.INIT('h1)
	) name7780 (
		_w13567_,
		_w13606_,
		_w13607_
	);
	LUT2 #(
		.INIT('h1)
	) name7781 (
		_w13568_,
		_w13567_,
		_w13608_
	);
	LUT4 #(
		.INIT('h0010)
	) name7782 (
		_w13568_,
		_w13569_,
		_w13571_,
		_w13567_,
		_w13609_
	);
	LUT4 #(
		.INIT('h0800)
	) name7783 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13610_
	);
	LUT2 #(
		.INIT('h1)
	) name7784 (
		_w13609_,
		_w13610_,
		_w13611_
	);
	LUT4 #(
		.INIT('h4000)
	) name7785 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13612_
	);
	LUT4 #(
		.INIT('h0122)
	) name7786 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13613_
	);
	LUT3 #(
		.INIT('h07)
	) name7787 (
		_w13567_,
		_w13612_,
		_w13613_,
		_w13614_
	);
	LUT4 #(
		.INIT('h4555)
	) name7788 (
		_w13566_,
		_w13607_,
		_w13611_,
		_w13614_,
		_w13615_
	);
	LUT4 #(
		.INIT('h9fe2)
	) name7789 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13616_
	);
	LUT4 #(
		.INIT('h0900)
	) name7790 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13617_
	);
	LUT4 #(
		.INIT('h0501)
	) name7791 (
		_w13567_,
		_w13566_,
		_w13617_,
		_w13616_,
		_w13618_
	);
	LUT3 #(
		.INIT('h51)
	) name7792 (
		_w13568_,
		_w13570_,
		_w13571_,
		_w13619_
	);
	LUT4 #(
		.INIT('hb300)
	) name7793 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13566_,
		_w13620_
	);
	LUT3 #(
		.INIT('h04)
	) name7794 (
		_w13568_,
		_w13569_,
		_w13571_,
		_w13621_
	);
	LUT4 #(
		.INIT('h0004)
	) name7795 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13622_
	);
	LUT4 #(
		.INIT('hdf00)
	) name7796 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13567_,
		_w13623_
	);
	LUT4 #(
		.INIT('h0b00)
	) name7797 (
		_w13619_,
		_w13620_,
		_w13622_,
		_w13623_,
		_w13624_
	);
	LUT2 #(
		.INIT('h1)
	) name7798 (
		_w13618_,
		_w13624_,
		_w13625_
	);
	LUT3 #(
		.INIT('h56)
	) name7799 (
		\u2_L1_reg[2]/NET0131 ,
		_w13615_,
		_w13625_,
		_w13626_
	);
	LUT4 #(
		.INIT('hd79b)
	) name7800 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13627_
	);
	LUT4 #(
		.INIT('h0040)
	) name7801 (
		_w13444_,
		_w13446_,
		_w13448_,
		_w13445_,
		_w13628_
	);
	LUT4 #(
		.INIT('h0031)
	) name7802 (
		_w13444_,
		_w13458_,
		_w13627_,
		_w13628_,
		_w13629_
	);
	LUT2 #(
		.INIT('h1)
	) name7803 (
		_w13443_,
		_w13629_,
		_w13630_
	);
	LUT4 #(
		.INIT('hebef)
	) name7804 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13631_
	);
	LUT3 #(
		.INIT('h01)
	) name7805 (
		_w13446_,
		_w13448_,
		_w13445_,
		_w13632_
	);
	LUT4 #(
		.INIT('hff8a)
	) name7806 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13633_
	);
	LUT4 #(
		.INIT('h3210)
	) name7807 (
		_w13443_,
		_w13632_,
		_w13631_,
		_w13633_,
		_w13634_
	);
	LUT4 #(
		.INIT('h0f77)
	) name7808 (
		_w13444_,
		_w13446_,
		_w13447_,
		_w13445_,
		_w13635_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name7809 (
		_w13448_,
		_w13443_,
		_w13469_,
		_w13635_,
		_w13636_
	);
	LUT4 #(
		.INIT('h82a8)
	) name7810 (
		_w13444_,
		_w13446_,
		_w13448_,
		_w13447_,
		_w13637_
	);
	LUT4 #(
		.INIT('h1551)
	) name7811 (
		_w13444_,
		_w13446_,
		_w13448_,
		_w13447_,
		_w13638_
	);
	LUT3 #(
		.INIT('h02)
	) name7812 (
		_w13445_,
		_w13638_,
		_w13637_,
		_w13639_
	);
	LUT4 #(
		.INIT('h000e)
	) name7813 (
		_w13444_,
		_w13634_,
		_w13636_,
		_w13639_,
		_w13640_
	);
	LUT3 #(
		.INIT('h65)
	) name7814 (
		\u2_L1_reg[4]/NET0131 ,
		_w13630_,
		_w13640_,
		_w13641_
	);
	LUT4 #(
		.INIT('hbbdb)
	) name7815 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13642_
	);
	LUT4 #(
		.INIT('h7dff)
	) name7816 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13643_
	);
	LUT4 #(
		.INIT('hefe7)
	) name7817 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13644_
	);
	LUT4 #(
		.INIT('hc480)
	) name7818 (
		_w13533_,
		_w13643_,
		_w13644_,
		_w13642_,
		_w13645_
	);
	LUT2 #(
		.INIT('h2)
	) name7819 (
		_w13542_,
		_w13645_,
		_w13646_
	);
	LUT4 #(
		.INIT('hf3d9)
	) name7820 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13647_
	);
	LUT2 #(
		.INIT('h2)
	) name7821 (
		_w13533_,
		_w13647_,
		_w13648_
	);
	LUT3 #(
		.INIT('h08)
	) name7822 (
		_w13531_,
		_w13532_,
		_w13535_,
		_w13649_
	);
	LUT2 #(
		.INIT('h1)
	) name7823 (
		_w13535_,
		_w13533_,
		_w13650_
	);
	LUT4 #(
		.INIT('h0008)
	) name7824 (
		_w13530_,
		_w13531_,
		_w13535_,
		_w13533_,
		_w13651_
	);
	LUT4 #(
		.INIT('h0002)
	) name7825 (
		_w13540_,
		_w13549_,
		_w13651_,
		_w13649_,
		_w13652_
	);
	LUT3 #(
		.INIT('h45)
	) name7826 (
		_w13542_,
		_w13648_,
		_w13652_,
		_w13653_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name7827 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13654_
	);
	LUT2 #(
		.INIT('h1)
	) name7828 (
		_w13533_,
		_w13654_,
		_w13655_
	);
	LUT3 #(
		.INIT('h23)
	) name7829 (
		_w13535_,
		_w13544_,
		_w13554_,
		_w13656_
	);
	LUT2 #(
		.INIT('h4)
	) name7830 (
		_w13655_,
		_w13656_,
		_w13657_
	);
	LUT4 #(
		.INIT('h5655)
	) name7831 (
		\u2_L1_reg[10]/NET0131 ,
		_w13653_,
		_w13646_,
		_w13657_,
		_w13658_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name7832 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13659_
	);
	LUT4 #(
		.INIT('hfbe5)
	) name7833 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13660_
	);
	LUT4 #(
		.INIT('h0515)
	) name7834 (
		_w13567_,
		_w13566_,
		_w13659_,
		_w13660_,
		_w13661_
	);
	LUT3 #(
		.INIT('h14)
	) name7835 (
		_w13568_,
		_w13570_,
		_w13571_,
		_w13662_
	);
	LUT4 #(
		.INIT('haa8a)
	) name7836 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13663_
	);
	LUT3 #(
		.INIT('h02)
	) name7837 (
		_w13567_,
		_w13663_,
		_w13662_,
		_w13664_
	);
	LUT2 #(
		.INIT('h8)
	) name7838 (
		_w13569_,
		_w13567_,
		_w13665_
	);
	LUT3 #(
		.INIT('hc4)
	) name7839 (
		_w13568_,
		_w13570_,
		_w13571_,
		_w13666_
	);
	LUT2 #(
		.INIT('h8)
	) name7840 (
		_w13665_,
		_w13666_,
		_w13667_
	);
	LUT3 #(
		.INIT('h10)
	) name7841 (
		_w13569_,
		_w13570_,
		_w13571_,
		_w13668_
	);
	LUT3 #(
		.INIT('h45)
	) name7842 (
		_w13566_,
		_w13608_,
		_w13668_,
		_w13669_
	);
	LUT3 #(
		.INIT('h10)
	) name7843 (
		_w13667_,
		_w13664_,
		_w13669_,
		_w13670_
	);
	LUT3 #(
		.INIT('h01)
	) name7844 (
		_w13568_,
		_w13569_,
		_w13571_,
		_w13671_
	);
	LUT4 #(
		.INIT('hdf00)
	) name7845 (
		_w13569_,
		_w13570_,
		_w13571_,
		_w13567_,
		_w13672_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name7846 (
		_w13577_,
		_w13621_,
		_w13671_,
		_w13672_,
		_w13673_
	);
	LUT4 #(
		.INIT('h0002)
	) name7847 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w13674_
	);
	LUT4 #(
		.INIT('h0002)
	) name7848 (
		_w13566_,
		_w13609_,
		_w13610_,
		_w13674_,
		_w13675_
	);
	LUT3 #(
		.INIT('h20)
	) name7849 (
		_w13659_,
		_w13673_,
		_w13675_,
		_w13676_
	);
	LUT4 #(
		.INIT('h999a)
	) name7850 (
		\u2_L1_reg[13]/NET0131 ,
		_w13661_,
		_w13670_,
		_w13676_,
		_w13677_
	);
	LUT4 #(
		.INIT('h02a0)
	) name7851 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13678_
	);
	LUT4 #(
		.INIT('h0100)
	) name7852 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13475_,
		_w13679_
	);
	LUT4 #(
		.INIT('h4000)
	) name7853 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13680_
	);
	LUT4 #(
		.INIT('h0040)
	) name7854 (
		_w13477_,
		_w13478_,
		_w13479_,
		_w13475_,
		_w13681_
	);
	LUT4 #(
		.INIT('h0002)
	) name7855 (
		_w13474_,
		_w13680_,
		_w13679_,
		_w13681_,
		_w13682_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name7856 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13683_
	);
	LUT4 #(
		.INIT('h5b59)
	) name7857 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13684_
	);
	LUT4 #(
		.INIT('h0010)
	) name7858 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13685_
	);
	LUT4 #(
		.INIT('h0501)
	) name7859 (
		_w13474_,
		_w13475_,
		_w13685_,
		_w13684_,
		_w13686_
	);
	LUT3 #(
		.INIT('h0b)
	) name7860 (
		_w13678_,
		_w13682_,
		_w13686_,
		_w13687_
	);
	LUT4 #(
		.INIT('h0009)
	) name7861 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13688_
	);
	LUT4 #(
		.INIT('h3010)
	) name7862 (
		_w13474_,
		_w13477_,
		_w13476_,
		_w13479_,
		_w13689_
	);
	LUT4 #(
		.INIT('h0200)
	) name7863 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13690_
	);
	LUT4 #(
		.INIT('h0001)
	) name7864 (
		_w13475_,
		_w13690_,
		_w13688_,
		_w13689_,
		_w13691_
	);
	LUT4 #(
		.INIT('h0004)
	) name7865 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13692_
	);
	LUT3 #(
		.INIT('h04)
	) name7866 (
		_w13496_,
		_w13475_,
		_w13692_,
		_w13693_
	);
	LUT2 #(
		.INIT('h1)
	) name7867 (
		_w13691_,
		_w13693_,
		_w13694_
	);
	LUT3 #(
		.INIT('h56)
	) name7868 (
		\u2_L1_reg[15]/NET0131 ,
		_w13687_,
		_w13694_,
		_w13695_
	);
	LUT4 #(
		.INIT('hc963)
	) name7869 (
		decrypt_pad,
		\u2_R1_reg[20]/NET0131 ,
		\u2_uk_K_r1_reg[44]/P0001 ,
		\u2_uk_K_r1_reg[50]/NET0131 ,
		_w13696_
	);
	LUT4 #(
		.INIT('hc963)
	) name7870 (
		decrypt_pad,
		\u2_R1_reg[19]/NET0131 ,
		\u2_uk_K_r1_reg[29]/NET0131 ,
		\u2_uk_K_r1_reg[35]/NET0131 ,
		_w13697_
	);
	LUT4 #(
		.INIT('hc963)
	) name7871 (
		decrypt_pad,
		\u2_R1_reg[18]/NET0131 ,
		\u2_uk_K_r1_reg[42]/NET0131 ,
		\u2_uk_K_r1_reg[52]/NET0131 ,
		_w13698_
	);
	LUT4 #(
		.INIT('hc693)
	) name7872 (
		decrypt_pad,
		\u2_R1_reg[17]/NET0131 ,
		\u2_uk_K_r1_reg[30]/NET0131 ,
		\u2_uk_K_r1_reg[52]/NET0131 ,
		_w13699_
	);
	LUT4 #(
		.INIT('hc963)
	) name7873 (
		decrypt_pad,
		\u2_R1_reg[21]/NET0131 ,
		\u2_uk_K_r1_reg[14]/NET0131 ,
		\u2_uk_K_r1_reg[51]/NET0131 ,
		_w13700_
	);
	LUT4 #(
		.INIT('hc963)
	) name7874 (
		decrypt_pad,
		\u2_R1_reg[16]/NET0131 ,
		\u2_uk_K_r1_reg[2]/NET0131 ,
		\u2_uk_K_r1_reg[8]/NET0131 ,
		_w13701_
	);
	LUT3 #(
		.INIT('h80)
	) name7875 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13702_
	);
	LUT4 #(
		.INIT('h0080)
	) name7876 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13703_
	);
	LUT3 #(
		.INIT('h40)
	) name7877 (
		_w13700_,
		_w13699_,
		_w13698_,
		_w13704_
	);
	LUT4 #(
		.INIT('h0004)
	) name7878 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13705_
	);
	LUT4 #(
		.INIT('had79)
	) name7879 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13706_
	);
	LUT2 #(
		.INIT('h1)
	) name7880 (
		_w13697_,
		_w13706_,
		_w13707_
	);
	LUT4 #(
		.INIT('h228a)
	) name7881 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13708_
	);
	LUT3 #(
		.INIT('hb0)
	) name7882 (
		_w13700_,
		_w13701_,
		_w13697_,
		_w13709_
	);
	LUT4 #(
		.INIT('h0800)
	) name7883 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13710_
	);
	LUT4 #(
		.INIT('hf7ef)
	) name7884 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13711_
	);
	LUT4 #(
		.INIT('hef00)
	) name7885 (
		_w13708_,
		_w13704_,
		_w13709_,
		_w13711_,
		_w13712_
	);
	LUT3 #(
		.INIT('h45)
	) name7886 (
		_w13696_,
		_w13707_,
		_w13712_,
		_w13713_
	);
	LUT4 #(
		.INIT('h9d35)
	) name7887 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13714_
	);
	LUT2 #(
		.INIT('h4)
	) name7888 (
		_w13714_,
		_w13697_,
		_w13715_
	);
	LUT4 #(
		.INIT('h0020)
	) name7889 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13697_,
		_w13716_
	);
	LUT4 #(
		.INIT('hffde)
	) name7890 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13697_,
		_w13717_
	);
	LUT2 #(
		.INIT('h1)
	) name7891 (
		_w13698_,
		_w13717_,
		_w13718_
	);
	LUT3 #(
		.INIT('hc4)
	) name7892 (
		_w13699_,
		_w13698_,
		_w13697_,
		_w13719_
	);
	LUT4 #(
		.INIT('h8808)
	) name7893 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13720_
	);
	LUT4 #(
		.INIT('h0440)
	) name7894 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13721_
	);
	LUT3 #(
		.INIT('h0b)
	) name7895 (
		_w13719_,
		_w13720_,
		_w13721_,
		_w13722_
	);
	LUT4 #(
		.INIT('hef00)
	) name7896 (
		_w13715_,
		_w13718_,
		_w13722_,
		_w13696_,
		_w13723_
	);
	LUT4 #(
		.INIT('h0040)
	) name7897 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13724_
	);
	LUT4 #(
		.INIT('hfebf)
	) name7898 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13725_
	);
	LUT4 #(
		.INIT('h0200)
	) name7899 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13726_
	);
	LUT4 #(
		.INIT('hedff)
	) name7900 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13727_
	);
	LUT3 #(
		.INIT('hd8)
	) name7901 (
		_w13697_,
		_w13725_,
		_w13727_,
		_w13728_
	);
	LUT4 #(
		.INIT('h5655)
	) name7902 (
		\u2_L1_reg[14]/NET0131 ,
		_w13723_,
		_w13713_,
		_w13728_,
		_w13729_
	);
	LUT3 #(
		.INIT('h04)
	) name7903 (
		_w13444_,
		_w13446_,
		_w13447_,
		_w13730_
	);
	LUT4 #(
		.INIT('hfb00)
	) name7904 (
		_w13448_,
		_w13447_,
		_w13445_,
		_w13443_,
		_w13731_
	);
	LUT3 #(
		.INIT('h10)
	) name7905 (
		_w13468_,
		_w13730_,
		_w13731_,
		_w13732_
	);
	LUT4 #(
		.INIT('hfb5b)
	) name7906 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13733_
	);
	LUT4 #(
		.INIT('h4100)
	) name7907 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13734_
	);
	LUT3 #(
		.INIT('h0d)
	) name7908 (
		_w13444_,
		_w13733_,
		_w13734_,
		_w13735_
	);
	LUT4 #(
		.INIT('h45e5)
	) name7909 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13736_
	);
	LUT2 #(
		.INIT('h2)
	) name7910 (
		_w13444_,
		_w13736_,
		_w13737_
	);
	LUT4 #(
		.INIT('h1001)
	) name7911 (
		_w13444_,
		_w13446_,
		_w13448_,
		_w13447_,
		_w13738_
	);
	LUT4 #(
		.INIT('h8000)
	) name7912 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13445_,
		_w13739_
	);
	LUT3 #(
		.INIT('h01)
	) name7913 (
		_w13443_,
		_w13739_,
		_w13738_,
		_w13740_
	);
	LUT4 #(
		.INIT('h7077)
	) name7914 (
		_w13732_,
		_w13735_,
		_w13737_,
		_w13740_,
		_w13741_
	);
	LUT3 #(
		.INIT('hd7)
	) name7915 (
		_w13446_,
		_w13448_,
		_w13447_,
		_w13742_
	);
	LUT4 #(
		.INIT('h5f4e)
	) name7916 (
		_w13444_,
		_w13445_,
		_w13468_,
		_w13742_,
		_w13743_
	);
	LUT3 #(
		.INIT('h65)
	) name7917 (
		\u2_L1_reg[19]/NET0131 ,
		_w13741_,
		_w13743_,
		_w13744_
	);
	LUT4 #(
		.INIT('h00fb)
	) name7918 (
		_w13478_,
		_w13476_,
		_w13479_,
		_w13475_,
		_w13745_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7919 (
		_w13477_,
		_w13476_,
		_w13479_,
		_w13475_,
		_w13746_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name7920 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13747_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7921 (
		_w13680_,
		_w13745_,
		_w13746_,
		_w13747_,
		_w13748_
	);
	LUT4 #(
		.INIT('h2100)
	) name7922 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13749_
	);
	LUT3 #(
		.INIT('h02)
	) name7923 (
		_w13474_,
		_w13692_,
		_w13749_,
		_w13750_
	);
	LUT2 #(
		.INIT('h4)
	) name7924 (
		_w13748_,
		_w13750_,
		_w13751_
	);
	LUT2 #(
		.INIT('h2)
	) name7925 (
		_w13478_,
		_w13475_,
		_w13752_
	);
	LUT3 #(
		.INIT('h73)
	) name7926 (
		_w13477_,
		_w13478_,
		_w13475_,
		_w13753_
	);
	LUT2 #(
		.INIT('h2)
	) name7927 (
		_w13482_,
		_w13753_,
		_w13754_
	);
	LUT3 #(
		.INIT('h51)
	) name7928 (
		_w13477_,
		_w13478_,
		_w13475_,
		_w13755_
	);
	LUT3 #(
		.INIT('h31)
	) name7929 (
		_w13483_,
		_w13480_,
		_w13755_,
		_w13756_
	);
	LUT4 #(
		.INIT('h8fdf)
	) name7930 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13757_
	);
	LUT2 #(
		.INIT('h2)
	) name7931 (
		_w13475_,
		_w13757_,
		_w13758_
	);
	LUT4 #(
		.INIT('h0002)
	) name7932 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13475_,
		_w13759_
	);
	LUT3 #(
		.INIT('h01)
	) name7933 (
		_w13474_,
		_w13492_,
		_w13759_,
		_w13760_
	);
	LUT4 #(
		.INIT('h1000)
	) name7934 (
		_w13758_,
		_w13754_,
		_w13760_,
		_w13756_,
		_w13761_
	);
	LUT4 #(
		.INIT('h0100)
	) name7935 (
		_w13477_,
		_w13476_,
		_w13479_,
		_w13475_,
		_w13762_
	);
	LUT3 #(
		.INIT('h13)
	) name7936 (
		_w13485_,
		_w13762_,
		_w13752_,
		_w13763_
	);
	LUT4 #(
		.INIT('ha955)
	) name7937 (
		\u2_L1_reg[21]/NET0131 ,
		_w13751_,
		_w13761_,
		_w13763_,
		_w13764_
	);
	LUT4 #(
		.INIT('h5545)
	) name7938 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13765_
	);
	LUT4 #(
		.INIT('h004c)
	) name7939 (
		_w13531_,
		_w13532_,
		_w13535_,
		_w13533_,
		_w13766_
	);
	LUT2 #(
		.INIT('h4)
	) name7940 (
		_w13765_,
		_w13766_,
		_w13767_
	);
	LUT3 #(
		.INIT('h51)
	) name7941 (
		_w13530_,
		_w13531_,
		_w13535_,
		_w13768_
	);
	LUT4 #(
		.INIT('h4000)
	) name7942 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13769_
	);
	LUT4 #(
		.INIT('hbcff)
	) name7943 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13770_
	);
	LUT3 #(
		.INIT('hd0)
	) name7944 (
		_w13550_,
		_w13768_,
		_w13770_,
		_w13771_
	);
	LUT3 #(
		.INIT('h8a)
	) name7945 (
		_w13542_,
		_w13767_,
		_w13771_,
		_w13772_
	);
	LUT4 #(
		.INIT('h084c)
	) name7946 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13773_
	);
	LUT4 #(
		.INIT('h0400)
	) name7947 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13774_
	);
	LUT4 #(
		.INIT('hfcb8)
	) name7948 (
		_w13539_,
		_w13533_,
		_w13773_,
		_w13774_,
		_w13775_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name7949 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13776_
	);
	LUT3 #(
		.INIT('h45)
	) name7950 (
		_w13542_,
		_w13775_,
		_w13776_,
		_w13777_
	);
	LUT4 #(
		.INIT('h6dff)
	) name7951 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13778_
	);
	LUT2 #(
		.INIT('h2)
	) name7952 (
		_w13533_,
		_w13778_,
		_w13779_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name7953 (
		_w13535_,
		_w13533_,
		_w13549_,
		_w13769_,
		_w13780_
	);
	LUT2 #(
		.INIT('h4)
	) name7954 (
		_w13779_,
		_w13780_,
		_w13781_
	);
	LUT4 #(
		.INIT('h5655)
	) name7955 (
		\u2_L1_reg[1]/NET0131 ,
		_w13777_,
		_w13772_,
		_w13781_,
		_w13782_
	);
	LUT4 #(
		.INIT('hf9ff)
	) name7956 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13783_
	);
	LUT3 #(
		.INIT('hf9)
	) name7957 (
		_w13414_,
		_w13415_,
		_w13413_,
		_w13784_
	);
	LUT4 #(
		.INIT('h0010)
	) name7958 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13785_
	);
	LUT4 #(
		.INIT('h0400)
	) name7959 (
		_w13411_,
		_w13784_,
		_w13785_,
		_w13783_,
		_w13786_
	);
	LUT4 #(
		.INIT('hf700)
	) name7960 (
		_w13414_,
		_w13415_,
		_w13413_,
		_w13411_,
		_w13787_
	);
	LUT2 #(
		.INIT('h4)
	) name7961 (
		_w13422_,
		_w13787_,
		_w13788_
	);
	LUT4 #(
		.INIT('h002a)
	) name7962 (
		_w13410_,
		_w13438_,
		_w13428_,
		_w13522_,
		_w13789_
	);
	LUT3 #(
		.INIT('he0)
	) name7963 (
		_w13786_,
		_w13788_,
		_w13789_,
		_w13790_
	);
	LUT4 #(
		.INIT('hfd00)
	) name7964 (
		_w13414_,
		_w13415_,
		_w13413_,
		_w13411_,
		_w13791_
	);
	LUT4 #(
		.INIT('h13ff)
	) name7965 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13792_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name7966 (
		_w13411_,
		_w13785_,
		_w13791_,
		_w13792_,
		_w13793_
	);
	LUT3 #(
		.INIT('h7e)
	) name7967 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13794_
	);
	LUT3 #(
		.INIT('h10)
	) name7968 (
		_w13410_,
		_w13419_,
		_w13794_,
		_w13795_
	);
	LUT2 #(
		.INIT('h4)
	) name7969 (
		_w13793_,
		_w13795_,
		_w13796_
	);
	LUT4 #(
		.INIT('h5100)
	) name7970 (
		_w13412_,
		_w13415_,
		_w13413_,
		_w13411_,
		_w13797_
	);
	LUT3 #(
		.INIT('h08)
	) name7971 (
		_w13412_,
		_w13414_,
		_w13411_,
		_w13798_
	);
	LUT4 #(
		.INIT('h153f)
	) name7972 (
		_w13423_,
		_w13432_,
		_w13797_,
		_w13798_,
		_w13799_
	);
	LUT4 #(
		.INIT('h56aa)
	) name7973 (
		\u2_L1_reg[23]/NET0131 ,
		_w13790_,
		_w13796_,
		_w13799_,
		_w13800_
	);
	LUT4 #(
		.INIT('h6c78)
	) name7974 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13801_
	);
	LUT4 #(
		.INIT('hf7c7)
	) name7975 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13802_
	);
	LUT4 #(
		.INIT('hbf5f)
	) name7976 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13803_
	);
	LUT4 #(
		.INIT('hd800)
	) name7977 (
		_w13697_,
		_w13801_,
		_w13802_,
		_w13803_,
		_w13804_
	);
	LUT2 #(
		.INIT('h2)
	) name7978 (
		_w13696_,
		_w13804_,
		_w13805_
	);
	LUT4 #(
		.INIT('hbefd)
	) name7979 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13806_
	);
	LUT2 #(
		.INIT('h2)
	) name7980 (
		_w13697_,
		_w13806_,
		_w13807_
	);
	LUT4 #(
		.INIT('hf351)
	) name7981 (
		_w13701_,
		_w13699_,
		_w13698_,
		_w13697_,
		_w13808_
	);
	LUT3 #(
		.INIT('h51)
	) name7982 (
		_w13700_,
		_w13699_,
		_w13697_,
		_w13809_
	);
	LUT3 #(
		.INIT('h70)
	) name7983 (
		_w13700_,
		_w13698_,
		_w13697_,
		_w13810_
	);
	LUT3 #(
		.INIT('h41)
	) name7984 (
		_w13701_,
		_w13699_,
		_w13698_,
		_w13811_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name7985 (
		_w13808_,
		_w13809_,
		_w13810_,
		_w13811_,
		_w13812_
	);
	LUT4 #(
		.INIT('h0020)
	) name7986 (
		_w13701_,
		_w13699_,
		_w13698_,
		_w13697_,
		_w13813_
	);
	LUT2 #(
		.INIT('h1)
	) name7987 (
		_w13703_,
		_w13813_,
		_w13814_
	);
	LUT4 #(
		.INIT('h0e00)
	) name7988 (
		_w13696_,
		_w13812_,
		_w13807_,
		_w13814_,
		_w13815_
	);
	LUT3 #(
		.INIT('h65)
	) name7989 (
		\u2_L1_reg[25]/NET0131 ,
		_w13805_,
		_w13815_,
		_w13816_
	);
	LUT4 #(
		.INIT('h9cee)
	) name7990 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13817_
	);
	LUT2 #(
		.INIT('h1)
	) name7991 (
		_w13548_,
		_w13817_,
		_w13818_
	);
	LUT4 #(
		.INIT('h7775)
	) name7992 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13819_
	);
	LUT3 #(
		.INIT('h0d)
	) name7993 (
		_w13531_,
		_w13535_,
		_w13533_,
		_w13820_
	);
	LUT3 #(
		.INIT('h8a)
	) name7994 (
		_w13542_,
		_w13819_,
		_w13820_,
		_w13821_
	);
	LUT2 #(
		.INIT('h4)
	) name7995 (
		_w13818_,
		_w13821_,
		_w13822_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name7996 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13535_,
		_w13823_
	);
	LUT2 #(
		.INIT('h1)
	) name7997 (
		_w13533_,
		_w13823_,
		_w13824_
	);
	LUT4 #(
		.INIT('h00fd)
	) name7998 (
		_w13531_,
		_w13532_,
		_w13535_,
		_w13542_,
		_w13825_
	);
	LUT3 #(
		.INIT('hd0)
	) name7999 (
		_w13543_,
		_w13551_,
		_w13825_,
		_w13826_
	);
	LUT3 #(
		.INIT('h20)
	) name8000 (
		_w13556_,
		_w13824_,
		_w13826_,
		_w13827_
	);
	LUT3 #(
		.INIT('h6b)
	) name8001 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13828_
	);
	LUT2 #(
		.INIT('h8)
	) name8002 (
		_w13530_,
		_w13533_,
		_w13829_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name8003 (
		_w13557_,
		_w13650_,
		_w13828_,
		_w13829_,
		_w13830_
	);
	LUT4 #(
		.INIT('ha955)
	) name8004 (
		\u2_L1_reg[26]/NET0131 ,
		_w13822_,
		_w13827_,
		_w13830_,
		_w13831_
	);
	LUT4 #(
		.INIT('hd7d2)
	) name8005 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13832_
	);
	LUT2 #(
		.INIT('h1)
	) name8006 (
		_w13475_,
		_w13832_,
		_w13833_
	);
	LUT3 #(
		.INIT('hb0)
	) name8007 (
		_w13478_,
		_w13476_,
		_w13475_,
		_w13834_
	);
	LUT4 #(
		.INIT('he7bb)
	) name8008 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13835_
	);
	LUT3 #(
		.INIT('hb0)
	) name8009 (
		_w13683_,
		_w13834_,
		_w13835_,
		_w13836_
	);
	LUT3 #(
		.INIT('h8a)
	) name8010 (
		_w13474_,
		_w13833_,
		_w13836_,
		_w13837_
	);
	LUT4 #(
		.INIT('hce44)
	) name8011 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13838_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8012 (
		_w13477_,
		_w13478_,
		_w13479_,
		_w13475_,
		_w13839_
	);
	LUT2 #(
		.INIT('h4)
	) name8013 (
		_w13838_,
		_w13839_,
		_w13840_
	);
	LUT4 #(
		.INIT('h0080)
	) name8014 (
		_w13478_,
		_w13476_,
		_w13479_,
		_w13475_,
		_w13841_
	);
	LUT3 #(
		.INIT('h01)
	) name8015 (
		_w13493_,
		_w13759_,
		_w13841_,
		_w13842_
	);
	LUT4 #(
		.INIT('h1000)
	) name8016 (
		_w13477_,
		_w13478_,
		_w13479_,
		_w13475_,
		_w13843_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name8017 (
		_w13477_,
		_w13478_,
		_w13476_,
		_w13479_,
		_w13844_
	);
	LUT3 #(
		.INIT('h32)
	) name8018 (
		_w13475_,
		_w13843_,
		_w13844_,
		_w13845_
	);
	LUT4 #(
		.INIT('hba00)
	) name8019 (
		_w13474_,
		_w13840_,
		_w13842_,
		_w13845_,
		_w13846_
	);
	LUT3 #(
		.INIT('h65)
	) name8020 (
		\u2_L1_reg[27]/NET0131 ,
		_w13837_,
		_w13846_,
		_w13847_
	);
	LUT3 #(
		.INIT('h40)
	) name8021 (
		_w13384_,
		_w13385_,
		_w13386_,
		_w13848_
	);
	LUT4 #(
		.INIT('hdee3)
	) name8022 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13849_
	);
	LUT2 #(
		.INIT('h1)
	) name8023 (
		_w13393_,
		_w13849_,
		_w13850_
	);
	LUT3 #(
		.INIT('h08)
	) name8024 (
		_w13383_,
		_w13385_,
		_w13386_,
		_w13851_
	);
	LUT4 #(
		.INIT('hbbfc)
	) name8025 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13852_
	);
	LUT4 #(
		.INIT('h1f13)
	) name8026 (
		_w13384_,
		_w13393_,
		_w13851_,
		_w13852_,
		_w13853_
	);
	LUT3 #(
		.INIT('h8a)
	) name8027 (
		_w13391_,
		_w13850_,
		_w13853_,
		_w13854_
	);
	LUT3 #(
		.INIT('h04)
	) name8028 (
		_w13383_,
		_w13385_,
		_w13386_,
		_w13855_
	);
	LUT2 #(
		.INIT('h6)
	) name8029 (
		_w13384_,
		_w13386_,
		_w13856_
	);
	LUT4 #(
		.INIT('hab89)
	) name8030 (
		_w13393_,
		_w13855_,
		_w13856_,
		_w13848_,
		_w13857_
	);
	LUT4 #(
		.INIT('h7db7)
	) name8031 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13858_
	);
	LUT4 #(
		.INIT('h00a2)
	) name8032 (
		_w13384_,
		_w13385_,
		_w13386_,
		_w13393_,
		_w13859_
	);
	LUT4 #(
		.INIT('h0777)
	) name8033 (
		_w13388_,
		_w13393_,
		_w13397_,
		_w13859_,
		_w13860_
	);
	LUT4 #(
		.INIT('hba00)
	) name8034 (
		_w13391_,
		_w13857_,
		_w13858_,
		_w13860_,
		_w13861_
	);
	LUT3 #(
		.INIT('h65)
	) name8035 (
		\u2_L1_reg[32]/NET0131 ,
		_w13854_,
		_w13861_,
		_w13862_
	);
	LUT4 #(
		.INIT('hc963)
	) name8036 (
		decrypt_pad,
		\u2_R1_reg[12]/NET0131 ,
		\u2_uk_K_r1_reg[13]/NET0131 ,
		\u2_uk_K_r1_reg[46]/NET0131 ,
		_w13863_
	);
	LUT4 #(
		.INIT('hc963)
	) name8037 (
		decrypt_pad,
		\u2_R1_reg[13]/NET0131 ,
		\u2_uk_K_r1_reg[26]/NET0131 ,
		\u2_uk_K_r1_reg[34]/NET0131 ,
		_w13864_
	);
	LUT4 #(
		.INIT('hc963)
	) name8038 (
		decrypt_pad,
		\u2_R1_reg[8]/NET0131 ,
		\u2_uk_K_r1_reg[17]/NET0131 ,
		\u2_uk_K_r1_reg[25]/NET0131 ,
		_w13865_
	);
	LUT2 #(
		.INIT('h6)
	) name8039 (
		_w13864_,
		_w13865_,
		_w13866_
	);
	LUT4 #(
		.INIT('hc963)
	) name8040 (
		decrypt_pad,
		\u2_R1_reg[9]/NET0131 ,
		\u2_uk_K_r1_reg[46]/NET0131 ,
		\u2_uk_K_r1_reg[54]/NET0131 ,
		_w13867_
	);
	LUT4 #(
		.INIT('hc963)
	) name8041 (
		decrypt_pad,
		\u2_R1_reg[10]/NET0131 ,
		\u2_uk_K_r1_reg[54]/NET0131 ,
		\u2_uk_K_r1_reg[5]/NET0131 ,
		_w13868_
	);
	LUT4 #(
		.INIT('h2100)
	) name8042 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13869_
	);
	LUT3 #(
		.INIT('h08)
	) name8043 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13870_
	);
	LUT4 #(
		.INIT('hc963)
	) name8044 (
		decrypt_pad,
		\u2_R1_reg[11]/P0001 ,
		\u2_uk_K_r1_reg[55]/NET0131 ,
		\u2_uk_K_r1_reg[6]/NET0131 ,
		_w13871_
	);
	LUT2 #(
		.INIT('h2)
	) name8045 (
		_w13868_,
		_w13871_,
		_w13872_
	);
	LUT3 #(
		.INIT('h40)
	) name8046 (
		_w13864_,
		_w13867_,
		_w13868_,
		_w13873_
	);
	LUT4 #(
		.INIT('h4000)
	) name8047 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13874_
	);
	LUT4 #(
		.INIT('h0007)
	) name8048 (
		_w13870_,
		_w13872_,
		_w13874_,
		_w13869_,
		_w13875_
	);
	LUT2 #(
		.INIT('h8)
	) name8049 (
		_w13864_,
		_w13871_,
		_w13876_
	);
	LUT3 #(
		.INIT('h46)
	) name8050 (
		_w13864_,
		_w13865_,
		_w13871_,
		_w13877_
	);
	LUT2 #(
		.INIT('h1)
	) name8051 (
		_w13867_,
		_w13868_,
		_w13878_
	);
	LUT2 #(
		.INIT('h8)
	) name8052 (
		_w13878_,
		_w13877_,
		_w13879_
	);
	LUT3 #(
		.INIT('hed)
	) name8053 (
		_w13867_,
		_w13868_,
		_w13877_,
		_w13880_
	);
	LUT3 #(
		.INIT('h15)
	) name8054 (
		_w13863_,
		_w13875_,
		_w13880_,
		_w13881_
	);
	LUT4 #(
		.INIT('h959d)
	) name8055 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13882_
	);
	LUT4 #(
		.INIT('h0001)
	) name8056 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13883_
	);
	LUT4 #(
		.INIT('hddfe)
	) name8057 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13884_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8058 (
		_w13882_,
		_w13863_,
		_w13884_,
		_w13871_,
		_w13885_
	);
	LUT2 #(
		.INIT('h8)
	) name8059 (
		_w13868_,
		_w13863_,
		_w13886_
	);
	LUT3 #(
		.INIT('h04)
	) name8060 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13887_
	);
	LUT2 #(
		.INIT('h2)
	) name8061 (
		_w13863_,
		_w13871_,
		_w13888_
	);
	LUT3 #(
		.INIT('h80)
	) name8062 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13889_
	);
	LUT4 #(
		.INIT('h6f67)
	) name8063 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13890_
	);
	LUT4 #(
		.INIT('h7707)
	) name8064 (
		_w13886_,
		_w13887_,
		_w13888_,
		_w13890_,
		_w13891_
	);
	LUT2 #(
		.INIT('h4)
	) name8065 (
		_w13885_,
		_w13891_,
		_w13892_
	);
	LUT3 #(
		.INIT('h65)
	) name8066 (
		\u2_L1_reg[6]/NET0131 ,
		_w13881_,
		_w13892_,
		_w13893_
	);
	LUT3 #(
		.INIT('h28)
	) name8067 (
		_w13384_,
		_w13385_,
		_w13386_,
		_w13894_
	);
	LUT4 #(
		.INIT('h2880)
	) name8068 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13895_
	);
	LUT4 #(
		.INIT('h5004)
	) name8069 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13896_
	);
	LUT2 #(
		.INIT('h2)
	) name8070 (
		_w13393_,
		_w13896_,
		_w13897_
	);
	LUT3 #(
		.INIT('h09)
	) name8071 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13898_
	);
	LUT4 #(
		.INIT('h00f7)
	) name8072 (
		_w13383_,
		_w13385_,
		_w13386_,
		_w13393_,
		_w13899_
	);
	LUT3 #(
		.INIT('h10)
	) name8073 (
		_w13894_,
		_w13898_,
		_w13899_,
		_w13900_
	);
	LUT4 #(
		.INIT('h888a)
	) name8074 (
		_w13391_,
		_w13895_,
		_w13897_,
		_w13900_,
		_w13901_
	);
	LUT4 #(
		.INIT('h5150)
	) name8075 (
		_w13391_,
		_w13393_,
		_w13398_,
		_w13896_,
		_w13902_
	);
	LUT4 #(
		.INIT('h7885)
	) name8076 (
		_w13383_,
		_w13384_,
		_w13385_,
		_w13386_,
		_w13903_
	);
	LUT4 #(
		.INIT('h00c4)
	) name8077 (
		_w13391_,
		_w13393_,
		_w13398_,
		_w13903_,
		_w13904_
	);
	LUT2 #(
		.INIT('h4)
	) name8078 (
		_w13393_,
		_w13895_,
		_w13905_
	);
	LUT3 #(
		.INIT('h01)
	) name8079 (
		_w13904_,
		_w13905_,
		_w13902_,
		_w13906_
	);
	LUT3 #(
		.INIT('h65)
	) name8080 (
		\u2_L1_reg[7]/NET0131 ,
		_w13901_,
		_w13906_,
		_w13907_
	);
	LUT3 #(
		.INIT('h02)
	) name8081 (
		_w13697_,
		_w13702_,
		_w13705_,
		_w13908_
	);
	LUT4 #(
		.INIT('h2022)
	) name8082 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13909_
	);
	LUT4 #(
		.INIT('h00f7)
	) name8083 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13697_,
		_w13910_
	);
	LUT2 #(
		.INIT('h4)
	) name8084 (
		_w13909_,
		_w13910_,
		_w13911_
	);
	LUT4 #(
		.INIT('hbecf)
	) name8085 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13912_
	);
	LUT4 #(
		.INIT('h0155)
	) name8086 (
		_w13696_,
		_w13908_,
		_w13911_,
		_w13912_,
		_w13913_
	);
	LUT4 #(
		.INIT('h0001)
	) name8087 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13914_
	);
	LUT4 #(
		.INIT('hf7f6)
	) name8088 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13915_
	);
	LUT3 #(
		.INIT('h02)
	) name8089 (
		_w13701_,
		_w13698_,
		_w13697_,
		_w13916_
	);
	LUT4 #(
		.INIT('h00c4)
	) name8090 (
		_w13697_,
		_w13727_,
		_w13915_,
		_w13916_,
		_w13917_
	);
	LUT4 #(
		.INIT('haddf)
	) name8091 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13918_
	);
	LUT4 #(
		.INIT('haf23)
	) name8092 (
		_w13700_,
		_w13697_,
		_w13813_,
		_w13918_,
		_w13919_
	);
	LUT3 #(
		.INIT('hd0)
	) name8093 (
		_w13696_,
		_w13917_,
		_w13919_,
		_w13920_
	);
	LUT3 #(
		.INIT('h65)
	) name8094 (
		\u2_L1_reg[8]/NET0131 ,
		_w13913_,
		_w13920_,
		_w13921_
	);
	LUT4 #(
		.INIT('hf700)
	) name8095 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13922_
	);
	LUT4 #(
		.INIT('h0400)
	) name8096 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13871_,
		_w13923_
	);
	LUT4 #(
		.INIT('h006d)
	) name8097 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13924_
	);
	LUT3 #(
		.INIT('h45)
	) name8098 (
		_w13922_,
		_w13923_,
		_w13924_,
		_w13925_
	);
	LUT4 #(
		.INIT('h0100)
	) name8099 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13926_
	);
	LUT3 #(
		.INIT('h14)
	) name8100 (
		_w13864_,
		_w13865_,
		_w13868_,
		_w13927_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8101 (
		_w13871_,
		_w13874_,
		_w13926_,
		_w13927_,
		_w13928_
	);
	LUT3 #(
		.INIT('ha8)
	) name8102 (
		_w13863_,
		_w13925_,
		_w13928_,
		_w13929_
	);
	LUT3 #(
		.INIT('h40)
	) name8103 (
		_w13867_,
		_w13865_,
		_w13868_,
		_w13930_
	);
	LUT4 #(
		.INIT('h00bf)
	) name8104 (
		_w13867_,
		_w13865_,
		_w13868_,
		_w13871_,
		_w13931_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8105 (
		_w13871_,
		_w13874_,
		_w13926_,
		_w13931_,
		_w13932_
	);
	LUT4 #(
		.INIT('h7d78)
	) name8106 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13933_
	);
	LUT3 #(
		.INIT('he0)
	) name8107 (
		_w13864_,
		_w13865_,
		_w13871_,
		_w13934_
	);
	LUT4 #(
		.INIT('h6800)
	) name8108 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13871_,
		_w13935_
	);
	LUT4 #(
		.INIT('h0504)
	) name8109 (
		_w13883_,
		_w13871_,
		_w13935_,
		_w13933_,
		_w13936_
	);
	LUT3 #(
		.INIT('h32)
	) name8110 (
		_w13863_,
		_w13932_,
		_w13936_,
		_w13937_
	);
	LUT3 #(
		.INIT('h65)
	) name8111 (
		\u2_L1_reg[16]/NET0131 ,
		_w13929_,
		_w13937_,
		_w13938_
	);
	LUT2 #(
		.INIT('h4)
	) name8112 (
		_w13868_,
		_w13871_,
		_w13939_
	);
	LUT3 #(
		.INIT('h31)
	) name8113 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13940_
	);
	LUT2 #(
		.INIT('h8)
	) name8114 (
		_w13939_,
		_w13940_,
		_w13941_
	);
	LUT3 #(
		.INIT('h0e)
	) name8115 (
		_w13867_,
		_w13868_,
		_w13871_,
		_w13942_
	);
	LUT3 #(
		.INIT('hb0)
	) name8116 (
		_w13867_,
		_w13865_,
		_w13868_,
		_w13943_
	);
	LUT4 #(
		.INIT('h23af)
	) name8117 (
		_w13866_,
		_w13934_,
		_w13942_,
		_w13943_,
		_w13944_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8118 (
		_w13863_,
		_w13879_,
		_w13941_,
		_w13944_,
		_w13945_
	);
	LUT4 #(
		.INIT('hcaf1)
	) name8119 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13946_
	);
	LUT4 #(
		.INIT('h1000)
	) name8120 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13947_
	);
	LUT4 #(
		.INIT('h5504)
	) name8121 (
		_w13863_,
		_w13871_,
		_w13946_,
		_w13947_,
		_w13948_
	);
	LUT4 #(
		.INIT('h0021)
	) name8122 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13949_
	);
	LUT4 #(
		.INIT('hb59e)
	) name8123 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13950_
	);
	LUT2 #(
		.INIT('h1)
	) name8124 (
		_w13863_,
		_w13871_,
		_w13951_
	);
	LUT2 #(
		.INIT('h4)
	) name8125 (
		_w13950_,
		_w13951_,
		_w13952_
	);
	LUT3 #(
		.INIT('he7)
	) name8126 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13953_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name8127 (
		_w13868_,
		_w13871_,
		_w13889_,
		_w13953_,
		_w13954_
	);
	LUT3 #(
		.INIT('h10)
	) name8128 (
		_w13948_,
		_w13952_,
		_w13954_,
		_w13955_
	);
	LUT3 #(
		.INIT('h65)
	) name8129 (
		\u2_L1_reg[24]/NET0131 ,
		_w13945_,
		_w13955_,
		_w13956_
	);
	LUT4 #(
		.INIT('hfae5)
	) name8130 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13957_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name8131 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13958_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name8132 (
		_w13863_,
		_w13873_,
		_w13957_,
		_w13958_,
		_w13959_
	);
	LUT2 #(
		.INIT('h2)
	) name8133 (
		_w13871_,
		_w13959_,
		_w13960_
	);
	LUT4 #(
		.INIT('h0200)
	) name8134 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13961_
	);
	LUT3 #(
		.INIT('h0e)
	) name8135 (
		_w13867_,
		_w13865_,
		_w13871_,
		_w13962_
	);
	LUT4 #(
		.INIT('h0015)
	) name8136 (
		_w13949_,
		_w13958_,
		_w13962_,
		_w13961_,
		_w13963_
	);
	LUT2 #(
		.INIT('h1)
	) name8137 (
		_w13863_,
		_w13963_,
		_w13964_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name8138 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13868_,
		_w13965_
	);
	LUT2 #(
		.INIT('h2)
	) name8139 (
		_w13888_,
		_w13965_,
		_w13966_
	);
	LUT3 #(
		.INIT('h4c)
	) name8140 (
		_w13864_,
		_w13867_,
		_w13865_,
		_w13967_
	);
	LUT2 #(
		.INIT('h8)
	) name8141 (
		_w13886_,
		_w13967_,
		_w13968_
	);
	LUT4 #(
		.INIT('h0040)
	) name8142 (
		_w13864_,
		_w13867_,
		_w13868_,
		_w13871_,
		_w13969_
	);
	LUT3 #(
		.INIT('h07)
	) name8143 (
		_w13876_,
		_w13930_,
		_w13969_,
		_w13970_
	);
	LUT3 #(
		.INIT('h10)
	) name8144 (
		_w13966_,
		_w13968_,
		_w13970_,
		_w13971_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name8145 (
		\u2_L1_reg[30]/NET0131 ,
		_w13960_,
		_w13964_,
		_w13971_,
		_w13972_
	);
	LUT3 #(
		.INIT('hc4)
	) name8146 (
		_w13700_,
		_w13701_,
		_w13698_,
		_w13973_
	);
	LUT4 #(
		.INIT('hdc00)
	) name8147 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13697_,
		_w13974_
	);
	LUT2 #(
		.INIT('h4)
	) name8148 (
		_w13973_,
		_w13974_,
		_w13975_
	);
	LUT4 #(
		.INIT('h0400)
	) name8149 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13976_
	);
	LUT4 #(
		.INIT('h0004)
	) name8150 (
		_w13716_,
		_w13696_,
		_w13703_,
		_w13976_,
		_w13977_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name8151 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13978_
	);
	LUT2 #(
		.INIT('h2)
	) name8152 (
		_w13697_,
		_w13978_,
		_w13979_
	);
	LUT3 #(
		.INIT('hb0)
	) name8153 (
		_w13699_,
		_w13698_,
		_w13697_,
		_w13980_
	);
	LUT4 #(
		.INIT('h44e6)
	) name8154 (
		_w13700_,
		_w13701_,
		_w13699_,
		_w13698_,
		_w13981_
	);
	LUT3 #(
		.INIT('h54)
	) name8155 (
		_w13696_,
		_w13980_,
		_w13981_,
		_w13982_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8156 (
		_w13975_,
		_w13977_,
		_w13979_,
		_w13982_,
		_w13983_
	);
	LUT3 #(
		.INIT('h02)
	) name8157 (
		_w13697_,
		_w13705_,
		_w13726_,
		_w13984_
	);
	LUT4 #(
		.INIT('h0001)
	) name8158 (
		_w13697_,
		_w13710_,
		_w13724_,
		_w13914_,
		_w13985_
	);
	LUT2 #(
		.INIT('h1)
	) name8159 (
		_w13984_,
		_w13985_,
		_w13986_
	);
	LUT3 #(
		.INIT('h56)
	) name8160 (
		\u2_L1_reg[3]/NET0131 ,
		_w13983_,
		_w13986_,
		_w13987_
	);
	LUT4 #(
		.INIT('h4000)
	) name8161 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13988_
	);
	LUT3 #(
		.INIT('he6)
	) name8162 (
		_w13414_,
		_w13415_,
		_w13413_,
		_w13989_
	);
	LUT4 #(
		.INIT('h00e6)
	) name8163 (
		_w13414_,
		_w13415_,
		_w13413_,
		_w13411_,
		_w13990_
	);
	LUT3 #(
		.INIT('hc7)
	) name8164 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13991_
	);
	LUT4 #(
		.INIT('h3230)
	) name8165 (
		_w13791_,
		_w13988_,
		_w13990_,
		_w13991_,
		_w13992_
	);
	LUT2 #(
		.INIT('h1)
	) name8166 (
		_w13410_,
		_w13992_,
		_w13993_
	);
	LUT4 #(
		.INIT('h2882)
	) name8167 (
		_w13410_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13994_
	);
	LUT4 #(
		.INIT('h4554)
	) name8168 (
		_w13410_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13995_
	);
	LUT3 #(
		.INIT('h02)
	) name8169 (
		_w13412_,
		_w13995_,
		_w13994_,
		_w13996_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name8170 (
		_w13410_,
		_w13424_,
		_w13525_,
		_w13989_,
		_w13997_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name8171 (
		_w13412_,
		_w13414_,
		_w13415_,
		_w13413_,
		_w13998_
	);
	LUT2 #(
		.INIT('h1)
	) name8172 (
		_w13411_,
		_w13998_,
		_w13999_
	);
	LUT3 #(
		.INIT('h01)
	) name8173 (
		_w13997_,
		_w13999_,
		_w13996_,
		_w14000_
	);
	LUT3 #(
		.INIT('h65)
	) name8174 (
		\u2_L1_reg[9]/NET0131 ,
		_w13993_,
		_w14000_,
		_w14001_
	);
	LUT4 #(
		.INIT('h1a00)
	) name8175 (
		_w13568_,
		_w13570_,
		_w13571_,
		_w13567_,
		_w14002_
	);
	LUT4 #(
		.INIT('hcfaf)
	) name8176 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w14003_
	);
	LUT4 #(
		.INIT('h0032)
	) name8177 (
		_w13567_,
		_w13622_,
		_w14003_,
		_w14002_,
		_w14004_
	);
	LUT4 #(
		.INIT('hbf6e)
	) name8178 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w14005_
	);
	LUT4 #(
		.INIT('h8000)
	) name8179 (
		_w13568_,
		_w13570_,
		_w13571_,
		_w13567_,
		_w14006_
	);
	LUT4 #(
		.INIT('h0109)
	) name8180 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13567_,
		_w14007_
	);
	LUT3 #(
		.INIT('h10)
	) name8181 (
		_w14006_,
		_w14007_,
		_w14005_,
		_w14008_
	);
	LUT4 #(
		.INIT('h0020)
	) name8182 (
		_w13568_,
		_w13570_,
		_w13571_,
		_w13567_,
		_w14009_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name8183 (
		_w13568_,
		_w13569_,
		_w13570_,
		_w13571_,
		_w14010_
	);
	LUT3 #(
		.INIT('h31)
	) name8184 (
		_w13567_,
		_w14009_,
		_w14010_,
		_w14011_
	);
	LUT4 #(
		.INIT('hd800)
	) name8185 (
		_w13566_,
		_w14004_,
		_w14008_,
		_w14011_,
		_w14012_
	);
	LUT2 #(
		.INIT('h9)
	) name8186 (
		\u2_L1_reg[18]/P0001 ,
		_w14012_,
		_w14013_
	);
	LUT4 #(
		.INIT('hc963)
	) name8187 (
		decrypt_pad,
		\u2_R0_reg[23]/NET0131 ,
		\u2_uk_K_r0_reg[16]/NET0131 ,
		\u2_uk_K_r0_reg[50]/NET0131 ,
		_w14014_
	);
	LUT4 #(
		.INIT('hc963)
	) name8188 (
		decrypt_pad,
		\u2_R0_reg[22]/NET0131 ,
		\u2_uk_K_r0_reg[31]/NET0131 ,
		\u2_uk_K_r0_reg[37]/NET0131 ,
		_w14015_
	);
	LUT4 #(
		.INIT('hc693)
	) name8189 (
		decrypt_pad,
		\u2_R0_reg[20]/NET0131 ,
		\u2_uk_K_r0_reg[0]/NET0131 ,
		\u2_uk_K_r0_reg[21]/NET0131 ,
		_w14016_
	);
	LUT4 #(
		.INIT('hc693)
	) name8190 (
		decrypt_pad,
		\u2_R0_reg[25]/NET0131 ,
		\u2_uk_K_r0_reg[16]/NET0131 ,
		\u2_uk_K_r0_reg[37]/NET0131 ,
		_w14017_
	);
	LUT4 #(
		.INIT('hc693)
	) name8191 (
		decrypt_pad,
		\u2_R0_reg[21]/NET0131 ,
		\u2_uk_K_r0_reg[15]/NET0131 ,
		\u2_uk_K_r0_reg[36]/NET0131 ,
		_w14018_
	);
	LUT3 #(
		.INIT('h20)
	) name8192 (
		_w14016_,
		_w14018_,
		_w14017_,
		_w14019_
	);
	LUT4 #(
		.INIT('h168a)
	) name8193 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14020_
	);
	LUT2 #(
		.INIT('h1)
	) name8194 (
		_w14014_,
		_w14020_,
		_w14021_
	);
	LUT4 #(
		.INIT('hc693)
	) name8195 (
		decrypt_pad,
		\u2_R0_reg[24]/NET0131 ,
		\u2_uk_K_r0_reg[21]/NET0131 ,
		\u2_uk_K_r0_reg[42]/NET0131 ,
		_w14022_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name8196 (
		_w14014_,
		_w14015_,
		_w14016_,
		_w14018_,
		_w14023_
	);
	LUT4 #(
		.INIT('h0004)
	) name8197 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14024_
	);
	LUT4 #(
		.INIT('h3ffb)
	) name8198 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14025_
	);
	LUT3 #(
		.INIT('h2a)
	) name8199 (
		_w14022_,
		_w14023_,
		_w14025_,
		_w14026_
	);
	LUT2 #(
		.INIT('h4)
	) name8200 (
		_w14021_,
		_w14026_,
		_w14027_
	);
	LUT4 #(
		.INIT('h0040)
	) name8201 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14028_
	);
	LUT4 #(
		.INIT('h0800)
	) name8202 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14029_
	);
	LUT4 #(
		.INIT('h0200)
	) name8203 (
		_w14014_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14030_
	);
	LUT3 #(
		.INIT('h01)
	) name8204 (
		_w14029_,
		_w14030_,
		_w14028_,
		_w14031_
	);
	LUT4 #(
		.INIT('h1400)
	) name8205 (
		_w14014_,
		_w14015_,
		_w14016_,
		_w14018_,
		_w14032_
	);
	LUT4 #(
		.INIT('h0010)
	) name8206 (
		_w14014_,
		_w14015_,
		_w14016_,
		_w14017_,
		_w14033_
	);
	LUT2 #(
		.INIT('h8)
	) name8207 (
		_w14014_,
		_w14015_,
		_w14034_
	);
	LUT4 #(
		.INIT('hfd7d)
	) name8208 (
		_w14014_,
		_w14015_,
		_w14016_,
		_w14018_,
		_w14035_
	);
	LUT3 #(
		.INIT('h10)
	) name8209 (
		_w14032_,
		_w14033_,
		_w14035_,
		_w14036_
	);
	LUT3 #(
		.INIT('h15)
	) name8210 (
		_w14022_,
		_w14031_,
		_w14036_,
		_w14037_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name8211 (
		_w14014_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14038_
	);
	LUT2 #(
		.INIT('h1)
	) name8212 (
		_w14015_,
		_w14038_,
		_w14039_
	);
	LUT4 #(
		.INIT('h0010)
	) name8213 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14040_
	);
	LUT4 #(
		.INIT('h77ef)
	) name8214 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14041_
	);
	LUT3 #(
		.INIT('h01)
	) name8215 (
		_w14016_,
		_w14018_,
		_w14017_,
		_w14042_
	);
	LUT4 #(
		.INIT('he4f5)
	) name8216 (
		_w14014_,
		_w14015_,
		_w14041_,
		_w14042_,
		_w14043_
	);
	LUT2 #(
		.INIT('h4)
	) name8217 (
		_w14039_,
		_w14043_,
		_w14044_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name8218 (
		\u2_L0_reg[11]/NET0131 ,
		_w14037_,
		_w14027_,
		_w14044_,
		_w14045_
	);
	LUT4 #(
		.INIT('hc963)
	) name8219 (
		decrypt_pad,
		\u2_R0_reg[26]/NET0131 ,
		\u2_uk_K_r0_reg[29]/NET0131 ,
		\u2_uk_K_r0_reg[8]/NET0131 ,
		_w14046_
	);
	LUT4 #(
		.INIT('hc693)
	) name8220 (
		decrypt_pad,
		\u2_R0_reg[25]/NET0131 ,
		\u2_uk_K_r0_reg[23]/NET0131 ,
		\u2_uk_K_r0_reg[44]/NET0131 ,
		_w14047_
	);
	LUT4 #(
		.INIT('hc693)
	) name8221 (
		decrypt_pad,
		\u2_R0_reg[24]/NET0131 ,
		\u2_uk_K_r0_reg[43]/NET0131 ,
		\u2_uk_K_r0_reg[9]/NET0131 ,
		_w14048_
	);
	LUT4 #(
		.INIT('hc963)
	) name8222 (
		decrypt_pad,
		\u2_R0_reg[29]/NET0131 ,
		\u2_uk_K_r0_reg[45]/NET0131 ,
		\u2_uk_K_r0_reg[51]/NET0131 ,
		_w14049_
	);
	LUT2 #(
		.INIT('h4)
	) name8223 (
		_w14048_,
		_w14049_,
		_w14050_
	);
	LUT4 #(
		.INIT('h0200)
	) name8224 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14051_
	);
	LUT4 #(
		.INIT('h0008)
	) name8225 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14052_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name8226 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14053_
	);
	LUT4 #(
		.INIT('hc693)
	) name8227 (
		decrypt_pad,
		\u2_R0_reg[28]/NET0131 ,
		\u2_uk_K_r0_reg[28]/NET0131 ,
		\u2_uk_K_r0_reg[49]/NET0131 ,
		_w14054_
	);
	LUT4 #(
		.INIT('h9cfc)
	) name8228 (
		_w14046_,
		_w14047_,
		_w14049_,
		_w14054_,
		_w14055_
	);
	LUT4 #(
		.INIT('hc693)
	) name8229 (
		decrypt_pad,
		\u2_R0_reg[27]/NET0131 ,
		\u2_uk_K_r0_reg[45]/NET0131 ,
		\u2_uk_K_r0_reg[7]/NET0131 ,
		_w14056_
	);
	LUT4 #(
		.INIT('h3b00)
	) name8230 (
		_w14048_,
		_w14053_,
		_w14055_,
		_w14056_,
		_w14057_
	);
	LUT2 #(
		.INIT('h4)
	) name8231 (
		_w14047_,
		_w14056_,
		_w14058_
	);
	LUT4 #(
		.INIT('heef2)
	) name8232 (
		_w14046_,
		_w14047_,
		_w14049_,
		_w14056_,
		_w14059_
	);
	LUT2 #(
		.INIT('h6)
	) name8233 (
		_w14046_,
		_w14048_,
		_w14060_
	);
	LUT4 #(
		.INIT('h0002)
	) name8234 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14061_
	);
	LUT4 #(
		.INIT('h5afd)
	) name8235 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14062_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name8236 (
		_w14048_,
		_w14058_,
		_w14059_,
		_w14062_,
		_w14063_
	);
	LUT4 #(
		.INIT('h1000)
	) name8237 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14064_
	);
	LUT4 #(
		.INIT('he3ff)
	) name8238 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14065_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name8239 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14066_
	);
	LUT3 #(
		.INIT('he0)
	) name8240 (
		_w14056_,
		_w14065_,
		_w14066_,
		_w14067_
	);
	LUT4 #(
		.INIT('h0100)
	) name8241 (
		_w14046_,
		_w14047_,
		_w14049_,
		_w14056_,
		_w14068_
	);
	LUT4 #(
		.INIT('h0084)
	) name8242 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14056_,
		_w14069_
	);
	LUT2 #(
		.INIT('h1)
	) name8243 (
		_w14068_,
		_w14069_,
		_w14070_
	);
	LUT4 #(
		.INIT('he400)
	) name8244 (
		_w14054_,
		_w14063_,
		_w14067_,
		_w14070_,
		_w14071_
	);
	LUT3 #(
		.INIT('h65)
	) name8245 (
		\u2_L0_reg[22]/NET0131 ,
		_w14057_,
		_w14071_,
		_w14072_
	);
	LUT4 #(
		.INIT('hc963)
	) name8246 (
		decrypt_pad,
		\u2_R0_reg[4]/NET0131 ,
		\u2_uk_K_r0_reg[20]/NET0131 ,
		\u2_uk_K_r0_reg[24]/P0001 ,
		_w14073_
	);
	LUT4 #(
		.INIT('hc963)
	) name8247 (
		decrypt_pad,
		\u2_R0_reg[3]/NET0131 ,
		\u2_uk_K_r0_reg[10]/NET0131 ,
		\u2_uk_K_r0_reg[46]/NET0131 ,
		_w14074_
	);
	LUT4 #(
		.INIT('hc693)
	) name8248 (
		decrypt_pad,
		\u2_R0_reg[2]/NET0131 ,
		\u2_uk_K_r0_reg[12]/NET0131 ,
		\u2_uk_K_r0_reg[33]/NET0131 ,
		_w14075_
	);
	LUT4 #(
		.INIT('hc693)
	) name8249 (
		decrypt_pad,
		\u2_R0_reg[32]/NET0131 ,
		\u2_uk_K_r0_reg[33]/NET0131 ,
		\u2_uk_K_r0_reg[54]/NET0131 ,
		_w14076_
	);
	LUT4 #(
		.INIT('hc963)
	) name8250 (
		decrypt_pad,
		\u2_R0_reg[1]/NET0131 ,
		\u2_uk_K_r0_reg[18]/NET0131 ,
		\u2_uk_K_r0_reg[54]/NET0131 ,
		_w14077_
	);
	LUT4 #(
		.INIT('hc693)
	) name8251 (
		decrypt_pad,
		\u2_R0_reg[5]/NET0131 ,
		\u2_uk_K_r0_reg[27]/NET0131 ,
		\u2_uk_K_r0_reg[48]/NET0131 ,
		_w14078_
	);
	LUT4 #(
		.INIT('hfdba)
	) name8252 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14079_
	);
	LUT2 #(
		.INIT('h1)
	) name8253 (
		_w14074_,
		_w14079_,
		_w14080_
	);
	LUT2 #(
		.INIT('h2)
	) name8254 (
		_w14078_,
		_w14076_,
		_w14081_
	);
	LUT4 #(
		.INIT('h0800)
	) name8255 (
		_w14075_,
		_w14078_,
		_w14076_,
		_w14074_,
		_w14082_
	);
	LUT4 #(
		.INIT('hf6fe)
	) name8256 (
		_w14075_,
		_w14078_,
		_w14076_,
		_w14074_,
		_w14083_
	);
	LUT2 #(
		.INIT('h2)
	) name8257 (
		_w14077_,
		_w14083_,
		_w14084_
	);
	LUT4 #(
		.INIT('h0800)
	) name8258 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14085_
	);
	LUT2 #(
		.INIT('h8)
	) name8259 (
		_w14078_,
		_w14076_,
		_w14086_
	);
	LUT2 #(
		.INIT('h4)
	) name8260 (
		_w14075_,
		_w14074_,
		_w14087_
	);
	LUT3 #(
		.INIT('hae)
	) name8261 (
		_w14075_,
		_w14077_,
		_w14074_,
		_w14088_
	);
	LUT4 #(
		.INIT('h7707)
	) name8262 (
		_w14085_,
		_w14074_,
		_w14086_,
		_w14088_,
		_w14089_
	);
	LUT4 #(
		.INIT('h5455)
	) name8263 (
		_w14073_,
		_w14080_,
		_w14084_,
		_w14089_,
		_w14090_
	);
	LUT3 #(
		.INIT('h02)
	) name8264 (
		_w14075_,
		_w14078_,
		_w14076_,
		_w14091_
	);
	LUT4 #(
		.INIT('hcfc5)
	) name8265 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14092_
	);
	LUT2 #(
		.INIT('h2)
	) name8266 (
		_w14074_,
		_w14092_,
		_w14093_
	);
	LUT3 #(
		.INIT('h8c)
	) name8267 (
		_w14075_,
		_w14077_,
		_w14074_,
		_w14094_
	);
	LUT4 #(
		.INIT('h0100)
	) name8268 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14095_
	);
	LUT2 #(
		.INIT('h2)
	) name8269 (
		_w14076_,
		_w14074_,
		_w14096_
	);
	LUT4 #(
		.INIT('h02c2)
	) name8270 (
		_w14075_,
		_w14077_,
		_w14076_,
		_w14074_,
		_w14097_
	);
	LUT4 #(
		.INIT('h0301)
	) name8271 (
		_w14081_,
		_w14095_,
		_w14097_,
		_w14094_,
		_w14098_
	);
	LUT2 #(
		.INIT('h4)
	) name8272 (
		_w14077_,
		_w14074_,
		_w14099_
	);
	LUT3 #(
		.INIT('had)
	) name8273 (
		_w14075_,
		_w14078_,
		_w14076_,
		_w14100_
	);
	LUT3 #(
		.INIT('h80)
	) name8274 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14101_
	);
	LUT4 #(
		.INIT('h7bdb)
	) name8275 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14102_
	);
	LUT4 #(
		.INIT('hfbc8)
	) name8276 (
		_w14077_,
		_w14074_,
		_w14100_,
		_w14102_,
		_w14103_
	);
	LUT4 #(
		.INIT('h7500)
	) name8277 (
		_w14073_,
		_w14093_,
		_w14098_,
		_w14103_,
		_w14104_
	);
	LUT3 #(
		.INIT('h65)
	) name8278 (
		\u2_L0_reg[31]/NET0131 ,
		_w14090_,
		_w14104_,
		_w14105_
	);
	LUT4 #(
		.INIT('hc693)
	) name8279 (
		decrypt_pad,
		\u2_R0_reg[13]/NET0131 ,
		\u2_uk_K_r0_reg[41]/NET0131 ,
		\u2_uk_K_r0_reg[5]/NET0131 ,
		_w14106_
	);
	LUT4 #(
		.INIT('hc963)
	) name8280 (
		decrypt_pad,
		\u2_R0_reg[12]/NET0131 ,
		\u2_uk_K_r0_reg[11]/NET0131 ,
		\u2_uk_K_r0_reg[47]/NET0131 ,
		_w14107_
	);
	LUT2 #(
		.INIT('h2)
	) name8281 (
		_w14106_,
		_w14107_,
		_w14108_
	);
	LUT4 #(
		.INIT('hc693)
	) name8282 (
		decrypt_pad,
		\u2_R0_reg[15]/NET0131 ,
		\u2_uk_K_r0_reg[18]/NET0131 ,
		\u2_uk_K_r0_reg[39]/NET0131 ,
		_w14109_
	);
	LUT4 #(
		.INIT('hc693)
	) name8283 (
		decrypt_pad,
		\u2_R0_reg[14]/NET0131 ,
		\u2_uk_K_r0_reg[10]/NET0131 ,
		\u2_uk_K_r0_reg[6]/NET0131 ,
		_w14110_
	);
	LUT4 #(
		.INIT('h0006)
	) name8284 (
		_w14106_,
		_w14107_,
		_w14109_,
		_w14110_,
		_w14111_
	);
	LUT2 #(
		.INIT('h4)
	) name8285 (
		_w14106_,
		_w14109_,
		_w14112_
	);
	LUT4 #(
		.INIT('hc963)
	) name8286 (
		decrypt_pad,
		\u2_R0_reg[17]/NET0131 ,
		\u2_uk_K_r0_reg[27]/NET0131 ,
		\u2_uk_K_r0_reg[6]/NET0131 ,
		_w14113_
	);
	LUT4 #(
		.INIT('h0400)
	) name8287 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14109_,
		_w14114_
	);
	LUT2 #(
		.INIT('h8)
	) name8288 (
		_w14106_,
		_w14109_,
		_w14115_
	);
	LUT4 #(
		.INIT('h2000)
	) name8289 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14109_,
		_w14116_
	);
	LUT4 #(
		.INIT('hc693)
	) name8290 (
		decrypt_pad,
		\u2_R0_reg[16]/NET0131 ,
		\u2_uk_K_r0_reg[26]/NET0131 ,
		\u2_uk_K_r0_reg[47]/NET0131 ,
		_w14117_
	);
	LUT4 #(
		.INIT('h0100)
	) name8291 (
		_w14116_,
		_w14114_,
		_w14111_,
		_w14117_,
		_w14118_
	);
	LUT3 #(
		.INIT('h01)
	) name8292 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14119_
	);
	LUT4 #(
		.INIT('h0001)
	) name8293 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14109_,
		_w14120_
	);
	LUT4 #(
		.INIT('h0008)
	) name8294 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14121_
	);
	LUT4 #(
		.INIT('h7ff7)
	) name8295 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14122_
	);
	LUT3 #(
		.INIT('h70)
	) name8296 (
		_w14120_,
		_w14110_,
		_w14122_,
		_w14123_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8297 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14109_,
		_w14124_
	);
	LUT4 #(
		.INIT('h7e00)
	) name8298 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14109_,
		_w14125_
	);
	LUT3 #(
		.INIT('h40)
	) name8299 (
		_w14113_,
		_w14107_,
		_w14110_,
		_w14126_
	);
	LUT3 #(
		.INIT('h0b)
	) name8300 (
		_w14106_,
		_w14113_,
		_w14109_,
		_w14127_
	);
	LUT3 #(
		.INIT('h45)
	) name8301 (
		_w14125_,
		_w14126_,
		_w14127_,
		_w14128_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name8302 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14129_
	);
	LUT4 #(
		.INIT('h0040)
	) name8303 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14130_
	);
	LUT4 #(
		.INIT('h2000)
	) name8304 (
		_w14106_,
		_w14107_,
		_w14109_,
		_w14110_,
		_w14131_
	);
	LUT4 #(
		.INIT('h0004)
	) name8305 (
		_w14117_,
		_w14129_,
		_w14131_,
		_w14130_,
		_w14132_
	);
	LUT4 #(
		.INIT('h7077)
	) name8306 (
		_w14118_,
		_w14123_,
		_w14128_,
		_w14132_,
		_w14133_
	);
	LUT3 #(
		.INIT('hbe)
	) name8307 (
		_w14113_,
		_w14107_,
		_w14110_,
		_w14134_
	);
	LUT2 #(
		.INIT('h2)
	) name8308 (
		_w14112_,
		_w14134_,
		_w14135_
	);
	LUT3 #(
		.INIT('h04)
	) name8309 (
		_w14113_,
		_w14107_,
		_w14110_,
		_w14136_
	);
	LUT3 #(
		.INIT('h02)
	) name8310 (
		_w14113_,
		_w14109_,
		_w14110_,
		_w14137_
	);
	LUT4 #(
		.INIT('h135f)
	) name8311 (
		_w14115_,
		_w14108_,
		_w14136_,
		_w14137_,
		_w14138_
	);
	LUT2 #(
		.INIT('h4)
	) name8312 (
		_w14135_,
		_w14138_,
		_w14139_
	);
	LUT3 #(
		.INIT('h65)
	) name8313 (
		\u2_L0_reg[20]/NET0131 ,
		_w14133_,
		_w14139_,
		_w14140_
	);
	LUT4 #(
		.INIT('h3fd2)
	) name8314 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14141_
	);
	LUT4 #(
		.INIT('hab6f)
	) name8315 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14142_
	);
	LUT4 #(
		.INIT('h0200)
	) name8316 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14143_
	);
	LUT4 #(
		.INIT('h00e4)
	) name8317 (
		_w14014_,
		_w14142_,
		_w14141_,
		_w14143_,
		_w14144_
	);
	LUT2 #(
		.INIT('h1)
	) name8318 (
		_w14022_,
		_w14144_,
		_w14145_
	);
	LUT4 #(
		.INIT('hcf6f)
	) name8319 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14146_
	);
	LUT2 #(
		.INIT('h2)
	) name8320 (
		_w14014_,
		_w14146_,
		_w14147_
	);
	LUT4 #(
		.INIT('h0102)
	) name8321 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14148_
	);
	LUT4 #(
		.INIT('h77dc)
	) name8322 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14149_
	);
	LUT4 #(
		.INIT('h0302)
	) name8323 (
		_w14014_,
		_w14033_,
		_w14029_,
		_w14149_,
		_w14150_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8324 (
		_w14022_,
		_w14147_,
		_w14148_,
		_w14150_,
		_w14151_
	);
	LUT4 #(
		.INIT('h2000)
	) name8325 (
		_w14014_,
		_w14015_,
		_w14018_,
		_w14017_,
		_w14152_
	);
	LUT2 #(
		.INIT('h1)
	) name8326 (
		_w14024_,
		_w14152_,
		_w14153_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name8327 (
		\u2_L0_reg[29]/NET0131 ,
		_w14151_,
		_w14145_,
		_w14153_,
		_w14154_
	);
	LUT4 #(
		.INIT('he63f)
	) name8328 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14155_
	);
	LUT2 #(
		.INIT('h2)
	) name8329 (
		_w14014_,
		_w14155_,
		_w14156_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name8330 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14157_
	);
	LUT4 #(
		.INIT('h1000)
	) name8331 (
		_w14014_,
		_w14015_,
		_w14016_,
		_w14017_,
		_w14158_
	);
	LUT4 #(
		.INIT('h0032)
	) name8332 (
		_w14014_,
		_w14024_,
		_w14157_,
		_w14158_,
		_w14159_
	);
	LUT3 #(
		.INIT('h45)
	) name8333 (
		_w14022_,
		_w14156_,
		_w14159_,
		_w14160_
	);
	LUT4 #(
		.INIT('heeae)
	) name8334 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14161_
	);
	LUT2 #(
		.INIT('h1)
	) name8335 (
		_w14014_,
		_w14161_,
		_w14162_
	);
	LUT3 #(
		.INIT('h80)
	) name8336 (
		_w14015_,
		_w14018_,
		_w14017_,
		_w14163_
	);
	LUT4 #(
		.INIT('h2000)
	) name8337 (
		_w14014_,
		_w14015_,
		_w14016_,
		_w14017_,
		_w14164_
	);
	LUT3 #(
		.INIT('h01)
	) name8338 (
		_w14040_,
		_w14163_,
		_w14164_,
		_w14165_
	);
	LUT3 #(
		.INIT('hb6)
	) name8339 (
		_w14016_,
		_w14018_,
		_w14017_,
		_w14166_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name8340 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14167_
	);
	LUT4 #(
		.INIT('h4445)
	) name8341 (
		_w14014_,
		_w14015_,
		_w14016_,
		_w14017_,
		_w14168_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name8342 (
		_w14034_,
		_w14166_,
		_w14167_,
		_w14168_,
		_w14169_
	);
	LUT4 #(
		.INIT('h7500)
	) name8343 (
		_w14022_,
		_w14162_,
		_w14165_,
		_w14169_,
		_w14170_
	);
	LUT3 #(
		.INIT('h65)
	) name8344 (
		\u2_L0_reg[4]/NET0131 ,
		_w14160_,
		_w14170_,
		_w14171_
	);
	LUT4 #(
		.INIT('hc963)
	) name8345 (
		decrypt_pad,
		\u2_R0_reg[32]/NET0131 ,
		\u2_uk_K_r0_reg[14]/NET0131 ,
		\u2_uk_K_r0_reg[52]/P0001 ,
		_w14172_
	);
	LUT4 #(
		.INIT('hc693)
	) name8346 (
		decrypt_pad,
		\u2_R0_reg[31]/P0001 ,
		\u2_uk_K_r0_reg[42]/NET0131 ,
		\u2_uk_K_r0_reg[8]/NET0131 ,
		_w14173_
	);
	LUT4 #(
		.INIT('hc963)
	) name8347 (
		decrypt_pad,
		\u2_R0_reg[28]/NET0131 ,
		\u2_uk_K_r0_reg[23]/NET0131 ,
		\u2_uk_K_r0_reg[2]/NET0131 ,
		_w14174_
	);
	LUT4 #(
		.INIT('hc693)
	) name8348 (
		decrypt_pad,
		\u2_R0_reg[29]/NET0131 ,
		\u2_uk_K_r0_reg[29]/NET0131 ,
		\u2_uk_K_r0_reg[50]/NET0131 ,
		_w14175_
	);
	LUT4 #(
		.INIT('hc693)
	) name8349 (
		decrypt_pad,
		\u2_R0_reg[1]/NET0131 ,
		\u2_uk_K_r0_reg[14]/NET0131 ,
		\u2_uk_K_r0_reg[35]/NET0131 ,
		_w14176_
	);
	LUT4 #(
		.INIT('hc693)
	) name8350 (
		decrypt_pad,
		\u2_R0_reg[30]/NET0131 ,
		\u2_uk_K_r0_reg[30]/NET0131 ,
		\u2_uk_K_r0_reg[51]/NET0131 ,
		_w14177_
	);
	LUT4 #(
		.INIT('h1000)
	) name8351 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14178_
	);
	LUT4 #(
		.INIT('hebfb)
	) name8352 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14179_
	);
	LUT2 #(
		.INIT('h2)
	) name8353 (
		_w14174_,
		_w14177_,
		_w14180_
	);
	LUT2 #(
		.INIT('h4)
	) name8354 (
		_w14174_,
		_w14177_,
		_w14181_
	);
	LUT4 #(
		.INIT('h7407)
	) name8355 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14182_
	);
	LUT3 #(
		.INIT('h08)
	) name8356 (
		_w14175_,
		_w14174_,
		_w14177_,
		_w14183_
	);
	LUT4 #(
		.INIT('h0020)
	) name8357 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14184_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name8358 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14185_
	);
	LUT4 #(
		.INIT('he400)
	) name8359 (
		_w14173_,
		_w14182_,
		_w14179_,
		_w14185_,
		_w14186_
	);
	LUT2 #(
		.INIT('h1)
	) name8360 (
		_w14172_,
		_w14186_,
		_w14187_
	);
	LUT4 #(
		.INIT('hcf45)
	) name8361 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14188_
	);
	LUT4 #(
		.INIT('h22d2)
	) name8362 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14189_
	);
	LUT4 #(
		.INIT('h0001)
	) name8363 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14190_
	);
	LUT4 #(
		.INIT('h0400)
	) name8364 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14191_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name8365 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14192_
	);
	LUT4 #(
		.INIT('h1f00)
	) name8366 (
		_w14172_,
		_w14188_,
		_w14189_,
		_w14192_,
		_w14193_
	);
	LUT4 #(
		.INIT('h0800)
	) name8367 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14194_
	);
	LUT2 #(
		.INIT('h8)
	) name8368 (
		_w14172_,
		_w14194_,
		_w14195_
	);
	LUT4 #(
		.INIT('h2002)
	) name8369 (
		_w14172_,
		_w14175_,
		_w14174_,
		_w14177_,
		_w14196_
	);
	LUT2 #(
		.INIT('h1)
	) name8370 (
		_w14196_,
		_w14184_,
		_w14197_
	);
	LUT4 #(
		.INIT('h5404)
	) name8371 (
		_w14195_,
		_w14197_,
		_w14173_,
		_w14193_,
		_w14198_
	);
	LUT3 #(
		.INIT('h9a)
	) name8372 (
		\u2_L0_reg[5]/NET0131 ,
		_w14187_,
		_w14198_,
		_w14199_
	);
	LUT4 #(
		.INIT('haf41)
	) name8373 (
		_w14106_,
		_w14113_,
		_w14109_,
		_w14110_,
		_w14200_
	);
	LUT2 #(
		.INIT('h2)
	) name8374 (
		_w14107_,
		_w14200_,
		_w14201_
	);
	LUT4 #(
		.INIT('h0020)
	) name8375 (
		_w14113_,
		_w14107_,
		_w14109_,
		_w14110_,
		_w14202_
	);
	LUT3 #(
		.INIT('h04)
	) name8376 (
		_w14120_,
		_w14129_,
		_w14202_,
		_w14203_
	);
	LUT3 #(
		.INIT('h45)
	) name8377 (
		_w14117_,
		_w14201_,
		_w14203_,
		_w14204_
	);
	LUT4 #(
		.INIT('hcfe7)
	) name8378 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14205_
	);
	LUT4 #(
		.INIT('h7bff)
	) name8379 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14206_
	);
	LUT4 #(
		.INIT('hfdbd)
	) name8380 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14207_
	);
	LUT4 #(
		.INIT('hc480)
	) name8381 (
		_w14109_,
		_w14206_,
		_w14207_,
		_w14205_,
		_w14208_
	);
	LUT4 #(
		.INIT('h7bfe)
	) name8382 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14209_
	);
	LUT2 #(
		.INIT('h1)
	) name8383 (
		_w14109_,
		_w14209_,
		_w14210_
	);
	LUT3 #(
		.INIT('h13)
	) name8384 (
		_w14115_,
		_w14131_,
		_w14136_,
		_w14211_
	);
	LUT4 #(
		.INIT('h0d00)
	) name8385 (
		_w14117_,
		_w14208_,
		_w14210_,
		_w14211_,
		_w14212_
	);
	LUT3 #(
		.INIT('h65)
	) name8386 (
		\u2_L0_reg[10]/NET0131 ,
		_w14204_,
		_w14212_,
		_w14213_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name8387 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14214_
	);
	LUT2 #(
		.INIT('h2)
	) name8388 (
		_w14056_,
		_w14214_,
		_w14215_
	);
	LUT4 #(
		.INIT('h0400)
	) name8389 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14216_
	);
	LUT3 #(
		.INIT('h02)
	) name8390 (
		_w14054_,
		_w14064_,
		_w14216_,
		_w14217_
	);
	LUT2 #(
		.INIT('h9)
	) name8391 (
		_w14048_,
		_w14049_,
		_w14218_
	);
	LUT4 #(
		.INIT('h2022)
	) name8392 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14056_,
		_w14219_
	);
	LUT3 #(
		.INIT('h45)
	) name8393 (
		_w14052_,
		_w14218_,
		_w14219_,
		_w14220_
	);
	LUT3 #(
		.INIT('h40)
	) name8394 (
		_w14215_,
		_w14217_,
		_w14220_,
		_w14221_
	);
	LUT3 #(
		.INIT('h47)
	) name8395 (
		_w14046_,
		_w14047_,
		_w14056_,
		_w14222_
	);
	LUT3 #(
		.INIT('h04)
	) name8396 (
		_w14046_,
		_w14048_,
		_w14049_,
		_w14223_
	);
	LUT4 #(
		.INIT('h0010)
	) name8397 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14224_
	);
	LUT4 #(
		.INIT('h0301)
	) name8398 (
		_w14050_,
		_w14054_,
		_w14224_,
		_w14222_,
		_w14225_
	);
	LUT2 #(
		.INIT('h6)
	) name8399 (
		_w14047_,
		_w14049_,
		_w14226_
	);
	LUT4 #(
		.INIT('h134c)
	) name8400 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14227_
	);
	LUT4 #(
		.INIT('h2006)
	) name8401 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14228_
	);
	LUT3 #(
		.INIT('h0e)
	) name8402 (
		_w14056_,
		_w14227_,
		_w14228_,
		_w14229_
	);
	LUT2 #(
		.INIT('h8)
	) name8403 (
		_w14225_,
		_w14229_,
		_w14230_
	);
	LUT3 #(
		.INIT('ha9)
	) name8404 (
		\u2_L0_reg[12]/NET0131 ,
		_w14221_,
		_w14230_,
		_w14231_
	);
	LUT4 #(
		.INIT('hc963)
	) name8405 (
		decrypt_pad,
		\u2_R0_reg[20]/NET0131 ,
		\u2_uk_K_r0_reg[30]/NET0131 ,
		\u2_uk_K_r0_reg[9]/NET0131 ,
		_w14232_
	);
	LUT4 #(
		.INIT('hc693)
	) name8406 (
		decrypt_pad,
		\u2_R0_reg[16]/NET0131 ,
		\u2_uk_K_r0_reg[22]/NET0131 ,
		\u2_uk_K_r0_reg[43]/NET0131 ,
		_w14233_
	);
	LUT4 #(
		.INIT('hc963)
	) name8407 (
		decrypt_pad,
		\u2_R0_reg[17]/NET0131 ,
		\u2_uk_K_r0_reg[38]/NET0131 ,
		\u2_uk_K_r0_reg[44]/NET0131 ,
		_w14234_
	);
	LUT4 #(
		.INIT('hc963)
	) name8408 (
		decrypt_pad,
		\u2_R0_reg[18]/NET0131 ,
		\u2_uk_K_r0_reg[28]/NET0131 ,
		\u2_uk_K_r0_reg[7]/NET0131 ,
		_w14235_
	);
	LUT4 #(
		.INIT('hc963)
	) name8409 (
		decrypt_pad,
		\u2_R0_reg[21]/NET0131 ,
		\u2_uk_K_r0_reg[0]/NET0131 ,
		\u2_uk_K_r0_reg[38]/NET0131 ,
		_w14236_
	);
	LUT3 #(
		.INIT('h2e)
	) name8410 (
		_w14233_,
		_w14236_,
		_w14235_,
		_w14237_
	);
	LUT4 #(
		.INIT('h2004)
	) name8411 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14238_
	);
	LUT4 #(
		.INIT('h1012)
	) name8412 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14239_
	);
	LUT4 #(
		.INIT('h0080)
	) name8413 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14240_
	);
	LUT4 #(
		.INIT('hc963)
	) name8414 (
		decrypt_pad,
		\u2_R0_reg[19]/NET0131 ,
		\u2_uk_K_r0_reg[15]/NET0131 ,
		\u2_uk_K_r0_reg[49]/NET0131 ,
		_w14241_
	);
	LUT4 #(
		.INIT('h00df)
	) name8415 (
		_w14234_,
		_w14236_,
		_w14235_,
		_w14241_,
		_w14242_
	);
	LUT3 #(
		.INIT('h10)
	) name8416 (
		_w14239_,
		_w14240_,
		_w14242_,
		_w14243_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8417 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14241_,
		_w14244_
	);
	LUT3 #(
		.INIT('h04)
	) name8418 (
		_w14233_,
		_w14234_,
		_w14235_,
		_w14245_
	);
	LUT4 #(
		.INIT('h5fbb)
	) name8419 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14246_
	);
	LUT2 #(
		.INIT('h8)
	) name8420 (
		_w14244_,
		_w14246_,
		_w14247_
	);
	LUT4 #(
		.INIT('h4445)
	) name8421 (
		_w14232_,
		_w14238_,
		_w14243_,
		_w14247_,
		_w14248_
	);
	LUT4 #(
		.INIT('ha747)
	) name8422 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14249_
	);
	LUT2 #(
		.INIT('h2)
	) name8423 (
		_w14241_,
		_w14249_,
		_w14250_
	);
	LUT2 #(
		.INIT('h1)
	) name8424 (
		_w14235_,
		_w14241_,
		_w14251_
	);
	LUT3 #(
		.INIT('hbe)
	) name8425 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14252_
	);
	LUT2 #(
		.INIT('h2)
	) name8426 (
		_w14251_,
		_w14252_,
		_w14253_
	);
	LUT3 #(
		.INIT('h80)
	) name8427 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14254_
	);
	LUT2 #(
		.INIT('h2)
	) name8428 (
		_w14235_,
		_w14241_,
		_w14255_
	);
	LUT4 #(
		.INIT('hfdd7)
	) name8429 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14256_
	);
	LUT3 #(
		.INIT('h70)
	) name8430 (
		_w14254_,
		_w14255_,
		_w14256_,
		_w14257_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8431 (
		_w14232_,
		_w14250_,
		_w14253_,
		_w14257_,
		_w14258_
	);
	LUT4 #(
		.INIT('hfef7)
	) name8432 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14259_
	);
	LUT4 #(
		.INIT('h1000)
	) name8433 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14260_
	);
	LUT4 #(
		.INIT('hebff)
	) name8434 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14261_
	);
	LUT3 #(
		.INIT('hd8)
	) name8435 (
		_w14241_,
		_w14259_,
		_w14261_,
		_w14262_
	);
	LUT4 #(
		.INIT('h5655)
	) name8436 (
		\u2_L0_reg[14]/NET0131 ,
		_w14258_,
		_w14248_,
		_w14262_,
		_w14263_
	);
	LUT4 #(
		.INIT('h1000)
	) name8437 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14264_
	);
	LUT4 #(
		.INIT('hef11)
	) name8438 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14265_
	);
	LUT4 #(
		.INIT('h00a1)
	) name8439 (
		_w14075_,
		_w14077_,
		_w14076_,
		_w14074_,
		_w14266_
	);
	LUT4 #(
		.INIT('h0400)
	) name8440 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14267_
	);
	LUT4 #(
		.INIT('h7b7f)
	) name8441 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14268_
	);
	LUT4 #(
		.INIT('h0d00)
	) name8442 (
		_w14074_,
		_w14265_,
		_w14266_,
		_w14268_,
		_w14269_
	);
	LUT4 #(
		.INIT('h0048)
	) name8443 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14270_
	);
	LUT4 #(
		.INIT('h4100)
	) name8444 (
		_w14073_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14271_
	);
	LUT3 #(
		.INIT('ha8)
	) name8445 (
		_w14074_,
		_w14270_,
		_w14271_,
		_w14272_
	);
	LUT4 #(
		.INIT('hccc8)
	) name8446 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14273_
	);
	LUT3 #(
		.INIT('h09)
	) name8447 (
		_w14078_,
		_w14076_,
		_w14074_,
		_w14274_
	);
	LUT4 #(
		.INIT('hf7df)
	) name8448 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14275_
	);
	LUT3 #(
		.INIT('hb0)
	) name8449 (
		_w14273_,
		_w14274_,
		_w14275_,
		_w14276_
	);
	LUT4 #(
		.INIT('h3210)
	) name8450 (
		_w14073_,
		_w14272_,
		_w14276_,
		_w14269_,
		_w14277_
	);
	LUT2 #(
		.INIT('h9)
	) name8451 (
		\u2_L0_reg[17]/NET0131 ,
		_w14277_,
		_w14278_
	);
	LUT4 #(
		.INIT('h7343)
	) name8452 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14279_
	);
	LUT2 #(
		.INIT('h2)
	) name8453 (
		_w14014_,
		_w14279_,
		_w14280_
	);
	LUT4 #(
		.INIT('h1001)
	) name8454 (
		_w14014_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14281_
	);
	LUT4 #(
		.INIT('h8000)
	) name8455 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14282_
	);
	LUT3 #(
		.INIT('h01)
	) name8456 (
		_w14022_,
		_w14282_,
		_w14281_,
		_w14283_
	);
	LUT4 #(
		.INIT('h2000)
	) name8457 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14284_
	);
	LUT3 #(
		.INIT('h04)
	) name8458 (
		_w14014_,
		_w14016_,
		_w14018_,
		_w14285_
	);
	LUT4 #(
		.INIT('haa8a)
	) name8459 (
		_w14022_,
		_w14015_,
		_w14018_,
		_w14017_,
		_w14286_
	);
	LUT3 #(
		.INIT('h10)
	) name8460 (
		_w14284_,
		_w14285_,
		_w14286_,
		_w14287_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name8461 (
		_w14015_,
		_w14016_,
		_w14018_,
		_w14017_,
		_w14288_
	);
	LUT3 #(
		.INIT('h31)
	) name8462 (
		_w14014_,
		_w14148_,
		_w14288_,
		_w14289_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name8463 (
		_w14280_,
		_w14283_,
		_w14287_,
		_w14289_,
		_w14290_
	);
	LUT4 #(
		.INIT('hefcc)
	) name8464 (
		_w14014_,
		_w14015_,
		_w14019_,
		_w14038_,
		_w14291_
	);
	LUT3 #(
		.INIT('h65)
	) name8465 (
		\u2_L0_reg[19]/NET0131 ,
		_w14290_,
		_w14291_,
		_w14292_
	);
	LUT3 #(
		.INIT('h40)
	) name8466 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14293_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name8467 (
		_w14113_,
		_w14107_,
		_w14109_,
		_w14110_,
		_w14294_
	);
	LUT4 #(
		.INIT('h1000)
	) name8468 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14295_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name8469 (
		_w14113_,
		_w14107_,
		_w14109_,
		_w14110_,
		_w14296_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8470 (
		_w14293_,
		_w14294_,
		_w14295_,
		_w14296_,
		_w14297_
	);
	LUT4 #(
		.INIT('h7fd7)
	) name8471 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14298_
	);
	LUT3 #(
		.INIT('h45)
	) name8472 (
		_w14117_,
		_w14297_,
		_w14298_,
		_w14299_
	);
	LUT3 #(
		.INIT('hd0)
	) name8473 (
		_w14113_,
		_w14107_,
		_w14110_,
		_w14300_
	);
	LUT4 #(
		.INIT('h008a)
	) name8474 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14109_,
		_w14301_
	);
	LUT4 #(
		.INIT('h2000)
	) name8475 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14302_
	);
	LUT4 #(
		.INIT('hdaff)
	) name8476 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14303_
	);
	LUT4 #(
		.INIT('h20aa)
	) name8477 (
		_w14117_,
		_w14300_,
		_w14301_,
		_w14303_,
		_w14304_
	);
	LUT4 #(
		.INIT('h79ff)
	) name8478 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14305_
	);
	LUT2 #(
		.INIT('h2)
	) name8479 (
		_w14109_,
		_w14305_,
		_w14306_
	);
	LUT4 #(
		.INIT('hbbab)
	) name8480 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14307_
	);
	LUT2 #(
		.INIT('h8)
	) name8481 (
		_w14109_,
		_w14117_,
		_w14308_
	);
	LUT2 #(
		.INIT('h4)
	) name8482 (
		_w14307_,
		_w14308_,
		_w14309_
	);
	LUT4 #(
		.INIT('hccdf)
	) name8483 (
		_w14119_,
		_w14109_,
		_w14110_,
		_w14302_,
		_w14310_
	);
	LUT4 #(
		.INIT('h0100)
	) name8484 (
		_w14306_,
		_w14309_,
		_w14304_,
		_w14310_,
		_w14311_
	);
	LUT3 #(
		.INIT('h65)
	) name8485 (
		\u2_L0_reg[1]/NET0131 ,
		_w14299_,
		_w14311_,
		_w14312_
	);
	LUT4 #(
		.INIT('h02a0)
	) name8486 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14313_
	);
	LUT4 #(
		.INIT('h0100)
	) name8487 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14173_,
		_w14314_
	);
	LUT4 #(
		.INIT('h4000)
	) name8488 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14315_
	);
	LUT4 #(
		.INIT('h0040)
	) name8489 (
		_w14175_,
		_w14176_,
		_w14177_,
		_w14173_,
		_w14316_
	);
	LUT4 #(
		.INIT('h0002)
	) name8490 (
		_w14172_,
		_w14315_,
		_w14314_,
		_w14316_,
		_w14317_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name8491 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14318_
	);
	LUT4 #(
		.INIT('h5b59)
	) name8492 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14319_
	);
	LUT4 #(
		.INIT('h0010)
	) name8493 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14320_
	);
	LUT4 #(
		.INIT('h0501)
	) name8494 (
		_w14172_,
		_w14173_,
		_w14320_,
		_w14319_,
		_w14321_
	);
	LUT3 #(
		.INIT('h0b)
	) name8495 (
		_w14313_,
		_w14317_,
		_w14321_,
		_w14322_
	);
	LUT4 #(
		.INIT('h0009)
	) name8496 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14323_
	);
	LUT4 #(
		.INIT('h3010)
	) name8497 (
		_w14172_,
		_w14175_,
		_w14174_,
		_w14177_,
		_w14324_
	);
	LUT4 #(
		.INIT('h0200)
	) name8498 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14325_
	);
	LUT4 #(
		.INIT('h0001)
	) name8499 (
		_w14173_,
		_w14325_,
		_w14323_,
		_w14324_,
		_w14326_
	);
	LUT4 #(
		.INIT('h0004)
	) name8500 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14327_
	);
	LUT3 #(
		.INIT('h04)
	) name8501 (
		_w14194_,
		_w14173_,
		_w14327_,
		_w14328_
	);
	LUT2 #(
		.INIT('h1)
	) name8502 (
		_w14326_,
		_w14328_,
		_w14329_
	);
	LUT3 #(
		.INIT('h56)
	) name8503 (
		\u2_L0_reg[15]/NET0131 ,
		_w14322_,
		_w14329_,
		_w14330_
	);
	LUT4 #(
		.INIT('h00fb)
	) name8504 (
		_w14176_,
		_w14174_,
		_w14177_,
		_w14173_,
		_w14331_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8505 (
		_w14175_,
		_w14174_,
		_w14177_,
		_w14173_,
		_w14332_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name8506 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14333_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name8507 (
		_w14315_,
		_w14331_,
		_w14332_,
		_w14333_,
		_w14334_
	);
	LUT4 #(
		.INIT('h2100)
	) name8508 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14335_
	);
	LUT3 #(
		.INIT('h02)
	) name8509 (
		_w14172_,
		_w14327_,
		_w14335_,
		_w14336_
	);
	LUT2 #(
		.INIT('h4)
	) name8510 (
		_w14334_,
		_w14336_,
		_w14337_
	);
	LUT2 #(
		.INIT('h2)
	) name8511 (
		_w14176_,
		_w14173_,
		_w14338_
	);
	LUT3 #(
		.INIT('h73)
	) name8512 (
		_w14175_,
		_w14176_,
		_w14173_,
		_w14339_
	);
	LUT2 #(
		.INIT('h2)
	) name8513 (
		_w14180_,
		_w14339_,
		_w14340_
	);
	LUT3 #(
		.INIT('h51)
	) name8514 (
		_w14175_,
		_w14176_,
		_w14173_,
		_w14341_
	);
	LUT3 #(
		.INIT('h31)
	) name8515 (
		_w14181_,
		_w14178_,
		_w14341_,
		_w14342_
	);
	LUT4 #(
		.INIT('h8fdf)
	) name8516 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14343_
	);
	LUT2 #(
		.INIT('h2)
	) name8517 (
		_w14173_,
		_w14343_,
		_w14344_
	);
	LUT4 #(
		.INIT('h0002)
	) name8518 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14173_,
		_w14345_
	);
	LUT3 #(
		.INIT('h01)
	) name8519 (
		_w14172_,
		_w14190_,
		_w14345_,
		_w14346_
	);
	LUT4 #(
		.INIT('h1000)
	) name8520 (
		_w14344_,
		_w14340_,
		_w14346_,
		_w14342_,
		_w14347_
	);
	LUT4 #(
		.INIT('h0100)
	) name8521 (
		_w14175_,
		_w14174_,
		_w14177_,
		_w14173_,
		_w14348_
	);
	LUT3 #(
		.INIT('h13)
	) name8522 (
		_w14183_,
		_w14348_,
		_w14338_,
		_w14349_
	);
	LUT4 #(
		.INIT('ha955)
	) name8523 (
		\u2_L0_reg[21]/NET0131 ,
		_w14337_,
		_w14347_,
		_w14349_,
		_w14350_
	);
	LUT4 #(
		.INIT('h08c0)
	) name8524 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14351_
	);
	LUT4 #(
		.INIT('h00df)
	) name8525 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14241_,
		_w14352_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8526 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14241_,
		_w14353_
	);
	LUT4 #(
		.INIT('heaec)
	) name8527 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14354_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name8528 (
		_w14245_,
		_w14352_,
		_w14353_,
		_w14354_,
		_w14355_
	);
	LUT3 #(
		.INIT('ha8)
	) name8529 (
		_w14232_,
		_w14351_,
		_w14355_,
		_w14356_
	);
	LUT3 #(
		.INIT('h0e)
	) name8530 (
		_w14233_,
		_w14234_,
		_w14241_,
		_w14357_
	);
	LUT4 #(
		.INIT('h020f)
	) name8531 (
		_w14234_,
		_w14236_,
		_w14235_,
		_w14241_,
		_w14358_
	);
	LUT2 #(
		.INIT('h4)
	) name8532 (
		_w14357_,
		_w14358_,
		_w14359_
	);
	LUT4 #(
		.INIT('h4000)
	) name8533 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14360_
	);
	LUT3 #(
		.INIT('h31)
	) name8534 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14361_
	);
	LUT4 #(
		.INIT('h0073)
	) name8535 (
		_w14233_,
		_w14234_,
		_w14235_,
		_w14241_,
		_w14362_
	);
	LUT3 #(
		.INIT('h45)
	) name8536 (
		_w14360_,
		_w14361_,
		_w14362_,
		_w14363_
	);
	LUT4 #(
		.INIT('hf6ef)
	) name8537 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14364_
	);
	LUT4 #(
		.INIT('h0020)
	) name8538 (
		_w14233_,
		_w14234_,
		_w14235_,
		_w14241_,
		_w14365_
	);
	LUT4 #(
		.INIT('h0031)
	) name8539 (
		_w14241_,
		_w14240_,
		_w14364_,
		_w14365_,
		_w14366_
	);
	LUT4 #(
		.INIT('hba00)
	) name8540 (
		_w14232_,
		_w14359_,
		_w14363_,
		_w14366_,
		_w14367_
	);
	LUT3 #(
		.INIT('h65)
	) name8541 (
		\u2_L0_reg[25]/NET0131 ,
		_w14356_,
		_w14367_,
		_w14368_
	);
	LUT4 #(
		.INIT('h0092)
	) name8542 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14369_
	);
	LUT4 #(
		.INIT('heaee)
	) name8543 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14370_
	);
	LUT4 #(
		.INIT('h0504)
	) name8544 (
		_w14109_,
		_w14117_,
		_w14369_,
		_w14370_,
		_w14371_
	);
	LUT3 #(
		.INIT('h02)
	) name8545 (
		_w14109_,
		_w14121_,
		_w14130_,
		_w14372_
	);
	LUT2 #(
		.INIT('h1)
	) name8546 (
		_w14371_,
		_w14372_,
		_w14373_
	);
	LUT4 #(
		.INIT('h0004)
	) name8547 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14374_
	);
	LUT4 #(
		.INIT('h070f)
	) name8548 (
		_w14113_,
		_w14107_,
		_w14109_,
		_w14110_,
		_w14375_
	);
	LUT3 #(
		.INIT('h45)
	) name8549 (
		_w14124_,
		_w14374_,
		_w14375_,
		_w14376_
	);
	LUT4 #(
		.INIT('h2002)
	) name8550 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14377_
	);
	LUT2 #(
		.INIT('h1)
	) name8551 (
		_w14106_,
		_w14109_,
		_w14378_
	);
	LUT3 #(
		.INIT('h20)
	) name8552 (
		_w14113_,
		_w14107_,
		_w14110_,
		_w14379_
	);
	LUT4 #(
		.INIT('h2022)
	) name8553 (
		_w14117_,
		_w14377_,
		_w14378_,
		_w14379_,
		_w14380_
	);
	LUT2 #(
		.INIT('h8)
	) name8554 (
		_w14115_,
		_w14300_,
		_w14381_
	);
	LUT4 #(
		.INIT('hffa7)
	) name8555 (
		_w14106_,
		_w14113_,
		_w14107_,
		_w14110_,
		_w14382_
	);
	LUT3 #(
		.INIT('h10)
	) name8556 (
		_w14116_,
		_w14117_,
		_w14382_,
		_w14383_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8557 (
		_w14376_,
		_w14380_,
		_w14381_,
		_w14383_,
		_w14384_
	);
	LUT3 #(
		.INIT('h56)
	) name8558 (
		\u2_L0_reg[26]/NET0131 ,
		_w14373_,
		_w14384_,
		_w14385_
	);
	LUT4 #(
		.INIT('hc693)
	) name8559 (
		decrypt_pad,
		\u2_R0_reg[8]/NET0131 ,
		\u2_uk_K_r0_reg[25]/P0001 ,
		\u2_uk_K_r0_reg[46]/NET0131 ,
		_w14386_
	);
	LUT4 #(
		.INIT('hc693)
	) name8560 (
		decrypt_pad,
		\u2_R0_reg[7]/NET0131 ,
		\u2_uk_K_r0_reg[34]/NET0131 ,
		\u2_uk_K_r0_reg[55]/NET0131 ,
		_w14387_
	);
	LUT4 #(
		.INIT('hc693)
	) name8561 (
		decrypt_pad,
		\u2_R0_reg[6]/NET0131 ,
		\u2_uk_K_r0_reg[40]/NET0131 ,
		\u2_uk_K_r0_reg[4]/NET0131 ,
		_w14388_
	);
	LUT4 #(
		.INIT('hc693)
	) name8562 (
		decrypt_pad,
		\u2_R0_reg[4]/NET0131 ,
		\u2_uk_K_r0_reg[13]/NET0131 ,
		\u2_uk_K_r0_reg[34]/NET0131 ,
		_w14389_
	);
	LUT4 #(
		.INIT('hc963)
	) name8563 (
		decrypt_pad,
		\u2_R0_reg[9]/NET0131 ,
		\u2_uk_K_r0_reg[26]/NET0131 ,
		\u2_uk_K_r0_reg[5]/NET0131 ,
		_w14390_
	);
	LUT4 #(
		.INIT('hc963)
	) name8564 (
		decrypt_pad,
		\u2_R0_reg[5]/NET0131 ,
		\u2_uk_K_r0_reg[13]/NET0131 ,
		\u2_uk_K_r0_reg[17]/NET0131 ,
		_w14391_
	);
	LUT4 #(
		.INIT('h5a4f)
	) name8565 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14392_
	);
	LUT4 #(
		.INIT('hf5fc)
	) name8566 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14393_
	);
	LUT4 #(
		.INIT('hbf7b)
	) name8567 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14394_
	);
	LUT4 #(
		.INIT('hd800)
	) name8568 (
		_w14387_,
		_w14393_,
		_w14392_,
		_w14394_,
		_w14395_
	);
	LUT2 #(
		.INIT('h1)
	) name8569 (
		_w14386_,
		_w14395_,
		_w14396_
	);
	LUT4 #(
		.INIT('hfb7b)
	) name8570 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14397_
	);
	LUT2 #(
		.INIT('h1)
	) name8571 (
		_w14397_,
		_w14387_,
		_w14398_
	);
	LUT3 #(
		.INIT('h02)
	) name8572 (
		_w14391_,
		_w14389_,
		_w14390_,
		_w14399_
	);
	LUT4 #(
		.INIT('h5fa7)
	) name8573 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14400_
	);
	LUT2 #(
		.INIT('h2)
	) name8574 (
		_w14387_,
		_w14400_,
		_w14401_
	);
	LUT2 #(
		.INIT('h1)
	) name8575 (
		_w14387_,
		_w14393_,
		_w14402_
	);
	LUT4 #(
		.INIT('h0400)
	) name8576 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14403_
	);
	LUT3 #(
		.INIT('h0b)
	) name8577 (
		_w14391_,
		_w14390_,
		_w14387_,
		_w14404_
	);
	LUT2 #(
		.INIT('h4)
	) name8578 (
		_w14388_,
		_w14389_,
		_w14405_
	);
	LUT3 #(
		.INIT('h45)
	) name8579 (
		_w14403_,
		_w14404_,
		_w14405_,
		_w14406_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8580 (
		_w14386_,
		_w14401_,
		_w14402_,
		_w14406_,
		_w14407_
	);
	LUT4 #(
		.INIT('h5556)
	) name8581 (
		\u2_L0_reg[28]/NET0131 ,
		_w14398_,
		_w14407_,
		_w14396_,
		_w14408_
	);
	LUT4 #(
		.INIT('h0122)
	) name8582 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14409_
	);
	LUT4 #(
		.INIT('h0800)
	) name8583 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14410_
	);
	LUT4 #(
		.INIT('h0010)
	) name8584 (
		_w14391_,
		_w14388_,
		_w14390_,
		_w14387_,
		_w14411_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name8585 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14412_
	);
	LUT4 #(
		.INIT('h00bf)
	) name8586 (
		_w14391_,
		_w14389_,
		_w14390_,
		_w14387_,
		_w14413_
	);
	LUT4 #(
		.INIT('h1011)
	) name8587 (
		_w14410_,
		_w14411_,
		_w14412_,
		_w14413_,
		_w14414_
	);
	LUT3 #(
		.INIT('h45)
	) name8588 (
		_w14386_,
		_w14409_,
		_w14414_,
		_w14415_
	);
	LUT4 #(
		.INIT('h2010)
	) name8589 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14416_
	);
	LUT4 #(
		.INIT('ha200)
	) name8590 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14387_,
		_w14417_
	);
	LUT3 #(
		.INIT('ha8)
	) name8591 (
		_w14386_,
		_w14416_,
		_w14417_,
		_w14418_
	);
	LUT3 #(
		.INIT('h04)
	) name8592 (
		_w14391_,
		_w14388_,
		_w14390_,
		_w14419_
	);
	LUT4 #(
		.INIT('h0004)
	) name8593 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14420_
	);
	LUT4 #(
		.INIT('h4000)
	) name8594 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14421_
	);
	LUT4 #(
		.INIT('hdf00)
	) name8595 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14387_,
		_w14422_
	);
	LUT4 #(
		.INIT('h0b00)
	) name8596 (
		_w14386_,
		_w14421_,
		_w14420_,
		_w14422_,
		_w14423_
	);
	LUT4 #(
		.INIT('hbff2)
	) name8597 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14424_
	);
	LUT4 #(
		.INIT('h0900)
	) name8598 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14425_
	);
	LUT4 #(
		.INIT('h0051)
	) name8599 (
		_w14387_,
		_w14386_,
		_w14424_,
		_w14425_,
		_w14426_
	);
	LUT3 #(
		.INIT('h54)
	) name8600 (
		_w14418_,
		_w14423_,
		_w14426_,
		_w14427_
	);
	LUT3 #(
		.INIT('h65)
	) name8601 (
		\u2_L0_reg[2]/NET0131 ,
		_w14415_,
		_w14427_,
		_w14428_
	);
	LUT4 #(
		.INIT('h0002)
	) name8602 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14429_
	);
	LUT4 #(
		.INIT('h4050)
	) name8603 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14430_
	);
	LUT4 #(
		.INIT('hf351)
	) name8604 (
		_w14352_,
		_w14353_,
		_w14429_,
		_w14430_,
		_w14431_
	);
	LUT4 #(
		.INIT('hf6bb)
	) name8605 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14432_
	);
	LUT3 #(
		.INIT('h45)
	) name8606 (
		_w14232_,
		_w14431_,
		_w14432_,
		_w14433_
	);
	LUT4 #(
		.INIT('h0200)
	) name8607 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14434_
	);
	LUT4 #(
		.INIT('hf3bf)
	) name8608 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14435_
	);
	LUT4 #(
		.INIT('hd8fa)
	) name8609 (
		_w14241_,
		_w14260_,
		_w14434_,
		_w14435_,
		_w14436_
	);
	LUT4 #(
		.INIT('hdfde)
	) name8610 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14437_
	);
	LUT3 #(
		.INIT('h02)
	) name8611 (
		_w14233_,
		_w14235_,
		_w14241_,
		_w14438_
	);
	LUT4 #(
		.INIT('h00c4)
	) name8612 (
		_w14241_,
		_w14261_,
		_w14437_,
		_w14438_,
		_w14439_
	);
	LUT3 #(
		.INIT('h31)
	) name8613 (
		_w14232_,
		_w14436_,
		_w14439_,
		_w14440_
	);
	LUT3 #(
		.INIT('h65)
	) name8614 (
		\u2_L0_reg[8]/NET0131 ,
		_w14433_,
		_w14440_,
		_w14441_
	);
	LUT3 #(
		.INIT('h01)
	) name8615 (
		_w14391_,
		_w14388_,
		_w14390_,
		_w14442_
	);
	LUT4 #(
		.INIT('hdf00)
	) name8616 (
		_w14388_,
		_w14389_,
		_w14390_,
		_w14387_,
		_w14443_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8617 (
		_w14419_,
		_w14413_,
		_w14442_,
		_w14443_,
		_w14444_
	);
	LUT4 #(
		.INIT('h0002)
	) name8618 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14445_
	);
	LUT4 #(
		.INIT('h0002)
	) name8619 (
		_w14386_,
		_w14410_,
		_w14411_,
		_w14445_,
		_w14446_
	);
	LUT4 #(
		.INIT('h0600)
	) name8620 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14447_
	);
	LUT4 #(
		.INIT('h0010)
	) name8621 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14448_
	);
	LUT2 #(
		.INIT('h1)
	) name8622 (
		_w14387_,
		_w14386_,
		_w14449_
	);
	LUT4 #(
		.INIT('h0100)
	) name8623 (
		_w14399_,
		_w14448_,
		_w14447_,
		_w14449_,
		_w14450_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name8624 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14451_
	);
	LUT4 #(
		.INIT('hf400)
	) name8625 (
		_w14444_,
		_w14446_,
		_w14450_,
		_w14451_,
		_w14452_
	);
	LUT4 #(
		.INIT('h1321)
	) name8626 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14453_
	);
	LUT4 #(
		.INIT('hc044)
	) name8627 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14454_
	);
	LUT2 #(
		.INIT('h2)
	) name8628 (
		_w14387_,
		_w14386_,
		_w14455_
	);
	LUT3 #(
		.INIT('h10)
	) name8629 (
		_w14453_,
		_w14454_,
		_w14455_,
		_w14456_
	);
	LUT3 #(
		.INIT('h56)
	) name8630 (
		\u2_L0_reg[13]/NET0131 ,
		_w14452_,
		_w14456_,
		_w14457_
	);
	LUT4 #(
		.INIT('hf73f)
	) name8631 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14458_
	);
	LUT2 #(
		.INIT('h2)
	) name8632 (
		_w14074_,
		_w14458_,
		_w14459_
	);
	LUT3 #(
		.INIT('h07)
	) name8633 (
		_w14091_,
		_w14099_,
		_w14264_,
		_w14460_
	);
	LUT3 #(
		.INIT('h8a)
	) name8634 (
		_w14073_,
		_w14459_,
		_w14460_,
		_w14461_
	);
	LUT4 #(
		.INIT('h7bef)
	) name8635 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14462_
	);
	LUT2 #(
		.INIT('h1)
	) name8636 (
		_w14074_,
		_w14462_,
		_w14463_
	);
	LUT3 #(
		.INIT('h01)
	) name8637 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14464_
	);
	LUT3 #(
		.INIT('h01)
	) name8638 (
		_w14082_,
		_w14101_,
		_w14464_,
		_w14465_
	);
	LUT3 #(
		.INIT('h02)
	) name8639 (
		_w14077_,
		_w14078_,
		_w14076_,
		_w14466_
	);
	LUT4 #(
		.INIT('h0200)
	) name8640 (
		_w14077_,
		_w14078_,
		_w14076_,
		_w14074_,
		_w14467_
	);
	LUT3 #(
		.INIT('hec)
	) name8641 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14468_
	);
	LUT3 #(
		.INIT('h13)
	) name8642 (
		_w14096_,
		_w14467_,
		_w14468_,
		_w14469_
	);
	LUT3 #(
		.INIT('had)
	) name8643 (
		_w14077_,
		_w14078_,
		_w14076_,
		_w14470_
	);
	LUT4 #(
		.INIT('hfdc3)
	) name8644 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14471_
	);
	LUT2 #(
		.INIT('h2)
	) name8645 (
		_w14073_,
		_w14074_,
		_w14472_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name8646 (
		_w14087_,
		_w14470_,
		_w14471_,
		_w14472_,
		_w14473_
	);
	LUT4 #(
		.INIT('hea00)
	) name8647 (
		_w14073_,
		_w14465_,
		_w14469_,
		_w14473_,
		_w14474_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name8648 (
		\u2_L0_reg[23]/NET0131 ,
		_w14463_,
		_w14461_,
		_w14474_,
		_w14475_
	);
	LUT4 #(
		.INIT('hd7d2)
	) name8649 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14476_
	);
	LUT2 #(
		.INIT('h1)
	) name8650 (
		_w14173_,
		_w14476_,
		_w14477_
	);
	LUT3 #(
		.INIT('hb0)
	) name8651 (
		_w14176_,
		_w14174_,
		_w14173_,
		_w14478_
	);
	LUT4 #(
		.INIT('he7bb)
	) name8652 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14479_
	);
	LUT3 #(
		.INIT('hb0)
	) name8653 (
		_w14318_,
		_w14478_,
		_w14479_,
		_w14480_
	);
	LUT3 #(
		.INIT('h8a)
	) name8654 (
		_w14172_,
		_w14477_,
		_w14480_,
		_w14481_
	);
	LUT4 #(
		.INIT('hce44)
	) name8655 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14482_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8656 (
		_w14175_,
		_w14176_,
		_w14177_,
		_w14173_,
		_w14483_
	);
	LUT2 #(
		.INIT('h4)
	) name8657 (
		_w14482_,
		_w14483_,
		_w14484_
	);
	LUT4 #(
		.INIT('h0080)
	) name8658 (
		_w14176_,
		_w14174_,
		_w14177_,
		_w14173_,
		_w14485_
	);
	LUT3 #(
		.INIT('h01)
	) name8659 (
		_w14191_,
		_w14345_,
		_w14485_,
		_w14486_
	);
	LUT4 #(
		.INIT('h1000)
	) name8660 (
		_w14175_,
		_w14176_,
		_w14177_,
		_w14173_,
		_w14487_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name8661 (
		_w14175_,
		_w14176_,
		_w14174_,
		_w14177_,
		_w14488_
	);
	LUT3 #(
		.INIT('h32)
	) name8662 (
		_w14173_,
		_w14487_,
		_w14488_,
		_w14489_
	);
	LUT4 #(
		.INIT('hba00)
	) name8663 (
		_w14172_,
		_w14484_,
		_w14486_,
		_w14489_,
		_w14490_
	);
	LUT3 #(
		.INIT('h65)
	) name8664 (
		\u2_L0_reg[27]/NET0131 ,
		_w14481_,
		_w14490_,
		_w14491_
	);
	LUT3 #(
		.INIT('h40)
	) name8665 (
		_w14047_,
		_w14048_,
		_w14049_,
		_w14492_
	);
	LUT4 #(
		.INIT('hdee3)
	) name8666 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14493_
	);
	LUT2 #(
		.INIT('h1)
	) name8667 (
		_w14056_,
		_w14493_,
		_w14494_
	);
	LUT3 #(
		.INIT('h08)
	) name8668 (
		_w14046_,
		_w14048_,
		_w14049_,
		_w14495_
	);
	LUT4 #(
		.INIT('hbbfc)
	) name8669 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14496_
	);
	LUT4 #(
		.INIT('h1f13)
	) name8670 (
		_w14047_,
		_w14056_,
		_w14495_,
		_w14496_,
		_w14497_
	);
	LUT3 #(
		.INIT('h8a)
	) name8671 (
		_w14054_,
		_w14494_,
		_w14497_,
		_w14498_
	);
	LUT4 #(
		.INIT('hab89)
	) name8672 (
		_w14056_,
		_w14223_,
		_w14226_,
		_w14492_,
		_w14499_
	);
	LUT4 #(
		.INIT('h7db7)
	) name8673 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14500_
	);
	LUT4 #(
		.INIT('h00a2)
	) name8674 (
		_w14047_,
		_w14048_,
		_w14049_,
		_w14056_,
		_w14501_
	);
	LUT4 #(
		.INIT('h0777)
	) name8675 (
		_w14051_,
		_w14056_,
		_w14060_,
		_w14501_,
		_w14502_
	);
	LUT4 #(
		.INIT('hba00)
	) name8676 (
		_w14054_,
		_w14499_,
		_w14500_,
		_w14502_,
		_w14503_
	);
	LUT3 #(
		.INIT('h65)
	) name8677 (
		\u2_L0_reg[32]/NET0131 ,
		_w14498_,
		_w14503_,
		_w14504_
	);
	LUT3 #(
		.INIT('h04)
	) name8678 (
		_w14233_,
		_w14236_,
		_w14235_,
		_w14505_
	);
	LUT4 #(
		.INIT('hf700)
	) name8679 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14241_,
		_w14506_
	);
	LUT4 #(
		.INIT('h7077)
	) name8680 (
		_w14237_,
		_w14352_,
		_w14505_,
		_w14506_,
		_w14507_
	);
	LUT4 #(
		.INIT('h3100)
	) name8681 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14508_
	);
	LUT2 #(
		.INIT('h1)
	) name8682 (
		_w14232_,
		_w14508_,
		_w14509_
	);
	LUT4 #(
		.INIT('hfb5b)
	) name8683 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14510_
	);
	LUT2 #(
		.INIT('h2)
	) name8684 (
		_w14241_,
		_w14510_,
		_w14511_
	);
	LUT4 #(
		.INIT('h0040)
	) name8685 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14241_,
		_w14512_
	);
	LUT4 #(
		.INIT('h0002)
	) name8686 (
		_w14232_,
		_w14240_,
		_w14434_,
		_w14512_,
		_w14513_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8687 (
		_w14507_,
		_w14509_,
		_w14511_,
		_w14513_,
		_w14514_
	);
	LUT3 #(
		.INIT('h02)
	) name8688 (
		_w14241_,
		_w14260_,
		_w14429_,
		_w14515_
	);
	LUT4 #(
		.INIT('hfff6)
	) name8689 (
		_w14233_,
		_w14234_,
		_w14236_,
		_w14235_,
		_w14516_
	);
	LUT3 #(
		.INIT('he0)
	) name8690 (
		_w14251_,
		_w14352_,
		_w14516_,
		_w14517_
	);
	LUT2 #(
		.INIT('h1)
	) name8691 (
		_w14515_,
		_w14517_,
		_w14518_
	);
	LUT3 #(
		.INIT('h56)
	) name8692 (
		\u2_L0_reg[3]/NET0131 ,
		_w14514_,
		_w14518_,
		_w14519_
	);
	LUT4 #(
		.INIT('hc693)
	) name8693 (
		decrypt_pad,
		\u2_R0_reg[11]/P0001 ,
		\u2_uk_K_r0_reg[20]/NET0131 ,
		\u2_uk_K_r0_reg[41]/NET0131 ,
		_w14520_
	);
	LUT4 #(
		.INIT('hc963)
	) name8694 (
		decrypt_pad,
		\u2_R0_reg[12]/NET0131 ,
		\u2_uk_K_r0_reg[24]/P0001 ,
		\u2_uk_K_r0_reg[3]/NET0131 ,
		_w14521_
	);
	LUT4 #(
		.INIT('hc963)
	) name8695 (
		decrypt_pad,
		\u2_R0_reg[13]/NET0131 ,
		\u2_uk_K_r0_reg[12]/NET0131 ,
		\u2_uk_K_r0_reg[48]/NET0131 ,
		_w14522_
	);
	LUT4 #(
		.INIT('hc693)
	) name8696 (
		decrypt_pad,
		\u2_R0_reg[9]/NET0131 ,
		\u2_uk_K_r0_reg[11]/NET0131 ,
		\u2_uk_K_r0_reg[32]/NET0131 ,
		_w14523_
	);
	LUT4 #(
		.INIT('hc693)
	) name8697 (
		decrypt_pad,
		\u2_R0_reg[8]/NET0131 ,
		\u2_uk_K_r0_reg[39]/NET0131 ,
		\u2_uk_K_r0_reg[3]/NET0131 ,
		_w14524_
	);
	LUT2 #(
		.INIT('h6)
	) name8698 (
		_w14522_,
		_w14524_,
		_w14525_
	);
	LUT4 #(
		.INIT('hc693)
	) name8699 (
		decrypt_pad,
		\u2_R0_reg[10]/NET0131 ,
		\u2_uk_K_r0_reg[19]/NET0131 ,
		\u2_uk_K_r0_reg[40]/NET0131 ,
		_w14526_
	);
	LUT4 #(
		.INIT('hc733)
	) name8700 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14527_
	);
	LUT2 #(
		.INIT('h1)
	) name8701 (
		_w14526_,
		_w14523_,
		_w14528_
	);
	LUT4 #(
		.INIT('h0001)
	) name8702 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14529_
	);
	LUT4 #(
		.INIT('hff76)
	) name8703 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14530_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8704 (
		_w14521_,
		_w14520_,
		_w14527_,
		_w14530_,
		_w14531_
	);
	LUT3 #(
		.INIT('h20)
	) name8705 (
		_w14522_,
		_w14524_,
		_w14523_,
		_w14532_
	);
	LUT2 #(
		.INIT('h2)
	) name8706 (
		_w14526_,
		_w14520_,
		_w14533_
	);
	LUT4 #(
		.INIT('h2000)
	) name8707 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14534_
	);
	LUT4 #(
		.INIT('hdf7d)
	) name8708 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14535_
	);
	LUT3 #(
		.INIT('h70)
	) name8709 (
		_w14532_,
		_w14533_,
		_w14535_,
		_w14536_
	);
	LUT2 #(
		.INIT('h8)
	) name8710 (
		_w14522_,
		_w14520_,
		_w14537_
	);
	LUT3 #(
		.INIT('h46)
	) name8711 (
		_w14522_,
		_w14524_,
		_w14520_,
		_w14538_
	);
	LUT2 #(
		.INIT('h8)
	) name8712 (
		_w14538_,
		_w14528_,
		_w14539_
	);
	LUT3 #(
		.INIT('heb)
	) name8713 (
		_w14526_,
		_w14523_,
		_w14538_,
		_w14540_
	);
	LUT2 #(
		.INIT('h8)
	) name8714 (
		_w14521_,
		_w14526_,
		_w14541_
	);
	LUT3 #(
		.INIT('h10)
	) name8715 (
		_w14522_,
		_w14524_,
		_w14523_,
		_w14542_
	);
	LUT2 #(
		.INIT('h2)
	) name8716 (
		_w14521_,
		_w14520_,
		_w14543_
	);
	LUT3 #(
		.INIT('h80)
	) name8717 (
		_w14522_,
		_w14524_,
		_w14523_,
		_w14544_
	);
	LUT4 #(
		.INIT('h3bcf)
	) name8718 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14545_
	);
	LUT4 #(
		.INIT('h7707)
	) name8719 (
		_w14541_,
		_w14542_,
		_w14543_,
		_w14545_,
		_w14546_
	);
	LUT4 #(
		.INIT('hea00)
	) name8720 (
		_w14521_,
		_w14536_,
		_w14540_,
		_w14546_,
		_w14547_
	);
	LUT3 #(
		.INIT('h65)
	) name8721 (
		\u2_L0_reg[6]/NET0131 ,
		_w14531_,
		_w14547_,
		_w14548_
	);
	LUT3 #(
		.INIT('h28)
	) name8722 (
		_w14047_,
		_w14048_,
		_w14049_,
		_w14549_
	);
	LUT4 #(
		.INIT('h2880)
	) name8723 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14550_
	);
	LUT4 #(
		.INIT('h5004)
	) name8724 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14551_
	);
	LUT2 #(
		.INIT('h2)
	) name8725 (
		_w14056_,
		_w14551_,
		_w14552_
	);
	LUT3 #(
		.INIT('h09)
	) name8726 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14553_
	);
	LUT4 #(
		.INIT('h00f7)
	) name8727 (
		_w14046_,
		_w14048_,
		_w14049_,
		_w14056_,
		_w14554_
	);
	LUT3 #(
		.INIT('h10)
	) name8728 (
		_w14549_,
		_w14553_,
		_w14554_,
		_w14555_
	);
	LUT4 #(
		.INIT('h888a)
	) name8729 (
		_w14054_,
		_w14550_,
		_w14552_,
		_w14555_,
		_w14556_
	);
	LUT4 #(
		.INIT('h5150)
	) name8730 (
		_w14054_,
		_w14056_,
		_w14061_,
		_w14551_,
		_w14557_
	);
	LUT4 #(
		.INIT('h7885)
	) name8731 (
		_w14046_,
		_w14047_,
		_w14048_,
		_w14049_,
		_w14558_
	);
	LUT4 #(
		.INIT('h00c4)
	) name8732 (
		_w14054_,
		_w14056_,
		_w14061_,
		_w14558_,
		_w14559_
	);
	LUT2 #(
		.INIT('h4)
	) name8733 (
		_w14056_,
		_w14550_,
		_w14560_
	);
	LUT3 #(
		.INIT('h01)
	) name8734 (
		_w14559_,
		_w14560_,
		_w14557_,
		_w14561_
	);
	LUT3 #(
		.INIT('h65)
	) name8735 (
		\u2_L0_reg[7]/NET0131 ,
		_w14556_,
		_w14561_,
		_w14562_
	);
	LUT4 #(
		.INIT('h0002)
	) name8736 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14563_
	);
	LUT3 #(
		.INIT('h12)
	) name8737 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14564_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8738 (
		_w14520_,
		_w14534_,
		_w14563_,
		_w14564_,
		_w14565_
	);
	LUT3 #(
		.INIT('h0d)
	) name8739 (
		_w14522_,
		_w14524_,
		_w14523_,
		_w14566_
	);
	LUT3 #(
		.INIT('h70)
	) name8740 (
		_w14522_,
		_w14524_,
		_w14523_,
		_w14567_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name8741 (
		_w14522_,
		_w14524_,
		_w14523_,
		_w14520_,
		_w14568_
	);
	LUT4 #(
		.INIT('hf7ef)
	) name8742 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14569_
	);
	LUT3 #(
		.INIT('he0)
	) name8743 (
		_w14526_,
		_w14568_,
		_w14569_,
		_w14570_
	);
	LUT3 #(
		.INIT('h8a)
	) name8744 (
		_w14521_,
		_w14565_,
		_w14570_,
		_w14571_
	);
	LUT3 #(
		.INIT('h08)
	) name8745 (
		_w14526_,
		_w14524_,
		_w14523_,
		_w14572_
	);
	LUT4 #(
		.INIT('h00f7)
	) name8746 (
		_w14526_,
		_w14524_,
		_w14523_,
		_w14520_,
		_w14573_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name8747 (
		_w14520_,
		_w14534_,
		_w14573_,
		_w14563_,
		_w14574_
	);
	LUT4 #(
		.INIT('h3ef2)
	) name8748 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14575_
	);
	LUT3 #(
		.INIT('he0)
	) name8749 (
		_w14522_,
		_w14524_,
		_w14520_,
		_w14576_
	);
	LUT4 #(
		.INIT('h6800)
	) name8750 (
		_w14522_,
		_w14524_,
		_w14523_,
		_w14520_,
		_w14577_
	);
	LUT4 #(
		.INIT('h0302)
	) name8751 (
		_w14520_,
		_w14529_,
		_w14577_,
		_w14575_,
		_w14578_
	);
	LUT3 #(
		.INIT('h32)
	) name8752 (
		_w14521_,
		_w14574_,
		_w14578_,
		_w14579_
	);
	LUT3 #(
		.INIT('h65)
	) name8753 (
		\u2_L0_reg[16]/NET0131 ,
		_w14571_,
		_w14579_,
		_w14580_
	);
	LUT4 #(
		.INIT('hf859)
	) name8754 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14581_
	);
	LUT4 #(
		.INIT('h0020)
	) name8755 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14582_
	);
	LUT4 #(
		.INIT('h5504)
	) name8756 (
		_w14521_,
		_w14520_,
		_w14581_,
		_w14582_,
		_w14583_
	);
	LUT4 #(
		.INIT('hc7b6)
	) name8757 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14584_
	);
	LUT3 #(
		.INIT('h54)
	) name8758 (
		_w14521_,
		_w14520_,
		_w14584_,
		_w14585_
	);
	LUT2 #(
		.INIT('h4)
	) name8759 (
		_w14526_,
		_w14520_,
		_w14586_
	);
	LUT3 #(
		.INIT('h2a)
	) name8760 (
		_w14521_,
		_w14566_,
		_w14586_,
		_w14587_
	);
	LUT3 #(
		.INIT('ha2)
	) name8761 (
		_w14526_,
		_w14524_,
		_w14523_,
		_w14588_
	);
	LUT3 #(
		.INIT('h0e)
	) name8762 (
		_w14526_,
		_w14523_,
		_w14520_,
		_w14589_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name8763 (
		_w14525_,
		_w14576_,
		_w14588_,
		_w14589_,
		_w14590_
	);
	LUT4 #(
		.INIT('h2333)
	) name8764 (
		_w14539_,
		_w14585_,
		_w14587_,
		_w14590_,
		_w14591_
	);
	LUT3 #(
		.INIT('hdb)
	) name8765 (
		_w14522_,
		_w14524_,
		_w14523_,
		_w14592_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name8766 (
		_w14526_,
		_w14520_,
		_w14544_,
		_w14592_,
		_w14593_
	);
	LUT4 #(
		.INIT('h5655)
	) name8767 (
		\u2_L0_reg[24]/NET0131 ,
		_w14591_,
		_w14583_,
		_w14593_,
		_w14594_
	);
	LUT4 #(
		.INIT('hf9e9)
	) name8768 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14595_
	);
	LUT3 #(
		.INIT('h20)
	) name8769 (
		_w14526_,
		_w14522_,
		_w14523_,
		_w14596_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name8770 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14597_
	);
	LUT4 #(
		.INIT('hddd8)
	) name8771 (
		_w14521_,
		_w14595_,
		_w14597_,
		_w14596_,
		_w14598_
	);
	LUT2 #(
		.INIT('h2)
	) name8772 (
		_w14520_,
		_w14598_,
		_w14599_
	);
	LUT3 #(
		.INIT('h0e)
	) name8773 (
		_w14524_,
		_w14523_,
		_w14520_,
		_w14600_
	);
	LUT4 #(
		.INIT('hffb6)
	) name8774 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14601_
	);
	LUT4 #(
		.INIT('h4055)
	) name8775 (
		_w14521_,
		_w14597_,
		_w14600_,
		_w14601_,
		_w14602_
	);
	LUT4 #(
		.INIT('h5c5f)
	) name8776 (
		_w14526_,
		_w14522_,
		_w14524_,
		_w14523_,
		_w14603_
	);
	LUT2 #(
		.INIT('h2)
	) name8777 (
		_w14543_,
		_w14603_,
		_w14604_
	);
	LUT2 #(
		.INIT('h8)
	) name8778 (
		_w14541_,
		_w14567_,
		_w14605_
	);
	LUT4 #(
		.INIT('h0020)
	) name8779 (
		_w14526_,
		_w14522_,
		_w14523_,
		_w14520_,
		_w14606_
	);
	LUT3 #(
		.INIT('h07)
	) name8780 (
		_w14537_,
		_w14572_,
		_w14606_,
		_w14607_
	);
	LUT4 #(
		.INIT('h0100)
	) name8781 (
		_w14602_,
		_w14604_,
		_w14605_,
		_w14607_,
		_w14608_
	);
	LUT3 #(
		.INIT('h9a)
	) name8782 (
		\u2_L0_reg[30]/NET0131 ,
		_w14599_,
		_w14608_,
		_w14609_
	);
	LUT4 #(
		.INIT('h8228)
	) name8783 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14610_
	);
	LUT3 #(
		.INIT('he6)
	) name8784 (
		_w14077_,
		_w14078_,
		_w14076_,
		_w14611_
	);
	LUT4 #(
		.INIT('h0031)
	) name8785 (
		_w14087_,
		_w14267_,
		_w14611_,
		_w14610_,
		_w14612_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name8786 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14613_
	);
	LUT2 #(
		.INIT('h1)
	) name8787 (
		_w14074_,
		_w14613_,
		_w14614_
	);
	LUT4 #(
		.INIT('h00e6)
	) name8788 (
		_w14077_,
		_w14078_,
		_w14076_,
		_w14074_,
		_w14615_
	);
	LUT4 #(
		.INIT('hc700)
	) name8789 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14074_,
		_w14616_
	);
	LUT4 #(
		.INIT('h9ffd)
	) name8790 (
		_w14075_,
		_w14077_,
		_w14078_,
		_w14076_,
		_w14617_
	);
	LUT4 #(
		.INIT('hdc00)
	) name8791 (
		_w14466_,
		_w14615_,
		_w14616_,
		_w14617_,
		_w14618_
	);
	LUT4 #(
		.INIT('h3210)
	) name8792 (
		_w14073_,
		_w14614_,
		_w14618_,
		_w14612_,
		_w14619_
	);
	LUT2 #(
		.INIT('h9)
	) name8793 (
		\u2_L0_reg[9]/NET0131 ,
		_w14619_,
		_w14620_
	);
	LUT4 #(
		.INIT('h1a00)
	) name8794 (
		_w14391_,
		_w14389_,
		_w14390_,
		_w14387_,
		_w14621_
	);
	LUT4 #(
		.INIT('hcfaf)
	) name8795 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14622_
	);
	LUT4 #(
		.INIT('h0032)
	) name8796 (
		_w14387_,
		_w14420_,
		_w14622_,
		_w14621_,
		_w14623_
	);
	LUT4 #(
		.INIT('hbf6e)
	) name8797 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14624_
	);
	LUT4 #(
		.INIT('h8000)
	) name8798 (
		_w14391_,
		_w14389_,
		_w14390_,
		_w14387_,
		_w14625_
	);
	LUT4 #(
		.INIT('h0109)
	) name8799 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14387_,
		_w14626_
	);
	LUT3 #(
		.INIT('h10)
	) name8800 (
		_w14625_,
		_w14626_,
		_w14624_,
		_w14627_
	);
	LUT4 #(
		.INIT('h0020)
	) name8801 (
		_w14391_,
		_w14389_,
		_w14390_,
		_w14387_,
		_w14628_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name8802 (
		_w14391_,
		_w14388_,
		_w14389_,
		_w14390_,
		_w14629_
	);
	LUT3 #(
		.INIT('h31)
	) name8803 (
		_w14387_,
		_w14628_,
		_w14629_,
		_w14630_
	);
	LUT4 #(
		.INIT('hd800)
	) name8804 (
		_w14386_,
		_w14623_,
		_w14627_,
		_w14630_,
		_w14631_
	);
	LUT2 #(
		.INIT('h9)
	) name8805 (
		\u2_L0_reg[18]/P0001 ,
		_w14631_,
		_w14632_
	);
	LUT4 #(
		.INIT('hc693)
	) name8806 (
		decrypt_pad,
		\u1_R1_reg[20]/NET0131 ,
		\u1_uk_K_r1_reg[44]/P0001 ,
		\u1_uk_K_r1_reg[50]/NET0131 ,
		_w14633_
	);
	LUT4 #(
		.INIT('hc693)
	) name8807 (
		decrypt_pad,
		\u1_R1_reg[19]/NET0131 ,
		\u1_uk_K_r1_reg[29]/NET0131 ,
		\u1_uk_K_r1_reg[35]/NET0131 ,
		_w14634_
	);
	LUT4 #(
		.INIT('hc693)
	) name8808 (
		decrypt_pad,
		\u1_R1_reg[18]/NET0131 ,
		\u1_uk_K_r1_reg[42]/NET0131 ,
		\u1_uk_K_r1_reg[52]/NET0131 ,
		_w14635_
	);
	LUT4 #(
		.INIT('hc693)
	) name8809 (
		decrypt_pad,
		\u1_R1_reg[16]/NET0131 ,
		\u1_uk_K_r1_reg[2]/NET0131 ,
		\u1_uk_K_r1_reg[8]/NET0131 ,
		_w14636_
	);
	LUT4 #(
		.INIT('hc693)
	) name8810 (
		decrypt_pad,
		\u1_R1_reg[21]/NET0131 ,
		\u1_uk_K_r1_reg[14]/NET0131 ,
		\u1_uk_K_r1_reg[51]/NET0131 ,
		_w14637_
	);
	LUT4 #(
		.INIT('hc963)
	) name8811 (
		decrypt_pad,
		\u1_R1_reg[17]/NET0131 ,
		\u1_uk_K_r1_reg[30]/NET0131 ,
		\u1_uk_K_r1_reg[52]/NET0131 ,
		_w14638_
	);
	LUT4 #(
		.INIT('h3ed0)
	) name8812 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w14639_
	);
	LUT4 #(
		.INIT('hf3af)
	) name8813 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w14640_
	);
	LUT4 #(
		.INIT('h9fbf)
	) name8814 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w14641_
	);
	LUT4 #(
		.INIT('hd800)
	) name8815 (
		_w14634_,
		_w14639_,
		_w14640_,
		_w14641_,
		_w14642_
	);
	LUT2 #(
		.INIT('h2)
	) name8816 (
		_w14633_,
		_w14642_,
		_w14643_
	);
	LUT4 #(
		.INIT('hdff9)
	) name8817 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w14644_
	);
	LUT2 #(
		.INIT('h2)
	) name8818 (
		_w14634_,
		_w14644_,
		_w14645_
	);
	LUT4 #(
		.INIT('hfc5f)
	) name8819 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w14646_
	);
	LUT2 #(
		.INIT('h4)
	) name8820 (
		_w14637_,
		_w14634_,
		_w14647_
	);
	LUT3 #(
		.INIT('hb0)
	) name8821 (
		_w14637_,
		_w14638_,
		_w14634_,
		_w14648_
	);
	LUT4 #(
		.INIT('h5051)
	) name8822 (
		_w14635_,
		_w14638_,
		_w14634_,
		_w14636_,
		_w14649_
	);
	LUT4 #(
		.INIT('he0ee)
	) name8823 (
		_w14646_,
		_w14647_,
		_w14648_,
		_w14649_,
		_w14650_
	);
	LUT4 #(
		.INIT('h0200)
	) name8824 (
		_w14635_,
		_w14638_,
		_w14634_,
		_w14636_,
		_w14651_
	);
	LUT4 #(
		.INIT('h4000)
	) name8825 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w14652_
	);
	LUT2 #(
		.INIT('h1)
	) name8826 (
		_w14651_,
		_w14652_,
		_w14653_
	);
	LUT4 #(
		.INIT('h0e00)
	) name8827 (
		_w14633_,
		_w14650_,
		_w14645_,
		_w14653_,
		_w14654_
	);
	LUT3 #(
		.INIT('h65)
	) name8828 (
		\u1_L1_reg[25]/NET0131 ,
		_w14643_,
		_w14654_,
		_w14655_
	);
	LUT4 #(
		.INIT('hc693)
	) name8829 (
		decrypt_pad,
		\u2_desIn_r_reg[25]/NET0131 ,
		\u2_key_r_reg[35]/P0001 ,
		\u2_key_r_reg[42]/P0001 ,
		_w14656_
	);
	LUT4 #(
		.INIT('hc963)
	) name8830 (
		decrypt_pad,
		\u2_desIn_r_reg[17]/NET0131 ,
		\u2_key_r_reg[0]/NET0131 ,
		\u2_key_r_reg[52]/NET0131 ,
		_w14657_
	);
	LUT4 #(
		.INIT('hc693)
	) name8831 (
		decrypt_pad,
		\u2_desIn_r_reg[9]/NET0131 ,
		\u2_key_r_reg[15]/NET0131 ,
		\u2_key_r_reg[22]/NET0131 ,
		_w14658_
	);
	LUT4 #(
		.INIT('hc693)
	) name8832 (
		decrypt_pad,
		\u2_desIn_r_reg[33]/NET0131 ,
		\u2_key_r_reg[31]/NET0131 ,
		\u2_key_r_reg[38]/NET0131 ,
		_w14659_
	);
	LUT4 #(
		.INIT('hc963)
	) name8833 (
		decrypt_pad,
		\u2_desIn_r_reg[59]/NET0131 ,
		\u2_key_r_reg[2]/NET0131 ,
		\u2_key_r_reg[50]/NET0131 ,
		_w14660_
	);
	LUT4 #(
		.INIT('hc693)
	) name8834 (
		decrypt_pad,
		\u2_desIn_r_reg[1]/NET0131 ,
		\u2_key_r_reg[30]/NET0131 ,
		\u2_key_r_reg[37]/NET0131 ,
		_w14661_
	);
	LUT4 #(
		.INIT('h0008)
	) name8835 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14662_
	);
	LUT2 #(
		.INIT('h2)
	) name8836 (
		_w14659_,
		_w14660_,
		_w14663_
	);
	LUT4 #(
		.INIT('hddf7)
	) name8837 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14664_
	);
	LUT2 #(
		.INIT('h1)
	) name8838 (
		_w14657_,
		_w14664_,
		_w14665_
	);
	LUT3 #(
		.INIT('hd3)
	) name8839 (
		_w14659_,
		_w14658_,
		_w14661_,
		_w14666_
	);
	LUT2 #(
		.INIT('h8)
	) name8840 (
		_w14660_,
		_w14657_,
		_w14667_
	);
	LUT4 #(
		.INIT('h0020)
	) name8841 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14668_
	);
	LUT4 #(
		.INIT('hffde)
	) name8842 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14669_
	);
	LUT3 #(
		.INIT('hb0)
	) name8843 (
		_w14666_,
		_w14667_,
		_w14669_,
		_w14670_
	);
	LUT3 #(
		.INIT('h8a)
	) name8844 (
		_w14656_,
		_w14665_,
		_w14670_,
		_w14671_
	);
	LUT4 #(
		.INIT('h0010)
	) name8845 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14672_
	);
	LUT3 #(
		.INIT('hca)
	) name8846 (
		_w14659_,
		_w14661_,
		_w14657_,
		_w14673_
	);
	LUT3 #(
		.INIT('ha2)
	) name8847 (
		_w14660_,
		_w14658_,
		_w14661_,
		_w14674_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8848 (
		_w14657_,
		_w14672_,
		_w14673_,
		_w14674_,
		_w14675_
	);
	LUT3 #(
		.INIT('h40)
	) name8849 (
		_w14660_,
		_w14658_,
		_w14661_,
		_w14676_
	);
	LUT4 #(
		.INIT('h1000)
	) name8850 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14677_
	);
	LUT4 #(
		.INIT('hefdf)
	) name8851 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14678_
	);
	LUT4 #(
		.INIT('hef9a)
	) name8852 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14679_
	);
	LUT4 #(
		.INIT('hf351)
	) name8853 (
		_w14659_,
		_w14661_,
		_w14657_,
		_w14656_,
		_w14680_
	);
	LUT4 #(
		.INIT('h9099)
	) name8854 (
		_w14660_,
		_w14658_,
		_w14661_,
		_w14657_,
		_w14681_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name8855 (
		_w14679_,
		_w14657_,
		_w14680_,
		_w14681_,
		_w14682_
	);
	LUT3 #(
		.INIT('he0)
	) name8856 (
		_w14656_,
		_w14675_,
		_w14682_,
		_w14683_
	);
	LUT3 #(
		.INIT('h65)
	) name8857 (
		\u2_desIn_r_reg[42]/NET0131 ,
		_w14671_,
		_w14683_,
		_w14684_
	);
	LUT4 #(
		.INIT('hc963)
	) name8858 (
		decrypt_pad,
		\u2_desIn_r_reg[23]/NET0131 ,
		\u2_key_r_reg[3]/NET0131 ,
		\u2_key_r_reg[53]/NET0131 ,
		_w14685_
	);
	LUT4 #(
		.INIT('hc963)
	) name8859 (
		decrypt_pad,
		\u2_desIn_r_reg[7]/NET0131 ,
		\u2_key_r_reg[11]/NET0131 ,
		\u2_key_r_reg[4]/NET0131 ,
		_w14686_
	);
	LUT4 #(
		.INIT('hc693)
	) name8860 (
		decrypt_pad,
		\u2_desIn_r_reg[39]/NET0131 ,
		\u2_key_r_reg[34]/NET0131 ,
		\u2_key_r_reg[41]/NET0131 ,
		_w14687_
	);
	LUT4 #(
		.INIT('hc693)
	) name8861 (
		decrypt_pad,
		\u2_desIn_r_reg[15]/NET0131 ,
		\u2_key_r_reg[19]/NET0131 ,
		\u2_key_r_reg[26]/NET0131 ,
		_w14688_
	);
	LUT4 #(
		.INIT('hc693)
	) name8862 (
		decrypt_pad,
		\u2_desIn_r_reg[57]/NET0131 ,
		\u2_key_r_reg[40]/NET0131 ,
		\u2_key_r_reg[47]/NET0131 ,
		_w14689_
	);
	LUT4 #(
		.INIT('hf0dd)
	) name8863 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14690_
	);
	LUT2 #(
		.INIT('h2)
	) name8864 (
		_w14685_,
		_w14690_,
		_w14691_
	);
	LUT2 #(
		.INIT('h9)
	) name8865 (
		_w14688_,
		_w14689_,
		_w14692_
	);
	LUT2 #(
		.INIT('h8)
	) name8866 (
		_w14689_,
		_w14687_,
		_w14693_
	);
	LUT4 #(
		.INIT('h0206)
	) name8867 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14694_
	);
	LUT2 #(
		.INIT('h4)
	) name8868 (
		_w14689_,
		_w14687_,
		_w14695_
	);
	LUT2 #(
		.INIT('h4)
	) name8869 (
		_w14688_,
		_w14685_,
		_w14696_
	);
	LUT3 #(
		.INIT('hb0)
	) name8870 (
		_w14688_,
		_w14685_,
		_w14686_,
		_w14697_
	);
	LUT4 #(
		.INIT('hc963)
	) name8871 (
		decrypt_pad,
		\u2_desIn_r_reg[31]/NET0131 ,
		\u2_key_r_reg[13]/NET0131 ,
		\u2_key_r_reg[6]/NET0131 ,
		_w14698_
	);
	LUT4 #(
		.INIT('hdf00)
	) name8872 (
		_w14689_,
		_w14685_,
		_w14686_,
		_w14698_,
		_w14699_
	);
	LUT4 #(
		.INIT('h0d00)
	) name8873 (
		_w14695_,
		_w14697_,
		_w14694_,
		_w14699_,
		_w14700_
	);
	LUT2 #(
		.INIT('h4)
	) name8874 (
		_w14691_,
		_w14700_,
		_w14701_
	);
	LUT3 #(
		.INIT('h20)
	) name8875 (
		_w14688_,
		_w14689_,
		_w14685_,
		_w14702_
	);
	LUT4 #(
		.INIT('h2000)
	) name8876 (
		_w14688_,
		_w14689_,
		_w14685_,
		_w14687_,
		_w14703_
	);
	LUT4 #(
		.INIT('hdfee)
	) name8877 (
		_w14688_,
		_w14689_,
		_w14685_,
		_w14687_,
		_w14704_
	);
	LUT2 #(
		.INIT('h2)
	) name8878 (
		_w14686_,
		_w14704_,
		_w14705_
	);
	LUT2 #(
		.INIT('h1)
	) name8879 (
		_w14686_,
		_w14687_,
		_w14706_
	);
	LUT4 #(
		.INIT('haaa2)
	) name8880 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14707_
	);
	LUT3 #(
		.INIT('h0b)
	) name8881 (
		_w14688_,
		_w14689_,
		_w14685_,
		_w14708_
	);
	LUT3 #(
		.INIT('h10)
	) name8882 (
		_w14689_,
		_w14686_,
		_w14687_,
		_w14709_
	);
	LUT3 #(
		.INIT('h02)
	) name8883 (
		_w14708_,
		_w14707_,
		_w14709_,
		_w14710_
	);
	LUT4 #(
		.INIT('h0080)
	) name8884 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14711_
	);
	LUT2 #(
		.INIT('h8)
	) name8885 (
		_w14685_,
		_w14711_,
		_w14712_
	);
	LUT2 #(
		.INIT('h1)
	) name8886 (
		_w14688_,
		_w14686_,
		_w14713_
	);
	LUT3 #(
		.INIT('hba)
	) name8887 (
		_w14688_,
		_w14685_,
		_w14686_,
		_w14714_
	);
	LUT3 #(
		.INIT('h51)
	) name8888 (
		_w14698_,
		_w14693_,
		_w14714_,
		_w14715_
	);
	LUT4 #(
		.INIT('h0100)
	) name8889 (
		_w14705_,
		_w14712_,
		_w14710_,
		_w14715_,
		_w14716_
	);
	LUT4 #(
		.INIT('h28aa)
	) name8890 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14717_
	);
	LUT4 #(
		.INIT('h2232)
	) name8891 (
		_w14688_,
		_w14685_,
		_w14686_,
		_w14687_,
		_w14718_
	);
	LUT2 #(
		.INIT('h4)
	) name8892 (
		_w14717_,
		_w14718_,
		_w14719_
	);
	LUT4 #(
		.INIT('h0040)
	) name8893 (
		_w14688_,
		_w14689_,
		_w14685_,
		_w14686_,
		_w14720_
	);
	LUT3 #(
		.INIT('h07)
	) name8894 (
		_w14702_,
		_w14706_,
		_w14720_,
		_w14721_
	);
	LUT2 #(
		.INIT('h4)
	) name8895 (
		_w14719_,
		_w14721_,
		_w14722_
	);
	LUT4 #(
		.INIT('ha955)
	) name8896 (
		\u2_desIn_r_reg[48]/NET0131 ,
		_w14701_,
		_w14716_,
		_w14722_,
		_w14723_
	);
	LUT4 #(
		.INIT('hc693)
	) name8897 (
		decrypt_pad,
		\u2_desIn_r_reg[59]/NET0131 ,
		\u2_key_r_reg[28]/NET0131 ,
		\u2_key_r_reg[35]/P0001 ,
		_w14724_
	);
	LUT4 #(
		.INIT('hc693)
	) name8898 (
		decrypt_pad,
		\u2_desIn_r_reg[51]/NET0131 ,
		\u2_key_r_reg[2]/NET0131 ,
		\u2_key_r_reg[9]/NET0131 ,
		_w14725_
	);
	LUT4 #(
		.INIT('hc693)
	) name8899 (
		decrypt_pad,
		\u2_desIn_r_reg[43]/NET0131 ,
		\u2_key_r_reg[44]/NET0131 ,
		\u2_key_r_reg[51]/NET0131 ,
		_w14726_
	);
	LUT4 #(
		.INIT('hc963)
	) name8900 (
		decrypt_pad,
		\u2_desIn_r_reg[27]/NET0131 ,
		\u2_key_r_reg[14]/NET0131 ,
		\u2_key_r_reg[7]/NET0131 ,
		_w14727_
	);
	LUT4 #(
		.INIT('hc693)
	) name8901 (
		decrypt_pad,
		\u2_desIn_r_reg[35]/NET0131 ,
		\u2_key_r_reg[22]/NET0131 ,
		\u2_key_r_reg[29]/NET0131 ,
		_w14728_
	);
	LUT4 #(
		.INIT('h4555)
	) name8902 (
		_w14725_,
		_w14727_,
		_w14728_,
		_w14726_,
		_w14729_
	);
	LUT4 #(
		.INIT('h4515)
	) name8903 (
		_w14725_,
		_w14727_,
		_w14728_,
		_w14726_,
		_w14730_
	);
	LUT4 #(
		.INIT('hc693)
	) name8904 (
		decrypt_pad,
		\u2_desIn_r_reg[1]/NET0131 ,
		\u2_key_r_reg[23]/NET0131 ,
		\u2_key_r_reg[30]/NET0131 ,
		_w14731_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8905 (
		_w14725_,
		_w14727_,
		_w14728_,
		_w14731_,
		_w14732_
	);
	LUT3 #(
		.INIT('hda)
	) name8906 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14733_
	);
	LUT3 #(
		.INIT('h13)
	) name8907 (
		_w14732_,
		_w14730_,
		_w14733_,
		_w14734_
	);
	LUT2 #(
		.INIT('h2)
	) name8908 (
		_w14727_,
		_w14731_,
		_w14735_
	);
	LUT3 #(
		.INIT('hf2)
	) name8909 (
		_w14725_,
		_w14728_,
		_w14726_,
		_w14736_
	);
	LUT3 #(
		.INIT('h80)
	) name8910 (
		_w14727_,
		_w14726_,
		_w14731_,
		_w14737_
	);
	LUT4 #(
		.INIT('h2000)
	) name8911 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14738_
	);
	LUT3 #(
		.INIT('h0d)
	) name8912 (
		_w14735_,
		_w14736_,
		_w14738_,
		_w14739_
	);
	LUT3 #(
		.INIT('h45)
	) name8913 (
		_w14724_,
		_w14734_,
		_w14739_,
		_w14740_
	);
	LUT4 #(
		.INIT('h0002)
	) name8914 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14741_
	);
	LUT4 #(
		.INIT('h37bd)
	) name8915 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14742_
	);
	LUT2 #(
		.INIT('h2)
	) name8916 (
		_w14725_,
		_w14742_,
		_w14743_
	);
	LUT4 #(
		.INIT('h090f)
	) name8917 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14744_
	);
	LUT3 #(
		.INIT('h02)
	) name8918 (
		_w14729_,
		_w14737_,
		_w14744_,
		_w14745_
	);
	LUT3 #(
		.INIT('ha8)
	) name8919 (
		_w14724_,
		_w14743_,
		_w14745_,
		_w14746_
	);
	LUT4 #(
		.INIT('h5515)
	) name8920 (
		_w14725_,
		_w14727_,
		_w14728_,
		_w14731_,
		_w14747_
	);
	LUT3 #(
		.INIT('h01)
	) name8921 (
		_w14726_,
		_w14732_,
		_w14747_,
		_w14748_
	);
	LUT4 #(
		.INIT('h0004)
	) name8922 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14749_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name8923 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14750_
	);
	LUT3 #(
		.INIT('h01)
	) name8924 (
		_w14727_,
		_w14728_,
		_w14731_,
		_w14751_
	);
	LUT4 #(
		.INIT('he4f5)
	) name8925 (
		_w14725_,
		_w14726_,
		_w14750_,
		_w14751_,
		_w14752_
	);
	LUT2 #(
		.INIT('h4)
	) name8926 (
		_w14748_,
		_w14752_,
		_w14753_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name8927 (
		\u2_desIn_r_reg[20]/NET0131 ,
		_w14746_,
		_w14740_,
		_w14753_,
		_w14754_
	);
	LUT4 #(
		.INIT('hc693)
	) name8928 (
		decrypt_pad,
		\u2_desIn_r_reg[3]/NET0131 ,
		\u2_key_r_reg[13]/NET0131 ,
		\u2_key_r_reg[20]/NET0131 ,
		_w14755_
	);
	LUT4 #(
		.INIT('hc963)
	) name8929 (
		decrypt_pad,
		\u2_desIn_r_reg[29]/NET0131 ,
		\u2_key_r_reg[4]/NET0131 ,
		\u2_key_r_reg[54]/NET0131 ,
		_w14756_
	);
	LUT4 #(
		.INIT('hc693)
	) name8930 (
		decrypt_pad,
		\u2_desIn_r_reg[37]/NET0131 ,
		\u2_key_r_reg[48]/NET0131 ,
		\u2_key_r_reg[55]/NET0131 ,
		_w14757_
	);
	LUT4 #(
		.INIT('hc693)
	) name8931 (
		decrypt_pad,
		\u2_desIn_r_reg[53]/NET0131 ,
		\u2_key_r_reg[25]/NET0131 ,
		\u2_key_r_reg[32]/NET0131 ,
		_w14758_
	);
	LUT4 #(
		.INIT('h7e00)
	) name8932 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14758_,
		_w14759_
	);
	LUT4 #(
		.INIT('hc693)
	) name8933 (
		decrypt_pad,
		\u2_desIn_r_reg[45]/NET0131 ,
		\u2_key_r_reg[17]/NET0131 ,
		\u2_key_r_reg[24]/NET0131 ,
		_w14760_
	);
	LUT3 #(
		.INIT('h40)
	) name8934 (
		_w14755_,
		_w14756_,
		_w14760_,
		_w14761_
	);
	LUT3 #(
		.INIT('h0d)
	) name8935 (
		_w14755_,
		_w14757_,
		_w14758_,
		_w14762_
	);
	LUT3 #(
		.INIT('h45)
	) name8936 (
		_w14759_,
		_w14761_,
		_w14762_,
		_w14763_
	);
	LUT3 #(
		.INIT('h01)
	) name8937 (
		_w14755_,
		_w14756_,
		_w14760_,
		_w14764_
	);
	LUT4 #(
		.INIT('heffe)
	) name8938 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14765_
	);
	LUT4 #(
		.INIT('h0008)
	) name8939 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14766_
	);
	LUT4 #(
		.INIT('hc693)
	) name8940 (
		decrypt_pad,
		\u2_desIn_r_reg[61]/NET0131 ,
		\u2_key_r_reg[33]/NET0131 ,
		\u2_key_r_reg[40]/NET0131 ,
		_w14767_
	);
	LUT3 #(
		.INIT('h80)
	) name8941 (
		_w14757_,
		_w14760_,
		_w14758_,
		_w14768_
	);
	LUT4 #(
		.INIT('h4000)
	) name8942 (
		_w14756_,
		_w14757_,
		_w14760_,
		_w14758_,
		_w14769_
	);
	LUT4 #(
		.INIT('h0002)
	) name8943 (
		_w14765_,
		_w14767_,
		_w14769_,
		_w14766_,
		_w14770_
	);
	LUT2 #(
		.INIT('h4)
	) name8944 (
		_w14763_,
		_w14770_,
		_w14771_
	);
	LUT4 #(
		.INIT('h8000)
	) name8945 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14772_
	);
	LUT2 #(
		.INIT('h1)
	) name8946 (
		_w14757_,
		_w14758_,
		_w14773_
	);
	LUT4 #(
		.INIT('h0001)
	) name8947 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14758_,
		_w14774_
	);
	LUT2 #(
		.INIT('h4)
	) name8948 (
		_w14757_,
		_w14758_,
		_w14775_
	);
	LUT2 #(
		.INIT('h2)
	) name8949 (
		_w14755_,
		_w14756_,
		_w14776_
	);
	LUT4 #(
		.INIT('h0200)
	) name8950 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14758_,
		_w14777_
	);
	LUT4 #(
		.INIT('h040c)
	) name8951 (
		_w14760_,
		_w14767_,
		_w14777_,
		_w14774_,
		_w14778_
	);
	LUT4 #(
		.INIT('h4000)
	) name8952 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14758_,
		_w14779_
	);
	LUT4 #(
		.INIT('h0020)
	) name8953 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14780_
	);
	LUT2 #(
		.INIT('h1)
	) name8954 (
		_w14779_,
		_w14780_,
		_w14781_
	);
	LUT3 #(
		.INIT('hf9)
	) name8955 (
		_w14756_,
		_w14757_,
		_w14760_,
		_w14782_
	);
	LUT4 #(
		.INIT('h0006)
	) name8956 (
		_w14756_,
		_w14757_,
		_w14760_,
		_w14758_,
		_w14783_
	);
	LUT3 #(
		.INIT('h01)
	) name8957 (
		_w14779_,
		_w14780_,
		_w14783_,
		_w14784_
	);
	LUT3 #(
		.INIT('h40)
	) name8958 (
		_w14772_,
		_w14778_,
		_w14784_,
		_w14785_
	);
	LUT2 #(
		.INIT('h4)
	) name8959 (
		_w14758_,
		_w14780_,
		_w14786_
	);
	LUT3 #(
		.INIT('hbe)
	) name8960 (
		_w14755_,
		_w14756_,
		_w14760_,
		_w14787_
	);
	LUT4 #(
		.INIT('haf23)
	) name8961 (
		_w14760_,
		_w14775_,
		_w14779_,
		_w14787_,
		_w14788_
	);
	LUT2 #(
		.INIT('h4)
	) name8962 (
		_w14786_,
		_w14788_,
		_w14789_
	);
	LUT4 #(
		.INIT('ha955)
	) name8963 (
		\u2_desIn_r_reg[26]/NET0131 ,
		_w14771_,
		_w14785_,
		_w14789_,
		_w14790_
	);
	LUT4 #(
		.INIT('hbbdb)
	) name8964 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14791_
	);
	LUT4 #(
		.INIT('h7dff)
	) name8965 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14792_
	);
	LUT4 #(
		.INIT('hefe7)
	) name8966 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14793_
	);
	LUT4 #(
		.INIT('hc480)
	) name8967 (
		_w14758_,
		_w14792_,
		_w14793_,
		_w14791_,
		_w14794_
	);
	LUT2 #(
		.INIT('h2)
	) name8968 (
		_w14767_,
		_w14794_,
		_w14795_
	);
	LUT4 #(
		.INIT('hf3d9)
	) name8969 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14796_
	);
	LUT2 #(
		.INIT('h2)
	) name8970 (
		_w14758_,
		_w14796_,
		_w14797_
	);
	LUT3 #(
		.INIT('h08)
	) name8971 (
		_w14756_,
		_w14757_,
		_w14760_,
		_w14798_
	);
	LUT2 #(
		.INIT('h1)
	) name8972 (
		_w14760_,
		_w14758_,
		_w14799_
	);
	LUT4 #(
		.INIT('h0008)
	) name8973 (
		_w14755_,
		_w14756_,
		_w14760_,
		_w14758_,
		_w14800_
	);
	LUT4 #(
		.INIT('h0002)
	) name8974 (
		_w14765_,
		_w14774_,
		_w14800_,
		_w14798_,
		_w14801_
	);
	LUT3 #(
		.INIT('h45)
	) name8975 (
		_w14767_,
		_w14797_,
		_w14801_,
		_w14802_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name8976 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14803_
	);
	LUT2 #(
		.INIT('h1)
	) name8977 (
		_w14758_,
		_w14803_,
		_w14804_
	);
	LUT3 #(
		.INIT('h23)
	) name8978 (
		_w14760_,
		_w14769_,
		_w14779_,
		_w14805_
	);
	LUT2 #(
		.INIT('h4)
	) name8979 (
		_w14804_,
		_w14805_,
		_w14806_
	);
	LUT4 #(
		.INIT('h5655)
	) name8980 (
		\u2_desIn_r_reg[12]/NET0131 ,
		_w14802_,
		_w14795_,
		_w14806_,
		_w14807_
	);
	LUT4 #(
		.INIT('h33fe)
	) name8981 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14808_
	);
	LUT2 #(
		.INIT('h2)
	) name8982 (
		_w14657_,
		_w14808_,
		_w14809_
	);
	LUT4 #(
		.INIT('h0200)
	) name8983 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14810_
	);
	LUT3 #(
		.INIT('h04)
	) name8984 (
		_w14677_,
		_w14656_,
		_w14810_,
		_w14811_
	);
	LUT2 #(
		.INIT('h9)
	) name8985 (
		_w14659_,
		_w14660_,
		_w14812_
	);
	LUT4 #(
		.INIT('h080c)
	) name8986 (
		_w14660_,
		_w14658_,
		_w14661_,
		_w14657_,
		_w14813_
	);
	LUT3 #(
		.INIT('h45)
	) name8987 (
		_w14662_,
		_w14812_,
		_w14813_,
		_w14814_
	);
	LUT3 #(
		.INIT('h40)
	) name8988 (
		_w14809_,
		_w14811_,
		_w14814_,
		_w14815_
	);
	LUT4 #(
		.INIT('h0004)
	) name8989 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14816_
	);
	LUT4 #(
		.INIT('h00f7)
	) name8990 (
		_w14660_,
		_w14658_,
		_w14657_,
		_w14656_,
		_w14817_
	);
	LUT2 #(
		.INIT('h4)
	) name8991 (
		_w14816_,
		_w14817_,
		_w14818_
	);
	LUT4 #(
		.INIT('hfe6f)
	) name8992 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w14819_
	);
	LUT3 #(
		.INIT('h47)
	) name8993 (
		_w14658_,
		_w14661_,
		_w14657_,
		_w14820_
	);
	LUT3 #(
		.INIT('h09)
	) name8994 (
		_w14659_,
		_w14661_,
		_w14657_,
		_w14821_
	);
	LUT4 #(
		.INIT('h0d00)
	) name8995 (
		_w14663_,
		_w14820_,
		_w14821_,
		_w14819_,
		_w14822_
	);
	LUT2 #(
		.INIT('h8)
	) name8996 (
		_w14818_,
		_w14822_,
		_w14823_
	);
	LUT3 #(
		.INIT('ha9)
	) name8997 (
		\u2_desIn_r_reg[28]/NET0131 ,
		_w14815_,
		_w14823_,
		_w14824_
	);
	LUT4 #(
		.INIT('hc693)
	) name8998 (
		decrypt_pad,
		\u2_desIn_r_reg[27]/NET0131 ,
		\u2_key_r_reg[16]/NET0131 ,
		\u2_key_r_reg[23]/NET0131 ,
		_w14825_
	);
	LUT4 #(
		.INIT('hc693)
	) name8999 (
		decrypt_pad,
		\u2_desIn_r_reg[11]/NET0131 ,
		\u2_key_r_reg[14]/NET0131 ,
		\u2_key_r_reg[21]/NET0131 ,
		_w14826_
	);
	LUT4 #(
		.INIT('hc693)
	) name9000 (
		decrypt_pad,
		\u2_desIn_r_reg[19]/NET0131 ,
		\u2_key_r_reg[1]/NET0131 ,
		\u2_key_r_reg[8]/NET0131 ,
		_w14827_
	);
	LUT4 #(
		.INIT('hc693)
	) name9001 (
		decrypt_pad,
		\u2_desIn_r_reg[35]/NET0131 ,
		\u2_key_r_reg[45]/NET0131 ,
		\u2_key_r_reg[52]/NET0131 ,
		_w14828_
	);
	LUT4 #(
		.INIT('hc693)
	) name9002 (
		decrypt_pad,
		\u2_desIn_r_reg[61]/NET0131 ,
		\u2_key_r_reg[29]/NET0131 ,
		\u2_key_r_reg[36]/NET0131 ,
		_w14829_
	);
	LUT4 #(
		.INIT('hc963)
	) name9003 (
		decrypt_pad,
		\u2_desIn_r_reg[3]/NET0131 ,
		\u2_key_r_reg[31]/NET0131 ,
		\u2_key_r_reg[51]/NET0131 ,
		_w14830_
	);
	LUT4 #(
		.INIT('h0020)
	) name9004 (
		_w14828_,
		_w14829_,
		_w14830_,
		_w14827_,
		_w14831_
	);
	LUT4 #(
		.INIT('hb796)
	) name9005 (
		_w14828_,
		_w14829_,
		_w14830_,
		_w14827_,
		_w14832_
	);
	LUT2 #(
		.INIT('h1)
	) name9006 (
		_w14826_,
		_w14832_,
		_w14833_
	);
	LUT4 #(
		.INIT('h93d5)
	) name9007 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14834_
	);
	LUT2 #(
		.INIT('h2)
	) name9008 (
		_w14827_,
		_w14834_,
		_w14835_
	);
	LUT3 #(
		.INIT('h80)
	) name9009 (
		_w14828_,
		_w14829_,
		_w14830_,
		_w14836_
	);
	LUT2 #(
		.INIT('h2)
	) name9010 (
		_w14826_,
		_w14827_,
		_w14837_
	);
	LUT4 #(
		.INIT('h0040)
	) name9011 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14838_
	);
	LUT3 #(
		.INIT('h07)
	) name9012 (
		_w14836_,
		_w14837_,
		_w14838_,
		_w14839_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9013 (
		_w14825_,
		_w14835_,
		_w14833_,
		_w14839_,
		_w14840_
	);
	LUT4 #(
		.INIT('h0180)
	) name9014 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14841_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9015 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14827_,
		_w14842_
	);
	LUT4 #(
		.INIT('hfcee)
	) name9016 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14843_
	);
	LUT2 #(
		.INIT('h8)
	) name9017 (
		_w14842_,
		_w14843_,
		_w14844_
	);
	LUT3 #(
		.INIT('h02)
	) name9018 (
		_w14828_,
		_w14829_,
		_w14830_,
		_w14845_
	);
	LUT4 #(
		.INIT('h00bf)
	) name9019 (
		_w14828_,
		_w14826_,
		_w14830_,
		_w14827_,
		_w14846_
	);
	LUT4 #(
		.INIT('h0004)
	) name9020 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14847_
	);
	LUT4 #(
		.INIT('h0800)
	) name9021 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14848_
	);
	LUT4 #(
		.INIT('hf7fb)
	) name9022 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14849_
	);
	LUT3 #(
		.INIT('h40)
	) name9023 (
		_w14845_,
		_w14846_,
		_w14849_,
		_w14850_
	);
	LUT4 #(
		.INIT('h00ab)
	) name9024 (
		_w14841_,
		_w14844_,
		_w14850_,
		_w14825_,
		_w14851_
	);
	LUT4 #(
		.INIT('h0400)
	) name9025 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14852_
	);
	LUT4 #(
		.INIT('hfbef)
	) name9026 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14853_
	);
	LUT4 #(
		.INIT('h0020)
	) name9027 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14854_
	);
	LUT4 #(
		.INIT('hefdf)
	) name9028 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w14855_
	);
	LUT3 #(
		.INIT('hd8)
	) name9029 (
		_w14827_,
		_w14853_,
		_w14855_,
		_w14856_
	);
	LUT4 #(
		.INIT('h5655)
	) name9030 (
		\u2_desIn_r_reg[44]/NET0131 ,
		_w14851_,
		_w14840_,
		_w14856_,
		_w14857_
	);
	LUT4 #(
		.INIT('hc693)
	) name9031 (
		decrypt_pad,
		\u2_desIn_r_reg[7]/NET0131 ,
		\u2_key_r_reg[21]/NET0131 ,
		\u2_key_r_reg[28]/NET0131 ,
		_w14858_
	);
	LUT4 #(
		.INIT('hc693)
	) name9032 (
		decrypt_pad,
		\u2_desIn_r_reg[41]/NET0131 ,
		\u2_key_r_reg[37]/NET0131 ,
		\u2_key_r_reg[44]/NET0131 ,
		_w14859_
	);
	LUT4 #(
		.INIT('hc963)
	) name9033 (
		decrypt_pad,
		\u2_desIn_r_reg[25]/NET0131 ,
		\u2_key_r_reg[16]/NET0131 ,
		\u2_key_r_reg[9]/NET0131 ,
		_w14860_
	);
	LUT4 #(
		.INIT('hc693)
	) name9034 (
		decrypt_pad,
		\u2_desIn_r_reg[33]/NET0131 ,
		\u2_key_r_reg[36]/NET0131 ,
		\u2_key_r_reg[43]/NET0131 ,
		_w14861_
	);
	LUT4 #(
		.INIT('hc963)
	) name9035 (
		decrypt_pad,
		\u2_desIn_r_reg[49]/NET0131 ,
		\u2_key_r_reg[1]/NET0131 ,
		\u2_key_r_reg[49]/NET0131 ,
		_w14862_
	);
	LUT3 #(
		.INIT('h10)
	) name9036 (
		_w14862_,
		_w14861_,
		_w14859_,
		_w14863_
	);
	LUT4 #(
		.INIT('hf2ff)
	) name9037 (
		_w14862_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14864_
	);
	LUT2 #(
		.INIT('h2)
	) name9038 (
		_w14858_,
		_w14864_,
		_w14865_
	);
	LUT3 #(
		.INIT('he3)
	) name9039 (
		_w14858_,
		_w14860_,
		_w14859_,
		_w14866_
	);
	LUT4 #(
		.INIT('h10c0)
	) name9040 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14867_
	);
	LUT4 #(
		.INIT('hc693)
	) name9041 (
		decrypt_pad,
		\u2_desIn_r_reg[57]/NET0131 ,
		\u2_key_r_reg[0]/NET0131 ,
		\u2_key_r_reg[7]/NET0131 ,
		_w14868_
	);
	LUT2 #(
		.INIT('h2)
	) name9042 (
		_w14862_,
		_w14861_,
		_w14869_
	);
	LUT4 #(
		.INIT('h0002)
	) name9043 (
		_w14862_,
		_w14858_,
		_w14860_,
		_w14861_,
		_w14870_
	);
	LUT3 #(
		.INIT('h02)
	) name9044 (
		_w14868_,
		_w14867_,
		_w14870_,
		_w14871_
	);
	LUT4 #(
		.INIT('h3d2d)
	) name9045 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14872_
	);
	LUT4 #(
		.INIT('h0004)
	) name9046 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14873_
	);
	LUT4 #(
		.INIT('h0301)
	) name9047 (
		_w14862_,
		_w14868_,
		_w14873_,
		_w14872_,
		_w14874_
	);
	LUT3 #(
		.INIT('h0b)
	) name9048 (
		_w14865_,
		_w14871_,
		_w14874_,
		_w14875_
	);
	LUT2 #(
		.INIT('h6)
	) name9049 (
		_w14861_,
		_w14859_,
		_w14876_
	);
	LUT4 #(
		.INIT('h1001)
	) name9050 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14877_
	);
	LUT4 #(
		.INIT('h0020)
	) name9051 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14878_
	);
	LUT4 #(
		.INIT('h2022)
	) name9052 (
		_w14860_,
		_w14861_,
		_w14859_,
		_w14868_,
		_w14879_
	);
	LUT4 #(
		.INIT('h5554)
	) name9053 (
		_w14862_,
		_w14878_,
		_w14877_,
		_w14879_,
		_w14880_
	);
	LUT3 #(
		.INIT('h08)
	) name9054 (
		_w14862_,
		_w14858_,
		_w14860_,
		_w14881_
	);
	LUT2 #(
		.INIT('h4)
	) name9055 (
		_w14876_,
		_w14881_,
		_w14882_
	);
	LUT2 #(
		.INIT('h1)
	) name9056 (
		_w14880_,
		_w14882_,
		_w14883_
	);
	LUT3 #(
		.INIT('h65)
	) name9057 (
		\u2_desIn_r_reg[52]/NET0131 ,
		_w14875_,
		_w14883_,
		_w14884_
	);
	LUT4 #(
		.INIT('h4010)
	) name9058 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14885_
	);
	LUT3 #(
		.INIT('h02)
	) name9059 (
		_w14728_,
		_w14726_,
		_w14731_,
		_w14886_
	);
	LUT4 #(
		.INIT('he6f7)
	) name9060 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14887_
	);
	LUT4 #(
		.INIT('h0031)
	) name9061 (
		_w14725_,
		_w14886_,
		_w14887_,
		_w14885_,
		_w14888_
	);
	LUT2 #(
		.INIT('h2)
	) name9062 (
		_w14724_,
		_w14888_,
		_w14889_
	);
	LUT4 #(
		.INIT('h1001)
	) name9063 (
		_w14725_,
		_w14727_,
		_w14728_,
		_w14731_,
		_w14890_
	);
	LUT4 #(
		.INIT('h8000)
	) name9064 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14891_
	);
	LUT4 #(
		.INIT('h5d19)
	) name9065 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14892_
	);
	LUT4 #(
		.INIT('h0031)
	) name9066 (
		_w14725_,
		_w14891_,
		_w14892_,
		_w14890_,
		_w14893_
	);
	LUT4 #(
		.INIT('hb8bb)
	) name9067 (
		_w14725_,
		_w14727_,
		_w14726_,
		_w14731_,
		_w14894_
	);
	LUT4 #(
		.INIT('h0400)
	) name9068 (
		_w14725_,
		_w14727_,
		_w14726_,
		_w14731_,
		_w14895_
	);
	LUT4 #(
		.INIT('h0032)
	) name9069 (
		_w14724_,
		_w14728_,
		_w14895_,
		_w14894_,
		_w14896_
	);
	LUT4 #(
		.INIT('h0032)
	) name9070 (
		_w14724_,
		_w14748_,
		_w14893_,
		_w14896_,
		_w14897_
	);
	LUT3 #(
		.INIT('h65)
	) name9071 (
		\u2_desIn_r_reg[18]/NET0131 ,
		_w14889_,
		_w14897_,
		_w14898_
	);
	LUT4 #(
		.INIT('h0400)
	) name9072 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14899_
	);
	LUT4 #(
		.INIT('hc9cd)
	) name9073 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14900_
	);
	LUT4 #(
		.INIT('h0809)
	) name9074 (
		_w14688_,
		_w14689_,
		_w14685_,
		_w14686_,
		_w14901_
	);
	LUT4 #(
		.INIT('h0040)
	) name9075 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14902_
	);
	LUT4 #(
		.INIT('h5fbf)
	) name9076 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14903_
	);
	LUT4 #(
		.INIT('h0d00)
	) name9077 (
		_w14685_,
		_w14900_,
		_w14901_,
		_w14903_,
		_w14904_
	);
	LUT4 #(
		.INIT('hf3ec)
	) name9078 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14905_
	);
	LUT4 #(
		.INIT('h0280)
	) name9079 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14906_
	);
	LUT3 #(
		.INIT('h0e)
	) name9080 (
		_w14685_,
		_w14905_,
		_w14906_,
		_w14907_
	);
	LUT4 #(
		.INIT('h1020)
	) name9081 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w14908_
	);
	LUT4 #(
		.INIT('h0082)
	) name9082 (
		_w14689_,
		_w14686_,
		_w14687_,
		_w14698_,
		_w14909_
	);
	LUT3 #(
		.INIT('ha8)
	) name9083 (
		_w14685_,
		_w14908_,
		_w14909_,
		_w14910_
	);
	LUT4 #(
		.INIT('h0e04)
	) name9084 (
		_w14698_,
		_w14907_,
		_w14910_,
		_w14904_,
		_w14911_
	);
	LUT2 #(
		.INIT('h9)
	) name9085 (
		\u2_desIn_r_reg[2]/NET0131 ,
		_w14911_,
		_w14912_
	);
	LUT4 #(
		.INIT('h5545)
	) name9086 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14913_
	);
	LUT4 #(
		.INIT('h004c)
	) name9087 (
		_w14756_,
		_w14757_,
		_w14760_,
		_w14758_,
		_w14914_
	);
	LUT2 #(
		.INIT('h4)
	) name9088 (
		_w14913_,
		_w14914_,
		_w14915_
	);
	LUT3 #(
		.INIT('h51)
	) name9089 (
		_w14755_,
		_w14756_,
		_w14760_,
		_w14916_
	);
	LUT4 #(
		.INIT('h4000)
	) name9090 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14917_
	);
	LUT4 #(
		.INIT('hbcff)
	) name9091 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14918_
	);
	LUT3 #(
		.INIT('hd0)
	) name9092 (
		_w14775_,
		_w14916_,
		_w14918_,
		_w14919_
	);
	LUT3 #(
		.INIT('h8a)
	) name9093 (
		_w14767_,
		_w14915_,
		_w14919_,
		_w14920_
	);
	LUT4 #(
		.INIT('h084c)
	) name9094 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14921_
	);
	LUT4 #(
		.INIT('h0400)
	) name9095 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14922_
	);
	LUT4 #(
		.INIT('hfcb8)
	) name9096 (
		_w14764_,
		_w14758_,
		_w14921_,
		_w14922_,
		_w14923_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name9097 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14924_
	);
	LUT3 #(
		.INIT('h45)
	) name9098 (
		_w14767_,
		_w14923_,
		_w14924_,
		_w14925_
	);
	LUT4 #(
		.INIT('h6dff)
	) name9099 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14926_
	);
	LUT2 #(
		.INIT('h2)
	) name9100 (
		_w14758_,
		_w14926_,
		_w14927_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name9101 (
		_w14760_,
		_w14758_,
		_w14774_,
		_w14917_,
		_w14928_
	);
	LUT2 #(
		.INIT('h4)
	) name9102 (
		_w14927_,
		_w14928_,
		_w14929_
	);
	LUT4 #(
		.INIT('h5655)
	) name9103 (
		\u2_desIn_r_reg[6]/NET0131 ,
		_w14925_,
		_w14920_,
		_w14929_,
		_w14930_
	);
	LUT2 #(
		.INIT('h4)
	) name9104 (
		_w14862_,
		_w14861_,
		_w14931_
	);
	LUT4 #(
		.INIT('h0100)
	) name9105 (
		_w14862_,
		_w14858_,
		_w14860_,
		_w14861_,
		_w14932_
	);
	LUT4 #(
		.INIT('h0400)
	) name9106 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14933_
	);
	LUT3 #(
		.INIT('h01)
	) name9107 (
		_w14868_,
		_w14933_,
		_w14932_,
		_w14934_
	);
	LUT3 #(
		.INIT('h01)
	) name9108 (
		_w14860_,
		_w14861_,
		_w14859_,
		_w14935_
	);
	LUT4 #(
		.INIT('h0001)
	) name9109 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14936_
	);
	LUT3 #(
		.INIT('h08)
	) name9110 (
		_w14858_,
		_w14860_,
		_w14859_,
		_w14937_
	);
	LUT3 #(
		.INIT('h0b)
	) name9111 (
		_w14869_,
		_w14937_,
		_w14936_,
		_w14938_
	);
	LUT4 #(
		.INIT('hb3bf)
	) name9112 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14939_
	);
	LUT4 #(
		.INIT('h0bff)
	) name9113 (
		_w14862_,
		_w14858_,
		_w14861_,
		_w14859_,
		_w14940_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name9114 (
		_w14862_,
		_w14860_,
		_w14939_,
		_w14940_,
		_w14941_
	);
	LUT3 #(
		.INIT('h80)
	) name9115 (
		_w14934_,
		_w14938_,
		_w14941_,
		_w14942_
	);
	LUT4 #(
		.INIT('h0844)
	) name9116 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14943_
	);
	LUT3 #(
		.INIT('h02)
	) name9117 (
		_w14858_,
		_w14861_,
		_w14859_,
		_w14944_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name9118 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14945_
	);
	LUT4 #(
		.INIT('he4ee)
	) name9119 (
		_w14862_,
		_w14943_,
		_w14944_,
		_w14945_,
		_w14946_
	);
	LUT4 #(
		.INIT('h4100)
	) name9120 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14947_
	);
	LUT4 #(
		.INIT('h0002)
	) name9121 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14948_
	);
	LUT3 #(
		.INIT('h02)
	) name9122 (
		_w14868_,
		_w14948_,
		_w14947_,
		_w14949_
	);
	LUT2 #(
		.INIT('h4)
	) name9123 (
		_w14946_,
		_w14949_,
		_w14950_
	);
	LUT4 #(
		.INIT('h0002)
	) name9124 (
		_w14862_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w14951_
	);
	LUT3 #(
		.INIT('h15)
	) name9125 (
		_w14951_,
		_w14931_,
		_w14937_,
		_w14952_
	);
	LUT4 #(
		.INIT('ha955)
	) name9126 (
		\u2_desIn_r_reg[34]/NET0131 ,
		_w14942_,
		_w14950_,
		_w14952_,
		_w14953_
	);
	LUT4 #(
		.INIT('h9cee)
	) name9127 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14954_
	);
	LUT2 #(
		.INIT('h1)
	) name9128 (
		_w14773_,
		_w14954_,
		_w14955_
	);
	LUT4 #(
		.INIT('h7775)
	) name9129 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14956_
	);
	LUT3 #(
		.INIT('h0d)
	) name9130 (
		_w14756_,
		_w14760_,
		_w14758_,
		_w14957_
	);
	LUT3 #(
		.INIT('h8a)
	) name9131 (
		_w14767_,
		_w14956_,
		_w14957_,
		_w14958_
	);
	LUT2 #(
		.INIT('h4)
	) name9132 (
		_w14955_,
		_w14958_,
		_w14959_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name9133 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14760_,
		_w14960_
	);
	LUT2 #(
		.INIT('h1)
	) name9134 (
		_w14758_,
		_w14960_,
		_w14961_
	);
	LUT4 #(
		.INIT('h00fd)
	) name9135 (
		_w14756_,
		_w14757_,
		_w14760_,
		_w14767_,
		_w14962_
	);
	LUT3 #(
		.INIT('hd0)
	) name9136 (
		_w14768_,
		_w14776_,
		_w14962_,
		_w14963_
	);
	LUT3 #(
		.INIT('h20)
	) name9137 (
		_w14781_,
		_w14961_,
		_w14963_,
		_w14964_
	);
	LUT3 #(
		.INIT('h6b)
	) name9138 (
		_w14755_,
		_w14756_,
		_w14757_,
		_w14965_
	);
	LUT2 #(
		.INIT('h8)
	) name9139 (
		_w14755_,
		_w14758_,
		_w14966_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name9140 (
		_w14782_,
		_w14799_,
		_w14965_,
		_w14966_,
		_w14967_
	);
	LUT4 #(
		.INIT('ha955)
	) name9141 (
		\u2_desIn_r_reg[8]/NET0131 ,
		_w14959_,
		_w14964_,
		_w14967_,
		_w14968_
	);
	LUT4 #(
		.INIT('hc693)
	) name9142 (
		decrypt_pad,
		\u2_desIn_r_reg[63]/NET0131 ,
		\u2_key_r_reg[32]/NET0131 ,
		\u2_key_r_reg[39]/P0001 ,
		_w14969_
	);
	LUT4 #(
		.INIT('hc693)
	) name9143 (
		decrypt_pad,
		\u2_desIn_r_reg[55]/NET0131 ,
		\u2_key_r_reg[41]/NET0131 ,
		\u2_key_r_reg[48]/NET0131 ,
		_w14970_
	);
	LUT4 #(
		.INIT('hc693)
	) name9144 (
		decrypt_pad,
		\u2_desIn_r_reg[47]/NET0131 ,
		\u2_key_r_reg[47]/NET0131 ,
		\u2_key_r_reg[54]/NET0131 ,
		_w14971_
	);
	LUT4 #(
		.INIT('hc693)
	) name9145 (
		decrypt_pad,
		\u2_desIn_r_reg[31]/NET0131 ,
		\u2_key_r_reg[20]/NET0131 ,
		\u2_key_r_reg[27]/NET0131 ,
		_w14972_
	);
	LUT4 #(
		.INIT('hc693)
	) name9146 (
		decrypt_pad,
		\u2_desIn_r_reg[5]/NET0131 ,
		\u2_key_r_reg[12]/NET0131 ,
		\u2_key_r_reg[19]/NET0131 ,
		_w14973_
	);
	LUT4 #(
		.INIT('hc693)
	) name9147 (
		decrypt_pad,
		\u2_desIn_r_reg[39]/NET0131 ,
		\u2_key_r_reg[24]/NET0131 ,
		\u2_key_r_reg[6]/NET0131 ,
		_w14974_
	);
	LUT4 #(
		.INIT('h5a4f)
	) name9148 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w14975_
	);
	LUT4 #(
		.INIT('hf5fc)
	) name9149 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w14976_
	);
	LUT4 #(
		.INIT('hbf7b)
	) name9150 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w14977_
	);
	LUT4 #(
		.INIT('hd800)
	) name9151 (
		_w14970_,
		_w14976_,
		_w14975_,
		_w14977_,
		_w14978_
	);
	LUT2 #(
		.INIT('h1)
	) name9152 (
		_w14969_,
		_w14978_,
		_w14979_
	);
	LUT4 #(
		.INIT('hfb7b)
	) name9153 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w14980_
	);
	LUT2 #(
		.INIT('h1)
	) name9154 (
		_w14980_,
		_w14970_,
		_w14981_
	);
	LUT3 #(
		.INIT('h02)
	) name9155 (
		_w14974_,
		_w14972_,
		_w14973_,
		_w14982_
	);
	LUT4 #(
		.INIT('h5fa7)
	) name9156 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w14983_
	);
	LUT2 #(
		.INIT('h2)
	) name9157 (
		_w14970_,
		_w14983_,
		_w14984_
	);
	LUT2 #(
		.INIT('h1)
	) name9158 (
		_w14970_,
		_w14976_,
		_w14985_
	);
	LUT4 #(
		.INIT('h0400)
	) name9159 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w14986_
	);
	LUT3 #(
		.INIT('h0b)
	) name9160 (
		_w14974_,
		_w14973_,
		_w14970_,
		_w14987_
	);
	LUT2 #(
		.INIT('h4)
	) name9161 (
		_w14971_,
		_w14972_,
		_w14988_
	);
	LUT3 #(
		.INIT('h45)
	) name9162 (
		_w14986_,
		_w14987_,
		_w14988_,
		_w14989_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9163 (
		_w14969_,
		_w14984_,
		_w14985_,
		_w14989_,
		_w14990_
	);
	LUT4 #(
		.INIT('h5556)
	) name9164 (
		\u2_desIn_r_reg[24]/NET0131 ,
		_w14981_,
		_w14990_,
		_w14979_,
		_w14991_
	);
	LUT4 #(
		.INIT('h779c)
	) name9165 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14992_
	);
	LUT4 #(
		.INIT('h0e04)
	) name9166 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14993_
	);
	LUT4 #(
		.INIT('hf17b)
	) name9167 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14994_
	);
	LUT4 #(
		.INIT('h1000)
	) name9168 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14995_
	);
	LUT4 #(
		.INIT('h00e4)
	) name9169 (
		_w14725_,
		_w14994_,
		_w14992_,
		_w14995_,
		_w14996_
	);
	LUT2 #(
		.INIT('h1)
	) name9170 (
		_w14724_,
		_w14996_,
		_w14997_
	);
	LUT4 #(
		.INIT('hbb7b)
	) name9171 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w14998_
	);
	LUT2 #(
		.INIT('h2)
	) name9172 (
		_w14725_,
		_w14998_,
		_w14999_
	);
	LUT3 #(
		.INIT('h48)
	) name9173 (
		_w14727_,
		_w14726_,
		_w14731_,
		_w15000_
	);
	LUT4 #(
		.INIT('h888a)
	) name9174 (
		_w14725_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w15001_
	);
	LUT3 #(
		.INIT('h01)
	) name9175 (
		_w14993_,
		_w15001_,
		_w15000_,
		_w15002_
	);
	LUT4 #(
		.INIT('h0800)
	) name9176 (
		_w14725_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w15003_
	);
	LUT2 #(
		.INIT('h1)
	) name9177 (
		_w14741_,
		_w15003_,
		_w15004_
	);
	LUT4 #(
		.INIT('h5700)
	) name9178 (
		_w14724_,
		_w14999_,
		_w15002_,
		_w15004_,
		_w15005_
	);
	LUT3 #(
		.INIT('h9a)
	) name9179 (
		\u2_desIn_r_reg[32]/NET0131 ,
		_w14997_,
		_w15005_,
		_w15006_
	);
	LUT4 #(
		.INIT('h0122)
	) name9180 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15007_
	);
	LUT4 #(
		.INIT('h0800)
	) name9181 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15008_
	);
	LUT4 #(
		.INIT('h0010)
	) name9182 (
		_w14974_,
		_w14971_,
		_w14973_,
		_w14970_,
		_w15009_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name9183 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15010_
	);
	LUT4 #(
		.INIT('h00bf)
	) name9184 (
		_w14974_,
		_w14972_,
		_w14973_,
		_w14970_,
		_w15011_
	);
	LUT4 #(
		.INIT('h1011)
	) name9185 (
		_w15008_,
		_w15009_,
		_w15010_,
		_w15011_,
		_w15012_
	);
	LUT3 #(
		.INIT('h45)
	) name9186 (
		_w14969_,
		_w15007_,
		_w15012_,
		_w15013_
	);
	LUT4 #(
		.INIT('h2010)
	) name9187 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15014_
	);
	LUT4 #(
		.INIT('ha200)
	) name9188 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14970_,
		_w15015_
	);
	LUT3 #(
		.INIT('ha8)
	) name9189 (
		_w14969_,
		_w15014_,
		_w15015_,
		_w15016_
	);
	LUT3 #(
		.INIT('h04)
	) name9190 (
		_w14974_,
		_w14971_,
		_w14973_,
		_w15017_
	);
	LUT4 #(
		.INIT('h0004)
	) name9191 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15018_
	);
	LUT4 #(
		.INIT('h4000)
	) name9192 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15019_
	);
	LUT4 #(
		.INIT('hdf00)
	) name9193 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14970_,
		_w15020_
	);
	LUT4 #(
		.INIT('h0b00)
	) name9194 (
		_w14969_,
		_w15019_,
		_w15018_,
		_w15020_,
		_w15021_
	);
	LUT4 #(
		.INIT('hbff2)
	) name9195 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15022_
	);
	LUT4 #(
		.INIT('h0900)
	) name9196 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15023_
	);
	LUT4 #(
		.INIT('h0051)
	) name9197 (
		_w14970_,
		_w14969_,
		_w15022_,
		_w15023_,
		_w15024_
	);
	LUT3 #(
		.INIT('h54)
	) name9198 (
		_w15016_,
		_w15021_,
		_w15024_,
		_w15025_
	);
	LUT3 #(
		.INIT('h65)
	) name9199 (
		\u2_desIn_r_reg[14]/NET0131 ,
		_w15013_,
		_w15025_,
		_w15026_
	);
	LUT4 #(
		.INIT('h67c8)
	) name9200 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15027_
	);
	LUT4 #(
		.INIT('hfc77)
	) name9201 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15028_
	);
	LUT4 #(
		.INIT('hb5ff)
	) name9202 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15029_
	);
	LUT4 #(
		.INIT('hd800)
	) name9203 (
		_w14827_,
		_w15027_,
		_w15028_,
		_w15029_,
		_w15030_
	);
	LUT2 #(
		.INIT('h2)
	) name9204 (
		_w14825_,
		_w15030_,
		_w15031_
	);
	LUT4 #(
		.INIT('hbfed)
	) name9205 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15032_
	);
	LUT2 #(
		.INIT('h2)
	) name9206 (
		_w14827_,
		_w15032_,
		_w15033_
	);
	LUT4 #(
		.INIT('hcfbb)
	) name9207 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15034_
	);
	LUT2 #(
		.INIT('h4)
	) name9208 (
		_w14828_,
		_w14827_,
		_w15035_
	);
	LUT3 #(
		.INIT('hb0)
	) name9209 (
		_w14828_,
		_w14830_,
		_w14827_,
		_w15036_
	);
	LUT4 #(
		.INIT('h3301)
	) name9210 (
		_w14829_,
		_w14826_,
		_w14830_,
		_w14827_,
		_w15037_
	);
	LUT4 #(
		.INIT('he0ee)
	) name9211 (
		_w15034_,
		_w15035_,
		_w15036_,
		_w15037_,
		_w15038_
	);
	LUT4 #(
		.INIT('h0008)
	) name9212 (
		_w14829_,
		_w14826_,
		_w14830_,
		_w14827_,
		_w15039_
	);
	LUT2 #(
		.INIT('h1)
	) name9213 (
		_w14848_,
		_w15039_,
		_w15040_
	);
	LUT4 #(
		.INIT('h0e00)
	) name9214 (
		_w14825_,
		_w15038_,
		_w15033_,
		_w15040_,
		_w15041_
	);
	LUT3 #(
		.INIT('h65)
	) name9215 (
		\u2_desIn_r_reg[0]/NET0131 ,
		_w15031_,
		_w15041_,
		_w15042_
	);
	LUT3 #(
		.INIT('h80)
	) name9216 (
		_w14728_,
		_w14726_,
		_w14731_,
		_w15043_
	);
	LUT4 #(
		.INIT('h0800)
	) name9217 (
		_w14725_,
		_w14727_,
		_w14726_,
		_w14731_,
		_w15044_
	);
	LUT4 #(
		.INIT('h0002)
	) name9218 (
		_w14724_,
		_w14749_,
		_w15044_,
		_w15043_,
		_w15045_
	);
	LUT4 #(
		.INIT('hda77)
	) name9219 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w15046_
	);
	LUT2 #(
		.INIT('h2)
	) name9220 (
		_w14725_,
		_w15046_,
		_w15047_
	);
	LUT3 #(
		.INIT('h01)
	) name9221 (
		_w14724_,
		_w14741_,
		_w14895_,
		_w15048_
	);
	LUT3 #(
		.INIT('h45)
	) name9222 (
		_w15045_,
		_w15047_,
		_w15048_,
		_w15049_
	);
	LUT4 #(
		.INIT('hefbb)
	) name9223 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w15050_
	);
	LUT3 #(
		.INIT('h01)
	) name9224 (
		_w14727_,
		_w14726_,
		_w14731_,
		_w15051_
	);
	LUT4 #(
		.INIT('hfaf2)
	) name9225 (
		_w14727_,
		_w14728_,
		_w14726_,
		_w14731_,
		_w15052_
	);
	LUT4 #(
		.INIT('h3210)
	) name9226 (
		_w14724_,
		_w15051_,
		_w15050_,
		_w15052_,
		_w15053_
	);
	LUT4 #(
		.INIT('h1551)
	) name9227 (
		_w14725_,
		_w14727_,
		_w14728_,
		_w14731_,
		_w15054_
	);
	LUT4 #(
		.INIT('h8a28)
	) name9228 (
		_w14725_,
		_w14727_,
		_w14728_,
		_w14731_,
		_w15055_
	);
	LUT3 #(
		.INIT('h02)
	) name9229 (
		_w14726_,
		_w15055_,
		_w15054_,
		_w15056_
	);
	LUT3 #(
		.INIT('h0e)
	) name9230 (
		_w14725_,
		_w15053_,
		_w15056_,
		_w15057_
	);
	LUT3 #(
		.INIT('h65)
	) name9231 (
		\u2_desIn_r_reg[30]/NET0131 ,
		_w15049_,
		_w15057_,
		_w15058_
	);
	LUT4 #(
		.INIT('haaa2)
	) name9232 (
		_w14862_,
		_w14858_,
		_w14860_,
		_w14861_,
		_w15059_
	);
	LUT3 #(
		.INIT('h15)
	) name9233 (
		_w14862_,
		_w14858_,
		_w14861_,
		_w15060_
	);
	LUT4 #(
		.INIT('h45cf)
	) name9234 (
		_w14866_,
		_w14933_,
		_w15059_,
		_w15060_,
		_w15061_
	);
	LUT4 #(
		.INIT('h0040)
	) name9235 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15062_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name9236 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15063_
	);
	LUT3 #(
		.INIT('h45)
	) name9237 (
		_w14868_,
		_w15061_,
		_w15063_,
		_w15064_
	);
	LUT4 #(
		.INIT('h509c)
	) name9238 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15065_
	);
	LUT4 #(
		.INIT('h2000)
	) name9239 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15066_
	);
	LUT4 #(
		.INIT('h001b)
	) name9240 (
		_w14862_,
		_w14935_,
		_w15065_,
		_w15066_,
		_w15067_
	);
	LUT4 #(
		.INIT('h0200)
	) name9241 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15068_
	);
	LUT4 #(
		.INIT('h1008)
	) name9242 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15069_
	);
	LUT4 #(
		.INIT('hedf6)
	) name9243 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15070_
	);
	LUT2 #(
		.INIT('h2)
	) name9244 (
		_w14862_,
		_w15070_,
		_w15071_
	);
	LUT2 #(
		.INIT('h8)
	) name9245 (
		_w14860_,
		_w14868_,
		_w15072_
	);
	LUT4 #(
		.INIT('h23af)
	) name9246 (
		_w14862_,
		_w14863_,
		_w15062_,
		_w15072_,
		_w15073_
	);
	LUT4 #(
		.INIT('h0d00)
	) name9247 (
		_w14868_,
		_w15067_,
		_w15071_,
		_w15073_,
		_w15074_
	);
	LUT3 #(
		.INIT('h9a)
	) name9248 (
		\u2_desIn_r_reg[38]/NET0131 ,
		_w15064_,
		_w15074_,
		_w15075_
	);
	LUT3 #(
		.INIT('h01)
	) name9249 (
		_w14974_,
		_w14971_,
		_w14973_,
		_w15076_
	);
	LUT4 #(
		.INIT('hdf00)
	) name9250 (
		_w14971_,
		_w14972_,
		_w14973_,
		_w14970_,
		_w15077_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9251 (
		_w15017_,
		_w15011_,
		_w15076_,
		_w15077_,
		_w15078_
	);
	LUT4 #(
		.INIT('h0002)
	) name9252 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15079_
	);
	LUT4 #(
		.INIT('h0002)
	) name9253 (
		_w14969_,
		_w15008_,
		_w15009_,
		_w15079_,
		_w15080_
	);
	LUT4 #(
		.INIT('h0600)
	) name9254 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15081_
	);
	LUT4 #(
		.INIT('h0010)
	) name9255 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15082_
	);
	LUT2 #(
		.INIT('h1)
	) name9256 (
		_w14970_,
		_w14969_,
		_w15083_
	);
	LUT4 #(
		.INIT('h0100)
	) name9257 (
		_w14982_,
		_w15082_,
		_w15081_,
		_w15083_,
		_w15084_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name9258 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15085_
	);
	LUT4 #(
		.INIT('hf400)
	) name9259 (
		_w15078_,
		_w15080_,
		_w15084_,
		_w15085_,
		_w15086_
	);
	LUT4 #(
		.INIT('h1321)
	) name9260 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15087_
	);
	LUT4 #(
		.INIT('hc044)
	) name9261 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15088_
	);
	LUT2 #(
		.INIT('h2)
	) name9262 (
		_w14970_,
		_w14969_,
		_w15089_
	);
	LUT3 #(
		.INIT('h10)
	) name9263 (
		_w15087_,
		_w15088_,
		_w15089_,
		_w15090_
	);
	LUT3 #(
		.INIT('h56)
	) name9264 (
		\u2_desIn_r_reg[36]/NET0131 ,
		_w15086_,
		_w15090_,
		_w15091_
	);
	LUT4 #(
		.INIT('hcf7f)
	) name9265 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w15092_
	);
	LUT2 #(
		.INIT('h2)
	) name9266 (
		_w14685_,
		_w15092_,
		_w15093_
	);
	LUT3 #(
		.INIT('h07)
	) name9267 (
		_w14702_,
		_w14706_,
		_w14899_,
		_w15094_
	);
	LUT3 #(
		.INIT('h8a)
	) name9268 (
		_w14698_,
		_w15093_,
		_w15094_,
		_w15095_
	);
	LUT4 #(
		.INIT('h007f)
	) name9269 (
		_w14689_,
		_w14686_,
		_w14687_,
		_w14698_,
		_w15096_
	);
	LUT4 #(
		.INIT('h8008)
	) name9270 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w15097_
	);
	LUT4 #(
		.INIT('h1400)
	) name9271 (
		_w14689_,
		_w14686_,
		_w14687_,
		_w14698_,
		_w15098_
	);
	LUT4 #(
		.INIT('h0140)
	) name9272 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w15099_
	);
	LUT4 #(
		.INIT('h1011)
	) name9273 (
		_w15098_,
		_w15099_,
		_w15096_,
		_w15097_,
		_w15100_
	);
	LUT2 #(
		.INIT('h1)
	) name9274 (
		_w14685_,
		_w15100_,
		_w15101_
	);
	LUT3 #(
		.INIT('hd9)
	) name9275 (
		_w14689_,
		_w14686_,
		_w14687_,
		_w15102_
	);
	LUT2 #(
		.INIT('h2)
	) name9276 (
		_w14696_,
		_w15102_,
		_w15103_
	);
	LUT3 #(
		.INIT('h7e)
	) name9277 (
		_w14688_,
		_w14686_,
		_w14687_,
		_w15104_
	);
	LUT2 #(
		.INIT('h4)
	) name9278 (
		_w14703_,
		_w15104_,
		_w15105_
	);
	LUT4 #(
		.INIT('h0040)
	) name9279 (
		_w14689_,
		_w14685_,
		_w14686_,
		_w14687_,
		_w15106_
	);
	LUT4 #(
		.INIT('h2220)
	) name9280 (
		_w14689_,
		_w14685_,
		_w14686_,
		_w14687_,
		_w15107_
	);
	LUT3 #(
		.INIT('h23)
	) name9281 (
		_w14713_,
		_w15106_,
		_w15107_,
		_w15108_
	);
	LUT4 #(
		.INIT('h3222)
	) name9282 (
		_w14698_,
		_w15103_,
		_w15105_,
		_w15108_,
		_w15109_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name9283 (
		\u2_desIn_r_reg[50]/NET0131 ,
		_w15101_,
		_w15095_,
		_w15109_,
		_w15110_
	);
	LUT4 #(
		.INIT('hb5ae)
	) name9284 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15111_
	);
	LUT2 #(
		.INIT('h2)
	) name9285 (
		_w14657_,
		_w15111_,
		_w15112_
	);
	LUT4 #(
		.INIT('h4000)
	) name9286 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15113_
	);
	LUT4 #(
		.INIT('hee70)
	) name9287 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15114_
	);
	LUT4 #(
		.INIT('h0009)
	) name9288 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15115_
	);
	LUT4 #(
		.INIT('h3332)
	) name9289 (
		_w14657_,
		_w15113_,
		_w15115_,
		_w15114_,
		_w15116_
	);
	LUT3 #(
		.INIT('h8a)
	) name9290 (
		_w14656_,
		_w15112_,
		_w15116_,
		_w15117_
	);
	LUT4 #(
		.INIT('h0800)
	) name9291 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15118_
	);
	LUT4 #(
		.INIT('h00bf)
	) name9292 (
		_w14660_,
		_w14658_,
		_w14661_,
		_w14657_,
		_w15119_
	);
	LUT4 #(
		.INIT('hafac)
	) name9293 (
		_w14668_,
		_w14676_,
		_w14657_,
		_w15118_,
		_w15120_
	);
	LUT3 #(
		.INIT('h04)
	) name9294 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w15121_
	);
	LUT4 #(
		.INIT('hfb73)
	) name9295 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15122_
	);
	LUT3 #(
		.INIT('ha2)
	) name9296 (
		_w14678_,
		_w14657_,
		_w15122_,
		_w15123_
	);
	LUT4 #(
		.INIT('h8400)
	) name9297 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15124_
	);
	LUT3 #(
		.INIT('h0d)
	) name9298 (
		_w14821_,
		_w15121_,
		_w15124_,
		_w15125_
	);
	LUT4 #(
		.INIT('h3222)
	) name9299 (
		_w14656_,
		_w15120_,
		_w15123_,
		_w15125_,
		_w15126_
	);
	LUT3 #(
		.INIT('h65)
	) name9300 (
		\u2_desIn_r_reg[56]/NET0131 ,
		_w15117_,
		_w15126_,
		_w15127_
	);
	LUT4 #(
		.INIT('hc693)
	) name9301 (
		decrypt_pad,
		\u2_desIn_r_reg[29]/NET0131 ,
		\u2_key_r_reg[10]/NET0131 ,
		\u2_key_r_reg[17]/NET0131 ,
		_w15128_
	);
	LUT4 #(
		.INIT('hc693)
	) name9302 (
		decrypt_pad,
		\u2_desIn_r_reg[37]/NET0131 ,
		\u2_key_r_reg[55]/NET0131 ,
		\u2_key_r_reg[5]/NET0131 ,
		_w15129_
	);
	LUT4 #(
		.INIT('hc693)
	) name9303 (
		decrypt_pad,
		\u2_desIn_r_reg[63]/NET0131 ,
		\u2_key_r_reg[46]/NET0131 ,
		\u2_key_r_reg[53]/NET0131 ,
		_w15130_
	);
	LUT2 #(
		.INIT('h6)
	) name9304 (
		_w15129_,
		_w15130_,
		_w15131_
	);
	LUT4 #(
		.INIT('hc693)
	) name9305 (
		decrypt_pad,
		\u2_desIn_r_reg[5]/NET0131 ,
		\u2_key_r_reg[18]/NET0131 ,
		\u2_key_r_reg[25]/NET0131 ,
		_w15132_
	);
	LUT4 #(
		.INIT('hc693)
	) name9306 (
		decrypt_pad,
		\u2_desIn_r_reg[13]/NET0131 ,
		\u2_key_r_reg[26]/NET0131 ,
		\u2_key_r_reg[33]/NET0131 ,
		_w15133_
	);
	LUT4 #(
		.INIT('h2100)
	) name9307 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15134_
	);
	LUT3 #(
		.INIT('h08)
	) name9308 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15135_
	);
	LUT4 #(
		.INIT('hc693)
	) name9309 (
		decrypt_pad,
		\u2_desIn_r_reg[21]/NET0131 ,
		\u2_key_r_reg[27]/NET0131 ,
		\u2_key_r_reg[34]/NET0131 ,
		_w15136_
	);
	LUT2 #(
		.INIT('h2)
	) name9310 (
		_w15133_,
		_w15136_,
		_w15137_
	);
	LUT3 #(
		.INIT('h40)
	) name9311 (
		_w15129_,
		_w15132_,
		_w15133_,
		_w15138_
	);
	LUT4 #(
		.INIT('h4000)
	) name9312 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15139_
	);
	LUT4 #(
		.INIT('h0007)
	) name9313 (
		_w15135_,
		_w15137_,
		_w15139_,
		_w15134_,
		_w15140_
	);
	LUT2 #(
		.INIT('h8)
	) name9314 (
		_w15129_,
		_w15136_,
		_w15141_
	);
	LUT3 #(
		.INIT('h46)
	) name9315 (
		_w15129_,
		_w15130_,
		_w15136_,
		_w15142_
	);
	LUT2 #(
		.INIT('h1)
	) name9316 (
		_w15132_,
		_w15133_,
		_w15143_
	);
	LUT2 #(
		.INIT('h8)
	) name9317 (
		_w15143_,
		_w15142_,
		_w15144_
	);
	LUT3 #(
		.INIT('hed)
	) name9318 (
		_w15132_,
		_w15133_,
		_w15142_,
		_w15145_
	);
	LUT3 #(
		.INIT('h15)
	) name9319 (
		_w15128_,
		_w15140_,
		_w15145_,
		_w15146_
	);
	LUT4 #(
		.INIT('h959d)
	) name9320 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15147_
	);
	LUT4 #(
		.INIT('h0001)
	) name9321 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15148_
	);
	LUT4 #(
		.INIT('hddfe)
	) name9322 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15149_
	);
	LUT4 #(
		.INIT('h4f00)
	) name9323 (
		_w15147_,
		_w15128_,
		_w15149_,
		_w15136_,
		_w15150_
	);
	LUT2 #(
		.INIT('h8)
	) name9324 (
		_w15133_,
		_w15128_,
		_w15151_
	);
	LUT3 #(
		.INIT('h04)
	) name9325 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15152_
	);
	LUT2 #(
		.INIT('h2)
	) name9326 (
		_w15128_,
		_w15136_,
		_w15153_
	);
	LUT3 #(
		.INIT('h80)
	) name9327 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15154_
	);
	LUT4 #(
		.INIT('h6f67)
	) name9328 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15155_
	);
	LUT4 #(
		.INIT('h7707)
	) name9329 (
		_w15151_,
		_w15152_,
		_w15153_,
		_w15155_,
		_w15156_
	);
	LUT2 #(
		.INIT('h4)
	) name9330 (
		_w15150_,
		_w15156_,
		_w15157_
	);
	LUT3 #(
		.INIT('h65)
	) name9331 (
		\u2_desIn_r_reg[46]/NET0131 ,
		_w15146_,
		_w15157_,
		_w15158_
	);
	LUT3 #(
		.INIT('h60)
	) name9332 (
		_w14659_,
		_w14660_,
		_w14661_,
		_w15159_
	);
	LUT4 #(
		.INIT('h6080)
	) name9333 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15160_
	);
	LUT4 #(
		.INIT('h0908)
	) name9334 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15161_
	);
	LUT2 #(
		.INIT('h2)
	) name9335 (
		_w14657_,
		_w15161_,
		_w15162_
	);
	LUT4 #(
		.INIT('hbfbc)
	) name9336 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15163_
	);
	LUT3 #(
		.INIT('h20)
	) name9337 (
		_w15119_,
		_w15159_,
		_w15163_,
		_w15164_
	);
	LUT4 #(
		.INIT('h888a)
	) name9338 (
		_w14656_,
		_w15160_,
		_w15162_,
		_w15164_,
		_w15165_
	);
	LUT2 #(
		.INIT('h2)
	) name9339 (
		_w14656_,
		_w14672_,
		_w15166_
	);
	LUT4 #(
		.INIT('h0989)
	) name9340 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15167_
	);
	LUT4 #(
		.INIT('h6000)
	) name9341 (
		_w14659_,
		_w14660_,
		_w14658_,
		_w14661_,
		_w15168_
	);
	LUT3 #(
		.INIT('h02)
	) name9342 (
		_w14657_,
		_w15168_,
		_w15167_,
		_w15169_
	);
	LUT2 #(
		.INIT('h4)
	) name9343 (
		_w14657_,
		_w15160_,
		_w15170_
	);
	LUT4 #(
		.INIT('h3130)
	) name9344 (
		_w14657_,
		_w14656_,
		_w14672_,
		_w15161_,
		_w15171_
	);
	LUT4 #(
		.INIT('h1011)
	) name9345 (
		_w15170_,
		_w15171_,
		_w15166_,
		_w15169_,
		_w15172_
	);
	LUT3 #(
		.INIT('h65)
	) name9346 (
		\u2_desIn_r_reg[54]/NET0131 ,
		_w15165_,
		_w15172_,
		_w15173_
	);
	LUT4 #(
		.INIT('hdd75)
	) name9347 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15174_
	);
	LUT4 #(
		.INIT('h77fb)
	) name9348 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15175_
	);
	LUT4 #(
		.INIT('hbcef)
	) name9349 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15176_
	);
	LUT4 #(
		.INIT('hd800)
	) name9350 (
		_w14827_,
		_w15175_,
		_w15174_,
		_w15176_,
		_w15177_
	);
	LUT4 #(
		.INIT('h0001)
	) name9351 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15178_
	);
	LUT4 #(
		.INIT('hff76)
	) name9352 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15179_
	);
	LUT3 #(
		.INIT('h02)
	) name9353 (
		_w14829_,
		_w14826_,
		_w14827_,
		_w15180_
	);
	LUT4 #(
		.INIT('h00c4)
	) name9354 (
		_w14827_,
		_w14855_,
		_w15179_,
		_w15180_,
		_w15181_
	);
	LUT4 #(
		.INIT('hadff)
	) name9355 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15182_
	);
	LUT4 #(
		.INIT('he4ee)
	) name9356 (
		_w14827_,
		_w14838_,
		_w14854_,
		_w15182_,
		_w15183_
	);
	LUT4 #(
		.INIT('h0d08)
	) name9357 (
		_w14825_,
		_w15181_,
		_w15183_,
		_w15177_,
		_w15184_
	);
	LUT2 #(
		.INIT('h9)
	) name9358 (
		\u2_desIn_r_reg[62]/NET0131 ,
		_w15184_,
		_w15185_
	);
	LUT4 #(
		.INIT('hf700)
	) name9359 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15186_
	);
	LUT4 #(
		.INIT('h0400)
	) name9360 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15136_,
		_w15187_
	);
	LUT4 #(
		.INIT('h006d)
	) name9361 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15188_
	);
	LUT3 #(
		.INIT('h45)
	) name9362 (
		_w15186_,
		_w15187_,
		_w15188_,
		_w15189_
	);
	LUT4 #(
		.INIT('h0100)
	) name9363 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15190_
	);
	LUT3 #(
		.INIT('h14)
	) name9364 (
		_w15129_,
		_w15130_,
		_w15133_,
		_w15191_
	);
	LUT4 #(
		.INIT('hfd00)
	) name9365 (
		_w15136_,
		_w15139_,
		_w15190_,
		_w15191_,
		_w15192_
	);
	LUT3 #(
		.INIT('ha8)
	) name9366 (
		_w15128_,
		_w15189_,
		_w15192_,
		_w15193_
	);
	LUT3 #(
		.INIT('h40)
	) name9367 (
		_w15132_,
		_w15130_,
		_w15133_,
		_w15194_
	);
	LUT4 #(
		.INIT('h00bf)
	) name9368 (
		_w15132_,
		_w15130_,
		_w15133_,
		_w15136_,
		_w15195_
	);
	LUT4 #(
		.INIT('h00fd)
	) name9369 (
		_w15136_,
		_w15139_,
		_w15190_,
		_w15195_,
		_w15196_
	);
	LUT4 #(
		.INIT('h7d78)
	) name9370 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15197_
	);
	LUT3 #(
		.INIT('he0)
	) name9371 (
		_w15129_,
		_w15130_,
		_w15136_,
		_w15198_
	);
	LUT4 #(
		.INIT('h6800)
	) name9372 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15136_,
		_w15199_
	);
	LUT4 #(
		.INIT('h0504)
	) name9373 (
		_w15148_,
		_w15136_,
		_w15199_,
		_w15197_,
		_w15200_
	);
	LUT3 #(
		.INIT('h32)
	) name9374 (
		_w15128_,
		_w15196_,
		_w15200_,
		_w15201_
	);
	LUT3 #(
		.INIT('h65)
	) name9375 (
		\u2_desIn_r_reg[60]/NET0131 ,
		_w15193_,
		_w15201_,
		_w15202_
	);
	LUT2 #(
		.INIT('h4)
	) name9376 (
		_w15133_,
		_w15136_,
		_w15203_
	);
	LUT3 #(
		.INIT('h31)
	) name9377 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15204_
	);
	LUT2 #(
		.INIT('h8)
	) name9378 (
		_w15203_,
		_w15204_,
		_w15205_
	);
	LUT3 #(
		.INIT('h0e)
	) name9379 (
		_w15132_,
		_w15133_,
		_w15136_,
		_w15206_
	);
	LUT3 #(
		.INIT('hb0)
	) name9380 (
		_w15132_,
		_w15130_,
		_w15133_,
		_w15207_
	);
	LUT4 #(
		.INIT('h23af)
	) name9381 (
		_w15131_,
		_w15198_,
		_w15206_,
		_w15207_,
		_w15208_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9382 (
		_w15128_,
		_w15144_,
		_w15205_,
		_w15208_,
		_w15209_
	);
	LUT4 #(
		.INIT('hcaf1)
	) name9383 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15210_
	);
	LUT4 #(
		.INIT('h1000)
	) name9384 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15211_
	);
	LUT4 #(
		.INIT('h5504)
	) name9385 (
		_w15128_,
		_w15136_,
		_w15210_,
		_w15211_,
		_w15212_
	);
	LUT4 #(
		.INIT('h0021)
	) name9386 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15213_
	);
	LUT4 #(
		.INIT('hb59e)
	) name9387 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15214_
	);
	LUT2 #(
		.INIT('h1)
	) name9388 (
		_w15128_,
		_w15136_,
		_w15215_
	);
	LUT2 #(
		.INIT('h4)
	) name9389 (
		_w15214_,
		_w15215_,
		_w15216_
	);
	LUT3 #(
		.INIT('he7)
	) name9390 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15217_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name9391 (
		_w15133_,
		_w15136_,
		_w15154_,
		_w15217_,
		_w15218_
	);
	LUT3 #(
		.INIT('h10)
	) name9392 (
		_w15212_,
		_w15216_,
		_w15218_,
		_w15219_
	);
	LUT3 #(
		.INIT('h65)
	) name9393 (
		\u2_desIn_r_reg[58]/NET0131 ,
		_w15209_,
		_w15219_,
		_w15220_
	);
	LUT4 #(
		.INIT('h8090)
	) name9394 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15221_
	);
	LUT3 #(
		.INIT('h9f)
	) name9395 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w15222_
	);
	LUT4 #(
		.INIT('he4f5)
	) name9396 (
		_w14862_,
		_w14935_,
		_w15221_,
		_w15222_,
		_w15223_
	);
	LUT4 #(
		.INIT('hdbf5)
	) name9397 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15224_
	);
	LUT3 #(
		.INIT('h8a)
	) name9398 (
		_w14868_,
		_w15223_,
		_w15224_,
		_w15225_
	);
	LUT4 #(
		.INIT('hba0a)
	) name9399 (
		_w14858_,
		_w14860_,
		_w14861_,
		_w14859_,
		_w15226_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9400 (
		_w14862_,
		_w14858_,
		_w14861_,
		_w14859_,
		_w15227_
	);
	LUT2 #(
		.INIT('h4)
	) name9401 (
		_w15226_,
		_w15227_,
		_w15228_
	);
	LUT4 #(
		.INIT('h4000)
	) name9402 (
		_w14862_,
		_w14858_,
		_w14860_,
		_w14859_,
		_w15229_
	);
	LUT3 #(
		.INIT('h01)
	) name9403 (
		_w14932_,
		_w15068_,
		_w15229_,
		_w15230_
	);
	LUT4 #(
		.INIT('h0200)
	) name9404 (
		_w14862_,
		_w14858_,
		_w14861_,
		_w14859_,
		_w15231_
	);
	LUT4 #(
		.INIT('h00ab)
	) name9405 (
		_w14862_,
		_w15062_,
		_w15069_,
		_w15231_,
		_w15232_
	);
	LUT4 #(
		.INIT('hba00)
	) name9406 (
		_w14868_,
		_w15228_,
		_w15230_,
		_w15232_,
		_w15233_
	);
	LUT3 #(
		.INIT('h65)
	) name9407 (
		\u2_desIn_r_reg[16]/NET0131 ,
		_w15225_,
		_w15233_,
		_w15234_
	);
	LUT4 #(
		.INIT('hfae5)
	) name9408 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15235_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name9409 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15236_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name9410 (
		_w15128_,
		_w15138_,
		_w15235_,
		_w15236_,
		_w15237_
	);
	LUT2 #(
		.INIT('h2)
	) name9411 (
		_w15136_,
		_w15237_,
		_w15238_
	);
	LUT4 #(
		.INIT('h0200)
	) name9412 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15239_
	);
	LUT3 #(
		.INIT('h0e)
	) name9413 (
		_w15132_,
		_w15130_,
		_w15136_,
		_w15240_
	);
	LUT4 #(
		.INIT('h0015)
	) name9414 (
		_w15213_,
		_w15236_,
		_w15240_,
		_w15239_,
		_w15241_
	);
	LUT2 #(
		.INIT('h1)
	) name9415 (
		_w15128_,
		_w15241_,
		_w15242_
	);
	LUT4 #(
		.INIT('h0bfb)
	) name9416 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15133_,
		_w15243_
	);
	LUT2 #(
		.INIT('h2)
	) name9417 (
		_w15153_,
		_w15243_,
		_w15244_
	);
	LUT3 #(
		.INIT('h4c)
	) name9418 (
		_w15129_,
		_w15132_,
		_w15130_,
		_w15245_
	);
	LUT2 #(
		.INIT('h8)
	) name9419 (
		_w15151_,
		_w15245_,
		_w15246_
	);
	LUT4 #(
		.INIT('h0040)
	) name9420 (
		_w15129_,
		_w15132_,
		_w15133_,
		_w15136_,
		_w15247_
	);
	LUT3 #(
		.INIT('h07)
	) name9421 (
		_w15141_,
		_w15194_,
		_w15247_,
		_w15248_
	);
	LUT3 #(
		.INIT('h10)
	) name9422 (
		_w15244_,
		_w15246_,
		_w15248_,
		_w15249_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name9423 (
		\u2_desIn_r_reg[40]/NET0131 ,
		_w15238_,
		_w15242_,
		_w15249_,
		_w15250_
	);
	LUT3 #(
		.INIT('h04)
	) name9424 (
		_w14848_,
		_w14825_,
		_w14838_,
		_w15251_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name9425 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15252_
	);
	LUT3 #(
		.INIT('hb0)
	) name9426 (
		_w14828_,
		_w14829_,
		_w14827_,
		_w15253_
	);
	LUT3 #(
		.INIT('h45)
	) name9427 (
		_w14831_,
		_w15252_,
		_w15253_,
		_w15254_
	);
	LUT4 #(
		.INIT('hb9fd)
	) name9428 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15255_
	);
	LUT2 #(
		.INIT('h2)
	) name9429 (
		_w14827_,
		_w15255_,
		_w15256_
	);
	LUT3 #(
		.INIT('hd0)
	) name9430 (
		_w14826_,
		_w14830_,
		_w14827_,
		_w15257_
	);
	LUT4 #(
		.INIT('h4e46)
	) name9431 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15258_
	);
	LUT3 #(
		.INIT('h54)
	) name9432 (
		_w14825_,
		_w15257_,
		_w15258_,
		_w15259_
	);
	LUT4 #(
		.INIT('h7077)
	) name9433 (
		_w15251_,
		_w15254_,
		_w15256_,
		_w15259_,
		_w15260_
	);
	LUT3 #(
		.INIT('h02)
	) name9434 (
		_w14827_,
		_w14847_,
		_w14854_,
		_w15261_
	);
	LUT4 #(
		.INIT('h0080)
	) name9435 (
		_w14828_,
		_w14829_,
		_w14826_,
		_w14830_,
		_w15262_
	);
	LUT4 #(
		.INIT('h0001)
	) name9436 (
		_w14827_,
		_w14852_,
		_w15178_,
		_w15262_,
		_w15263_
	);
	LUT2 #(
		.INIT('h1)
	) name9437 (
		_w15261_,
		_w15263_,
		_w15264_
	);
	LUT3 #(
		.INIT('h56)
	) name9438 (
		\u2_desIn_r_reg[22]/NET0131 ,
		_w15260_,
		_w15264_,
		_w15265_
	);
	LUT4 #(
		.INIT('h0802)
	) name9439 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w15266_
	);
	LUT4 #(
		.INIT('h4000)
	) name9440 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w15267_
	);
	LUT3 #(
		.INIT('h01)
	) name9441 (
		_w14698_,
		_w15266_,
		_w15267_,
		_w15268_
	);
	LUT3 #(
		.INIT('hbc)
	) name9442 (
		_w14689_,
		_w14686_,
		_w14687_,
		_w15269_
	);
	LUT4 #(
		.INIT('h1003)
	) name9443 (
		_w14689_,
		_w14685_,
		_w14686_,
		_w14687_,
		_w15270_
	);
	LUT4 #(
		.INIT('hf04f)
	) name9444 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w15271_
	);
	LUT3 #(
		.INIT('h31)
	) name9445 (
		_w14685_,
		_w15270_,
		_w15271_,
		_w15272_
	);
	LUT4 #(
		.INIT('h8228)
	) name9446 (
		_w14688_,
		_w14689_,
		_w14686_,
		_w14687_,
		_w15273_
	);
	LUT4 #(
		.INIT('h0c04)
	) name9447 (
		_w14696_,
		_w14698_,
		_w14902_,
		_w15269_,
		_w15274_
	);
	LUT4 #(
		.INIT('h7077)
	) name9448 (
		_w15268_,
		_w15272_,
		_w15273_,
		_w15274_,
		_w15275_
	);
	LUT3 #(
		.INIT('h40)
	) name9449 (
		_w14685_,
		_w14686_,
		_w14687_,
		_w15276_
	);
	LUT2 #(
		.INIT('h4)
	) name9450 (
		_w14692_,
		_w15276_,
		_w15277_
	);
	LUT3 #(
		.INIT('h56)
	) name9451 (
		\u2_desIn_r_reg[4]/NET0131 ,
		_w15275_,
		_w15277_,
		_w15278_
	);
	LUT4 #(
		.INIT('h1a00)
	) name9452 (
		_w14974_,
		_w14972_,
		_w14973_,
		_w14970_,
		_w15279_
	);
	LUT4 #(
		.INIT('hcfaf)
	) name9453 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15280_
	);
	LUT4 #(
		.INIT('h0032)
	) name9454 (
		_w14970_,
		_w15018_,
		_w15280_,
		_w15279_,
		_w15281_
	);
	LUT4 #(
		.INIT('hbf6e)
	) name9455 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15282_
	);
	LUT4 #(
		.INIT('h8000)
	) name9456 (
		_w14974_,
		_w14972_,
		_w14973_,
		_w14970_,
		_w15283_
	);
	LUT4 #(
		.INIT('h0109)
	) name9457 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14970_,
		_w15284_
	);
	LUT3 #(
		.INIT('h10)
	) name9458 (
		_w15283_,
		_w15284_,
		_w15282_,
		_w15285_
	);
	LUT4 #(
		.INIT('h0020)
	) name9459 (
		_w14974_,
		_w14972_,
		_w14973_,
		_w14970_,
		_w15286_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name9460 (
		_w14974_,
		_w14971_,
		_w14972_,
		_w14973_,
		_w15287_
	);
	LUT3 #(
		.INIT('h31)
	) name9461 (
		_w14970_,
		_w15286_,
		_w15287_,
		_w15288_
	);
	LUT4 #(
		.INIT('hd800)
	) name9462 (
		_w14969_,
		_w15281_,
		_w15285_,
		_w15288_,
		_w15289_
	);
	LUT2 #(
		.INIT('h9)
	) name9463 (
		\u2_desIn_r_reg[10]/P0001 ,
		_w15289_,
		_w15290_
	);
	LUT4 #(
		.INIT('hc963)
	) name9464 (
		decrypt_pad,
		\u1_R14_reg[31]/P0001 ,
		\u1_uk_K_r14_reg[1]/NET0131 ,
		\u1_uk_K_r14_reg[49]/NET0131 ,
		_w15291_
	);
	LUT4 #(
		.INIT('hc693)
	) name9465 (
		decrypt_pad,
		\u1_R14_reg[29]/NET0131 ,
		\u1_uk_K_r14_reg[36]/NET0131 ,
		\u1_uk_K_r14_reg[43]/NET0131 ,
		_w15292_
	);
	LUT4 #(
		.INIT('hc693)
	) name9466 (
		decrypt_pad,
		\u1_R14_reg[1]/NET0131 ,
		\u1_uk_K_r14_reg[21]/NET0131 ,
		\u1_uk_K_r14_reg[28]/NET0131 ,
		_w15293_
	);
	LUT4 #(
		.INIT('hc693)
	) name9467 (
		decrypt_pad,
		\u1_R14_reg[30]/NET0131 ,
		\u1_uk_K_r14_reg[37]/NET0131 ,
		\u1_uk_K_r14_reg[44]/NET0131 ,
		_w15294_
	);
	LUT4 #(
		.INIT('hc963)
	) name9468 (
		decrypt_pad,
		\u1_R14_reg[28]/NET0131 ,
		\u1_uk_K_r14_reg[16]/NET0131 ,
		\u1_uk_K_r14_reg[9]/NET0131 ,
		_w15295_
	);
	LUT4 #(
		.INIT('h5b59)
	) name9469 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w15296_
	);
	LUT2 #(
		.INIT('h2)
	) name9470 (
		_w15295_,
		_w15294_,
		_w15297_
	);
	LUT4 #(
		.INIT('h0010)
	) name9471 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w15298_
	);
	LUT4 #(
		.INIT('hc693)
	) name9472 (
		decrypt_pad,
		\u1_R14_reg[32]/NET0131 ,
		\u1_uk_K_r14_reg[0]/P0001 ,
		\u1_uk_K_r14_reg[7]/NET0131 ,
		_w15299_
	);
	LUT4 #(
		.INIT('h000d)
	) name9473 (
		_w15291_,
		_w15296_,
		_w15298_,
		_w15299_,
		_w15300_
	);
	LUT2 #(
		.INIT('h2)
	) name9474 (
		_w15292_,
		_w15294_,
		_w15301_
	);
	LUT4 #(
		.INIT('hf700)
	) name9475 (
		_w15292_,
		_w15295_,
		_w15294_,
		_w15299_,
		_w15302_
	);
	LUT4 #(
		.INIT('h0002)
	) name9476 (
		_w15291_,
		_w15292_,
		_w15293_,
		_w15295_,
		_w15303_
	);
	LUT4 #(
		.INIT('h1000)
	) name9477 (
		_w15291_,
		_w15292_,
		_w15293_,
		_w15294_,
		_w15304_
	);
	LUT4 #(
		.INIT('h0200)
	) name9478 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w15305_
	);
	LUT4 #(
		.INIT('h4000)
	) name9479 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w15306_
	);
	LUT4 #(
		.INIT('hbdff)
	) name9480 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w15307_
	);
	LUT4 #(
		.INIT('h1000)
	) name9481 (
		_w15303_,
		_w15304_,
		_w15302_,
		_w15307_,
		_w15308_
	);
	LUT2 #(
		.INIT('h1)
	) name9482 (
		_w15300_,
		_w15308_,
		_w15309_
	);
	LUT4 #(
		.INIT('h4555)
	) name9483 (
		_w15291_,
		_w15292_,
		_w15295_,
		_w15294_,
		_w15310_
	);
	LUT3 #(
		.INIT('h01)
	) name9484 (
		_w15292_,
		_w15295_,
		_w15294_,
		_w15311_
	);
	LUT4 #(
		.INIT('h0001)
	) name9485 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w15312_
	);
	LUT4 #(
		.INIT('hfff6)
	) name9486 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w15313_
	);
	LUT3 #(
		.INIT('h40)
	) name9487 (
		_w15305_,
		_w15310_,
		_w15313_,
		_w15314_
	);
	LUT4 #(
		.INIT('h0004)
	) name9488 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w15315_
	);
	LUT4 #(
		.INIT('h0800)
	) name9489 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w15316_
	);
	LUT3 #(
		.INIT('h02)
	) name9490 (
		_w15291_,
		_w15316_,
		_w15315_,
		_w15317_
	);
	LUT4 #(
		.INIT('h0010)
	) name9491 (
		_w15291_,
		_w15292_,
		_w15295_,
		_w15299_,
		_w15318_
	);
	LUT3 #(
		.INIT('h0e)
	) name9492 (
		_w15314_,
		_w15317_,
		_w15318_,
		_w15319_
	);
	LUT3 #(
		.INIT('h65)
	) name9493 (
		\u1_L14_reg[15]/P0001 ,
		_w15309_,
		_w15319_,
		_w15320_
	);
	LUT4 #(
		.INIT('hc963)
	) name9494 (
		decrypt_pad,
		\u1_R14_reg[3]/NET0131 ,
		\u1_uk_K_r14_reg[3]/NET0131 ,
		\u1_uk_K_r14_reg[53]/NET0131 ,
		_w15321_
	);
	LUT4 #(
		.INIT('hc693)
	) name9495 (
		decrypt_pad,
		\u1_R14_reg[2]/NET0131 ,
		\u1_uk_K_r14_reg[19]/NET0131 ,
		\u1_uk_K_r14_reg[26]/NET0131 ,
		_w15322_
	);
	LUT4 #(
		.INIT('hc693)
	) name9496 (
		decrypt_pad,
		\u1_R14_reg[32]/NET0131 ,
		\u1_uk_K_r14_reg[40]/NET0131 ,
		\u1_uk_K_r14_reg[47]/NET0131 ,
		_w15323_
	);
	LUT4 #(
		.INIT('hc693)
	) name9497 (
		decrypt_pad,
		\u1_R14_reg[5]/NET0131 ,
		\u1_uk_K_r14_reg[34]/NET0131 ,
		\u1_uk_K_r14_reg[41]/NET0131 ,
		_w15324_
	);
	LUT4 #(
		.INIT('hc963)
	) name9498 (
		decrypt_pad,
		\u1_R14_reg[1]/NET0131 ,
		\u1_uk_K_r14_reg[11]/NET0131 ,
		\u1_uk_K_r14_reg[4]/NET0131 ,
		_w15325_
	);
	LUT2 #(
		.INIT('h1)
	) name9499 (
		_w15324_,
		_w15325_,
		_w15326_
	);
	LUT4 #(
		.INIT('h0200)
	) name9500 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w15327_
	);
	LUT2 #(
		.INIT('h1)
	) name9501 (
		_w15324_,
		_w15323_,
		_w15328_
	);
	LUT3 #(
		.INIT('h04)
	) name9502 (
		_w15324_,
		_w15325_,
		_w15323_,
		_w15329_
	);
	LUT4 #(
		.INIT('hfdc3)
	) name9503 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w15330_
	);
	LUT4 #(
		.INIT('hc963)
	) name9504 (
		decrypt_pad,
		\u1_R14_reg[4]/NET0131 ,
		\u1_uk_K_r14_reg[13]/NET0131 ,
		\u1_uk_K_r14_reg[6]/NET0131 ,
		_w15331_
	);
	LUT4 #(
		.INIT('h1000)
	) name9505 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w15332_
	);
	LUT4 #(
		.INIT('h6ffb)
	) name9506 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w15333_
	);
	LUT4 #(
		.INIT('h1055)
	) name9507 (
		_w15321_,
		_w15330_,
		_w15331_,
		_w15333_,
		_w15334_
	);
	LUT3 #(
		.INIT('h08)
	) name9508 (
		_w15321_,
		_w15322_,
		_w15323_,
		_w15335_
	);
	LUT4 #(
		.INIT('h4080)
	) name9509 (
		_w15321_,
		_w15322_,
		_w15324_,
		_w15323_,
		_w15336_
	);
	LUT4 #(
		.INIT('h0020)
	) name9510 (
		_w15321_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w15337_
	);
	LUT3 #(
		.INIT('h80)
	) name9511 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15338_
	);
	LUT4 #(
		.INIT('h007f)
	) name9512 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15331_,
		_w15339_
	);
	LUT3 #(
		.INIT('h01)
	) name9513 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15340_
	);
	LUT3 #(
		.INIT('h40)
	) name9514 (
		_w15321_,
		_w15325_,
		_w15323_,
		_w15341_
	);
	LUT4 #(
		.INIT('h0100)
	) name9515 (
		_w15340_,
		_w15337_,
		_w15341_,
		_w15339_,
		_w15342_
	);
	LUT4 #(
		.INIT('h2000)
	) name9516 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w15343_
	);
	LUT4 #(
		.INIT('hdf3f)
	) name9517 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w15344_
	);
	LUT2 #(
		.INIT('h2)
	) name9518 (
		_w15321_,
		_w15344_,
		_w15345_
	);
	LUT4 #(
		.INIT('h0400)
	) name9519 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w15346_
	);
	LUT4 #(
		.INIT('h004c)
	) name9520 (
		_w15326_,
		_w15331_,
		_w15335_,
		_w15346_,
		_w15347_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9521 (
		_w15336_,
		_w15342_,
		_w15345_,
		_w15347_,
		_w15348_
	);
	LUT4 #(
		.INIT('h0200)
	) name9522 (
		_w15321_,
		_w15322_,
		_w15325_,
		_w15323_,
		_w15349_
	);
	LUT2 #(
		.INIT('h2)
	) name9523 (
		_w15321_,
		_w15322_,
		_w15350_
	);
	LUT3 #(
		.INIT('h13)
	) name9524 (
		_w15329_,
		_w15349_,
		_w15350_,
		_w15351_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name9525 (
		\u1_L14_reg[23]/P0001 ,
		_w15334_,
		_w15348_,
		_w15351_,
		_w15352_
	);
	LUT4 #(
		.INIT('hc693)
	) name9526 (
		decrypt_pad,
		\u1_R14_reg[12]/NET0131 ,
		\u1_uk_K_r14_reg[10]/P0001 ,
		\u1_uk_K_r14_reg[17]/NET0131 ,
		_w15353_
	);
	LUT4 #(
		.INIT('hc693)
	) name9527 (
		decrypt_pad,
		\u1_R14_reg[10]/P0001 ,
		\u1_uk_K_r14_reg[26]/NET0131 ,
		\u1_uk_K_r14_reg[33]/NET0131 ,
		_w15354_
	);
	LUT4 #(
		.INIT('hc693)
	) name9528 (
		decrypt_pad,
		\u1_R14_reg[8]/NET0131 ,
		\u1_uk_K_r14_reg[46]/NET0131 ,
		\u1_uk_K_r14_reg[53]/NET0131 ,
		_w15355_
	);
	LUT4 #(
		.INIT('hc693)
	) name9529 (
		decrypt_pad,
		\u1_R14_reg[13]/NET0131 ,
		\u1_uk_K_r14_reg[55]/NET0131 ,
		\u1_uk_K_r14_reg[5]/NET0131 ,
		_w15356_
	);
	LUT3 #(
		.INIT('heb)
	) name9530 (
		_w15355_,
		_w15356_,
		_w15354_,
		_w15357_
	);
	LUT4 #(
		.INIT('hc693)
	) name9531 (
		decrypt_pad,
		\u1_R14_reg[9]/NET0131 ,
		\u1_uk_K_r14_reg[18]/NET0131 ,
		\u1_uk_K_r14_reg[25]/NET0131 ,
		_w15358_
	);
	LUT4 #(
		.INIT('h0004)
	) name9532 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w15359_
	);
	LUT4 #(
		.INIT('hc693)
	) name9533 (
		decrypt_pad,
		\u1_R14_reg[11]/P0001 ,
		\u1_uk_K_r14_reg[27]/NET0131 ,
		\u1_uk_K_r14_reg[34]/NET0131 ,
		_w15360_
	);
	LUT3 #(
		.INIT('h40)
	) name9534 (
		_w15359_,
		_w15357_,
		_w15360_,
		_w15361_
	);
	LUT3 #(
		.INIT('h02)
	) name9535 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15362_
	);
	LUT3 #(
		.INIT('h07)
	) name9536 (
		_w15355_,
		_w15354_,
		_w15360_,
		_w15363_
	);
	LUT2 #(
		.INIT('h4)
	) name9537 (
		_w15362_,
		_w15363_,
		_w15364_
	);
	LUT3 #(
		.INIT('ha8)
	) name9538 (
		_w15353_,
		_w15361_,
		_w15364_,
		_w15365_
	);
	LUT4 #(
		.INIT('hc400)
	) name9539 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w15366_
	);
	LUT4 #(
		.INIT('hfd00)
	) name9540 (
		_w15358_,
		_w15356_,
		_w15354_,
		_w15360_,
		_w15367_
	);
	LUT4 #(
		.INIT('h00c4)
	) name9541 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w15368_
	);
	LUT3 #(
		.INIT('h20)
	) name9542 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15369_
	);
	LUT4 #(
		.INIT('h00df)
	) name9543 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15360_,
		_w15370_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9544 (
		_w15366_,
		_w15367_,
		_w15368_,
		_w15370_,
		_w15371_
	);
	LUT2 #(
		.INIT('h6)
	) name9545 (
		_w15355_,
		_w15356_,
		_w15372_
	);
	LUT4 #(
		.INIT('h0041)
	) name9546 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w15373_
	);
	LUT2 #(
		.INIT('h4)
	) name9547 (
		_w15358_,
		_w15356_,
		_w15374_
	);
	LUT4 #(
		.INIT('h1000)
	) name9548 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w15375_
	);
	LUT3 #(
		.INIT('h01)
	) name9549 (
		_w15353_,
		_w15375_,
		_w15373_,
		_w15376_
	);
	LUT2 #(
		.INIT('h4)
	) name9550 (
		_w15371_,
		_w15376_,
		_w15377_
	);
	LUT3 #(
		.INIT('h80)
	) name9551 (
		_w15355_,
		_w15354_,
		_w15360_,
		_w15378_
	);
	LUT2 #(
		.INIT('h8)
	) name9552 (
		_w15374_,
		_w15378_,
		_w15379_
	);
	LUT2 #(
		.INIT('h2)
	) name9553 (
		_w15354_,
		_w15360_,
		_w15380_
	);
	LUT4 #(
		.INIT('h0020)
	) name9554 (
		_w15358_,
		_w15356_,
		_w15354_,
		_w15360_,
		_w15381_
	);
	LUT3 #(
		.INIT('h2a)
	) name9555 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15382_
	);
	LUT2 #(
		.INIT('h8)
	) name9556 (
		_w15353_,
		_w15354_,
		_w15383_
	);
	LUT3 #(
		.INIT('h15)
	) name9557 (
		_w15381_,
		_w15382_,
		_w15383_,
		_w15384_
	);
	LUT2 #(
		.INIT('h4)
	) name9558 (
		_w15379_,
		_w15384_,
		_w15385_
	);
	LUT4 #(
		.INIT('h56aa)
	) name9559 (
		\u1_L14_reg[30]/P0001 ,
		_w15365_,
		_w15377_,
		_w15385_,
		_w15386_
	);
	LUT4 #(
		.INIT('hc693)
	) name9560 (
		decrypt_pad,
		\u1_R14_reg[8]/NET0131 ,
		\u1_uk_K_r14_reg[32]/NET0131 ,
		\u1_uk_K_r14_reg[39]/P0001 ,
		_w15387_
	);
	LUT4 #(
		.INIT('hc693)
	) name9561 (
		decrypt_pad,
		\u1_R14_reg[4]/NET0131 ,
		\u1_uk_K_r14_reg[20]/NET0131 ,
		\u1_uk_K_r14_reg[27]/NET0131 ,
		_w15388_
	);
	LUT4 #(
		.INIT('hc693)
	) name9562 (
		decrypt_pad,
		\u1_R14_reg[9]/NET0131 ,
		\u1_uk_K_r14_reg[12]/NET0131 ,
		\u1_uk_K_r14_reg[19]/NET0131 ,
		_w15389_
	);
	LUT2 #(
		.INIT('h8)
	) name9563 (
		_w15388_,
		_w15389_,
		_w15390_
	);
	LUT4 #(
		.INIT('hc693)
	) name9564 (
		decrypt_pad,
		\u1_R14_reg[5]/NET0131 ,
		\u1_uk_K_r14_reg[24]/NET0131 ,
		\u1_uk_K_r14_reg[6]/NET0131 ,
		_w15391_
	);
	LUT4 #(
		.INIT('hc693)
	) name9565 (
		decrypt_pad,
		\u1_R14_reg[6]/NET0131 ,
		\u1_uk_K_r14_reg[47]/NET0131 ,
		\u1_uk_K_r14_reg[54]/NET0131 ,
		_w15392_
	);
	LUT4 #(
		.INIT('hc693)
	) name9566 (
		decrypt_pad,
		\u1_R14_reg[7]/P0001 ,
		\u1_uk_K_r14_reg[41]/NET0131 ,
		\u1_uk_K_r14_reg[48]/NET0131 ,
		_w15393_
	);
	LUT3 #(
		.INIT('h47)
	) name9567 (
		_w15393_,
		_w15391_,
		_w15392_,
		_w15394_
	);
	LUT3 #(
		.INIT('h51)
	) name9568 (
		_w15388_,
		_w15391_,
		_w15392_,
		_w15395_
	);
	LUT2 #(
		.INIT('h8)
	) name9569 (
		_w15388_,
		_w15392_,
		_w15396_
	);
	LUT4 #(
		.INIT('h2000)
	) name9570 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w15397_
	);
	LUT4 #(
		.INIT('hdffc)
	) name9571 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w15398_
	);
	LUT4 #(
		.INIT('h1d00)
	) name9572 (
		_w15390_,
		_w15394_,
		_w15395_,
		_w15398_,
		_w15399_
	);
	LUT4 #(
		.INIT('h0a20)
	) name9573 (
		_w15393_,
		_w15388_,
		_w15389_,
		_w15391_,
		_w15400_
	);
	LUT2 #(
		.INIT('h8)
	) name9574 (
		_w15389_,
		_w15392_,
		_w15401_
	);
	LUT4 #(
		.INIT('h4044)
	) name9575 (
		_w15393_,
		_w15388_,
		_w15389_,
		_w15391_,
		_w15402_
	);
	LUT4 #(
		.INIT('h0100)
	) name9576 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w15403_
	);
	LUT4 #(
		.INIT('h000b)
	) name9577 (
		_w15401_,
		_w15402_,
		_w15400_,
		_w15403_,
		_w15404_
	);
	LUT4 #(
		.INIT('h0010)
	) name9578 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w15405_
	);
	LUT4 #(
		.INIT('h77ef)
	) name9579 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w15406_
	);
	LUT4 #(
		.INIT('h1000)
	) name9580 (
		_w15393_,
		_w15388_,
		_w15389_,
		_w15391_,
		_w15407_
	);
	LUT3 #(
		.INIT('h0d)
	) name9581 (
		_w15393_,
		_w15406_,
		_w15407_,
		_w15408_
	);
	LUT4 #(
		.INIT('hd800)
	) name9582 (
		_w15387_,
		_w15404_,
		_w15399_,
		_w15408_,
		_w15409_
	);
	LUT2 #(
		.INIT('h9)
	) name9583 (
		\u1_L14_reg[18]/P0001 ,
		_w15409_,
		_w15410_
	);
	LUT4 #(
		.INIT('hc963)
	) name9584 (
		decrypt_pad,
		\u1_R13_reg[4]/NET0131 ,
		\u1_uk_K_r13_reg[20]/NET0131 ,
		\u1_uk_K_r13_reg[24]/NET0131 ,
		_w15411_
	);
	LUT4 #(
		.INIT('hc963)
	) name9585 (
		decrypt_pad,
		\u1_R13_reg[3]/NET0131 ,
		\u1_uk_K_r13_reg[10]/NET0131 ,
		\u1_uk_K_r13_reg[46]/NET0131 ,
		_w15412_
	);
	LUT4 #(
		.INIT('hc693)
	) name9586 (
		decrypt_pad,
		\u1_R13_reg[32]/NET0131 ,
		\u1_uk_K_r13_reg[33]/NET0131 ,
		\u1_uk_K_r13_reg[54]/NET0131 ,
		_w15413_
	);
	LUT4 #(
		.INIT('hc693)
	) name9587 (
		decrypt_pad,
		\u1_R13_reg[5]/NET0131 ,
		\u1_uk_K_r13_reg[27]/NET0131 ,
		\u1_uk_K_r13_reg[48]/NET0131 ,
		_w15414_
	);
	LUT4 #(
		.INIT('hc963)
	) name9588 (
		decrypt_pad,
		\u1_R13_reg[1]/NET0131 ,
		\u1_uk_K_r13_reg[18]/NET0131 ,
		\u1_uk_K_r13_reg[54]/NET0131 ,
		_w15415_
	);
	LUT4 #(
		.INIT('hc693)
	) name9589 (
		decrypt_pad,
		\u1_R13_reg[2]/NET0131 ,
		\u1_uk_K_r13_reg[12]/NET0131 ,
		\u1_uk_K_r13_reg[33]/NET0131 ,
		_w15416_
	);
	LUT4 #(
		.INIT('h2000)
	) name9590 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15417_
	);
	LUT2 #(
		.INIT('h4)
	) name9591 (
		_w15416_,
		_w15413_,
		_w15418_
	);
	LUT3 #(
		.INIT('hb0)
	) name9592 (
		_w15412_,
		_w15415_,
		_w15414_,
		_w15419_
	);
	LUT4 #(
		.INIT('h0777)
	) name9593 (
		_w15412_,
		_w15417_,
		_w15418_,
		_w15419_,
		_w15420_
	);
	LUT4 #(
		.INIT('h0080)
	) name9594 (
		_w15412_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15421_
	);
	LUT4 #(
		.INIT('hff7c)
	) name9595 (
		_w15412_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15422_
	);
	LUT2 #(
		.INIT('h2)
	) name9596 (
		_w15415_,
		_w15422_,
		_w15423_
	);
	LUT3 #(
		.INIT('h8c)
	) name9597 (
		_w15415_,
		_w15416_,
		_w15413_,
		_w15424_
	);
	LUT2 #(
		.INIT('h4)
	) name9598 (
		_w15415_,
		_w15414_,
		_w15425_
	);
	LUT3 #(
		.INIT('h45)
	) name9599 (
		_w15412_,
		_w15416_,
		_w15413_,
		_w15426_
	);
	LUT3 #(
		.INIT('h04)
	) name9600 (
		_w15425_,
		_w15426_,
		_w15424_,
		_w15427_
	);
	LUT4 #(
		.INIT('h5455)
	) name9601 (
		_w15411_,
		_w15423_,
		_w15427_,
		_w15420_,
		_w15428_
	);
	LUT3 #(
		.INIT('h04)
	) name9602 (
		_w15414_,
		_w15416_,
		_w15413_,
		_w15429_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name9603 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15430_
	);
	LUT2 #(
		.INIT('h2)
	) name9604 (
		_w15412_,
		_w15430_,
		_w15431_
	);
	LUT3 #(
		.INIT('h01)
	) name9605 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15432_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name9606 (
		_w15412_,
		_w15415_,
		_w15414_,
		_w15416_,
		_w15433_
	);
	LUT2 #(
		.INIT('h2)
	) name9607 (
		_w15412_,
		_w15416_,
		_w15434_
	);
	LUT3 #(
		.INIT('hc4)
	) name9608 (
		_w15412_,
		_w15415_,
		_w15416_,
		_w15435_
	);
	LUT3 #(
		.INIT('h0e)
	) name9609 (
		_w15414_,
		_w15416_,
		_w15413_,
		_w15436_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9610 (
		_w15433_,
		_w15413_,
		_w15435_,
		_w15436_,
		_w15437_
	);
	LUT3 #(
		.INIT('h80)
	) name9611 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15438_
	);
	LUT4 #(
		.INIT('h7dbd)
	) name9612 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15439_
	);
	LUT2 #(
		.INIT('h2)
	) name9613 (
		_w15412_,
		_w15415_,
		_w15440_
	);
	LUT3 #(
		.INIT('hcb)
	) name9614 (
		_w15414_,
		_w15416_,
		_w15413_,
		_w15441_
	);
	LUT4 #(
		.INIT('hfad8)
	) name9615 (
		_w15412_,
		_w15415_,
		_w15439_,
		_w15441_,
		_w15442_
	);
	LUT4 #(
		.INIT('h4f00)
	) name9616 (
		_w15431_,
		_w15437_,
		_w15411_,
		_w15442_,
		_w15443_
	);
	LUT3 #(
		.INIT('h65)
	) name9617 (
		\u1_L13_reg[31]/NET0131 ,
		_w15428_,
		_w15443_,
		_w15444_
	);
	LUT4 #(
		.INIT('hc693)
	) name9618 (
		decrypt_pad,
		\u1_R13_reg[28]/NET0131 ,
		\u1_uk_K_r13_reg[28]/NET0131 ,
		\u1_uk_K_r13_reg[49]/NET0131 ,
		_w15445_
	);
	LUT4 #(
		.INIT('hc693)
	) name9619 (
		decrypt_pad,
		\u1_R13_reg[27]/P0001 ,
		\u1_uk_K_r13_reg[45]/NET0131 ,
		\u1_uk_K_r13_reg[7]/NET0131 ,
		_w15446_
	);
	LUT4 #(
		.INIT('hc963)
	) name9620 (
		decrypt_pad,
		\u1_R13_reg[26]/NET0131 ,
		\u1_uk_K_r13_reg[29]/NET0131 ,
		\u1_uk_K_r13_reg[8]/NET0131 ,
		_w15447_
	);
	LUT4 #(
		.INIT('hc963)
	) name9621 (
		decrypt_pad,
		\u1_R13_reg[29]/NET0131 ,
		\u1_uk_K_r13_reg[45]/NET0131 ,
		\u1_uk_K_r13_reg[51]/NET0131 ,
		_w15448_
	);
	LUT4 #(
		.INIT('hc693)
	) name9622 (
		decrypt_pad,
		\u1_R13_reg[24]/NET0131 ,
		\u1_uk_K_r13_reg[43]/NET0131 ,
		\u1_uk_K_r13_reg[9]/NET0131 ,
		_w15449_
	);
	LUT4 #(
		.INIT('hc693)
	) name9623 (
		decrypt_pad,
		\u1_R13_reg[25]/NET0131 ,
		\u1_uk_K_r13_reg[23]/NET0131 ,
		\u1_uk_K_r13_reg[44]/NET0131 ,
		_w15450_
	);
	LUT4 #(
		.INIT('h1bef)
	) name9624 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15451_
	);
	LUT2 #(
		.INIT('h1)
	) name9625 (
		_w15446_,
		_w15451_,
		_w15452_
	);
	LUT4 #(
		.INIT('hefe5)
	) name9626 (
		_w15448_,
		_w15450_,
		_w15449_,
		_w15446_,
		_w15453_
	);
	LUT4 #(
		.INIT('h8008)
	) name9627 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15454_
	);
	LUT2 #(
		.INIT('h8)
	) name9628 (
		_w15449_,
		_w15446_,
		_w15455_
	);
	LUT4 #(
		.INIT('h1000)
	) name9629 (
		_w15450_,
		_w15447_,
		_w15449_,
		_w15446_,
		_w15456_
	);
	LUT4 #(
		.INIT('h0032)
	) name9630 (
		_w15447_,
		_w15454_,
		_w15453_,
		_w15456_,
		_w15457_
	);
	LUT3 #(
		.INIT('h45)
	) name9631 (
		_w15445_,
		_w15452_,
		_w15457_,
		_w15458_
	);
	LUT2 #(
		.INIT('h4)
	) name9632 (
		_w15450_,
		_w15447_,
		_w15459_
	);
	LUT3 #(
		.INIT('hc7)
	) name9633 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15460_
	);
	LUT4 #(
		.INIT('h0020)
	) name9634 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15461_
	);
	LUT4 #(
		.INIT('hffde)
	) name9635 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15462_
	);
	LUT4 #(
		.INIT('h08aa)
	) name9636 (
		_w15445_,
		_w15455_,
		_w15460_,
		_w15462_,
		_w15463_
	);
	LUT3 #(
		.INIT('h82)
	) name9637 (
		_w15450_,
		_w15447_,
		_w15449_,
		_w15464_
	);
	LUT4 #(
		.INIT('h0200)
	) name9638 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15465_
	);
	LUT4 #(
		.INIT('hfd77)
	) name9639 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15466_
	);
	LUT4 #(
		.INIT('h3032)
	) name9640 (
		_w15445_,
		_w15446_,
		_w15464_,
		_w15466_,
		_w15467_
	);
	LUT4 #(
		.INIT('h0060)
	) name9641 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15468_
	);
	LUT4 #(
		.INIT('hee9e)
	) name9642 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15469_
	);
	LUT2 #(
		.INIT('h2)
	) name9643 (
		_w15446_,
		_w15469_,
		_w15470_
	);
	LUT3 #(
		.INIT('h01)
	) name9644 (
		_w15467_,
		_w15470_,
		_w15463_,
		_w15471_
	);
	LUT3 #(
		.INIT('h65)
	) name9645 (
		\u1_L13_reg[22]/NET0131 ,
		_w15458_,
		_w15471_,
		_w15472_
	);
	LUT4 #(
		.INIT('hc963)
	) name9646 (
		decrypt_pad,
		\u1_R13_reg[23]/P0001 ,
		\u1_uk_K_r13_reg[16]/NET0131 ,
		\u1_uk_K_r13_reg[50]/NET0131 ,
		_w15473_
	);
	LUT4 #(
		.INIT('hc963)
	) name9647 (
		decrypt_pad,
		\u1_R13_reg[22]/NET0131 ,
		\u1_uk_K_r13_reg[31]/NET0131 ,
		\u1_uk_K_r13_reg[37]/NET0131 ,
		_w15474_
	);
	LUT4 #(
		.INIT('hc693)
	) name9648 (
		decrypt_pad,
		\u1_R13_reg[20]/NET0131 ,
		\u1_uk_K_r13_reg[0]/NET0131 ,
		\u1_uk_K_r13_reg[21]/NET0131 ,
		_w15475_
	);
	LUT4 #(
		.INIT('hc693)
	) name9649 (
		decrypt_pad,
		\u1_R13_reg[21]/NET0131 ,
		\u1_uk_K_r13_reg[15]/NET0131 ,
		\u1_uk_K_r13_reg[36]/NET0131 ,
		_w15476_
	);
	LUT4 #(
		.INIT('hc693)
	) name9650 (
		decrypt_pad,
		\u1_R13_reg[25]/NET0131 ,
		\u1_uk_K_r13_reg[16]/NET0131 ,
		\u1_uk_K_r13_reg[37]/NET0131 ,
		_w15477_
	);
	LUT2 #(
		.INIT('h4)
	) name9651 (
		_w15476_,
		_w15477_,
		_w15478_
	);
	LUT4 #(
		.INIT('h16b0)
	) name9652 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15479_
	);
	LUT4 #(
		.INIT('hc693)
	) name9653 (
		decrypt_pad,
		\u1_R13_reg[24]/NET0131 ,
		\u1_uk_K_r13_reg[21]/NET0131 ,
		\u1_uk_K_r13_reg[42]/NET0131 ,
		_w15480_
	);
	LUT4 #(
		.INIT('hc842)
	) name9654 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15481_
	);
	LUT4 #(
		.INIT('hc480)
	) name9655 (
		_w15473_,
		_w15480_,
		_w15481_,
		_w15479_,
		_w15482_
	);
	LUT2 #(
		.INIT('h1)
	) name9656 (
		_w15473_,
		_w15474_,
		_w15483_
	);
	LUT3 #(
		.INIT('h02)
	) name9657 (
		_w15475_,
		_w15473_,
		_w15474_,
		_w15484_
	);
	LUT4 #(
		.INIT('hff75)
	) name9658 (
		_w15475_,
		_w15476_,
		_w15473_,
		_w15474_,
		_w15485_
	);
	LUT2 #(
		.INIT('h1)
	) name9659 (
		_w15477_,
		_w15485_,
		_w15486_
	);
	LUT4 #(
		.INIT('h0408)
	) name9660 (
		_w15475_,
		_w15476_,
		_w15473_,
		_w15474_,
		_w15487_
	);
	LUT3 #(
		.INIT('h04)
	) name9661 (
		_w15475_,
		_w15473_,
		_w15474_,
		_w15488_
	);
	LUT3 #(
		.INIT('h13)
	) name9662 (
		_w15475_,
		_w15473_,
		_w15477_,
		_w15489_
	);
	LUT4 #(
		.INIT('h3020)
	) name9663 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15490_
	);
	LUT4 #(
		.INIT('h0045)
	) name9664 (
		_w15488_,
		_w15489_,
		_w15490_,
		_w15487_,
		_w15491_
	);
	LUT3 #(
		.INIT('h45)
	) name9665 (
		_w15480_,
		_w15486_,
		_w15491_,
		_w15492_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name9666 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15493_
	);
	LUT4 #(
		.INIT('h8c0c)
	) name9667 (
		_w15475_,
		_w15473_,
		_w15474_,
		_w15477_,
		_w15494_
	);
	LUT2 #(
		.INIT('h4)
	) name9668 (
		_w15493_,
		_w15494_,
		_w15495_
	);
	LUT3 #(
		.INIT('h0d)
	) name9669 (
		_w15475_,
		_w15476_,
		_w15473_,
		_w15496_
	);
	LUT4 #(
		.INIT('h000b)
	) name9670 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15497_
	);
	LUT4 #(
		.INIT('h0777)
	) name9671 (
		_w15496_,
		_w15497_,
		_w15478_,
		_w15488_,
		_w15498_
	);
	LUT2 #(
		.INIT('h4)
	) name9672 (
		_w15495_,
		_w15498_,
		_w15499_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name9673 (
		\u1_L13_reg[11]/NET0131 ,
		_w15492_,
		_w15482_,
		_w15499_,
		_w15500_
	);
	LUT4 #(
		.INIT('h2000)
	) name9674 (
		_w15475_,
		_w15474_,
		_w15477_,
		_w15480_,
		_w15501_
	);
	LUT3 #(
		.INIT('h08)
	) name9675 (
		_w15475_,
		_w15476_,
		_w15477_,
		_w15502_
	);
	LUT3 #(
		.INIT('h51)
	) name9676 (
		_w15475_,
		_w15476_,
		_w15477_,
		_w15503_
	);
	LUT4 #(
		.INIT('h4090)
	) name9677 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15504_
	);
	LUT3 #(
		.INIT('ha8)
	) name9678 (
		_w15473_,
		_w15501_,
		_w15504_,
		_w15505_
	);
	LUT3 #(
		.INIT('h80)
	) name9679 (
		_w15476_,
		_w15474_,
		_w15477_,
		_w15506_
	);
	LUT4 #(
		.INIT('hf0b0)
	) name9680 (
		_w15475_,
		_w15476_,
		_w15473_,
		_w15477_,
		_w15507_
	);
	LUT4 #(
		.INIT('h050d)
	) name9681 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15508_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9682 (
		_w15480_,
		_w15506_,
		_w15507_,
		_w15508_,
		_w15509_
	);
	LUT2 #(
		.INIT('h1)
	) name9683 (
		_w15505_,
		_w15509_,
		_w15510_
	);
	LUT3 #(
		.INIT('h10)
	) name9684 (
		_w15475_,
		_w15476_,
		_w15477_,
		_w15511_
	);
	LUT4 #(
		.INIT('h1000)
	) name9685 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15512_
	);
	LUT4 #(
		.INIT('hefbb)
	) name9686 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15513_
	);
	LUT4 #(
		.INIT('h8025)
	) name9687 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15514_
	);
	LUT4 #(
		.INIT('h5501)
	) name9688 (
		_w15473_,
		_w15480_,
		_w15513_,
		_w15514_,
		_w15515_
	);
	LUT4 #(
		.INIT('h0002)
	) name9689 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15516_
	);
	LUT4 #(
		.INIT('h3133)
	) name9690 (
		_w15475_,
		_w15473_,
		_w15474_,
		_w15477_,
		_w15517_
	);
	LUT4 #(
		.INIT('h2500)
	) name9691 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15518_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name9692 (
		_w15483_,
		_w15502_,
		_w15517_,
		_w15518_,
		_w15519_
	);
	LUT4 #(
		.INIT('h2223)
	) name9693 (
		_w15480_,
		_w15515_,
		_w15516_,
		_w15519_,
		_w15520_
	);
	LUT3 #(
		.INIT('h95)
	) name9694 (
		\u1_L13_reg[4]/NET0131 ,
		_w15510_,
		_w15520_,
		_w15521_
	);
	LUT4 #(
		.INIT('hbbec)
	) name9695 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15522_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name9696 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15523_
	);
	LUT4 #(
		.INIT('h0133)
	) name9697 (
		_w15412_,
		_w15411_,
		_w15522_,
		_w15523_,
		_w15524_
	);
	LUT4 #(
		.INIT('h0028)
	) name9698 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15525_
	);
	LUT4 #(
		.INIT('h0090)
	) name9699 (
		_w15415_,
		_w15414_,
		_w15413_,
		_w15411_,
		_w15526_
	);
	LUT3 #(
		.INIT('ha8)
	) name9700 (
		_w15412_,
		_w15525_,
		_w15526_,
		_w15527_
	);
	LUT4 #(
		.INIT('h0400)
	) name9701 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15528_
	);
	LUT4 #(
		.INIT('hfb05)
	) name9702 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15529_
	);
	LUT4 #(
		.INIT('h5001)
	) name9703 (
		_w15412_,
		_w15415_,
		_w15416_,
		_w15413_,
		_w15530_
	);
	LUT4 #(
		.INIT('h0200)
	) name9704 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15531_
	);
	LUT4 #(
		.INIT('h7d7f)
	) name9705 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15532_
	);
	LUT4 #(
		.INIT('h0d00)
	) name9706 (
		_w15412_,
		_w15529_,
		_w15530_,
		_w15532_,
		_w15533_
	);
	LUT4 #(
		.INIT('h0031)
	) name9707 (
		_w15411_,
		_w15527_,
		_w15533_,
		_w15524_,
		_w15534_
	);
	LUT2 #(
		.INIT('h9)
	) name9708 (
		\u1_L13_reg[17]/NET0131 ,
		_w15534_,
		_w15535_
	);
	LUT4 #(
		.INIT('hc693)
	) name9709 (
		decrypt_pad,
		\u1_R13_reg[15]/NET0131 ,
		\u1_uk_K_r13_reg[18]/NET0131 ,
		\u1_uk_K_r13_reg[39]/NET0131 ,
		_w15536_
	);
	LUT4 #(
		.INIT('hc693)
	) name9710 (
		decrypt_pad,
		\u1_R13_reg[14]/NET0131 ,
		\u1_uk_K_r13_reg[10]/NET0131 ,
		\u1_uk_K_r13_reg[6]/NET0131 ,
		_w15537_
	);
	LUT4 #(
		.INIT('hc963)
	) name9711 (
		decrypt_pad,
		\u1_R13_reg[12]/NET0131 ,
		\u1_uk_K_r13_reg[11]/NET0131 ,
		\u1_uk_K_r13_reg[47]/NET0131 ,
		_w15538_
	);
	LUT4 #(
		.INIT('hc693)
	) name9712 (
		decrypt_pad,
		\u1_R13_reg[13]/NET0131 ,
		\u1_uk_K_r13_reg[41]/NET0131 ,
		\u1_uk_K_r13_reg[5]/NET0131 ,
		_w15539_
	);
	LUT4 #(
		.INIT('h0012)
	) name9713 (
		_w15538_,
		_w15536_,
		_w15539_,
		_w15537_,
		_w15540_
	);
	LUT4 #(
		.INIT('hc963)
	) name9714 (
		decrypt_pad,
		\u1_R13_reg[17]/NET0131 ,
		\u1_uk_K_r13_reg[27]/NET0131 ,
		\u1_uk_K_r13_reg[6]/NET0131 ,
		_w15541_
	);
	LUT2 #(
		.INIT('h4)
	) name9715 (
		_w15538_,
		_w15541_,
		_w15542_
	);
	LUT4 #(
		.INIT('h0040)
	) name9716 (
		_w15538_,
		_w15541_,
		_w15536_,
		_w15539_,
		_w15543_
	);
	LUT2 #(
		.INIT('h8)
	) name9717 (
		_w15536_,
		_w15539_,
		_w15544_
	);
	LUT4 #(
		.INIT('h2000)
	) name9718 (
		_w15538_,
		_w15541_,
		_w15536_,
		_w15539_,
		_w15545_
	);
	LUT4 #(
		.INIT('hc693)
	) name9719 (
		decrypt_pad,
		\u1_R13_reg[16]/NET0131 ,
		\u1_uk_K_r13_reg[26]/NET0131 ,
		\u1_uk_K_r13_reg[47]/NET0131 ,
		_w15546_
	);
	LUT4 #(
		.INIT('h0004)
	) name9720 (
		_w15545_,
		_w15546_,
		_w15543_,
		_w15540_,
		_w15547_
	);
	LUT4 #(
		.INIT('h0001)
	) name9721 (
		_w15538_,
		_w15541_,
		_w15536_,
		_w15539_,
		_w15548_
	);
	LUT4 #(
		.INIT('h0040)
	) name9722 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15549_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name9723 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15550_
	);
	LUT3 #(
		.INIT('h70)
	) name9724 (
		_w15548_,
		_w15537_,
		_w15550_,
		_w15551_
	);
	LUT2 #(
		.INIT('h8)
	) name9725 (
		_w15547_,
		_w15551_,
		_w15552_
	);
	LUT4 #(
		.INIT('h0010)
	) name9726 (
		_w15538_,
		_w15541_,
		_w15536_,
		_w15539_,
		_w15553_
	);
	LUT4 #(
		.INIT('h8000)
	) name9727 (
		_w15538_,
		_w15541_,
		_w15536_,
		_w15539_,
		_w15554_
	);
	LUT3 #(
		.INIT('h01)
	) name9728 (
		_w15546_,
		_w15554_,
		_w15553_,
		_w15555_
	);
	LUT4 #(
		.INIT('h0008)
	) name9729 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15556_
	);
	LUT3 #(
		.INIT('h80)
	) name9730 (
		_w15536_,
		_w15539_,
		_w15537_,
		_w15557_
	);
	LUT4 #(
		.INIT('h4000)
	) name9731 (
		_w15538_,
		_w15536_,
		_w15539_,
		_w15537_,
		_w15558_
	);
	LUT2 #(
		.INIT('h1)
	) name9732 (
		_w15556_,
		_w15558_,
		_w15559_
	);
	LUT4 #(
		.INIT('h0001)
	) name9733 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15560_
	);
	LUT4 #(
		.INIT('heffe)
	) name9734 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15561_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name9735 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15562_
	);
	LUT3 #(
		.INIT('hc8)
	) name9736 (
		_w15536_,
		_w15561_,
		_w15562_,
		_w15563_
	);
	LUT3 #(
		.INIT('h80)
	) name9737 (
		_w15555_,
		_w15559_,
		_w15563_,
		_w15564_
	);
	LUT4 #(
		.INIT('h0200)
	) name9738 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15565_
	);
	LUT4 #(
		.INIT('heee4)
	) name9739 (
		_w15536_,
		_w15549_,
		_w15560_,
		_w15565_,
		_w15566_
	);
	LUT3 #(
		.INIT('h02)
	) name9740 (
		_w15538_,
		_w15541_,
		_w15537_,
		_w15567_
	);
	LUT2 #(
		.INIT('h8)
	) name9741 (
		_w15544_,
		_w15567_,
		_w15568_
	);
	LUT2 #(
		.INIT('h1)
	) name9742 (
		_w15566_,
		_w15568_,
		_w15569_
	);
	LUT4 #(
		.INIT('ha955)
	) name9743 (
		\u1_L13_reg[20]/NET0131 ,
		_w15552_,
		_w15564_,
		_w15569_,
		_w15570_
	);
	LUT4 #(
		.INIT('hc693)
	) name9744 (
		decrypt_pad,
		\u1_R13_reg[8]/NET0131 ,
		\u1_uk_K_r13_reg[25]/P0001 ,
		\u1_uk_K_r13_reg[46]/NET0131 ,
		_w15571_
	);
	LUT4 #(
		.INIT('hc693)
	) name9745 (
		decrypt_pad,
		\u1_R13_reg[6]/NET0131 ,
		\u1_uk_K_r13_reg[40]/NET0131 ,
		\u1_uk_K_r13_reg[4]/NET0131 ,
		_w15572_
	);
	LUT4 #(
		.INIT('hc693)
	) name9746 (
		decrypt_pad,
		\u1_R13_reg[4]/NET0131 ,
		\u1_uk_K_r13_reg[13]/NET0131 ,
		\u1_uk_K_r13_reg[34]/NET0131 ,
		_w15573_
	);
	LUT4 #(
		.INIT('hc963)
	) name9747 (
		decrypt_pad,
		\u1_R13_reg[5]/NET0131 ,
		\u1_uk_K_r13_reg[13]/NET0131 ,
		\u1_uk_K_r13_reg[17]/NET0131 ,
		_w15574_
	);
	LUT4 #(
		.INIT('hc963)
	) name9748 (
		decrypt_pad,
		\u1_R13_reg[9]/NET0131 ,
		\u1_uk_K_r13_reg[26]/NET0131 ,
		\u1_uk_K_r13_reg[5]/NET0131 ,
		_w15575_
	);
	LUT2 #(
		.INIT('h2)
	) name9749 (
		_w15574_,
		_w15575_,
		_w15576_
	);
	LUT4 #(
		.INIT('h0212)
	) name9750 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15577_
	);
	LUT4 #(
		.INIT('hc693)
	) name9751 (
		decrypt_pad,
		\u1_R13_reg[7]/NET0131 ,
		\u1_uk_K_r13_reg[34]/NET0131 ,
		\u1_uk_K_r13_reg[55]/NET0131 ,
		_w15578_
	);
	LUT2 #(
		.INIT('h1)
	) name9752 (
		_w15574_,
		_w15578_,
		_w15579_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name9753 (
		_w15574_,
		_w15572_,
		_w15573_,
		_w15578_,
		_w15580_
	);
	LUT3 #(
		.INIT('hb0)
	) name9754 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15581_
	);
	LUT4 #(
		.INIT('h73af)
	) name9755 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15582_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name9756 (
		_w15578_,
		_w15580_,
		_w15581_,
		_w15582_,
		_w15583_
	);
	LUT3 #(
		.INIT('h45)
	) name9757 (
		_w15571_,
		_w15577_,
		_w15583_,
		_w15584_
	);
	LUT4 #(
		.INIT('h4000)
	) name9758 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15585_
	);
	LUT4 #(
		.INIT('hbff2)
	) name9759 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15586_
	);
	LUT2 #(
		.INIT('h1)
	) name9760 (
		_w15578_,
		_w15586_,
		_w15587_
	);
	LUT4 #(
		.INIT('h0100)
	) name9761 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15588_
	);
	LUT4 #(
		.INIT('h2000)
	) name9762 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15589_
	);
	LUT4 #(
		.INIT('ha200)
	) name9763 (
		_w15574_,
		_w15572_,
		_w15573_,
		_w15578_,
		_w15590_
	);
	LUT3 #(
		.INIT('h01)
	) name9764 (
		_w15589_,
		_w15590_,
		_w15588_,
		_w15591_
	);
	LUT3 #(
		.INIT('h8a)
	) name9765 (
		_w15571_,
		_w15587_,
		_w15591_,
		_w15592_
	);
	LUT2 #(
		.INIT('h9)
	) name9766 (
		_w15574_,
		_w15572_,
		_w15593_
	);
	LUT3 #(
		.INIT('h02)
	) name9767 (
		_w15575_,
		_w15573_,
		_w15578_,
		_w15594_
	);
	LUT2 #(
		.INIT('h8)
	) name9768 (
		_w15593_,
		_w15594_,
		_w15595_
	);
	LUT3 #(
		.INIT('h04)
	) name9769 (
		_w15574_,
		_w15572_,
		_w15573_,
		_w15596_
	);
	LUT4 #(
		.INIT('h0004)
	) name9770 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15597_
	);
	LUT4 #(
		.INIT('hddfb)
	) name9771 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15598_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9772 (
		_w15578_,
		_w15571_,
		_w15585_,
		_w15598_,
		_w15599_
	);
	LUT2 #(
		.INIT('h1)
	) name9773 (
		_w15595_,
		_w15599_,
		_w15600_
	);
	LUT4 #(
		.INIT('h5655)
	) name9774 (
		\u1_L13_reg[2]/NET0131 ,
		_w15592_,
		_w15584_,
		_w15600_,
		_w15601_
	);
	LUT4 #(
		.INIT('h0484)
	) name9775 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15602_
	);
	LUT4 #(
		.INIT('h0043)
	) name9776 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15603_
	);
	LUT4 #(
		.INIT('h70d0)
	) name9777 (
		_w15475_,
		_w15476_,
		_w15473_,
		_w15477_,
		_w15604_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name9778 (
		_w15517_,
		_w15602_,
		_w15603_,
		_w15604_,
		_w15605_
	);
	LUT2 #(
		.INIT('h1)
	) name9779 (
		_w15480_,
		_w15512_,
		_w15606_
	);
	LUT4 #(
		.INIT('hbb7b)
	) name9780 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15607_
	);
	LUT2 #(
		.INIT('h2)
	) name9781 (
		_w15473_,
		_w15607_,
		_w15608_
	);
	LUT3 #(
		.INIT('h48)
	) name9782 (
		_w15475_,
		_w15474_,
		_w15477_,
		_w15609_
	);
	LUT4 #(
		.INIT('h0e04)
	) name9783 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15610_
	);
	LUT4 #(
		.INIT('h888c)
	) name9784 (
		_w15476_,
		_w15473_,
		_w15474_,
		_w15477_,
		_w15611_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9785 (
		_w15480_,
		_w15610_,
		_w15611_,
		_w15609_,
		_w15612_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9786 (
		_w15605_,
		_w15606_,
		_w15608_,
		_w15612_,
		_w15613_
	);
	LUT4 #(
		.INIT('h0800)
	) name9787 (
		_w15476_,
		_w15473_,
		_w15474_,
		_w15477_,
		_w15614_
	);
	LUT2 #(
		.INIT('h1)
	) name9788 (
		_w15516_,
		_w15614_,
		_w15615_
	);
	LUT3 #(
		.INIT('h9a)
	) name9789 (
		\u1_L13_reg[29]/NET0131 ,
		_w15613_,
		_w15615_,
		_w15616_
	);
	LUT4 #(
		.INIT('hc963)
	) name9790 (
		decrypt_pad,
		\u1_R13_reg[32]/NET0131 ,
		\u1_uk_K_r13_reg[14]/NET0131 ,
		\u1_uk_K_r13_reg[52]/P0001 ,
		_w15617_
	);
	LUT4 #(
		.INIT('hc693)
	) name9791 (
		decrypt_pad,
		\u1_R13_reg[31]/P0001 ,
		\u1_uk_K_r13_reg[42]/NET0131 ,
		\u1_uk_K_r13_reg[8]/NET0131 ,
		_w15618_
	);
	LUT4 #(
		.INIT('hc693)
	) name9792 (
		decrypt_pad,
		\u1_R13_reg[30]/NET0131 ,
		\u1_uk_K_r13_reg[30]/NET0131 ,
		\u1_uk_K_r13_reg[51]/NET0131 ,
		_w15619_
	);
	LUT4 #(
		.INIT('hc693)
	) name9793 (
		decrypt_pad,
		\u1_R13_reg[29]/NET0131 ,
		\u1_uk_K_r13_reg[29]/NET0131 ,
		\u1_uk_K_r13_reg[50]/NET0131 ,
		_w15620_
	);
	LUT4 #(
		.INIT('hc963)
	) name9794 (
		decrypt_pad,
		\u1_R13_reg[28]/NET0131 ,
		\u1_uk_K_r13_reg[23]/NET0131 ,
		\u1_uk_K_r13_reg[2]/NET0131 ,
		_w15621_
	);
	LUT4 #(
		.INIT('hc693)
	) name9795 (
		decrypt_pad,
		\u1_R13_reg[1]/NET0131 ,
		\u1_uk_K_r13_reg[14]/NET0131 ,
		\u1_uk_K_r13_reg[35]/NET0131 ,
		_w15622_
	);
	LUT2 #(
		.INIT('h8)
	) name9796 (
		_w15622_,
		_w15621_,
		_w15623_
	);
	LUT4 #(
		.INIT('ha6f3)
	) name9797 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15624_
	);
	LUT3 #(
		.INIT('h08)
	) name9798 (
		_w15619_,
		_w15620_,
		_w15621_,
		_w15625_
	);
	LUT4 #(
		.INIT('h0080)
	) name9799 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15626_
	);
	LUT3 #(
		.INIT('h01)
	) name9800 (
		_w15619_,
		_w15620_,
		_w15621_,
		_w15627_
	);
	LUT4 #(
		.INIT('h2031)
	) name9801 (
		_w15618_,
		_w15626_,
		_w15624_,
		_w15627_,
		_w15628_
	);
	LUT2 #(
		.INIT('h2)
	) name9802 (
		_w15617_,
		_w15628_,
		_w15629_
	);
	LUT4 #(
		.INIT('h0200)
	) name9803 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15630_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name9804 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15631_
	);
	LUT2 #(
		.INIT('h2)
	) name9805 (
		_w15618_,
		_w15631_,
		_w15632_
	);
	LUT2 #(
		.INIT('h1)
	) name9806 (
		_w15618_,
		_w15619_,
		_w15633_
	);
	LUT4 #(
		.INIT('heece)
	) name9807 (
		_w15618_,
		_w15619_,
		_w15620_,
		_w15622_,
		_w15634_
	);
	LUT2 #(
		.INIT('h4)
	) name9808 (
		_w15634_,
		_w15621_,
		_w15635_
	);
	LUT4 #(
		.INIT('h8000)
	) name9809 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15636_
	);
	LUT3 #(
		.INIT('h45)
	) name9810 (
		_w15618_,
		_w15622_,
		_w15621_,
		_w15637_
	);
	LUT3 #(
		.INIT('hca)
	) name9811 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15638_
	);
	LUT3 #(
		.INIT('h15)
	) name9812 (
		_w15636_,
		_w15637_,
		_w15638_,
		_w15639_
	);
	LUT4 #(
		.INIT('h00ef)
	) name9813 (
		_w15635_,
		_w15632_,
		_w15639_,
		_w15617_,
		_w15640_
	);
	LUT4 #(
		.INIT('h0008)
	) name9814 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15641_
	);
	LUT4 #(
		.INIT('heff7)
	) name9815 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15642_
	);
	LUT4 #(
		.INIT('h0020)
	) name9816 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15643_
	);
	LUT4 #(
		.INIT('h0001)
	) name9817 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15644_
	);
	LUT4 #(
		.INIT('hefd6)
	) name9818 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15645_
	);
	LUT2 #(
		.INIT('h2)
	) name9819 (
		_w15618_,
		_w15645_,
		_w15646_
	);
	LUT3 #(
		.INIT('h40)
	) name9820 (
		_w15620_,
		_w15621_,
		_w15617_,
		_w15647_
	);
	LUT3 #(
		.INIT('h20)
	) name9821 (
		_w15620_,
		_w15622_,
		_w15621_,
		_w15648_
	);
	LUT4 #(
		.INIT('haebf)
	) name9822 (
		_w15618_,
		_w15619_,
		_w15647_,
		_w15648_,
		_w15649_
	);
	LUT2 #(
		.INIT('h4)
	) name9823 (
		_w15646_,
		_w15649_,
		_w15650_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name9824 (
		\u1_L13_reg[5]/NET0131 ,
		_w15640_,
		_w15629_,
		_w15650_,
		_w15651_
	);
	LUT4 #(
		.INIT('h0800)
	) name9825 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15652_
	);
	LUT4 #(
		.INIT('hd7ff)
	) name9826 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15653_
	);
	LUT4 #(
		.INIT('hfeb5)
	) name9827 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15654_
	);
	LUT4 #(
		.INIT('h0515)
	) name9828 (
		_w15578_,
		_w15571_,
		_w15653_,
		_w15654_,
		_w15655_
	);
	LUT4 #(
		.INIT('h5404)
	) name9829 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15656_
	);
	LUT3 #(
		.INIT('h08)
	) name9830 (
		_w15572_,
		_w15575_,
		_w15573_,
		_w15657_
	);
	LUT3 #(
		.INIT('h01)
	) name9831 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15658_
	);
	LUT4 #(
		.INIT('heee4)
	) name9832 (
		_w15578_,
		_w15656_,
		_w15658_,
		_w15657_,
		_w15659_
	);
	LUT4 #(
		.INIT('h0002)
	) name9833 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15660_
	);
	LUT4 #(
		.INIT('h008a)
	) name9834 (
		_w15571_,
		_w15580_,
		_w15581_,
		_w15660_,
		_w15661_
	);
	LUT3 #(
		.INIT('h20)
	) name9835 (
		_w15653_,
		_w15659_,
		_w15661_,
		_w15662_
	);
	LUT3 #(
		.INIT('h8e)
	) name9836 (
		_w15574_,
		_w15575_,
		_w15573_,
		_w15663_
	);
	LUT4 #(
		.INIT('h0d00)
	) name9837 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15664_
	);
	LUT3 #(
		.INIT('h02)
	) name9838 (
		_w15578_,
		_w15664_,
		_w15663_,
		_w15665_
	);
	LUT3 #(
		.INIT('h80)
	) name9839 (
		_w15572_,
		_w15573_,
		_w15578_,
		_w15666_
	);
	LUT2 #(
		.INIT('h4)
	) name9840 (
		_w15576_,
		_w15666_,
		_w15667_
	);
	LUT3 #(
		.INIT('h04)
	) name9841 (
		_w15572_,
		_w15575_,
		_w15573_,
		_w15668_
	);
	LUT3 #(
		.INIT('h45)
	) name9842 (
		_w15571_,
		_w15579_,
		_w15668_,
		_w15669_
	);
	LUT3 #(
		.INIT('h10)
	) name9843 (
		_w15665_,
		_w15667_,
		_w15669_,
		_w15670_
	);
	LUT4 #(
		.INIT('h999a)
	) name9844 (
		\u1_L13_reg[13]/NET0131 ,
		_w15655_,
		_w15662_,
		_w15670_,
		_w15671_
	);
	LUT4 #(
		.INIT('hc963)
	) name9845 (
		decrypt_pad,
		\u1_R13_reg[19]/NET0131 ,
		\u1_uk_K_r13_reg[15]/NET0131 ,
		\u1_uk_K_r13_reg[49]/NET0131 ,
		_w15672_
	);
	LUT4 #(
		.INIT('hc693)
	) name9846 (
		decrypt_pad,
		\u1_R13_reg[16]/NET0131 ,
		\u1_uk_K_r13_reg[22]/NET0131 ,
		\u1_uk_K_r13_reg[43]/NET0131 ,
		_w15673_
	);
	LUT4 #(
		.INIT('hc963)
	) name9847 (
		decrypt_pad,
		\u1_R13_reg[21]/NET0131 ,
		\u1_uk_K_r13_reg[0]/NET0131 ,
		\u1_uk_K_r13_reg[38]/NET0131 ,
		_w15674_
	);
	LUT4 #(
		.INIT('hc963)
	) name9848 (
		decrypt_pad,
		\u1_R13_reg[17]/NET0131 ,
		\u1_uk_K_r13_reg[38]/NET0131 ,
		\u1_uk_K_r13_reg[44]/NET0131 ,
		_w15675_
	);
	LUT4 #(
		.INIT('hc963)
	) name9849 (
		decrypt_pad,
		\u1_R13_reg[18]/NET0131 ,
		\u1_uk_K_r13_reg[28]/NET0131 ,
		\u1_uk_K_r13_reg[7]/NET0131 ,
		_w15676_
	);
	LUT4 #(
		.INIT('h0080)
	) name9850 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15677_
	);
	LUT4 #(
		.INIT('h0002)
	) name9851 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15678_
	);
	LUT4 #(
		.INIT('hcb79)
	) name9852 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15679_
	);
	LUT4 #(
		.INIT('h76ae)
	) name9853 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15680_
	);
	LUT4 #(
		.INIT('h0800)
	) name9854 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15681_
	);
	LUT4 #(
		.INIT('hf7ef)
	) name9855 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15682_
	);
	LUT4 #(
		.INIT('he400)
	) name9856 (
		_w15672_,
		_w15679_,
		_w15680_,
		_w15682_,
		_w15683_
	);
	LUT4 #(
		.INIT('hc963)
	) name9857 (
		decrypt_pad,
		\u1_R13_reg[20]/NET0131 ,
		\u1_uk_K_r13_reg[30]/NET0131 ,
		\u1_uk_K_r13_reg[9]/NET0131 ,
		_w15684_
	);
	LUT2 #(
		.INIT('h1)
	) name9858 (
		_w15683_,
		_w15684_,
		_w15685_
	);
	LUT4 #(
		.INIT('h9b53)
	) name9859 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15686_
	);
	LUT2 #(
		.INIT('h2)
	) name9860 (
		_w15672_,
		_w15686_,
		_w15687_
	);
	LUT2 #(
		.INIT('h1)
	) name9861 (
		_w15672_,
		_w15676_,
		_w15688_
	);
	LUT3 #(
		.INIT('hbe)
	) name9862 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15689_
	);
	LUT2 #(
		.INIT('h2)
	) name9863 (
		_w15688_,
		_w15689_,
		_w15690_
	);
	LUT2 #(
		.INIT('h9)
	) name9864 (
		_w15675_,
		_w15676_,
		_w15691_
	);
	LUT4 #(
		.INIT('h0220)
	) name9865 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15692_
	);
	LUT4 #(
		.INIT('h40c0)
	) name9866 (
		_w15672_,
		_w15673_,
		_w15674_,
		_w15675_,
		_w15693_
	);
	LUT3 #(
		.INIT('h13)
	) name9867 (
		_w15691_,
		_w15692_,
		_w15693_,
		_w15694_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9868 (
		_w15684_,
		_w15687_,
		_w15690_,
		_w15694_,
		_w15695_
	);
	LUT4 #(
		.INIT('h0020)
	) name9869 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15696_
	);
	LUT4 #(
		.INIT('hfedf)
	) name9870 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15697_
	);
	LUT4 #(
		.INIT('h0400)
	) name9871 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15698_
	);
	LUT4 #(
		.INIT('hebff)
	) name9872 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15699_
	);
	LUT3 #(
		.INIT('hd8)
	) name9873 (
		_w15672_,
		_w15697_,
		_w15699_,
		_w15700_
	);
	LUT4 #(
		.INIT('h5655)
	) name9874 (
		\u1_L13_reg[14]/NET0131 ,
		_w15685_,
		_w15695_,
		_w15700_,
		_w15701_
	);
	LUT4 #(
		.INIT('h672f)
	) name9875 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15702_
	);
	LUT4 #(
		.INIT('h2000)
	) name9876 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15703_
	);
	LUT4 #(
		.INIT('hdaff)
	) name9877 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15704_
	);
	LUT4 #(
		.INIT('h0010)
	) name9878 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15705_
	);
	LUT4 #(
		.INIT('hf7ed)
	) name9879 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15706_
	);
	LUT4 #(
		.INIT('he400)
	) name9880 (
		_w15618_,
		_w15704_,
		_w15702_,
		_w15706_,
		_w15707_
	);
	LUT2 #(
		.INIT('h2)
	) name9881 (
		_w15617_,
		_w15707_,
		_w15708_
	);
	LUT4 #(
		.INIT('h0004)
	) name9882 (
		_w15618_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15709_
	);
	LUT3 #(
		.INIT('hce)
	) name9883 (
		_w15618_,
		_w15619_,
		_w15620_,
		_w15710_
	);
	LUT4 #(
		.INIT('h0031)
	) name9884 (
		_w15623_,
		_w15644_,
		_w15710_,
		_w15709_,
		_w15711_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name9885 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15712_
	);
	LUT2 #(
		.INIT('h2)
	) name9886 (
		_w15618_,
		_w15712_,
		_w15713_
	);
	LUT4 #(
		.INIT('h0040)
	) name9887 (
		_w15618_,
		_w15619_,
		_w15622_,
		_w15621_,
		_w15714_
	);
	LUT3 #(
		.INIT('h01)
	) name9888 (
		_w15630_,
		_w15625_,
		_w15714_,
		_w15715_
	);
	LUT4 #(
		.INIT('h4555)
	) name9889 (
		_w15617_,
		_w15713_,
		_w15715_,
		_w15711_,
		_w15716_
	);
	LUT4 #(
		.INIT('h0002)
	) name9890 (
		_w15618_,
		_w15619_,
		_w15620_,
		_w15621_,
		_w15717_
	);
	LUT3 #(
		.INIT('h80)
	) name9891 (
		_w15620_,
		_w15622_,
		_w15621_,
		_w15718_
	);
	LUT3 #(
		.INIT('h13)
	) name9892 (
		_w15633_,
		_w15717_,
		_w15718_,
		_w15719_
	);
	LUT4 #(
		.INIT('h5655)
	) name9893 (
		\u1_L13_reg[21]/NET0131 ,
		_w15716_,
		_w15708_,
		_w15719_,
		_w15720_
	);
	LUT4 #(
		.INIT('hf309)
	) name9894 (
		_w15541_,
		_w15536_,
		_w15539_,
		_w15537_,
		_w15721_
	);
	LUT2 #(
		.INIT('h2)
	) name9895 (
		_w15538_,
		_w15721_,
		_w15722_
	);
	LUT4 #(
		.INIT('h0040)
	) name9896 (
		_w15538_,
		_w15541_,
		_w15536_,
		_w15537_,
		_w15723_
	);
	LUT3 #(
		.INIT('h04)
	) name9897 (
		_w15548_,
		_w15561_,
		_w15723_,
		_w15724_
	);
	LUT3 #(
		.INIT('h45)
	) name9898 (
		_w15546_,
		_w15722_,
		_w15724_,
		_w15725_
	);
	LUT4 #(
		.INIT('h7bff)
	) name9899 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15726_
	);
	LUT4 #(
		.INIT('h2202)
	) name9900 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15727_
	);
	LUT3 #(
		.INIT('h01)
	) name9901 (
		_w15536_,
		_w15549_,
		_w15727_,
		_w15728_
	);
	LUT4 #(
		.INIT('he0f0)
	) name9902 (
		_w15538_,
		_w15541_,
		_w15536_,
		_w15539_,
		_w15729_
	);
	LUT2 #(
		.INIT('h4)
	) name9903 (
		_w15556_,
		_w15729_,
		_w15730_
	);
	LUT4 #(
		.INIT('h222a)
	) name9904 (
		_w15546_,
		_w15726_,
		_w15728_,
		_w15730_,
		_w15731_
	);
	LUT4 #(
		.INIT('h7bfe)
	) name9905 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15732_
	);
	LUT2 #(
		.INIT('h1)
	) name9906 (
		_w15536_,
		_w15732_,
		_w15733_
	);
	LUT3 #(
		.INIT('h13)
	) name9907 (
		_w15544_,
		_w15558_,
		_w15567_,
		_w15734_
	);
	LUT2 #(
		.INIT('h4)
	) name9908 (
		_w15733_,
		_w15734_,
		_w15735_
	);
	LUT4 #(
		.INIT('h5655)
	) name9909 (
		\u1_L13_reg[10]/NET0131 ,
		_w15731_,
		_w15725_,
		_w15735_,
		_w15736_
	);
	LUT4 #(
		.INIT('h0100)
	) name9910 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15737_
	);
	LUT3 #(
		.INIT('h08)
	) name9911 (
		_w15447_,
		_w15449_,
		_w15446_,
		_w15738_
	);
	LUT4 #(
		.INIT('h0004)
	) name9912 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15739_
	);
	LUT4 #(
		.INIT('h0001)
	) name9913 (
		_w15445_,
		_w15737_,
		_w15738_,
		_w15739_,
		_w15740_
	);
	LUT2 #(
		.INIT('h1)
	) name9914 (
		_w15450_,
		_w15446_,
		_w15741_
	);
	LUT4 #(
		.INIT('h00a2)
	) name9915 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15742_
	);
	LUT4 #(
		.INIT('h2010)
	) name9916 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15743_
	);
	LUT3 #(
		.INIT('h09)
	) name9917 (
		_w15448_,
		_w15450_,
		_w15446_,
		_w15744_
	);
	LUT4 #(
		.INIT('h1011)
	) name9918 (
		_w15743_,
		_w15744_,
		_w15741_,
		_w15742_,
		_w15745_
	);
	LUT3 #(
		.INIT('h08)
	) name9919 (
		_w15450_,
		_w15447_,
		_w15449_,
		_w15746_
	);
	LUT4 #(
		.INIT('h0040)
	) name9920 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15747_
	);
	LUT4 #(
		.INIT('h0008)
	) name9921 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15748_
	);
	LUT4 #(
		.INIT('h0002)
	) name9922 (
		_w15445_,
		_w15465_,
		_w15748_,
		_w15747_,
		_w15749_
	);
	LUT3 #(
		.INIT('hb9)
	) name9923 (
		_w15448_,
		_w15449_,
		_w15446_,
		_w15750_
	);
	LUT4 #(
		.INIT('h33fe)
	) name9924 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15751_
	);
	LUT4 #(
		.INIT('hf351)
	) name9925 (
		_w15446_,
		_w15459_,
		_w15750_,
		_w15751_,
		_w15752_
	);
	LUT4 #(
		.INIT('h0777)
	) name9926 (
		_w15740_,
		_w15745_,
		_w15749_,
		_w15752_,
		_w15753_
	);
	LUT2 #(
		.INIT('h6)
	) name9927 (
		\u1_L13_reg[12]/NET0131 ,
		_w15753_,
		_w15754_
	);
	LUT4 #(
		.INIT('h33cb)
	) name9928 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15755_
	);
	LUT4 #(
		.INIT('h0100)
	) name9929 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15756_
	);
	LUT4 #(
		.INIT('h3302)
	) name9930 (
		_w15618_,
		_w15617_,
		_w15755_,
		_w15756_,
		_w15757_
	);
	LUT3 #(
		.INIT('h40)
	) name9931 (
		_w15619_,
		_w15620_,
		_w15621_,
		_w15758_
	);
	LUT4 #(
		.INIT('h0400)
	) name9932 (
		_w15618_,
		_w15619_,
		_w15620_,
		_w15622_,
		_w15759_
	);
	LUT3 #(
		.INIT('h01)
	) name9933 (
		_w15641_,
		_w15758_,
		_w15759_,
		_w15760_
	);
	LUT4 #(
		.INIT('h0002)
	) name9934 (
		_w15618_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15761_
	);
	LUT2 #(
		.INIT('h1)
	) name9935 (
		_w15703_,
		_w15761_,
		_w15762_
	);
	LUT3 #(
		.INIT('h2a)
	) name9936 (
		_w15617_,
		_w15760_,
		_w15762_,
		_w15763_
	);
	LUT4 #(
		.INIT('h5155)
	) name9937 (
		_w15618_,
		_w15619_,
		_w15620_,
		_w15621_,
		_w15764_
	);
	LUT4 #(
		.INIT('h0040)
	) name9938 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15765_
	);
	LUT3 #(
		.INIT('h04)
	) name9939 (
		_w15620_,
		_w15621_,
		_w15617_,
		_w15766_
	);
	LUT4 #(
		.INIT('hfff6)
	) name9940 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15767_
	);
	LUT4 #(
		.INIT('h1000)
	) name9941 (
		_w15765_,
		_w15766_,
		_w15764_,
		_w15767_,
		_w15768_
	);
	LUT3 #(
		.INIT('h02)
	) name9942 (
		_w15618_,
		_w15626_,
		_w15705_,
		_w15769_
	);
	LUT2 #(
		.INIT('h1)
	) name9943 (
		_w15768_,
		_w15769_,
		_w15770_
	);
	LUT4 #(
		.INIT('h5556)
	) name9944 (
		\u1_L13_reg[15]/P0001 ,
		_w15757_,
		_w15763_,
		_w15770_,
		_w15771_
	);
	LUT4 #(
		.INIT('hf070)
	) name9945 (
		_w15475_,
		_w15476_,
		_w15473_,
		_w15474_,
		_w15772_
	);
	LUT3 #(
		.INIT('h45)
	) name9946 (
		_w15496_,
		_w15511_,
		_w15772_,
		_w15773_
	);
	LUT4 #(
		.INIT('h010c)
	) name9947 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15774_
	);
	LUT4 #(
		.INIT('h4010)
	) name9948 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15775_
	);
	LUT3 #(
		.INIT('h02)
	) name9949 (
		_w15480_,
		_w15775_,
		_w15774_,
		_w15776_
	);
	LUT4 #(
		.INIT('h0401)
	) name9950 (
		_w15475_,
		_w15476_,
		_w15473_,
		_w15477_,
		_w15777_
	);
	LUT4 #(
		.INIT('h8000)
	) name9951 (
		_w15475_,
		_w15476_,
		_w15474_,
		_w15477_,
		_w15778_
	);
	LUT4 #(
		.INIT('h0045)
	) name9952 (
		_w15480_,
		_w15503_,
		_w15772_,
		_w15778_,
		_w15779_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9953 (
		_w15773_,
		_w15776_,
		_w15777_,
		_w15779_,
		_w15780_
	);
	LUT4 #(
		.INIT('h99bf)
	) name9954 (
		_w15476_,
		_w15477_,
		_w15488_,
		_w15484_,
		_w15781_
	);
	LUT3 #(
		.INIT('h65)
	) name9955 (
		\u1_L13_reg[19]/P0001 ,
		_w15780_,
		_w15781_,
		_w15782_
	);
	LUT3 #(
		.INIT('h02)
	) name9956 (
		_w15538_,
		_w15539_,
		_w15537_,
		_w15783_
	);
	LUT4 #(
		.INIT('hf3f1)
	) name9957 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15784_
	);
	LUT4 #(
		.INIT('h6bff)
	) name9958 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15785_
	);
	LUT4 #(
		.INIT('h08aa)
	) name9959 (
		_w15536_,
		_w15546_,
		_w15784_,
		_w15785_,
		_w15786_
	);
	LUT3 #(
		.INIT('h01)
	) name9960 (
		_w15538_,
		_w15541_,
		_w15537_,
		_w15787_
	);
	LUT3 #(
		.INIT('h02)
	) name9961 (
		_w15536_,
		_w15565_,
		_w15787_,
		_w15788_
	);
	LUT4 #(
		.INIT('h0f07)
	) name9962 (
		_w15538_,
		_w15541_,
		_w15536_,
		_w15539_,
		_w15789_
	);
	LUT2 #(
		.INIT('h4)
	) name9963 (
		_w15567_,
		_w15789_,
		_w15790_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name9964 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15791_
	);
	LUT4 #(
		.INIT('h0155)
	) name9965 (
		_w15546_,
		_w15788_,
		_w15790_,
		_w15791_,
		_w15792_
	);
	LUT4 #(
		.INIT('hbf2f)
	) name9966 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15793_
	);
	LUT4 #(
		.INIT('h2500)
	) name9967 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15794_
	);
	LUT4 #(
		.INIT('hcc04)
	) name9968 (
		_w15536_,
		_w15546_,
		_w15793_,
		_w15794_,
		_w15795_
	);
	LUT2 #(
		.INIT('h1)
	) name9969 (
		_w15541_,
		_w15536_,
		_w15796_
	);
	LUT2 #(
		.INIT('h8)
	) name9970 (
		_w15794_,
		_w15796_,
		_w15797_
	);
	LUT2 #(
		.INIT('h1)
	) name9971 (
		_w15795_,
		_w15797_,
		_w15798_
	);
	LUT4 #(
		.INIT('h5655)
	) name9972 (
		\u1_L13_reg[1]/NET0131 ,
		_w15792_,
		_w15786_,
		_w15798_,
		_w15799_
	);
	LUT4 #(
		.INIT('h15ff)
	) name9973 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15800_
	);
	LUT2 #(
		.INIT('h1)
	) name9974 (
		_w15412_,
		_w15800_,
		_w15801_
	);
	LUT4 #(
		.INIT('h0008)
	) name9975 (
		_w15412_,
		_w15415_,
		_w15414_,
		_w15413_,
		_w15802_
	);
	LUT4 #(
		.INIT('h0001)
	) name9976 (
		_w15432_,
		_w15421_,
		_w15438_,
		_w15802_,
		_w15803_
	);
	LUT3 #(
		.INIT('h45)
	) name9977 (
		_w15411_,
		_w15801_,
		_w15803_,
		_w15804_
	);
	LUT4 #(
		.INIT('h007f)
	) name9978 (
		_w15415_,
		_w15414_,
		_w15413_,
		_w15411_,
		_w15805_
	);
	LUT4 #(
		.INIT('h9000)
	) name9979 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15806_
	);
	LUT4 #(
		.INIT('h0600)
	) name9980 (
		_w15415_,
		_w15414_,
		_w15413_,
		_w15411_,
		_w15807_
	);
	LUT4 #(
		.INIT('hfdfb)
	) name9981 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15808_
	);
	LUT4 #(
		.INIT('h4500)
	) name9982 (
		_w15807_,
		_w15805_,
		_w15806_,
		_w15808_,
		_w15809_
	);
	LUT2 #(
		.INIT('h1)
	) name9983 (
		_w15412_,
		_w15809_,
		_w15810_
	);
	LUT3 #(
		.INIT('had)
	) name9984 (
		_w15415_,
		_w15414_,
		_w15413_,
		_w15811_
	);
	LUT2 #(
		.INIT('h2)
	) name9985 (
		_w15434_,
		_w15811_,
		_w15812_
	);
	LUT3 #(
		.INIT('h28)
	) name9986 (
		_w15415_,
		_w15414_,
		_w15413_,
		_w15813_
	);
	LUT3 #(
		.INIT('ha8)
	) name9987 (
		_w15412_,
		_w15414_,
		_w15416_,
		_w15814_
	);
	LUT2 #(
		.INIT('h8)
	) name9988 (
		_w15813_,
		_w15814_,
		_w15815_
	);
	LUT3 #(
		.INIT('h07)
	) name9989 (
		_w15429_,
		_w15440_,
		_w15528_,
		_w15816_
	);
	LUT4 #(
		.INIT('h1311)
	) name9990 (
		_w15411_,
		_w15812_,
		_w15815_,
		_w15816_,
		_w15817_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name9991 (
		\u1_L13_reg[23]/P0001 ,
		_w15810_,
		_w15804_,
		_w15817_,
		_w15818_
	);
	LUT3 #(
		.INIT('h80)
	) name9992 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15819_
	);
	LUT4 #(
		.INIT('h6a78)
	) name9993 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15820_
	);
	LUT4 #(
		.INIT('hf7a7)
	) name9994 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15821_
	);
	LUT4 #(
		.INIT('hdf3f)
	) name9995 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15822_
	);
	LUT4 #(
		.INIT('hd800)
	) name9996 (
		_w15672_,
		_w15820_,
		_w15821_,
		_w15822_,
		_w15823_
	);
	LUT2 #(
		.INIT('h2)
	) name9997 (
		_w15684_,
		_w15823_,
		_w15824_
	);
	LUT3 #(
		.INIT('h8a)
	) name9998 (
		_w15672_,
		_w15674_,
		_w15675_,
		_w15825_
	);
	LUT4 #(
		.INIT('h00ab)
	) name9999 (
		_w15672_,
		_w15673_,
		_w15675_,
		_w15676_,
		_w15826_
	);
	LUT2 #(
		.INIT('h4)
	) name10000 (
		_w15825_,
		_w15826_,
		_w15827_
	);
	LUT4 #(
		.INIT('h0004)
	) name10001 (
		_w15672_,
		_w15673_,
		_w15674_,
		_w15675_,
		_w15828_
	);
	LUT2 #(
		.INIT('h2)
	) name10002 (
		_w15672_,
		_w15674_,
		_w15829_
	);
	LUT3 #(
		.INIT('h40)
	) name10003 (
		_w15673_,
		_w15675_,
		_w15676_,
		_w15830_
	);
	LUT3 #(
		.INIT('h45)
	) name10004 (
		_w15828_,
		_w15829_,
		_w15830_,
		_w15831_
	);
	LUT4 #(
		.INIT('hdefb)
	) name10005 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15832_
	);
	LUT4 #(
		.INIT('h0400)
	) name10006 (
		_w15672_,
		_w15673_,
		_w15675_,
		_w15676_,
		_w15833_
	);
	LUT4 #(
		.INIT('h0031)
	) name10007 (
		_w15672_,
		_w15677_,
		_w15832_,
		_w15833_,
		_w15834_
	);
	LUT4 #(
		.INIT('hba00)
	) name10008 (
		_w15684_,
		_w15827_,
		_w15831_,
		_w15834_,
		_w15835_
	);
	LUT3 #(
		.INIT('h65)
	) name10009 (
		\u1_L13_reg[25]/NET0131 ,
		_w15824_,
		_w15835_,
		_w15836_
	);
	LUT4 #(
		.INIT('h77fb)
	) name10010 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15837_
	);
	LUT3 #(
		.INIT('h32)
	) name10011 (
		_w15536_,
		_w15553_,
		_w15837_,
		_w15838_
	);
	LUT4 #(
		.INIT('h2010)
	) name10012 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15839_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name10013 (
		_w15538_,
		_w15541_,
		_w15536_,
		_w15539_,
		_w15840_
	);
	LUT3 #(
		.INIT('h31)
	) name10014 (
		_w15537_,
		_w15839_,
		_w15840_,
		_w15841_
	);
	LUT3 #(
		.INIT('h2a)
	) name10015 (
		_w15546_,
		_w15838_,
		_w15841_,
		_w15842_
	);
	LUT4 #(
		.INIT('hf8fc)
	) name10016 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15843_
	);
	LUT4 #(
		.INIT('h0092)
	) name10017 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15844_
	);
	LUT4 #(
		.INIT('h5501)
	) name10018 (
		_w15536_,
		_w15546_,
		_w15843_,
		_w15844_,
		_w15845_
	);
	LUT4 #(
		.INIT('hffb7)
	) name10019 (
		_w15538_,
		_w15541_,
		_w15539_,
		_w15537_,
		_w15846_
	);
	LUT2 #(
		.INIT('h2)
	) name10020 (
		_w15536_,
		_w15846_,
		_w15847_
	);
	LUT2 #(
		.INIT('h4)
	) name10021 (
		_w15542_,
		_w15557_,
		_w15848_
	);
	LUT3 #(
		.INIT('h01)
	) name10022 (
		_w15545_,
		_w15549_,
		_w15783_,
		_w15849_
	);
	LUT4 #(
		.INIT('h2322)
	) name10023 (
		_w15546_,
		_w15847_,
		_w15848_,
		_w15849_,
		_w15850_
	);
	LUT4 #(
		.INIT('h5655)
	) name10024 (
		\u1_L13_reg[26]/NET0131 ,
		_w15845_,
		_w15842_,
		_w15850_,
		_w15851_
	);
	LUT4 #(
		.INIT('h0008)
	) name10025 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15852_
	);
	LUT3 #(
		.INIT('h80)
	) name10026 (
		_w15574_,
		_w15575_,
		_w15573_,
		_w15853_
	);
	LUT3 #(
		.INIT('h10)
	) name10027 (
		_w15574_,
		_w15575_,
		_w15573_,
		_w15854_
	);
	LUT3 #(
		.INIT('hb0)
	) name10028 (
		_w15572_,
		_w15573_,
		_w15578_,
		_w15855_
	);
	LUT4 #(
		.INIT('h0100)
	) name10029 (
		_w15852_,
		_w15854_,
		_w15853_,
		_w15855_,
		_w15856_
	);
	LUT4 #(
		.INIT('h00a3)
	) name10030 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15857_
	);
	LUT4 #(
		.INIT('h00fb)
	) name10031 (
		_w15574_,
		_w15572_,
		_w15573_,
		_w15578_,
		_w15858_
	);
	LUT3 #(
		.INIT('h04)
	) name10032 (
		_w15652_,
		_w15858_,
		_w15857_,
		_w15859_
	);
	LUT4 #(
		.INIT('h1040)
	) name10033 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15860_
	);
	LUT2 #(
		.INIT('h2)
	) name10034 (
		_w15571_,
		_w15860_,
		_w15861_
	);
	LUT3 #(
		.INIT('he0)
	) name10035 (
		_w15856_,
		_w15859_,
		_w15861_,
		_w15862_
	);
	LUT4 #(
		.INIT('h54af)
	) name10036 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15863_
	);
	LUT4 #(
		.INIT('he4f5)
	) name10037 (
		_w15578_,
		_w15596_,
		_w15857_,
		_w15863_,
		_w15864_
	);
	LUT4 #(
		.INIT('h4804)
	) name10038 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w15865_
	);
	LUT2 #(
		.INIT('h1)
	) name10039 (
		_w15571_,
		_w15865_,
		_w15866_
	);
	LUT2 #(
		.INIT('h4)
	) name10040 (
		_w15864_,
		_w15866_,
		_w15867_
	);
	LUT3 #(
		.INIT('ha9)
	) name10041 (
		\u1_L13_reg[28]/NET0131 ,
		_w15862_,
		_w15867_,
		_w15868_
	);
	LUT3 #(
		.INIT('h02)
	) name10042 (
		_w15672_,
		_w15678_,
		_w15819_,
		_w15869_
	);
	LUT4 #(
		.INIT('h4044)
	) name10043 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15870_
	);
	LUT4 #(
		.INIT('h5515)
	) name10044 (
		_w15672_,
		_w15673_,
		_w15674_,
		_w15675_,
		_w15871_
	);
	LUT2 #(
		.INIT('h4)
	) name10045 (
		_w15870_,
		_w15871_,
		_w15872_
	);
	LUT4 #(
		.INIT('hdeaf)
	) name10046 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15873_
	);
	LUT4 #(
		.INIT('h0155)
	) name10047 (
		_w15684_,
		_w15869_,
		_w15872_,
		_w15873_,
		_w15874_
	);
	LUT4 #(
		.INIT('h0001)
	) name10048 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15875_
	);
	LUT4 #(
		.INIT('hf7f6)
	) name10049 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15876_
	);
	LUT3 #(
		.INIT('h04)
	) name10050 (
		_w15672_,
		_w15673_,
		_w15676_,
		_w15877_
	);
	LUT4 #(
		.INIT('h00c4)
	) name10051 (
		_w15672_,
		_w15699_,
		_w15876_,
		_w15877_,
		_w15878_
	);
	LUT4 #(
		.INIT('hcbbf)
	) name10052 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15879_
	);
	LUT4 #(
		.INIT('hcf45)
	) name10053 (
		_w15672_,
		_w15674_,
		_w15833_,
		_w15879_,
		_w15880_
	);
	LUT3 #(
		.INIT('hd0)
	) name10054 (
		_w15684_,
		_w15878_,
		_w15880_,
		_w15881_
	);
	LUT3 #(
		.INIT('h65)
	) name10055 (
		\u1_L13_reg[8]/NET0131 ,
		_w15874_,
		_w15881_,
		_w15882_
	);
	LUT4 #(
		.INIT('h9b99)
	) name10056 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15883_
	);
	LUT3 #(
		.INIT('h19)
	) name10057 (
		_w15415_,
		_w15414_,
		_w15413_,
		_w15884_
	);
	LUT4 #(
		.INIT('hb7ef)
	) name10058 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15885_
	);
	LUT4 #(
		.INIT('h8d00)
	) name10059 (
		_w15412_,
		_w15883_,
		_w15884_,
		_w15885_,
		_w15886_
	);
	LUT4 #(
		.INIT('hf77f)
	) name10060 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15887_
	);
	LUT2 #(
		.INIT('h1)
	) name10061 (
		_w15412_,
		_w15887_,
		_w15888_
	);
	LUT4 #(
		.INIT('h9060)
	) name10062 (
		_w15415_,
		_w15414_,
		_w15416_,
		_w15413_,
		_w15889_
	);
	LUT4 #(
		.INIT('h0013)
	) name10063 (
		_w15434_,
		_w15531_,
		_w15884_,
		_w15889_,
		_w15890_
	);
	LUT4 #(
		.INIT('h0e04)
	) name10064 (
		_w15411_,
		_w15886_,
		_w15888_,
		_w15890_,
		_w15891_
	);
	LUT2 #(
		.INIT('h9)
	) name10065 (
		\u1_L13_reg[9]/NET0131 ,
		_w15891_,
		_w15892_
	);
	LUT4 #(
		.INIT('hdeb9)
	) name10066 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15893_
	);
	LUT2 #(
		.INIT('h1)
	) name10067 (
		_w15446_,
		_w15893_,
		_w15894_
	);
	LUT3 #(
		.INIT('h40)
	) name10068 (
		_w15448_,
		_w15447_,
		_w15449_,
		_w15895_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name10069 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15896_
	);
	LUT4 #(
		.INIT('h1f13)
	) name10070 (
		_w15450_,
		_w15446_,
		_w15895_,
		_w15896_,
		_w15897_
	);
	LUT3 #(
		.INIT('h8a)
	) name10071 (
		_w15445_,
		_w15894_,
		_w15897_,
		_w15898_
	);
	LUT4 #(
		.INIT('h00f7)
	) name10072 (
		_w15450_,
		_w15447_,
		_w15449_,
		_w15446_,
		_w15899_
	);
	LUT4 #(
		.INIT('h0800)
	) name10073 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15900_
	);
	LUT4 #(
		.INIT('hddd8)
	) name10074 (
		_w15446_,
		_w15461_,
		_w15746_,
		_w15900_,
		_w15901_
	);
	LUT3 #(
		.INIT('h10)
	) name10075 (
		_w15448_,
		_w15447_,
		_w15449_,
		_w15902_
	);
	LUT2 #(
		.INIT('h2)
	) name10076 (
		_w15744_,
		_w15902_,
		_w15903_
	);
	LUT4 #(
		.INIT('h58ff)
	) name10077 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15904_
	);
	LUT3 #(
		.INIT('h54)
	) name10078 (
		_w15468_,
		_w15741_,
		_w15904_,
		_w15905_
	);
	LUT4 #(
		.INIT('h2322)
	) name10079 (
		_w15445_,
		_w15901_,
		_w15903_,
		_w15905_,
		_w15906_
	);
	LUT3 #(
		.INIT('h65)
	) name10080 (
		\u1_L13_reg[32]/NET0131 ,
		_w15898_,
		_w15906_,
		_w15907_
	);
	LUT4 #(
		.INIT('h3ffb)
	) name10081 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15908_
	);
	LUT4 #(
		.INIT('hf32e)
	) name10082 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15909_
	);
	LUT4 #(
		.INIT('hed6f)
	) name10083 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15910_
	);
	LUT4 #(
		.INIT('he400)
	) name10084 (
		_w15618_,
		_w15909_,
		_w15908_,
		_w15910_,
		_w15911_
	);
	LUT2 #(
		.INIT('h2)
	) name10085 (
		_w15617_,
		_w15911_,
		_w15912_
	);
	LUT4 #(
		.INIT('haa8a)
	) name10086 (
		_w15618_,
		_w15619_,
		_w15620_,
		_w15622_,
		_w15913_
	);
	LUT4 #(
		.INIT('h4f47)
	) name10087 (
		_w15619_,
		_w15620_,
		_w15622_,
		_w15621_,
		_w15914_
	);
	LUT2 #(
		.INIT('h8)
	) name10088 (
		_w15913_,
		_w15914_,
		_w15915_
	);
	LUT4 #(
		.INIT('h4000)
	) name10089 (
		_w15618_,
		_w15619_,
		_w15622_,
		_w15621_,
		_w15916_
	);
	LUT3 #(
		.INIT('h01)
	) name10090 (
		_w15643_,
		_w15709_,
		_w15916_,
		_w15917_
	);
	LUT3 #(
		.INIT('h45)
	) name10091 (
		_w15617_,
		_w15915_,
		_w15917_,
		_w15918_
	);
	LUT2 #(
		.INIT('h1)
	) name10092 (
		_w15618_,
		_w15642_,
		_w15919_
	);
	LUT4 #(
		.INIT('h0008)
	) name10093 (
		_w15618_,
		_w15619_,
		_w15620_,
		_w15622_,
		_w15920_
	);
	LUT3 #(
		.INIT('h07)
	) name10094 (
		_w15633_,
		_w15648_,
		_w15920_,
		_w15921_
	);
	LUT2 #(
		.INIT('h4)
	) name10095 (
		_w15919_,
		_w15921_,
		_w15922_
	);
	LUT4 #(
		.INIT('h5655)
	) name10096 (
		\u1_L13_reg[27]/NET0131 ,
		_w15918_,
		_w15912_,
		_w15922_,
		_w15923_
	);
	LUT3 #(
		.INIT('h2e)
	) name10097 (
		_w15673_,
		_w15674_,
		_w15676_,
		_w15924_
	);
	LUT3 #(
		.INIT('h04)
	) name10098 (
		_w15673_,
		_w15674_,
		_w15676_,
		_w15925_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name10099 (
		_w15672_,
		_w15673_,
		_w15674_,
		_w15675_,
		_w15926_
	);
	LUT4 #(
		.INIT('h7077)
	) name10100 (
		_w15871_,
		_w15924_,
		_w15925_,
		_w15926_,
		_w15927_
	);
	LUT4 #(
		.INIT('h0d00)
	) name10101 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15928_
	);
	LUT2 #(
		.INIT('h1)
	) name10102 (
		_w15684_,
		_w15928_,
		_w15929_
	);
	LUT4 #(
		.INIT('hef67)
	) name10103 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15930_
	);
	LUT2 #(
		.INIT('h2)
	) name10104 (
		_w15672_,
		_w15930_,
		_w15931_
	);
	LUT4 #(
		.INIT('h0200)
	) name10105 (
		_w15673_,
		_w15674_,
		_w15675_,
		_w15676_,
		_w15932_
	);
	LUT4 #(
		.INIT('h1000)
	) name10106 (
		_w15672_,
		_w15673_,
		_w15674_,
		_w15675_,
		_w15933_
	);
	LUT4 #(
		.INIT('h0004)
	) name10107 (
		_w15677_,
		_w15684_,
		_w15932_,
		_w15933_,
		_w15934_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name10108 (
		_w15927_,
		_w15929_,
		_w15931_,
		_w15934_,
		_w15935_
	);
	LUT3 #(
		.INIT('h02)
	) name10109 (
		_w15672_,
		_w15678_,
		_w15698_,
		_w15936_
	);
	LUT4 #(
		.INIT('h0001)
	) name10110 (
		_w15672_,
		_w15681_,
		_w15696_,
		_w15875_,
		_w15937_
	);
	LUT2 #(
		.INIT('h1)
	) name10111 (
		_w15936_,
		_w15937_,
		_w15938_
	);
	LUT3 #(
		.INIT('h56)
	) name10112 (
		\u1_L13_reg[3]/NET0131 ,
		_w15935_,
		_w15938_,
		_w15939_
	);
	LUT4 #(
		.INIT('hc693)
	) name10113 (
		decrypt_pad,
		\u1_R13_reg[11]/P0001 ,
		\u1_uk_K_r13_reg[20]/NET0131 ,
		\u1_uk_K_r13_reg[41]/NET0131 ,
		_w15940_
	);
	LUT4 #(
		.INIT('hc963)
	) name10114 (
		decrypt_pad,
		\u1_R13_reg[12]/NET0131 ,
		\u1_uk_K_r13_reg[24]/NET0131 ,
		\u1_uk_K_r13_reg[3]/NET0131 ,
		_w15941_
	);
	LUT4 #(
		.INIT('hc963)
	) name10115 (
		decrypt_pad,
		\u1_R13_reg[13]/NET0131 ,
		\u1_uk_K_r13_reg[12]/NET0131 ,
		\u1_uk_K_r13_reg[48]/NET0131 ,
		_w15942_
	);
	LUT4 #(
		.INIT('hc693)
	) name10116 (
		decrypt_pad,
		\u1_R13_reg[9]/NET0131 ,
		\u1_uk_K_r13_reg[11]/NET0131 ,
		\u1_uk_K_r13_reg[32]/NET0131 ,
		_w15943_
	);
	LUT4 #(
		.INIT('hc693)
	) name10117 (
		decrypt_pad,
		\u1_R13_reg[10]/NET0131 ,
		\u1_uk_K_r13_reg[19]/NET0131 ,
		\u1_uk_K_r13_reg[40]/NET0131 ,
		_w15944_
	);
	LUT4 #(
		.INIT('hc693)
	) name10118 (
		decrypt_pad,
		\u1_R13_reg[8]/NET0131 ,
		\u1_uk_K_r13_reg[39]/NET0131 ,
		\u1_uk_K_r13_reg[3]/NET0131 ,
		_w15945_
	);
	LUT4 #(
		.INIT('h95b5)
	) name10119 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w15946_
	);
	LUT2 #(
		.INIT('h1)
	) name10120 (
		_w15942_,
		_w15945_,
		_w15947_
	);
	LUT4 #(
		.INIT('h0001)
	) name10121 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w15948_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name10122 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w15949_
	);
	LUT4 #(
		.INIT('h08cc)
	) name10123 (
		_w15941_,
		_w15940_,
		_w15946_,
		_w15949_,
		_w15950_
	);
	LUT2 #(
		.INIT('h1)
	) name10124 (
		_w15943_,
		_w15944_,
		_w15951_
	);
	LUT2 #(
		.INIT('h6)
	) name10125 (
		_w15943_,
		_w15944_,
		_w15952_
	);
	LUT2 #(
		.INIT('h9)
	) name10126 (
		_w15942_,
		_w15945_,
		_w15953_
	);
	LUT3 #(
		.INIT('h46)
	) name10127 (
		_w15942_,
		_w15945_,
		_w15940_,
		_w15954_
	);
	LUT2 #(
		.INIT('h1)
	) name10128 (
		_w15952_,
		_w15954_,
		_w15955_
	);
	LUT4 #(
		.INIT('h383c)
	) name10129 (
		_w15945_,
		_w15943_,
		_w15944_,
		_w15940_,
		_w15956_
	);
	LUT3 #(
		.INIT('h45)
	) name10130 (
		_w15941_,
		_w15953_,
		_w15956_,
		_w15957_
	);
	LUT3 #(
		.INIT('h80)
	) name10131 (
		_w15943_,
		_w15944_,
		_w15941_,
		_w15958_
	);
	LUT3 #(
		.INIT('h51)
	) name10132 (
		_w15945_,
		_w15943_,
		_w15944_,
		_w15959_
	);
	LUT2 #(
		.INIT('h2)
	) name10133 (
		_w15941_,
		_w15940_,
		_w15960_
	);
	LUT4 #(
		.INIT('h0090)
	) name10134 (
		_w15942_,
		_w15943_,
		_w15941_,
		_w15940_,
		_w15961_
	);
	LUT4 #(
		.INIT('h7077)
	) name10135 (
		_w15947_,
		_w15958_,
		_w15959_,
		_w15961_,
		_w15962_
	);
	LUT4 #(
		.INIT('h4500)
	) name10136 (
		_w15950_,
		_w15955_,
		_w15957_,
		_w15962_,
		_w15963_
	);
	LUT2 #(
		.INIT('h9)
	) name10137 (
		\u1_L13_reg[6]/NET0131 ,
		_w15963_,
		_w15964_
	);
	LUT3 #(
		.INIT('h48)
	) name10138 (
		_w15448_,
		_w15450_,
		_w15449_,
		_w15965_
	);
	LUT4 #(
		.INIT('h4080)
	) name10139 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15966_
	);
	LUT4 #(
		.INIT('h9f7f)
	) name10140 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15967_
	);
	LUT3 #(
		.INIT('h21)
	) name10141 (
		_w15448_,
		_w15447_,
		_w15449_,
		_w15968_
	);
	LUT4 #(
		.INIT('h0a04)
	) name10142 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15969_
	);
	LUT2 #(
		.INIT('h2)
	) name10143 (
		_w15446_,
		_w15969_,
		_w15970_
	);
	LUT4 #(
		.INIT('haffc)
	) name10144 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15971_
	);
	LUT3 #(
		.INIT('h20)
	) name10145 (
		_w15899_,
		_w15965_,
		_w15971_,
		_w15972_
	);
	LUT4 #(
		.INIT('h222a)
	) name10146 (
		_w15445_,
		_w15967_,
		_w15970_,
		_w15972_,
		_w15973_
	);
	LUT4 #(
		.INIT('h0010)
	) name10147 (
		_w15448_,
		_w15450_,
		_w15447_,
		_w15449_,
		_w15974_
	);
	LUT4 #(
		.INIT('h5510)
	) name10148 (
		_w15445_,
		_w15446_,
		_w15969_,
		_w15974_,
		_w15975_
	);
	LUT2 #(
		.INIT('h1)
	) name10149 (
		_w15446_,
		_w15967_,
		_w15976_
	);
	LUT4 #(
		.INIT('hdf00)
	) name10150 (
		_w15448_,
		_w15450_,
		_w15449_,
		_w15446_,
		_w15977_
	);
	LUT4 #(
		.INIT('h3100)
	) name10151 (
		_w15445_,
		_w15968_,
		_w15974_,
		_w15977_,
		_w15978_
	);
	LUT4 #(
		.INIT('h0203)
	) name10152 (
		_w15966_,
		_w15976_,
		_w15975_,
		_w15978_,
		_w15979_
	);
	LUT3 #(
		.INIT('h65)
	) name10153 (
		\u1_L13_reg[7]/NET0131 ,
		_w15973_,
		_w15979_,
		_w15980_
	);
	LUT4 #(
		.INIT('heed9)
	) name10154 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w15981_
	);
	LUT3 #(
		.INIT('ha2)
	) name10155 (
		_w15941_,
		_w15940_,
		_w15981_,
		_w15982_
	);
	LUT4 #(
		.INIT('h8c00)
	) name10156 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w15983_
	);
	LUT3 #(
		.INIT('h04)
	) name10157 (
		_w15942_,
		_w15943_,
		_w15944_,
		_w15984_
	);
	LUT2 #(
		.INIT('h4)
	) name10158 (
		_w15941_,
		_w15940_,
		_w15985_
	);
	LUT3 #(
		.INIT('h10)
	) name10159 (
		_w15984_,
		_w15983_,
		_w15985_,
		_w15986_
	);
	LUT4 #(
		.INIT('h008c)
	) name10160 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w15987_
	);
	LUT4 #(
		.INIT('h00df)
	) name10161 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15940_,
		_w15988_
	);
	LUT2 #(
		.INIT('h4)
	) name10162 (
		_w15987_,
		_w15988_,
		_w15989_
	);
	LUT4 #(
		.INIT('hfdf6)
	) name10163 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w15990_
	);
	LUT4 #(
		.INIT('h0155)
	) name10164 (
		_w15982_,
		_w15986_,
		_w15989_,
		_w15990_,
		_w15991_
	);
	LUT4 #(
		.INIT('h23ef)
	) name10165 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w15992_
	);
	LUT2 #(
		.INIT('h2)
	) name10166 (
		_w15960_,
		_w15992_,
		_w15993_
	);
	LUT2 #(
		.INIT('h8)
	) name10167 (
		_w15944_,
		_w15940_,
		_w15994_
	);
	LUT2 #(
		.INIT('h8)
	) name10168 (
		_w15942_,
		_w15945_,
		_w15995_
	);
	LUT3 #(
		.INIT('h08)
	) name10169 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15996_
	);
	LUT2 #(
		.INIT('h8)
	) name10170 (
		_w15994_,
		_w15996_,
		_w15997_
	);
	LUT4 #(
		.INIT('h0040)
	) name10171 (
		_w15942_,
		_w15943_,
		_w15944_,
		_w15940_,
		_w15998_
	);
	LUT3 #(
		.INIT('h0d)
	) name10172 (
		_w15958_,
		_w15995_,
		_w15998_,
		_w15999_
	);
	LUT3 #(
		.INIT('h10)
	) name10173 (
		_w15993_,
		_w15997_,
		_w15999_,
		_w16000_
	);
	LUT3 #(
		.INIT('h9a)
	) name10174 (
		\u1_L13_reg[30]/NET0131 ,
		_w15991_,
		_w16000_,
		_w16001_
	);
	LUT3 #(
		.INIT('hbe)
	) name10175 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w16002_
	);
	LUT2 #(
		.INIT('h2)
	) name10176 (
		_w15994_,
		_w16002_,
		_w16003_
	);
	LUT4 #(
		.INIT('hdf00)
	) name10177 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w16004_
	);
	LUT3 #(
		.INIT('h80)
	) name10178 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w16005_
	);
	LUT3 #(
		.INIT('h7d)
	) name10179 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w16006_
	);
	LUT4 #(
		.INIT('h1000)
	) name10180 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15940_,
		_w16007_
	);
	LUT4 #(
		.INIT('h00fb)
	) name10181 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w16008_
	);
	LUT4 #(
		.INIT('h5155)
	) name10182 (
		_w16004_,
		_w16006_,
		_w16007_,
		_w16008_,
		_w16009_
	);
	LUT4 #(
		.INIT('he2bb)
	) name10183 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w16010_
	);
	LUT3 #(
		.INIT('ha8)
	) name10184 (
		_w15941_,
		_w15940_,
		_w16010_,
		_w16011_
	);
	LUT4 #(
		.INIT('h716c)
	) name10185 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w16012_
	);
	LUT2 #(
		.INIT('h1)
	) name10186 (
		_w15940_,
		_w16012_,
		_w16013_
	);
	LUT4 #(
		.INIT('h6800)
	) name10187 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15940_,
		_w16014_
	);
	LUT3 #(
		.INIT('h01)
	) name10188 (
		_w15941_,
		_w15948_,
		_w16014_,
		_w16015_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name10189 (
		_w16009_,
		_w16011_,
		_w16013_,
		_w16015_,
		_w16016_
	);
	LUT3 #(
		.INIT('h56)
	) name10190 (
		\u1_L13_reg[16]/NET0131 ,
		_w16003_,
		_w16016_,
		_w16017_
	);
	LUT4 #(
		.INIT('h2600)
	) name10191 (
		_w15574_,
		_w15575_,
		_w15573_,
		_w15578_,
		_w16018_
	);
	LUT4 #(
		.INIT('hcaff)
	) name10192 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w16019_
	);
	LUT4 #(
		.INIT('h0032)
	) name10193 (
		_w15578_,
		_w15597_,
		_w16019_,
		_w16018_,
		_w16020_
	);
	LUT4 #(
		.INIT('h0109)
	) name10194 (
		_w15574_,
		_w15572_,
		_w15573_,
		_w15578_,
		_w16021_
	);
	LUT2 #(
		.INIT('h2)
	) name10195 (
		_w15575_,
		_w15578_,
		_w16022_
	);
	LUT4 #(
		.INIT('ha800)
	) name10196 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w16023_
	);
	LUT4 #(
		.INIT('hbefe)
	) name10197 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w16024_
	);
	LUT4 #(
		.INIT('h0b00)
	) name10198 (
		_w16022_,
		_w16023_,
		_w16021_,
		_w16024_,
		_w16025_
	);
	LUT4 #(
		.INIT('h0008)
	) name10199 (
		_w15574_,
		_w15575_,
		_w15573_,
		_w15578_,
		_w16026_
	);
	LUT4 #(
		.INIT('h33f5)
	) name10200 (
		_w15574_,
		_w15572_,
		_w15575_,
		_w15573_,
		_w16027_
	);
	LUT3 #(
		.INIT('hd0)
	) name10201 (
		_w15572_,
		_w15575_,
		_w15578_,
		_w16028_
	);
	LUT3 #(
		.INIT('h45)
	) name10202 (
		_w16026_,
		_w16027_,
		_w16028_,
		_w16029_
	);
	LUT4 #(
		.INIT('hd800)
	) name10203 (
		_w15571_,
		_w16020_,
		_w16025_,
		_w16029_,
		_w16030_
	);
	LUT2 #(
		.INIT('h9)
	) name10204 (
		\u1_L13_reg[18]/P0001 ,
		_w16030_,
		_w16031_
	);
	LUT4 #(
		.INIT('he2cd)
	) name10205 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w16032_
	);
	LUT4 #(
		.INIT('h0400)
	) name10206 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w16033_
	);
	LUT4 #(
		.INIT('h5504)
	) name10207 (
		_w15941_,
		_w15940_,
		_w16032_,
		_w16033_,
		_w16034_
	);
	LUT2 #(
		.INIT('h8)
	) name10208 (
		_w15951_,
		_w15954_,
		_w16035_
	);
	LUT4 #(
		.INIT('h1dff)
	) name10209 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w16036_
	);
	LUT2 #(
		.INIT('h2)
	) name10210 (
		_w15940_,
		_w16036_,
		_w16037_
	);
	LUT3 #(
		.INIT('h0e)
	) name10211 (
		_w15943_,
		_w15944_,
		_w15940_,
		_w16038_
	);
	LUT2 #(
		.INIT('h4)
	) name10212 (
		_w15944_,
		_w15940_,
		_w16039_
	);
	LUT3 #(
		.INIT('h0d)
	) name10213 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w16040_
	);
	LUT4 #(
		.INIT('h0777)
	) name10214 (
		_w15953_,
		_w16038_,
		_w16039_,
		_w16040_,
		_w16041_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10215 (
		_w15941_,
		_w16037_,
		_w16035_,
		_w16041_,
		_w16042_
	);
	LUT4 #(
		.INIT('h9db6)
	) name10216 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w15944_,
		_w16043_
	);
	LUT2 #(
		.INIT('h1)
	) name10217 (
		_w15941_,
		_w15940_,
		_w16044_
	);
	LUT2 #(
		.INIT('h4)
	) name10218 (
		_w16043_,
		_w16044_,
		_w16045_
	);
	LUT3 #(
		.INIT('hdb)
	) name10219 (
		_w15942_,
		_w15945_,
		_w15943_,
		_w16046_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name10220 (
		_w15944_,
		_w15940_,
		_w16005_,
		_w16046_,
		_w16047_
	);
	LUT2 #(
		.INIT('h4)
	) name10221 (
		_w16045_,
		_w16047_,
		_w16048_
	);
	LUT4 #(
		.INIT('h5655)
	) name10222 (
		\u1_L13_reg[24]/NET0131 ,
		_w16042_,
		_w16034_,
		_w16048_,
		_w16049_
	);
	LUT4 #(
		.INIT('hc693)
	) name10223 (
		decrypt_pad,
		\u1_R12_reg[28]/NET0131 ,
		\u1_uk_K_r12_reg[14]/NET0131 ,
		\u1_uk_K_r12_reg[8]/NET0131 ,
		_w16050_
	);
	LUT4 #(
		.INIT('hc963)
	) name10224 (
		decrypt_pad,
		\u1_R12_reg[27]/NET0131 ,
		\u1_uk_K_r12_reg[21]/NET0131 ,
		\u1_uk_K_r12_reg[31]/NET0131 ,
		_w16051_
	);
	LUT4 #(
		.INIT('hc963)
	) name10225 (
		decrypt_pad,
		\u1_R12_reg[24]/NET0131 ,
		\u1_uk_K_r12_reg[23]/NET0131 ,
		\u1_uk_K_r12_reg[29]/NET0131 ,
		_w16052_
	);
	LUT4 #(
		.INIT('hc963)
	) name10226 (
		decrypt_pad,
		\u1_R12_reg[26]/NET0131 ,
		\u1_uk_K_r12_reg[43]/NET0131 ,
		\u1_uk_K_r12_reg[49]/NET0131 ,
		_w16053_
	);
	LUT4 #(
		.INIT('hc963)
	) name10227 (
		decrypt_pad,
		\u1_R12_reg[29]/NET0131 ,
		\u1_uk_K_r12_reg[0]/NET0131 ,
		\u1_uk_K_r12_reg[37]/NET0131 ,
		_w16054_
	);
	LUT4 #(
		.INIT('hc963)
	) name10228 (
		decrypt_pad,
		\u1_R12_reg[25]/NET0131 ,
		\u1_uk_K_r12_reg[31]/NET0131 ,
		\u1_uk_K_r12_reg[9]/NET0131 ,
		_w16055_
	);
	LUT4 #(
		.INIT('h0080)
	) name10229 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16056_
	);
	LUT4 #(
		.INIT('hf37f)
	) name10230 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16057_
	);
	LUT3 #(
		.INIT('h08)
	) name10231 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16058_
	);
	LUT4 #(
		.INIT('h0008)
	) name10232 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16059_
	);
	LUT4 #(
		.INIT('hdfd7)
	) name10233 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16060_
	);
	LUT4 #(
		.INIT('h0200)
	) name10234 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16061_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name10235 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16062_
	);
	LUT4 #(
		.INIT('he400)
	) name10236 (
		_w16051_,
		_w16060_,
		_w16057_,
		_w16062_,
		_w16063_
	);
	LUT2 #(
		.INIT('h2)
	) name10237 (
		_w16050_,
		_w16063_,
		_w16064_
	);
	LUT4 #(
		.INIT('h0100)
	) name10238 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16065_
	);
	LUT4 #(
		.INIT('h36bf)
	) name10239 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16066_
	);
	LUT2 #(
		.INIT('h1)
	) name10240 (
		_w16051_,
		_w16066_,
		_w16067_
	);
	LUT3 #(
		.INIT('h51)
	) name10241 (
		_w16051_,
		_w16054_,
		_w16052_,
		_w16068_
	);
	LUT4 #(
		.INIT('h005d)
	) name10242 (
		_w16051_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16069_
	);
	LUT3 #(
		.INIT('h04)
	) name10243 (
		_w16054_,
		_w16052_,
		_w16053_,
		_w16070_
	);
	LUT4 #(
		.INIT('h7fdb)
	) name10244 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16071_
	);
	LUT3 #(
		.INIT('hb0)
	) name10245 (
		_w16068_,
		_w16069_,
		_w16071_,
		_w16072_
	);
	LUT4 #(
		.INIT('h1000)
	) name10246 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16073_
	);
	LUT4 #(
		.INIT('he9fb)
	) name10247 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16074_
	);
	LUT4 #(
		.INIT('h0002)
	) name10248 (
		_w16051_,
		_w16054_,
		_w16055_,
		_w16053_,
		_w16075_
	);
	LUT4 #(
		.INIT('h4010)
	) name10249 (
		_w16051_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16076_
	);
	LUT4 #(
		.INIT('h000d)
	) name10250 (
		_w16051_,
		_w16074_,
		_w16075_,
		_w16076_,
		_w16077_
	);
	LUT4 #(
		.INIT('hba00)
	) name10251 (
		_w16050_,
		_w16067_,
		_w16072_,
		_w16077_,
		_w16078_
	);
	LUT3 #(
		.INIT('h65)
	) name10252 (
		\u1_L12_reg[22]/NET0131 ,
		_w16064_,
		_w16078_,
		_w16079_
	);
	LUT4 #(
		.INIT('hc693)
	) name10253 (
		decrypt_pad,
		\u1_R12_reg[4]/NET0131 ,
		\u1_uk_K_r12_reg[10]/P0001 ,
		\u1_uk_K_r12_reg[34]/NET0131 ,
		_w16080_
	);
	LUT4 #(
		.INIT('hc963)
	) name10254 (
		decrypt_pad,
		\u1_R12_reg[1]/NET0131 ,
		\u1_uk_K_r12_reg[32]/NET0131 ,
		\u1_uk_K_r12_reg[40]/NET0131 ,
		_w16081_
	);
	LUT4 #(
		.INIT('hc693)
	) name10255 (
		decrypt_pad,
		\u1_R12_reg[5]/NET0131 ,
		\u1_uk_K_r12_reg[13]/NET0131 ,
		\u1_uk_K_r12_reg[5]/NET0131 ,
		_w16082_
	);
	LUT4 #(
		.INIT('hc963)
	) name10256 (
		decrypt_pad,
		\u1_R12_reg[32]/NET0131 ,
		\u1_uk_K_r12_reg[11]/NET0131 ,
		\u1_uk_K_r12_reg[19]/NET0131 ,
		_w16083_
	);
	LUT4 #(
		.INIT('hc963)
	) name10257 (
		decrypt_pad,
		\u1_R12_reg[2]/NET0131 ,
		\u1_uk_K_r12_reg[47]/NET0131 ,
		\u1_uk_K_r12_reg[55]/NET0131 ,
		_w16084_
	);
	LUT4 #(
		.INIT('heff4)
	) name10258 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16085_
	);
	LUT4 #(
		.INIT('hc963)
	) name10259 (
		decrypt_pad,
		\u1_R12_reg[3]/NET0131 ,
		\u1_uk_K_r12_reg[24]/NET0131 ,
		\u1_uk_K_r12_reg[32]/NET0131 ,
		_w16086_
	);
	LUT2 #(
		.INIT('h1)
	) name10260 (
		_w16085_,
		_w16086_,
		_w16087_
	);
	LUT4 #(
		.INIT('hc040)
	) name10261 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16086_,
		_w16088_
	);
	LUT3 #(
		.INIT('h02)
	) name10262 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16089_
	);
	LUT4 #(
		.INIT('h00fd)
	) name10263 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16090_
	);
	LUT3 #(
		.INIT('h28)
	) name10264 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16091_
	);
	LUT4 #(
		.INIT('hd700)
	) name10265 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16092_
	);
	LUT2 #(
		.INIT('h2)
	) name10266 (
		_w16084_,
		_w16086_,
		_w16093_
	);
	LUT4 #(
		.INIT('h1011)
	) name10267 (
		_w16092_,
		_w16093_,
		_w16088_,
		_w16090_,
		_w16094_
	);
	LUT3 #(
		.INIT('h54)
	) name10268 (
		_w16080_,
		_w16087_,
		_w16094_,
		_w16095_
	);
	LUT3 #(
		.INIT('h10)
	) name10269 (
		_w16082_,
		_w16083_,
		_w16084_,
		_w16096_
	);
	LUT4 #(
		.INIT('hb8bb)
	) name10270 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16097_
	);
	LUT2 #(
		.INIT('h2)
	) name10271 (
		_w16086_,
		_w16097_,
		_w16098_
	);
	LUT4 #(
		.INIT('h0510)
	) name10272 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16099_
	);
	LUT2 #(
		.INIT('h2)
	) name10273 (
		_w16082_,
		_w16083_,
		_w16100_
	);
	LUT2 #(
		.INIT('h4)
	) name10274 (
		_w16084_,
		_w16086_,
		_w16101_
	);
	LUT3 #(
		.INIT('h8a)
	) name10275 (
		_w16081_,
		_w16084_,
		_w16086_,
		_w16102_
	);
	LUT3 #(
		.INIT('h08)
	) name10276 (
		_w16081_,
		_w16083_,
		_w16086_,
		_w16103_
	);
	LUT4 #(
		.INIT('h000d)
	) name10277 (
		_w16100_,
		_w16102_,
		_w16103_,
		_w16099_,
		_w16104_
	);
	LUT3 #(
		.INIT('h8a)
	) name10278 (
		_w16080_,
		_w16098_,
		_w16104_,
		_w16105_
	);
	LUT3 #(
		.INIT('h80)
	) name10279 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16106_
	);
	LUT4 #(
		.INIT('h7bdd)
	) name10280 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16107_
	);
	LUT2 #(
		.INIT('h1)
	) name10281 (
		_w16086_,
		_w16107_,
		_w16108_
	);
	LUT2 #(
		.INIT('h4)
	) name10282 (
		_w16081_,
		_w16086_,
		_w16109_
	);
	LUT4 #(
		.INIT('h0400)
	) name10283 (
		_w16081_,
		_w16083_,
		_w16084_,
		_w16086_,
		_w16110_
	);
	LUT3 #(
		.INIT('h07)
	) name10284 (
		_w16096_,
		_w16109_,
		_w16110_,
		_w16111_
	);
	LUT2 #(
		.INIT('h4)
	) name10285 (
		_w16108_,
		_w16111_,
		_w16112_
	);
	LUT4 #(
		.INIT('h5655)
	) name10286 (
		\u1_L12_reg[31]/NET0131 ,
		_w16095_,
		_w16105_,
		_w16112_,
		_w16113_
	);
	LUT4 #(
		.INIT('hc963)
	) name10287 (
		decrypt_pad,
		\u1_R12_reg[24]/NET0131 ,
		\u1_uk_K_r12_reg[1]/NET0131 ,
		\u1_uk_K_r12_reg[7]/P0001 ,
		_w16114_
	);
	LUT4 #(
		.INIT('hc963)
	) name10288 (
		decrypt_pad,
		\u1_R12_reg[23]/NET0131 ,
		\u1_uk_K_r12_reg[30]/NET0131 ,
		\u1_uk_K_r12_reg[36]/NET0131 ,
		_w16115_
	);
	LUT4 #(
		.INIT('hc693)
	) name10289 (
		decrypt_pad,
		\u1_R12_reg[21]/NET0131 ,
		\u1_uk_K_r12_reg[1]/NET0131 ,
		\u1_uk_K_r12_reg[50]/NET0131 ,
		_w16116_
	);
	LUT4 #(
		.INIT('hc963)
	) name10290 (
		decrypt_pad,
		\u1_R12_reg[20]/NET0131 ,
		\u1_uk_K_r12_reg[35]/NET0131 ,
		\u1_uk_K_r12_reg[45]/NET0131 ,
		_w16117_
	);
	LUT4 #(
		.INIT('hc693)
	) name10291 (
		decrypt_pad,
		\u1_R12_reg[25]/NET0131 ,
		\u1_uk_K_r12_reg[2]/NET0131 ,
		\u1_uk_K_r12_reg[51]/NET0131 ,
		_w16118_
	);
	LUT4 #(
		.INIT('hc693)
	) name10292 (
		decrypt_pad,
		\u1_R12_reg[22]/NET0131 ,
		\u1_uk_K_r12_reg[23]/NET0131 ,
		\u1_uk_K_r12_reg[45]/NET0131 ,
		_w16119_
	);
	LUT3 #(
		.INIT('h08)
	) name10293 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16120_
	);
	LUT4 #(
		.INIT('h0010)
	) name10294 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16121_
	);
	LUT4 #(
		.INIT('h37e7)
	) name10295 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16122_
	);
	LUT2 #(
		.INIT('h2)
	) name10296 (
		_w16115_,
		_w16122_,
		_w16123_
	);
	LUT2 #(
		.INIT('h1)
	) name10297 (
		_w16119_,
		_w16115_,
		_w16124_
	);
	LUT4 #(
		.INIT('h0400)
	) name10298 (
		_w16119_,
		_w16117_,
		_w16115_,
		_w16118_,
		_w16125_
	);
	LUT2 #(
		.INIT('h4)
	) name10299 (
		_w16116_,
		_w16125_,
		_w16126_
	);
	LUT3 #(
		.INIT('h15)
	) name10300 (
		_w16119_,
		_w16116_,
		_w16118_,
		_w16127_
	);
	LUT3 #(
		.INIT('h13)
	) name10301 (
		_w16117_,
		_w16115_,
		_w16118_,
		_w16128_
	);
	LUT3 #(
		.INIT('h10)
	) name10302 (
		_w16120_,
		_w16127_,
		_w16128_,
		_w16129_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10303 (
		_w16114_,
		_w16123_,
		_w16126_,
		_w16129_,
		_w16130_
	);
	LUT4 #(
		.INIT('h0048)
	) name10304 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16115_,
		_w16131_
	);
	LUT4 #(
		.INIT('h0004)
	) name10305 (
		_w16119_,
		_w16117_,
		_w16115_,
		_w16118_,
		_w16132_
	);
	LUT4 #(
		.INIT('h2000)
	) name10306 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16133_
	);
	LUT2 #(
		.INIT('h1)
	) name10307 (
		_w16132_,
		_w16133_,
		_w16134_
	);
	LUT3 #(
		.INIT('hb0)
	) name10308 (
		_w16119_,
		_w16117_,
		_w16115_,
		_w16135_
	);
	LUT4 #(
		.INIT('h2500)
	) name10309 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16115_,
		_w16136_
	);
	LUT4 #(
		.INIT('h1000)
	) name10310 (
		_w16116_,
		_w16117_,
		_w16115_,
		_w16118_,
		_w16137_
	);
	LUT4 #(
		.INIT('h0040)
	) name10311 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16138_
	);
	LUT3 #(
		.INIT('h01)
	) name10312 (
		_w16136_,
		_w16137_,
		_w16138_,
		_w16139_
	);
	LUT4 #(
		.INIT('h00bf)
	) name10313 (
		_w16131_,
		_w16134_,
		_w16139_,
		_w16114_,
		_w16140_
	);
	LUT4 #(
		.INIT('heff7)
	) name10314 (
		_w16116_,
		_w16117_,
		_w16115_,
		_w16118_,
		_w16141_
	);
	LUT2 #(
		.INIT('h1)
	) name10315 (
		_w16119_,
		_w16141_,
		_w16142_
	);
	LUT3 #(
		.INIT('h01)
	) name10316 (
		_w16116_,
		_w16117_,
		_w16118_,
		_w16143_
	);
	LUT4 #(
		.INIT('h0fbb)
	) name10317 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16144_
	);
	LUT4 #(
		.INIT('h3f15)
	) name10318 (
		_w16135_,
		_w16124_,
		_w16143_,
		_w16144_,
		_w16145_
	);
	LUT2 #(
		.INIT('h4)
	) name10319 (
		_w16142_,
		_w16145_,
		_w16146_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name10320 (
		\u1_L12_reg[11]/NET0131 ,
		_w16140_,
		_w16130_,
		_w16146_,
		_w16147_
	);
	LUT4 #(
		.INIT('hc963)
	) name10321 (
		decrypt_pad,
		\u1_R12_reg[13]/NET0131 ,
		\u1_uk_K_r12_reg[19]/NET0131 ,
		\u1_uk_K_r12_reg[27]/NET0131 ,
		_w16148_
	);
	LUT4 #(
		.INIT('hc963)
	) name10322 (
		decrypt_pad,
		\u1_R12_reg[12]/NET0131 ,
		\u1_uk_K_r12_reg[25]/NET0131 ,
		\u1_uk_K_r12_reg[33]/NET0131 ,
		_w16149_
	);
	LUT4 #(
		.INIT('hc693)
	) name10323 (
		decrypt_pad,
		\u1_R12_reg[17]/NET0131 ,
		\u1_uk_K_r12_reg[17]/NET0131 ,
		\u1_uk_K_r12_reg[41]/NET0131 ,
		_w16150_
	);
	LUT2 #(
		.INIT('h1)
	) name10324 (
		_w16149_,
		_w16150_,
		_w16151_
	);
	LUT4 #(
		.INIT('hc963)
	) name10325 (
		decrypt_pad,
		\u1_R12_reg[14]/NET0131 ,
		\u1_uk_K_r12_reg[20]/NET0131 ,
		\u1_uk_K_r12_reg[53]/NET0131 ,
		_w16152_
	);
	LUT4 #(
		.INIT('h0200)
	) name10326 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16153_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name10327 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16154_
	);
	LUT4 #(
		.INIT('hc693)
	) name10328 (
		decrypt_pad,
		\u1_R12_reg[15]/NET0131 ,
		\u1_uk_K_r12_reg[4]/NET0131 ,
		\u1_uk_K_r12_reg[53]/NET0131 ,
		_w16155_
	);
	LUT3 #(
		.INIT('h80)
	) name10329 (
		_w16148_,
		_w16155_,
		_w16152_,
		_w16156_
	);
	LUT4 #(
		.INIT('h0800)
	) name10330 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16152_,
		_w16157_
	);
	LUT2 #(
		.INIT('h2)
	) name10331 (
		_w16150_,
		_w16152_,
		_w16158_
	);
	LUT4 #(
		.INIT('h0040)
	) name10332 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16159_
	);
	LUT4 #(
		.INIT('hc693)
	) name10333 (
		decrypt_pad,
		\u1_R12_reg[16]/NET0131 ,
		\u1_uk_K_r12_reg[12]/NET0131 ,
		\u1_uk_K_r12_reg[4]/NET0131 ,
		_w16160_
	);
	LUT4 #(
		.INIT('h0002)
	) name10334 (
		_w16154_,
		_w16159_,
		_w16157_,
		_w16160_,
		_w16161_
	);
	LUT4 #(
		.INIT('ha3af)
	) name10335 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16162_
	);
	LUT4 #(
		.INIT('h8004)
	) name10336 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16150_,
		_w16163_
	);
	LUT3 #(
		.INIT('h0e)
	) name10337 (
		_w16155_,
		_w16162_,
		_w16163_,
		_w16164_
	);
	LUT2 #(
		.INIT('h8)
	) name10338 (
		_w16161_,
		_w16164_,
		_w16165_
	);
	LUT4 #(
		.INIT('h0080)
	) name10339 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16150_,
		_w16166_
	);
	LUT2 #(
		.INIT('h4)
	) name10340 (
		_w16149_,
		_w16150_,
		_w16167_
	);
	LUT3 #(
		.INIT('h20)
	) name10341 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16168_
	);
	LUT4 #(
		.INIT('h0020)
	) name10342 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16169_
	);
	LUT2 #(
		.INIT('h1)
	) name10343 (
		_w16166_,
		_w16169_,
		_w16170_
	);
	LUT2 #(
		.INIT('h1)
	) name10344 (
		_w16155_,
		_w16150_,
		_w16171_
	);
	LUT3 #(
		.INIT('h10)
	) name10345 (
		_w16148_,
		_w16149_,
		_w16152_,
		_w16172_
	);
	LUT2 #(
		.INIT('h8)
	) name10346 (
		_w16171_,
		_w16172_,
		_w16173_
	);
	LUT4 #(
		.INIT('h8000)
	) name10347 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16174_
	);
	LUT4 #(
		.INIT('h002a)
	) name10348 (
		_w16160_,
		_w16171_,
		_w16172_,
		_w16174_,
		_w16175_
	);
	LUT4 #(
		.INIT('h0012)
	) name10349 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16152_,
		_w16176_
	);
	LUT4 #(
		.INIT('h0400)
	) name10350 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16150_,
		_w16177_
	);
	LUT2 #(
		.INIT('h1)
	) name10351 (
		_w16176_,
		_w16177_,
		_w16178_
	);
	LUT3 #(
		.INIT('h80)
	) name10352 (
		_w16170_,
		_w16175_,
		_w16178_,
		_w16179_
	);
	LUT2 #(
		.INIT('h4)
	) name10353 (
		_w16148_,
		_w16155_,
		_w16180_
	);
	LUT3 #(
		.INIT('hde)
	) name10354 (
		_w16149_,
		_w16150_,
		_w16152_,
		_w16181_
	);
	LUT2 #(
		.INIT('h2)
	) name10355 (
		_w16180_,
		_w16181_,
		_w16182_
	);
	LUT4 #(
		.INIT('hcecf)
	) name10356 (
		_w16155_,
		_w16152_,
		_w16166_,
		_w16168_,
		_w16183_
	);
	LUT2 #(
		.INIT('h4)
	) name10357 (
		_w16182_,
		_w16183_,
		_w16184_
	);
	LUT4 #(
		.INIT('ha955)
	) name10358 (
		\u1_L12_reg[20]/NET0131 ,
		_w16165_,
		_w16179_,
		_w16184_,
		_w16185_
	);
	LUT4 #(
		.INIT('h0040)
	) name10359 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16186_
	);
	LUT4 #(
		.INIT('hf0b5)
	) name10360 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16187_
	);
	LUT4 #(
		.INIT('h00c1)
	) name10361 (
		_w16081_,
		_w16083_,
		_w16084_,
		_w16086_,
		_w16188_
	);
	LUT3 #(
		.INIT('h80)
	) name10362 (
		_w16081_,
		_w16082_,
		_w16084_,
		_w16189_
	);
	LUT4 #(
		.INIT('h0020)
	) name10363 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16190_
	);
	LUT4 #(
		.INIT('h77df)
	) name10364 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16191_
	);
	LUT4 #(
		.INIT('h0d00)
	) name10365 (
		_w16086_,
		_w16187_,
		_w16188_,
		_w16191_,
		_w16192_
	);
	LUT4 #(
		.INIT('hbebc)
	) name10366 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16193_
	);
	LUT3 #(
		.INIT('h6f)
	) name10367 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16194_
	);
	LUT4 #(
		.INIT('hdbff)
	) name10368 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16195_
	);
	LUT4 #(
		.INIT('he400)
	) name10369 (
		_w16086_,
		_w16193_,
		_w16194_,
		_w16195_,
		_w16196_
	);
	LUT4 #(
		.INIT('hfd00)
	) name10370 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16197_
	);
	LUT4 #(
		.INIT('h00f7)
	) name10371 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16198_
	);
	LUT3 #(
		.INIT('h02)
	) name10372 (
		_w16086_,
		_w16198_,
		_w16197_,
		_w16199_
	);
	LUT4 #(
		.INIT('h0e04)
	) name10373 (
		_w16080_,
		_w16196_,
		_w16199_,
		_w16192_,
		_w16200_
	);
	LUT2 #(
		.INIT('h9)
	) name10374 (
		\u1_L12_reg[17]/NET0131 ,
		_w16200_,
		_w16201_
	);
	LUT4 #(
		.INIT('h0800)
	) name10375 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16202_
	);
	LUT3 #(
		.INIT('h41)
	) name10376 (
		_w16051_,
		_w16054_,
		_w16055_,
		_w16203_
	);
	LUT4 #(
		.INIT('hbbe6)
	) name10377 (
		_w16051_,
		_w16054_,
		_w16052_,
		_w16055_,
		_w16204_
	);
	LUT2 #(
		.INIT('h4)
	) name10378 (
		_w16202_,
		_w16204_,
		_w16205_
	);
	LUT3 #(
		.INIT('h40)
	) name10379 (
		_w16051_,
		_w16052_,
		_w16053_,
		_w16206_
	);
	LUT4 #(
		.INIT('h2000)
	) name10380 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16207_
	);
	LUT4 #(
		.INIT('hfeeb)
	) name10381 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16208_
	);
	LUT4 #(
		.INIT('h0100)
	) name10382 (
		_w16050_,
		_w16207_,
		_w16206_,
		_w16208_,
		_w16209_
	);
	LUT4 #(
		.INIT('h0420)
	) name10383 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16210_
	);
	LUT4 #(
		.INIT('h0004)
	) name10384 (
		_w16073_,
		_w16050_,
		_w16059_,
		_w16210_,
		_w16211_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name10385 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16212_
	);
	LUT3 #(
		.INIT('hb1)
	) name10386 (
		_w16051_,
		_w16061_,
		_w16212_,
		_w16213_
	);
	LUT4 #(
		.INIT('h0777)
	) name10387 (
		_w16205_,
		_w16209_,
		_w16211_,
		_w16213_,
		_w16214_
	);
	LUT2 #(
		.INIT('h6)
	) name10388 (
		\u1_L12_reg[12]/NET0131 ,
		_w16214_,
		_w16215_
	);
	LUT4 #(
		.INIT('hc963)
	) name10389 (
		decrypt_pad,
		\u1_R12_reg[28]/NET0131 ,
		\u1_uk_K_r12_reg[37]/NET0131 ,
		\u1_uk_K_r12_reg[43]/NET0131 ,
		_w16216_
	);
	LUT4 #(
		.INIT('hc693)
	) name10390 (
		decrypt_pad,
		\u1_R12_reg[29]/NET0131 ,
		\u1_uk_K_r12_reg[15]/NET0131 ,
		\u1_uk_K_r12_reg[9]/NET0131 ,
		_w16217_
	);
	LUT2 #(
		.INIT('h2)
	) name10391 (
		_w16216_,
		_w16217_,
		_w16218_
	);
	LUT4 #(
		.INIT('hc693)
	) name10392 (
		decrypt_pad,
		\u1_R12_reg[1]/NET0131 ,
		\u1_uk_K_r12_reg[0]/NET0131 ,
		\u1_uk_K_r12_reg[49]/NET0131 ,
		_w16219_
	);
	LUT4 #(
		.INIT('hc693)
	) name10393 (
		decrypt_pad,
		\u1_R12_reg[30]/NET0131 ,
		\u1_uk_K_r12_reg[16]/NET0131 ,
		\u1_uk_K_r12_reg[38]/NET0131 ,
		_w16220_
	);
	LUT3 #(
		.INIT('h01)
	) name10394 (
		_w16216_,
		_w16217_,
		_w16220_,
		_w16221_
	);
	LUT4 #(
		.INIT('h0001)
	) name10395 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16222_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name10396 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16223_
	);
	LUT2 #(
		.INIT('h8)
	) name10397 (
		_w16217_,
		_w16219_,
		_w16224_
	);
	LUT4 #(
		.INIT('h0040)
	) name10398 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16225_
	);
	LUT4 #(
		.INIT('hc963)
	) name10399 (
		decrypt_pad,
		\u1_R12_reg[31]/NET0131 ,
		\u1_uk_K_r12_reg[22]/NET0131 ,
		\u1_uk_K_r12_reg[28]/NET0131 ,
		_w16226_
	);
	LUT2 #(
		.INIT('h8)
	) name10400 (
		_w16216_,
		_w16220_,
		_w16227_
	);
	LUT4 #(
		.INIT('h00df)
	) name10401 (
		_w16216_,
		_w16217_,
		_w16220_,
		_w16226_,
		_w16228_
	);
	LUT3 #(
		.INIT('h40)
	) name10402 (
		_w16225_,
		_w16223_,
		_w16228_,
		_w16229_
	);
	LUT4 #(
		.INIT('h1000)
	) name10403 (
		_w16218_,
		_w16225_,
		_w16223_,
		_w16228_,
		_w16230_
	);
	LUT4 #(
		.INIT('h0010)
	) name10404 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16231_
	);
	LUT4 #(
		.INIT('h4000)
	) name10405 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16232_
	);
	LUT4 #(
		.INIT('h6763)
	) name10406 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16233_
	);
	LUT4 #(
		.INIT('h0200)
	) name10407 (
		_w16226_,
		_w16231_,
		_w16232_,
		_w16233_,
		_w16234_
	);
	LUT4 #(
		.INIT('hc963)
	) name10408 (
		decrypt_pad,
		\u1_R12_reg[32]/NET0131 ,
		\u1_uk_K_r12_reg[28]/NET0131 ,
		\u1_uk_K_r12_reg[38]/NET0131 ,
		_w16235_
	);
	LUT2 #(
		.INIT('h2)
	) name10409 (
		_w16216_,
		_w16220_,
		_w16236_
	);
	LUT4 #(
		.INIT('h0002)
	) name10410 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16237_
	);
	LUT2 #(
		.INIT('h1)
	) name10411 (
		_w16235_,
		_w16237_,
		_w16238_
	);
	LUT3 #(
		.INIT('he0)
	) name10412 (
		_w16230_,
		_w16234_,
		_w16238_,
		_w16239_
	);
	LUT3 #(
		.INIT('h01)
	) name10413 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16240_
	);
	LUT4 #(
		.INIT('h0002)
	) name10414 (
		_w16226_,
		_w16231_,
		_w16232_,
		_w16240_,
		_w16241_
	);
	LUT3 #(
		.INIT('h08)
	) name10415 (
		_w16216_,
		_w16217_,
		_w16220_,
		_w16242_
	);
	LUT2 #(
		.INIT('h2)
	) name10416 (
		_w16219_,
		_w16226_,
		_w16243_
	);
	LUT4 #(
		.INIT('h0040)
	) name10417 (
		_w16217_,
		_w16219_,
		_w16220_,
		_w16226_,
		_w16244_
	);
	LUT4 #(
		.INIT('hdbff)
	) name10418 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16245_
	);
	LUT4 #(
		.INIT('h0200)
	) name10419 (
		_w16235_,
		_w16244_,
		_w16242_,
		_w16245_,
		_w16246_
	);
	LUT3 #(
		.INIT('he0)
	) name10420 (
		_w16229_,
		_w16241_,
		_w16246_,
		_w16247_
	);
	LUT3 #(
		.INIT('ha9)
	) name10421 (
		\u1_L12_reg[15]/P0001 ,
		_w16239_,
		_w16247_,
		_w16248_
	);
	LUT3 #(
		.INIT('h08)
	) name10422 (
		_w16148_,
		_w16149_,
		_w16152_,
		_w16249_
	);
	LUT3 #(
		.INIT('hc6)
	) name10423 (
		_w16148_,
		_w16149_,
		_w16152_,
		_w16250_
	);
	LUT4 #(
		.INIT('h3391)
	) name10424 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16251_
	);
	LUT3 #(
		.INIT('h31)
	) name10425 (
		_w16149_,
		_w16150_,
		_w16152_,
		_w16252_
	);
	LUT3 #(
		.INIT('h01)
	) name10426 (
		_w16180_,
		_w16252_,
		_w16251_,
		_w16253_
	);
	LUT3 #(
		.INIT('hb0)
	) name10427 (
		_w16148_,
		_w16149_,
		_w16152_,
		_w16254_
	);
	LUT4 #(
		.INIT('h0a02)
	) name10428 (
		_w16155_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16255_
	);
	LUT3 #(
		.INIT('h45)
	) name10429 (
		_w16160_,
		_w16254_,
		_w16255_,
		_w16256_
	);
	LUT4 #(
		.INIT('h0800)
	) name10430 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16257_
	);
	LUT2 #(
		.INIT('h2)
	) name10431 (
		_w16160_,
		_w16257_,
		_w16258_
	);
	LUT3 #(
		.INIT('h31)
	) name10432 (
		_w16180_,
		_w16172_,
		_w16252_,
		_w16259_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name10433 (
		_w16253_,
		_w16256_,
		_w16258_,
		_w16259_,
		_w16260_
	);
	LUT4 #(
		.INIT('hdf5d)
	) name10434 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16261_
	);
	LUT4 #(
		.INIT('h0501)
	) name10435 (
		_w16155_,
		_w16160_,
		_w16257_,
		_w16261_,
		_w16262_
	);
	LUT4 #(
		.INIT('h9000)
	) name10436 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16263_
	);
	LUT3 #(
		.INIT('h02)
	) name10437 (
		_w16155_,
		_w16153_,
		_w16263_,
		_w16264_
	);
	LUT3 #(
		.INIT('h54)
	) name10438 (
		_w16173_,
		_w16262_,
		_w16264_,
		_w16265_
	);
	LUT3 #(
		.INIT('h65)
	) name10439 (
		\u1_L12_reg[1]/NET0131 ,
		_w16260_,
		_w16265_,
		_w16266_
	);
	LUT4 #(
		.INIT('h378f)
	) name10440 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16267_
	);
	LUT4 #(
		.INIT('hdff5)
	) name10441 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16268_
	);
	LUT4 #(
		.INIT('hf6ef)
	) name10442 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16269_
	);
	LUT4 #(
		.INIT('he400)
	) name10443 (
		_w16226_,
		_w16268_,
		_w16267_,
		_w16269_,
		_w16270_
	);
	LUT2 #(
		.INIT('h2)
	) name10444 (
		_w16235_,
		_w16270_,
		_w16271_
	);
	LUT4 #(
		.INIT('hd5f7)
	) name10445 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16272_
	);
	LUT2 #(
		.INIT('h2)
	) name10446 (
		_w16226_,
		_w16272_,
		_w16273_
	);
	LUT2 #(
		.INIT('h9)
	) name10447 (
		_w16216_,
		_w16220_,
		_w16274_
	);
	LUT4 #(
		.INIT('h3b0b)
	) name10448 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16226_,
		_w16275_
	);
	LUT2 #(
		.INIT('h1)
	) name10449 (
		_w16274_,
		_w16275_,
		_w16276_
	);
	LUT4 #(
		.INIT('h0200)
	) name10450 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16277_
	);
	LUT4 #(
		.INIT('h0004)
	) name10451 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16226_,
		_w16278_
	);
	LUT3 #(
		.INIT('h01)
	) name10452 (
		_w16222_,
		_w16277_,
		_w16278_,
		_w16279_
	);
	LUT4 #(
		.INIT('h5455)
	) name10453 (
		_w16235_,
		_w16276_,
		_w16273_,
		_w16279_,
		_w16280_
	);
	LUT4 #(
		.INIT('h0100)
	) name10454 (
		_w16216_,
		_w16217_,
		_w16220_,
		_w16226_,
		_w16281_
	);
	LUT3 #(
		.INIT('h07)
	) name10455 (
		_w16243_,
		_w16242_,
		_w16281_,
		_w16282_
	);
	LUT4 #(
		.INIT('h5655)
	) name10456 (
		\u1_L12_reg[21]/NET0131 ,
		_w16280_,
		_w16271_,
		_w16282_,
		_w16283_
	);
	LUT3 #(
		.INIT('hb1)
	) name10457 (
		_w16148_,
		_w16155_,
		_w16152_,
		_w16284_
	);
	LUT4 #(
		.INIT('h0c04)
	) name10458 (
		_w16151_,
		_w16160_,
		_w16257_,
		_w16284_,
		_w16285_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name10459 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16150_,
		_w16286_
	);
	LUT4 #(
		.INIT('h3f2f)
	) name10460 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16287_
	);
	LUT3 #(
		.INIT('h51)
	) name10461 (
		_w16155_,
		_w16149_,
		_w16152_,
		_w16288_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name10462 (
		_w16152_,
		_w16286_,
		_w16287_,
		_w16288_,
		_w16289_
	);
	LUT2 #(
		.INIT('h8)
	) name10463 (
		_w16285_,
		_w16289_,
		_w16290_
	);
	LUT3 #(
		.INIT('h0b)
	) name10464 (
		_w16167_,
		_w16156_,
		_w16160_,
		_w16291_
	);
	LUT4 #(
		.INIT('h0100)
	) name10465 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16152_,
		_w16292_
	);
	LUT4 #(
		.INIT('hfa32)
	) name10466 (
		_w16155_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16293_
	);
	LUT3 #(
		.INIT('h32)
	) name10467 (
		_w16148_,
		_w16292_,
		_w16293_,
		_w16294_
	);
	LUT3 #(
		.INIT('h80)
	) name10468 (
		_w16170_,
		_w16291_,
		_w16294_,
		_w16295_
	);
	LUT4 #(
		.INIT('h8421)
	) name10469 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16150_,
		_w16296_
	);
	LUT4 #(
		.INIT('h13cc)
	) name10470 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16150_,
		_w16297_
	);
	LUT3 #(
		.INIT('h01)
	) name10471 (
		_w16152_,
		_w16297_,
		_w16296_,
		_w16298_
	);
	LUT4 #(
		.INIT('h55a9)
	) name10472 (
		\u1_L12_reg[26]/NET0131 ,
		_w16290_,
		_w16295_,
		_w16298_,
		_w16299_
	);
	LUT4 #(
		.INIT('h3fc6)
	) name10473 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16300_
	);
	LUT2 #(
		.INIT('h2)
	) name10474 (
		_w16115_,
		_w16300_,
		_w16301_
	);
	LUT4 #(
		.INIT('h0484)
	) name10475 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16302_
	);
	LUT4 #(
		.INIT('h0200)
	) name10476 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16303_
	);
	LUT4 #(
		.INIT('h0023)
	) name10477 (
		_w16115_,
		_w16125_,
		_w16302_,
		_w16303_,
		_w16304_
	);
	LUT3 #(
		.INIT('h45)
	) name10478 (
		_w16114_,
		_w16301_,
		_w16304_,
		_w16305_
	);
	LUT4 #(
		.INIT('hf37b)
	) name10479 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16306_
	);
	LUT2 #(
		.INIT('h2)
	) name10480 (
		_w16115_,
		_w16306_,
		_w16307_
	);
	LUT4 #(
		.INIT('h5ff4)
	) name10481 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16308_
	);
	LUT2 #(
		.INIT('h1)
	) name10482 (
		_w16115_,
		_w16308_,
		_w16309_
	);
	LUT4 #(
		.INIT('h0002)
	) name10483 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16310_
	);
	LUT4 #(
		.INIT('h0100)
	) name10484 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16311_
	);
	LUT4 #(
		.INIT('h0001)
	) name10485 (
		_w16132_,
		_w16133_,
		_w16311_,
		_w16310_,
		_w16312_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10486 (
		_w16114_,
		_w16309_,
		_w16307_,
		_w16312_,
		_w16313_
	);
	LUT4 #(
		.INIT('h4000)
	) name10487 (
		_w16119_,
		_w16116_,
		_w16115_,
		_w16118_,
		_w16314_
	);
	LUT2 #(
		.INIT('h1)
	) name10488 (
		_w16121_,
		_w16314_,
		_w16315_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name10489 (
		\u1_L12_reg[29]/NET0131 ,
		_w16313_,
		_w16305_,
		_w16315_,
		_w16316_
	);
	LUT4 #(
		.INIT('hc693)
	) name10490 (
		decrypt_pad,
		\u1_R12_reg[4]/NET0131 ,
		\u1_uk_K_r12_reg[24]/NET0131 ,
		\u1_uk_K_r12_reg[48]/NET0131 ,
		_w16317_
	);
	LUT4 #(
		.INIT('hc963)
	) name10491 (
		decrypt_pad,
		\u1_R12_reg[9]/NET0131 ,
		\u1_uk_K_r12_reg[40]/NET0131 ,
		\u1_uk_K_r12_reg[48]/NET0131 ,
		_w16318_
	);
	LUT4 #(
		.INIT('hc963)
	) name10492 (
		decrypt_pad,
		\u1_R12_reg[5]/NET0131 ,
		\u1_uk_K_r12_reg[27]/NET0131 ,
		\u1_uk_K_r12_reg[3]/NET0131 ,
		_w16319_
	);
	LUT3 #(
		.INIT('h59)
	) name10493 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16320_
	);
	LUT4 #(
		.INIT('hc963)
	) name10494 (
		decrypt_pad,
		\u1_R12_reg[6]/NET0131 ,
		\u1_uk_K_r12_reg[18]/NET0131 ,
		\u1_uk_K_r12_reg[26]/NET0131 ,
		_w16321_
	);
	LUT4 #(
		.INIT('hc963)
	) name10495 (
		decrypt_pad,
		\u1_R12_reg[7]/NET0131 ,
		\u1_uk_K_r12_reg[12]/NET0131 ,
		\u1_uk_K_r12_reg[20]/NET0131 ,
		_w16322_
	);
	LUT2 #(
		.INIT('h2)
	) name10496 (
		_w16321_,
		_w16322_,
		_w16323_
	);
	LUT2 #(
		.INIT('h4)
	) name10497 (
		_w16320_,
		_w16323_,
		_w16324_
	);
	LUT4 #(
		.INIT('h0034)
	) name10498 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16325_
	);
	LUT4 #(
		.INIT('hc693)
	) name10499 (
		decrypt_pad,
		\u1_R12_reg[8]/NET0131 ,
		\u1_uk_K_r12_reg[11]/NET0131 ,
		\u1_uk_K_r12_reg[3]/NET0131 ,
		_w16326_
	);
	LUT2 #(
		.INIT('h1)
	) name10500 (
		_w16325_,
		_w16326_,
		_w16327_
	);
	LUT4 #(
		.INIT('h0800)
	) name10501 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16328_
	);
	LUT2 #(
		.INIT('h8)
	) name10502 (
		_w16322_,
		_w16328_,
		_w16329_
	);
	LUT3 #(
		.INIT('h8c)
	) name10503 (
		_w16317_,
		_w16319_,
		_w16321_,
		_w16330_
	);
	LUT3 #(
		.INIT('hb0)
	) name10504 (
		_w16317_,
		_w16321_,
		_w16322_,
		_w16331_
	);
	LUT3 #(
		.INIT('h8a)
	) name10505 (
		_w16318_,
		_w16319_,
		_w16321_,
		_w16332_
	);
	LUT3 #(
		.INIT('h10)
	) name10506 (
		_w16331_,
		_w16330_,
		_w16332_,
		_w16333_
	);
	LUT4 #(
		.INIT('h0100)
	) name10507 (
		_w16324_,
		_w16329_,
		_w16333_,
		_w16327_,
		_w16334_
	);
	LUT4 #(
		.INIT('h0082)
	) name10508 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16335_
	);
	LUT4 #(
		.INIT('h8c00)
	) name10509 (
		_w16317_,
		_w16319_,
		_w16321_,
		_w16322_,
		_w16336_
	);
	LUT3 #(
		.INIT('h02)
	) name10510 (
		_w16326_,
		_w16336_,
		_w16335_,
		_w16337_
	);
	LUT2 #(
		.INIT('h2)
	) name10511 (
		_w16319_,
		_w16321_,
		_w16338_
	);
	LUT4 #(
		.INIT('he6ee)
	) name10512 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16339_
	);
	LUT4 #(
		.INIT('h4044)
	) name10513 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16340_
	);
	LUT4 #(
		.INIT('h3302)
	) name10514 (
		_w16326_,
		_w16338_,
		_w16339_,
		_w16340_,
		_w16341_
	);
	LUT4 #(
		.INIT('h0100)
	) name10515 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16342_
	);
	LUT2 #(
		.INIT('h2)
	) name10516 (
		_w16317_,
		_w16321_,
		_w16343_
	);
	LUT4 #(
		.INIT('hf700)
	) name10517 (
		_w16317_,
		_w16319_,
		_w16321_,
		_w16322_,
		_w16344_
	);
	LUT2 #(
		.INIT('h4)
	) name10518 (
		_w16342_,
		_w16344_,
		_w16345_
	);
	LUT3 #(
		.INIT('h0e)
	) name10519 (
		_w16322_,
		_w16341_,
		_w16345_,
		_w16346_
	);
	LUT4 #(
		.INIT('h55a9)
	) name10520 (
		\u1_L12_reg[2]/NET0131 ,
		_w16334_,
		_w16337_,
		_w16346_,
		_w16347_
	);
	LUT4 #(
		.INIT('hbfae)
	) name10521 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16348_
	);
	LUT4 #(
		.INIT('h2000)
	) name10522 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16349_
	);
	LUT4 #(
		.INIT('h00ef)
	) name10523 (
		_w16317_,
		_w16319_,
		_w16321_,
		_w16322_,
		_w16350_
	);
	LUT3 #(
		.INIT('h20)
	) name10524 (
		_w16348_,
		_w16349_,
		_w16350_,
		_w16351_
	);
	LUT3 #(
		.INIT('h10)
	) name10525 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16352_
	);
	LUT4 #(
		.INIT('h1000)
	) name10526 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16353_
	);
	LUT4 #(
		.INIT('h7d00)
	) name10527 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16322_,
		_w16354_
	);
	LUT2 #(
		.INIT('h4)
	) name10528 (
		_w16353_,
		_w16354_,
		_w16355_
	);
	LUT4 #(
		.INIT('h00f7)
	) name10529 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16322_,
		_w16356_
	);
	LUT4 #(
		.INIT('h0400)
	) name10530 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16357_
	);
	LUT4 #(
		.INIT('h00a2)
	) name10531 (
		_w16326_,
		_w16343_,
		_w16356_,
		_w16357_,
		_w16358_
	);
	LUT3 #(
		.INIT('he0)
	) name10532 (
		_w16351_,
		_w16355_,
		_w16358_,
		_w16359_
	);
	LUT2 #(
		.INIT('h8)
	) name10533 (
		_w16322_,
		_w16348_,
		_w16360_
	);
	LUT4 #(
		.INIT('h5b59)
	) name10534 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16361_
	);
	LUT3 #(
		.INIT('h40)
	) name10535 (
		_w16349_,
		_w16350_,
		_w16361_,
		_w16362_
	);
	LUT4 #(
		.INIT('h2900)
	) name10536 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16363_
	);
	LUT2 #(
		.INIT('h1)
	) name10537 (
		_w16326_,
		_w16363_,
		_w16364_
	);
	LUT3 #(
		.INIT('he0)
	) name10538 (
		_w16360_,
		_w16362_,
		_w16364_,
		_w16365_
	);
	LUT3 #(
		.INIT('ha9)
	) name10539 (
		\u1_L12_reg[28]/NET0131 ,
		_w16359_,
		_w16365_,
		_w16366_
	);
	LUT4 #(
		.INIT('h2777)
	) name10540 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16115_,
		_w16367_
	);
	LUT2 #(
		.INIT('h2)
	) name10541 (
		_w16118_,
		_w16367_,
		_w16368_
	);
	LUT4 #(
		.INIT('hfaba)
	) name10542 (
		_w16119_,
		_w16116_,
		_w16115_,
		_w16118_,
		_w16369_
	);
	LUT4 #(
		.INIT('h0004)
	) name10543 (
		_w16119_,
		_w16116_,
		_w16115_,
		_w16118_,
		_w16370_
	);
	LUT4 #(
		.INIT('h0c08)
	) name10544 (
		_w16117_,
		_w16114_,
		_w16370_,
		_w16369_,
		_w16371_
	);
	LUT2 #(
		.INIT('h4)
	) name10545 (
		_w16368_,
		_w16371_,
		_w16372_
	);
	LUT4 #(
		.INIT('hf070)
	) name10546 (
		_w16116_,
		_w16117_,
		_w16115_,
		_w16118_,
		_w16373_
	);
	LUT4 #(
		.INIT('h2500)
	) name10547 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16374_
	);
	LUT2 #(
		.INIT('h2)
	) name10548 (
		_w16373_,
		_w16374_,
		_w16375_
	);
	LUT3 #(
		.INIT('h02)
	) name10549 (
		_w16116_,
		_w16117_,
		_w16118_,
		_w16376_
	);
	LUT3 #(
		.INIT('h01)
	) name10550 (
		_w16115_,
		_w16303_,
		_w16376_,
		_w16377_
	);
	LUT3 #(
		.INIT('h01)
	) name10551 (
		_w16114_,
		_w16121_,
		_w16125_,
		_w16378_
	);
	LUT3 #(
		.INIT('he0)
	) name10552 (
		_w16375_,
		_w16377_,
		_w16378_,
		_w16379_
	);
	LUT4 #(
		.INIT('h0001)
	) name10553 (
		_w16119_,
		_w16117_,
		_w16115_,
		_w16118_,
		_w16380_
	);
	LUT4 #(
		.INIT('h070b)
	) name10554 (
		_w16116_,
		_w16117_,
		_w16115_,
		_w16118_,
		_w16381_
	);
	LUT4 #(
		.INIT('hd060)
	) name10555 (
		_w16116_,
		_w16117_,
		_w16115_,
		_w16118_,
		_w16382_
	);
	LUT4 #(
		.INIT('h3331)
	) name10556 (
		_w16119_,
		_w16380_,
		_w16382_,
		_w16381_,
		_w16383_
	);
	LUT4 #(
		.INIT('ha955)
	) name10557 (
		\u1_L12_reg[4]/NET0131 ,
		_w16372_,
		_w16379_,
		_w16383_,
		_w16384_
	);
	LUT3 #(
		.INIT('h14)
	) name10558 (
		_w16155_,
		_w16149_,
		_w16150_,
		_w16385_
	);
	LUT2 #(
		.INIT('h8)
	) name10559 (
		_w16250_,
		_w16385_,
		_w16386_
	);
	LUT4 #(
		.INIT('hfdbd)
	) name10560 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16387_
	);
	LUT3 #(
		.INIT('h31)
	) name10561 (
		_w16155_,
		_w16263_,
		_w16387_,
		_w16388_
	);
	LUT3 #(
		.INIT('h8a)
	) name10562 (
		_w16160_,
		_w16386_,
		_w16388_,
		_w16389_
	);
	LUT4 #(
		.INIT('h0040)
	) name10563 (
		_w16155_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16390_
	);
	LUT4 #(
		.INIT('h0001)
	) name10564 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16150_,
		_w16391_
	);
	LUT3 #(
		.INIT('h01)
	) name10565 (
		_w16249_,
		_w16391_,
		_w16390_,
		_w16392_
	);
	LUT3 #(
		.INIT('h40)
	) name10566 (
		_w16148_,
		_w16155_,
		_w16149_,
		_w16393_
	);
	LUT4 #(
		.INIT('h0020)
	) name10567 (
		_w16155_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16394_
	);
	LUT3 #(
		.INIT('h0b)
	) name10568 (
		_w16158_,
		_w16393_,
		_w16394_,
		_w16395_
	);
	LUT4 #(
		.INIT('h1333)
	) name10569 (
		_w16154_,
		_w16160_,
		_w16392_,
		_w16395_,
		_w16396_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name10570 (
		_w16148_,
		_w16149_,
		_w16150_,
		_w16152_,
		_w16397_
	);
	LUT2 #(
		.INIT('h1)
	) name10571 (
		_w16155_,
		_w16397_,
		_w16398_
	);
	LUT3 #(
		.INIT('h0b)
	) name10572 (
		_w16152_,
		_w16166_,
		_w16157_,
		_w16399_
	);
	LUT2 #(
		.INIT('h4)
	) name10573 (
		_w16398_,
		_w16399_,
		_w16400_
	);
	LUT4 #(
		.INIT('h5655)
	) name10574 (
		\u1_L12_reg[10]/NET0131 ,
		_w16396_,
		_w16389_,
		_w16400_,
		_w16401_
	);
	LUT4 #(
		.INIT('hc963)
	) name10575 (
		decrypt_pad,
		\u1_R12_reg[21]/NET0131 ,
		\u1_uk_K_r12_reg[14]/NET0131 ,
		\u1_uk_K_r12_reg[51]/NET0131 ,
		_w16402_
	);
	LUT4 #(
		.INIT('hc963)
	) name10576 (
		decrypt_pad,
		\u1_R12_reg[18]/NET0131 ,
		\u1_uk_K_r12_reg[42]/NET0131 ,
		\u1_uk_K_r12_reg[52]/NET0131 ,
		_w16403_
	);
	LUT4 #(
		.INIT('hc963)
	) name10577 (
		decrypt_pad,
		\u1_R12_reg[16]/NET0131 ,
		\u1_uk_K_r12_reg[2]/NET0131 ,
		\u1_uk_K_r12_reg[8]/NET0131 ,
		_w16404_
	);
	LUT4 #(
		.INIT('hc693)
	) name10578 (
		decrypt_pad,
		\u1_R12_reg[17]/NET0131 ,
		\u1_uk_K_r12_reg[30]/NET0131 ,
		\u1_uk_K_r12_reg[52]/NET0131 ,
		_w16405_
	);
	LUT4 #(
		.INIT('h0180)
	) name10579 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16406_
	);
	LUT3 #(
		.INIT('h02)
	) name10580 (
		_w16402_,
		_w16404_,
		_w16405_,
		_w16407_
	);
	LUT4 #(
		.INIT('hc963)
	) name10581 (
		decrypt_pad,
		\u1_R12_reg[19]/NET0131 ,
		\u1_uk_K_r12_reg[29]/NET0131 ,
		\u1_uk_K_r12_reg[35]/NET0131 ,
		_w16408_
	);
	LUT4 #(
		.INIT('h00bf)
	) name10582 (
		_w16402_,
		_w16403_,
		_w16405_,
		_w16408_,
		_w16409_
	);
	LUT4 #(
		.INIT('h0010)
	) name10583 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16410_
	);
	LUT4 #(
		.INIT('h2000)
	) name10584 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16411_
	);
	LUT4 #(
		.INIT('hdfef)
	) name10585 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16412_
	);
	LUT3 #(
		.INIT('h40)
	) name10586 (
		_w16407_,
		_w16409_,
		_w16412_,
		_w16413_
	);
	LUT4 #(
		.INIT('h7f00)
	) name10587 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16408_,
		_w16414_
	);
	LUT3 #(
		.INIT('h10)
	) name10588 (
		_w16403_,
		_w16404_,
		_w16405_,
		_w16415_
	);
	LUT4 #(
		.INIT('hfcfa)
	) name10589 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16416_
	);
	LUT2 #(
		.INIT('h8)
	) name10590 (
		_w16414_,
		_w16416_,
		_w16417_
	);
	LUT4 #(
		.INIT('hc963)
	) name10591 (
		decrypt_pad,
		\u1_R12_reg[20]/NET0131 ,
		\u1_uk_K_r12_reg[44]/P0001 ,
		\u1_uk_K_r12_reg[50]/NET0131 ,
		_w16418_
	);
	LUT4 #(
		.INIT('h00ab)
	) name10592 (
		_w16406_,
		_w16413_,
		_w16417_,
		_w16418_,
		_w16419_
	);
	LUT4 #(
		.INIT('h87d5)
	) name10593 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16420_
	);
	LUT2 #(
		.INIT('h2)
	) name10594 (
		_w16408_,
		_w16420_,
		_w16421_
	);
	LUT3 #(
		.INIT('h7c)
	) name10595 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16422_
	);
	LUT3 #(
		.INIT('h09)
	) name10596 (
		_w16402_,
		_w16405_,
		_w16408_,
		_w16423_
	);
	LUT4 #(
		.INIT('h0040)
	) name10597 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16424_
	);
	LUT4 #(
		.INIT('hef9f)
	) name10598 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16425_
	);
	LUT3 #(
		.INIT('hb0)
	) name10599 (
		_w16422_,
		_w16423_,
		_w16425_,
		_w16426_
	);
	LUT4 #(
		.INIT('h0408)
	) name10600 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16427_
	);
	LUT4 #(
		.INIT('h1000)
	) name10601 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16428_
	);
	LUT4 #(
		.INIT('heffb)
	) name10602 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16429_
	);
	LUT3 #(
		.INIT('hb1)
	) name10603 (
		_w16408_,
		_w16427_,
		_w16429_,
		_w16430_
	);
	LUT4 #(
		.INIT('h7500)
	) name10604 (
		_w16418_,
		_w16421_,
		_w16426_,
		_w16430_,
		_w16431_
	);
	LUT3 #(
		.INIT('h65)
	) name10605 (
		\u1_L12_reg[14]/NET0131 ,
		_w16419_,
		_w16431_,
		_w16432_
	);
	LUT4 #(
		.INIT('h5be0)
	) name10606 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16433_
	);
	LUT3 #(
		.INIT('h08)
	) name10607 (
		_w16402_,
		_w16404_,
		_w16405_,
		_w16434_
	);
	LUT4 #(
		.INIT('hfc5f)
	) name10608 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16435_
	);
	LUT4 #(
		.INIT('h9dff)
	) name10609 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16436_
	);
	LUT4 #(
		.INIT('hd800)
	) name10610 (
		_w16408_,
		_w16433_,
		_w16435_,
		_w16436_,
		_w16437_
	);
	LUT3 #(
		.INIT('hd0)
	) name10611 (
		_w16403_,
		_w16404_,
		_w16405_,
		_w16438_
	);
	LUT4 #(
		.INIT('h5f0b)
	) name10612 (
		_w16402_,
		_w16404_,
		_w16405_,
		_w16408_,
		_w16439_
	);
	LUT3 #(
		.INIT('h0e)
	) name10613 (
		_w16404_,
		_w16405_,
		_w16408_,
		_w16440_
	);
	LUT4 #(
		.INIT('h1033)
	) name10614 (
		_w16402_,
		_w16403_,
		_w16405_,
		_w16408_,
		_w16441_
	);
	LUT4 #(
		.INIT('he0ee)
	) name10615 (
		_w16438_,
		_w16439_,
		_w16440_,
		_w16441_,
		_w16442_
	);
	LUT4 #(
		.INIT('hbffb)
	) name10616 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16443_
	);
	LUT4 #(
		.INIT('hbff9)
	) name10617 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16444_
	);
	LUT4 #(
		.INIT('h0008)
	) name10618 (
		_w16403_,
		_w16404_,
		_w16405_,
		_w16408_,
		_w16445_
	);
	LUT4 #(
		.INIT('h0301)
	) name10619 (
		_w16408_,
		_w16411_,
		_w16445_,
		_w16444_,
		_w16446_
	);
	LUT4 #(
		.INIT('he400)
	) name10620 (
		_w16418_,
		_w16442_,
		_w16437_,
		_w16446_,
		_w16447_
	);
	LUT2 #(
		.INIT('h9)
	) name10621 (
		\u1_L12_reg[25]/NET0131 ,
		_w16447_,
		_w16448_
	);
	LUT3 #(
		.INIT('h01)
	) name10622 (
		_w16322_,
		_w16357_,
		_w16352_,
		_w16449_
	);
	LUT4 #(
		.INIT('h0002)
	) name10623 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16450_
	);
	LUT4 #(
		.INIT('h0040)
	) name10624 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16451_
	);
	LUT3 #(
		.INIT('h01)
	) name10625 (
		_w16326_,
		_w16450_,
		_w16451_,
		_w16452_
	);
	LUT2 #(
		.INIT('h8)
	) name10626 (
		_w16449_,
		_w16452_,
		_w16453_
	);
	LUT3 #(
		.INIT('h10)
	) name10627 (
		_w16318_,
		_w16319_,
		_w16321_,
		_w16454_
	);
	LUT3 #(
		.INIT('h40)
	) name10628 (
		_w16317_,
		_w16318_,
		_w16321_,
		_w16455_
	);
	LUT4 #(
		.INIT('hfe00)
	) name10629 (
		_w16318_,
		_w16319_,
		_w16321_,
		_w16322_,
		_w16456_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name10630 (
		_w16356_,
		_w16454_,
		_w16455_,
		_w16456_,
		_w16457_
	);
	LUT4 #(
		.INIT('h0010)
	) name10631 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16458_
	);
	LUT2 #(
		.INIT('h2)
	) name10632 (
		_w16326_,
		_w16458_,
		_w16459_
	);
	LUT3 #(
		.INIT('h10)
	) name10633 (
		_w16333_,
		_w16457_,
		_w16459_,
		_w16460_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name10634 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16461_
	);
	LUT4 #(
		.INIT('h002d)
	) name10635 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16462_
	);
	LUT4 #(
		.INIT('h8b00)
	) name10636 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16463_
	);
	LUT4 #(
		.INIT('h0002)
	) name10637 (
		_w16322_,
		_w16326_,
		_w16451_,
		_w16463_,
		_w16464_
	);
	LUT2 #(
		.INIT('h4)
	) name10638 (
		_w16462_,
		_w16464_,
		_w16465_
	);
	LUT4 #(
		.INIT('h001f)
	) name10639 (
		_w16453_,
		_w16460_,
		_w16461_,
		_w16465_,
		_w16466_
	);
	LUT2 #(
		.INIT('h9)
	) name10640 (
		\u1_L12_reg[13]/NET0131 ,
		_w16466_,
		_w16467_
	);
	LUT4 #(
		.INIT('hbf00)
	) name10641 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16115_,
		_w16468_
	);
	LUT3 #(
		.INIT('h31)
	) name10642 (
		_w16116_,
		_w16117_,
		_w16118_,
		_w16469_
	);
	LUT2 #(
		.INIT('h2)
	) name10643 (
		_w16468_,
		_w16469_,
		_w16470_
	);
	LUT4 #(
		.INIT('h0201)
	) name10644 (
		_w16116_,
		_w16117_,
		_w16115_,
		_w16118_,
		_w16471_
	);
	LUT4 #(
		.INIT('h8000)
	) name10645 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16472_
	);
	LUT3 #(
		.INIT('h01)
	) name10646 (
		_w16114_,
		_w16472_,
		_w16471_,
		_w16473_
	);
	LUT4 #(
		.INIT('h0802)
	) name10647 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16474_
	);
	LUT4 #(
		.INIT('h4030)
	) name10648 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16115_,
		_w16475_
	);
	LUT4 #(
		.INIT('hfebb)
	) name10649 (
		_w16119_,
		_w16116_,
		_w16117_,
		_w16118_,
		_w16476_
	);
	LUT4 #(
		.INIT('h0400)
	) name10650 (
		_w16137_,
		_w16114_,
		_w16475_,
		_w16476_,
		_w16477_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name10651 (
		_w16470_,
		_w16473_,
		_w16474_,
		_w16477_,
		_w16478_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name10652 (
		_w16119_,
		_w16116_,
		_w16125_,
		_w16141_,
		_w16479_
	);
	LUT3 #(
		.INIT('h65)
	) name10653 (
		\u1_L12_reg[19]/NET0131 ,
		_w16478_,
		_w16479_,
		_w16480_
	);
	LUT4 #(
		.INIT('he9f9)
	) name10654 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16481_
	);
	LUT4 #(
		.INIT('hffdb)
	) name10655 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16482_
	);
	LUT4 #(
		.INIT('h0233)
	) name10656 (
		_w16080_,
		_w16086_,
		_w16481_,
		_w16482_,
		_w16483_
	);
	LUT3 #(
		.INIT('he0)
	) name10657 (
		_w16082_,
		_w16084_,
		_w16086_,
		_w16484_
	);
	LUT2 #(
		.INIT('h8)
	) name10658 (
		_w16091_,
		_w16484_,
		_w16485_
	);
	LUT4 #(
		.INIT('h002a)
	) name10659 (
		_w16080_,
		_w16096_,
		_w16109_,
		_w16186_,
		_w16486_
	);
	LUT4 #(
		.INIT('h2000)
	) name10660 (
		_w16082_,
		_w16083_,
		_w16084_,
		_w16086_,
		_w16487_
	);
	LUT4 #(
		.INIT('h0080)
	) name10661 (
		_w16082_,
		_w16083_,
		_w16084_,
		_w16086_,
		_w16488_
	);
	LUT3 #(
		.INIT('h01)
	) name10662 (
		_w16081_,
		_w16082_,
		_w16084_,
		_w16489_
	);
	LUT4 #(
		.INIT('h0001)
	) name10663 (
		_w16189_,
		_w16487_,
		_w16488_,
		_w16489_,
		_w16490_
	);
	LUT4 #(
		.INIT('h0200)
	) name10664 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16086_,
		_w16491_
	);
	LUT4 #(
		.INIT('h5515)
	) name10665 (
		_w16080_,
		_w16081_,
		_w16083_,
		_w16086_,
		_w16492_
	);
	LUT2 #(
		.INIT('h4)
	) name10666 (
		_w16491_,
		_w16492_,
		_w16493_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name10667 (
		_w16485_,
		_w16486_,
		_w16490_,
		_w16493_,
		_w16494_
	);
	LUT2 #(
		.INIT('h8)
	) name10668 (
		_w16089_,
		_w16101_,
		_w16495_
	);
	LUT3 #(
		.INIT('h07)
	) name10669 (
		_w16093_,
		_w16106_,
		_w16110_,
		_w16496_
	);
	LUT2 #(
		.INIT('h4)
	) name10670 (
		_w16495_,
		_w16496_,
		_w16497_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name10671 (
		\u1_L12_reg[23]/P0001 ,
		_w16494_,
		_w16483_,
		_w16497_,
		_w16498_
	);
	LUT4 #(
		.INIT('h8084)
	) name10672 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16499_
	);
	LUT4 #(
		.INIT('h00fe)
	) name10673 (
		_w16216_,
		_w16217_,
		_w16220_,
		_w16226_,
		_w16500_
	);
	LUT3 #(
		.INIT('hb7)
	) name10674 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16501_
	);
	LUT4 #(
		.INIT('he4f5)
	) name10675 (
		_w16226_,
		_w16221_,
		_w16499_,
		_w16501_,
		_w16502_
	);
	LUT4 #(
		.INIT('hbdcf)
	) name10676 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16503_
	);
	LUT3 #(
		.INIT('h8a)
	) name10677 (
		_w16235_,
		_w16502_,
		_w16503_,
		_w16504_
	);
	LUT4 #(
		.INIT('hf430)
	) name10678 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16505_
	);
	LUT4 #(
		.INIT('hfd00)
	) name10679 (
		_w16217_,
		_w16219_,
		_w16220_,
		_w16226_,
		_w16506_
	);
	LUT2 #(
		.INIT('h4)
	) name10680 (
		_w16505_,
		_w16506_,
		_w16507_
	);
	LUT4 #(
		.INIT('h1000)
	) name10681 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16508_
	);
	LUT4 #(
		.INIT('h0080)
	) name10682 (
		_w16216_,
		_w16219_,
		_w16220_,
		_w16226_,
		_w16509_
	);
	LUT3 #(
		.INIT('h01)
	) name10683 (
		_w16278_,
		_w16508_,
		_w16509_,
		_w16510_
	);
	LUT4 #(
		.INIT('h1000)
	) name10684 (
		_w16217_,
		_w16219_,
		_w16220_,
		_w16226_,
		_w16511_
	);
	LUT4 #(
		.INIT('h0008)
	) name10685 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16512_
	);
	LUT4 #(
		.INIT('h0ac6)
	) name10686 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16513_
	);
	LUT4 #(
		.INIT('hf351)
	) name10687 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w16514_
	);
	LUT4 #(
		.INIT('h3332)
	) name10688 (
		_w16226_,
		_w16511_,
		_w16513_,
		_w16514_,
		_w16515_
	);
	LUT4 #(
		.INIT('hba00)
	) name10689 (
		_w16235_,
		_w16507_,
		_w16510_,
		_w16515_,
		_w16516_
	);
	LUT3 #(
		.INIT('h65)
	) name10690 (
		\u1_L12_reg[27]/NET0131 ,
		_w16504_,
		_w16516_,
		_w16517_
	);
	LUT3 #(
		.INIT('h40)
	) name10691 (
		_w16052_,
		_w16055_,
		_w16053_,
		_w16518_
	);
	LUT4 #(
		.INIT('h4555)
	) name10692 (
		_w16051_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16519_
	);
	LUT4 #(
		.INIT('hddd8)
	) name10693 (
		_w16051_,
		_w16061_,
		_w16056_,
		_w16518_,
		_w16520_
	);
	LUT4 #(
		.INIT('h1016)
	) name10694 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16521_
	);
	LUT3 #(
		.INIT('h01)
	) name10695 (
		_w16051_,
		_w16202_,
		_w16521_,
		_w16522_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10696 (
		_w16051_,
		_w16054_,
		_w16052_,
		_w16055_,
		_w16523_
	);
	LUT4 #(
		.INIT('hbb5f)
	) name10697 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16524_
	);
	LUT2 #(
		.INIT('h8)
	) name10698 (
		_w16523_,
		_w16524_,
		_w16525_
	);
	LUT4 #(
		.INIT('h4000)
	) name10699 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16526_
	);
	LUT2 #(
		.INIT('h2)
	) name10700 (
		_w16050_,
		_w16526_,
		_w16527_
	);
	LUT3 #(
		.INIT('he0)
	) name10701 (
		_w16522_,
		_w16525_,
		_w16527_,
		_w16528_
	);
	LUT4 #(
		.INIT('h0240)
	) name10702 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16529_
	);
	LUT4 #(
		.INIT('h9000)
	) name10703 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16530_
	);
	LUT3 #(
		.INIT('h01)
	) name10704 (
		_w16050_,
		_w16530_,
		_w16529_,
		_w16531_
	);
	LUT4 #(
		.INIT('h4457)
	) name10705 (
		_w16051_,
		_w16070_,
		_w16058_,
		_w16203_,
		_w16532_
	);
	LUT2 #(
		.INIT('h8)
	) name10706 (
		_w16531_,
		_w16532_,
		_w16533_
	);
	LUT4 #(
		.INIT('h6665)
	) name10707 (
		\u1_L12_reg[32]/NET0131 ,
		_w16520_,
		_w16528_,
		_w16533_,
		_w16534_
	);
	LUT4 #(
		.INIT('hc963)
	) name10708 (
		decrypt_pad,
		\u1_R12_reg[11]/NET0131 ,
		\u1_uk_K_r12_reg[55]/NET0131 ,
		\u1_uk_K_r12_reg[6]/NET0131 ,
		_w16535_
	);
	LUT4 #(
		.INIT('hc963)
	) name10709 (
		decrypt_pad,
		\u1_R12_reg[12]/NET0131 ,
		\u1_uk_K_r12_reg[13]/NET0131 ,
		\u1_uk_K_r12_reg[46]/NET0131 ,
		_w16536_
	);
	LUT4 #(
		.INIT('hc963)
	) name10710 (
		decrypt_pad,
		\u1_R12_reg[13]/NET0131 ,
		\u1_uk_K_r12_reg[26]/NET0131 ,
		\u1_uk_K_r12_reg[34]/NET0131 ,
		_w16537_
	);
	LUT4 #(
		.INIT('hc963)
	) name10711 (
		decrypt_pad,
		\u1_R12_reg[9]/NET0131 ,
		\u1_uk_K_r12_reg[46]/NET0131 ,
		\u1_uk_K_r12_reg[54]/NET0131 ,
		_w16538_
	);
	LUT4 #(
		.INIT('hc963)
	) name10712 (
		decrypt_pad,
		\u1_R12_reg[8]/NET0131 ,
		\u1_uk_K_r12_reg[17]/NET0131 ,
		\u1_uk_K_r12_reg[25]/NET0131 ,
		_w16539_
	);
	LUT2 #(
		.INIT('h1)
	) name10713 (
		_w16539_,
		_w16537_,
		_w16540_
	);
	LUT4 #(
		.INIT('hc963)
	) name10714 (
		decrypt_pad,
		\u1_R12_reg[10]/NET0131 ,
		\u1_uk_K_r12_reg[54]/NET0131 ,
		\u1_uk_K_r12_reg[5]/NET0131 ,
		_w16541_
	);
	LUT4 #(
		.INIT('h8acf)
	) name10715 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16542_
	);
	LUT4 #(
		.INIT('h93d3)
	) name10716 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16543_
	);
	LUT3 #(
		.INIT('hf2)
	) name10717 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16544_
	);
	LUT4 #(
		.INIT('h0c01)
	) name10718 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16545_
	);
	LUT4 #(
		.INIT('hcc08)
	) name10719 (
		_w16536_,
		_w16535_,
		_w16543_,
		_w16545_,
		_w16546_
	);
	LUT2 #(
		.INIT('h1)
	) name10720 (
		_w16538_,
		_w16541_,
		_w16547_
	);
	LUT2 #(
		.INIT('h8)
	) name10721 (
		_w16539_,
		_w16537_,
		_w16548_
	);
	LUT2 #(
		.INIT('h6)
	) name10722 (
		_w16539_,
		_w16537_,
		_w16549_
	);
	LUT4 #(
		.INIT('h0990)
	) name10723 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16550_
	);
	LUT2 #(
		.INIT('h4)
	) name10724 (
		_w16539_,
		_w16538_,
		_w16551_
	);
	LUT3 #(
		.INIT('h08)
	) name10725 (
		_w16537_,
		_w16541_,
		_w16535_,
		_w16552_
	);
	LUT3 #(
		.INIT('hc7)
	) name10726 (
		_w16537_,
		_w16541_,
		_w16535_,
		_w16553_
	);
	LUT2 #(
		.INIT('h2)
	) name10727 (
		_w16551_,
		_w16553_,
		_w16554_
	);
	LUT4 #(
		.INIT('h2000)
	) name10728 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16555_
	);
	LUT2 #(
		.INIT('h8)
	) name10729 (
		_w16537_,
		_w16535_,
		_w16556_
	);
	LUT4 #(
		.INIT('h0103)
	) name10730 (
		_w16537_,
		_w16538_,
		_w16541_,
		_w16535_,
		_w16557_
	);
	LUT3 #(
		.INIT('h15)
	) name10731 (
		_w16555_,
		_w16549_,
		_w16557_,
		_w16558_
	);
	LUT4 #(
		.INIT('h5455)
	) name10732 (
		_w16536_,
		_w16554_,
		_w16550_,
		_w16558_,
		_w16559_
	);
	LUT3 #(
		.INIT('h80)
	) name10733 (
		_w16538_,
		_w16541_,
		_w16536_,
		_w16560_
	);
	LUT2 #(
		.INIT('h8)
	) name10734 (
		_w16540_,
		_w16560_,
		_w16561_
	);
	LUT2 #(
		.INIT('h2)
	) name10735 (
		_w16536_,
		_w16535_,
		_w16562_
	);
	LUT3 #(
		.INIT('h80)
	) name10736 (
		_w16542_,
		_w16544_,
		_w16562_,
		_w16563_
	);
	LUT2 #(
		.INIT('h1)
	) name10737 (
		_w16561_,
		_w16563_,
		_w16564_
	);
	LUT4 #(
		.INIT('h5655)
	) name10738 (
		\u1_L12_reg[6]/NET0131 ,
		_w16559_,
		_w16546_,
		_w16564_,
		_w16565_
	);
	LUT3 #(
		.INIT('h60)
	) name10739 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16566_
	);
	LUT4 #(
		.INIT('h6000)
	) name10740 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16567_
	);
	LUT4 #(
		.INIT('h97ff)
	) name10741 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16568_
	);
	LUT4 #(
		.INIT('h0098)
	) name10742 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16569_
	);
	LUT2 #(
		.INIT('h2)
	) name10743 (
		_w16051_,
		_w16569_,
		_w16570_
	);
	LUT4 #(
		.INIT('hbbfc)
	) name10744 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16571_
	);
	LUT3 #(
		.INIT('h20)
	) name10745 (
		_w16519_,
		_w16566_,
		_w16571_,
		_w16572_
	);
	LUT4 #(
		.INIT('h222a)
	) name10746 (
		_w16050_,
		_w16568_,
		_w16570_,
		_w16572_,
		_w16573_
	);
	LUT4 #(
		.INIT('h0899)
	) name10747 (
		_w16054_,
		_w16052_,
		_w16055_,
		_w16053_,
		_w16574_
	);
	LUT4 #(
		.INIT('h3332)
	) name10748 (
		_w16050_,
		_w16065_,
		_w16567_,
		_w16574_,
		_w16575_
	);
	LUT4 #(
		.INIT('h3130)
	) name10749 (
		_w16051_,
		_w16050_,
		_w16065_,
		_w16569_,
		_w16576_
	);
	LUT4 #(
		.INIT('h00e4)
	) name10750 (
		_w16051_,
		_w16568_,
		_w16575_,
		_w16576_,
		_w16577_
	);
	LUT3 #(
		.INIT('h65)
	) name10751 (
		\u1_L12_reg[7]/NET0131 ,
		_w16573_,
		_w16577_,
		_w16578_
	);
	LUT4 #(
		.INIT('hf5fd)
	) name10752 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16579_
	);
	LUT4 #(
		.INIT('hb8bb)
	) name10753 (
		_w16410_,
		_w16408_,
		_w16434_,
		_w16579_,
		_w16580_
	);
	LUT4 #(
		.INIT('h8000)
	) name10754 (
		_w16402_,
		_w16404_,
		_w16405_,
		_w16408_,
		_w16581_
	);
	LUT3 #(
		.INIT('h04)
	) name10755 (
		_w16415_,
		_w16443_,
		_w16581_,
		_w16582_
	);
	LUT3 #(
		.INIT('h45)
	) name10756 (
		_w16418_,
		_w16580_,
		_w16582_,
		_w16583_
	);
	LUT4 #(
		.INIT('hff5e)
	) name10757 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16584_
	);
	LUT4 #(
		.INIT('h0008)
	) name10758 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16585_
	);
	LUT4 #(
		.INIT('hb9f7)
	) name10759 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16586_
	);
	LUT4 #(
		.INIT('h08aa)
	) name10760 (
		_w16408_,
		_w16418_,
		_w16584_,
		_w16586_,
		_w16587_
	);
	LUT2 #(
		.INIT('h8)
	) name10761 (
		_w16418_,
		_w16427_,
		_w16588_
	);
	LUT3 #(
		.INIT('h40)
	) name10762 (
		_w16403_,
		_w16404_,
		_w16418_,
		_w16589_
	);
	LUT3 #(
		.INIT('h54)
	) name10763 (
		_w16408_,
		_w16424_,
		_w16589_,
		_w16590_
	);
	LUT3 #(
		.INIT('h01)
	) name10764 (
		_w16587_,
		_w16588_,
		_w16590_,
		_w16591_
	);
	LUT3 #(
		.INIT('h65)
	) name10765 (
		\u1_L12_reg[8]/NET0131 ,
		_w16583_,
		_w16591_,
		_w16592_
	);
	LUT3 #(
		.INIT('h84)
	) name10766 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16593_
	);
	LUT4 #(
		.INIT('h0084)
	) name10767 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16535_,
		_w16594_
	);
	LUT3 #(
		.INIT('h01)
	) name10768 (
		_w16539_,
		_w16537_,
		_w16541_,
		_w16595_
	);
	LUT3 #(
		.INIT('h13)
	) name10769 (
		_w16538_,
		_w16536_,
		_w16535_,
		_w16596_
	);
	LUT3 #(
		.INIT('he0)
	) name10770 (
		_w16594_,
		_w16595_,
		_w16596_,
		_w16597_
	);
	LUT4 #(
		.INIT('h1000)
	) name10771 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16535_,
		_w16598_
	);
	LUT4 #(
		.INIT('h0222)
	) name10772 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16535_,
		_w16599_
	);
	LUT4 #(
		.INIT('h0001)
	) name10773 (
		_w16541_,
		_w16599_,
		_w16593_,
		_w16598_,
		_w16600_
	);
	LUT3 #(
		.INIT('h40)
	) name10774 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16601_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name10775 (
		_w16539_,
		_w16537_,
		_w16541_,
		_w16535_,
		_w16602_
	);
	LUT3 #(
		.INIT('h8a)
	) name10776 (
		_w16536_,
		_w16601_,
		_w16602_,
		_w16603_
	);
	LUT3 #(
		.INIT('h20)
	) name10777 (
		_w16539_,
		_w16538_,
		_w16541_,
		_w16604_
	);
	LUT4 #(
		.INIT('h0020)
	) name10778 (
		_w16539_,
		_w16538_,
		_w16541_,
		_w16535_,
		_w16605_
	);
	LUT4 #(
		.INIT('h00ec)
	) name10779 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16536_,
		_w16606_
	);
	LUT3 #(
		.INIT('h90)
	) name10780 (
		_w16539_,
		_w16538_,
		_w16541_,
		_w16607_
	);
	LUT4 #(
		.INIT('h7b00)
	) name10781 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16535_,
		_w16608_
	);
	LUT4 #(
		.INIT('h0155)
	) name10782 (
		_w16605_,
		_w16606_,
		_w16607_,
		_w16608_,
		_w16609_
	);
	LUT4 #(
		.INIT('h0b00)
	) name10783 (
		_w16600_,
		_w16603_,
		_w16597_,
		_w16609_,
		_w16610_
	);
	LUT2 #(
		.INIT('h9)
	) name10784 (
		\u1_L12_reg[16]/NET0131 ,
		_w16610_,
		_w16611_
	);
	LUT4 #(
		.INIT('h1bf4)
	) name10785 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16612_
	);
	LUT2 #(
		.INIT('h2)
	) name10786 (
		_w16535_,
		_w16612_,
		_w16613_
	);
	LUT4 #(
		.INIT('hfe3e)
	) name10787 (
		_w16535_,
		_w16547_,
		_w16549_,
		_w16556_,
		_w16614_
	);
	LUT3 #(
		.INIT('h8a)
	) name10788 (
		_w16536_,
		_w16613_,
		_w16614_,
		_w16615_
	);
	LUT4 #(
		.INIT('h0200)
	) name10789 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16616_
	);
	LUT3 #(
		.INIT('h14)
	) name10790 (
		_w16539_,
		_w16537_,
		_w16541_,
		_w16617_
	);
	LUT4 #(
		.INIT('h45cf)
	) name10791 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16618_
	);
	LUT4 #(
		.INIT('h448b)
	) name10792 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16619_
	);
	LUT3 #(
		.INIT('h70)
	) name10793 (
		_w16539_,
		_w16538_,
		_w16535_,
		_w16620_
	);
	LUT4 #(
		.INIT('h4544)
	) name10794 (
		_w16536_,
		_w16616_,
		_w16619_,
		_w16620_,
		_w16621_
	);
	LUT4 #(
		.INIT('h9bd6)
	) name10795 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16622_
	);
	LUT2 #(
		.INIT('h1)
	) name10796 (
		_w16536_,
		_w16535_,
		_w16623_
	);
	LUT2 #(
		.INIT('h4)
	) name10797 (
		_w16622_,
		_w16623_,
		_w16624_
	);
	LUT4 #(
		.INIT('h0600)
	) name10798 (
		_w16539_,
		_w16537_,
		_w16541_,
		_w16535_,
		_w16625_
	);
	LUT4 #(
		.INIT('h197f)
	) name10799 (
		_w16539_,
		_w16538_,
		_w16552_,
		_w16625_,
		_w16626_
	);
	LUT3 #(
		.INIT('h10)
	) name10800 (
		_w16621_,
		_w16624_,
		_w16626_,
		_w16627_
	);
	LUT3 #(
		.INIT('h65)
	) name10801 (
		\u1_L12_reg[24]/NET0131 ,
		_w16615_,
		_w16627_,
		_w16628_
	);
	LUT4 #(
		.INIT('h8a30)
	) name10802 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16629_
	);
	LUT2 #(
		.INIT('h1)
	) name10803 (
		_w16536_,
		_w16629_,
		_w16630_
	);
	LUT4 #(
		.INIT('h0002)
	) name10804 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16631_
	);
	LUT4 #(
		.INIT('hccc4)
	) name10805 (
		_w16536_,
		_w16535_,
		_w16617_,
		_w16631_,
		_w16632_
	);
	LUT2 #(
		.INIT('h4)
	) name10806 (
		_w16630_,
		_w16632_,
		_w16633_
	);
	LUT3 #(
		.INIT('h0e)
	) name10807 (
		_w16539_,
		_w16538_,
		_w16535_,
		_w16634_
	);
	LUT4 #(
		.INIT('hfbf6)
	) name10808 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16635_
	);
	LUT4 #(
		.INIT('h4055)
	) name10809 (
		_w16536_,
		_w16618_,
		_w16634_,
		_w16635_,
		_w16636_
	);
	LUT4 #(
		.INIT('h45ef)
	) name10810 (
		_w16539_,
		_w16537_,
		_w16538_,
		_w16541_,
		_w16637_
	);
	LUT2 #(
		.INIT('h2)
	) name10811 (
		_w16562_,
		_w16637_,
		_w16638_
	);
	LUT2 #(
		.INIT('h8)
	) name10812 (
		_w16556_,
		_w16604_,
		_w16639_
	);
	LUT4 #(
		.INIT('h0040)
	) name10813 (
		_w16537_,
		_w16538_,
		_w16541_,
		_w16535_,
		_w16640_
	);
	LUT3 #(
		.INIT('h0d)
	) name10814 (
		_w16560_,
		_w16548_,
		_w16640_,
		_w16641_
	);
	LUT4 #(
		.INIT('h0100)
	) name10815 (
		_w16636_,
		_w16638_,
		_w16639_,
		_w16641_,
		_w16642_
	);
	LUT3 #(
		.INIT('h9a)
	) name10816 (
		\u1_L12_reg[30]/NET0131 ,
		_w16633_,
		_w16642_,
		_w16643_
	);
	LUT4 #(
		.INIT('h99b9)
	) name10817 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16644_
	);
	LUT3 #(
		.INIT('he6)
	) name10818 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16645_
	);
	LUT4 #(
		.INIT('hbe7f)
	) name10819 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16646_
	);
	LUT4 #(
		.INIT('hd800)
	) name10820 (
		_w16086_,
		_w16644_,
		_w16645_,
		_w16646_,
		_w16647_
	);
	LUT4 #(
		.INIT('hf77f)
	) name10821 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16648_
	);
	LUT2 #(
		.INIT('h1)
	) name10822 (
		_w16086_,
		_w16648_,
		_w16649_
	);
	LUT4 #(
		.INIT('h9600)
	) name10823 (
		_w16081_,
		_w16082_,
		_w16083_,
		_w16084_,
		_w16650_
	);
	LUT4 #(
		.INIT('h0031)
	) name10824 (
		_w16101_,
		_w16190_,
		_w16645_,
		_w16650_,
		_w16651_
	);
	LUT4 #(
		.INIT('h0e04)
	) name10825 (
		_w16080_,
		_w16647_,
		_w16649_,
		_w16651_,
		_w16652_
	);
	LUT2 #(
		.INIT('h9)
	) name10826 (
		\u1_L12_reg[9]/NET0131 ,
		_w16652_,
		_w16653_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10827 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16654_
	);
	LUT3 #(
		.INIT('h02)
	) name10828 (
		_w16418_,
		_w16424_,
		_w16654_,
		_w16655_
	);
	LUT4 #(
		.INIT('h008c)
	) name10829 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16656_
	);
	LUT4 #(
		.INIT('h7252)
	) name10830 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16657_
	);
	LUT3 #(
		.INIT('h10)
	) name10831 (
		_w16418_,
		_w16656_,
		_w16657_,
		_w16658_
	);
	LUT4 #(
		.INIT('h0081)
	) name10832 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16659_
	);
	LUT3 #(
		.INIT('h01)
	) name10833 (
		_w16408_,
		_w16428_,
		_w16659_,
		_w16660_
	);
	LUT3 #(
		.INIT('he0)
	) name10834 (
		_w16655_,
		_w16658_,
		_w16660_,
		_w16661_
	);
	LUT4 #(
		.INIT('hdadf)
	) name10835 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16662_
	);
	LUT3 #(
		.INIT('h20)
	) name10836 (
		_w16418_,
		_w16424_,
		_w16662_,
		_w16663_
	);
	LUT4 #(
		.INIT('hadfd)
	) name10837 (
		_w16402_,
		_w16403_,
		_w16404_,
		_w16405_,
		_w16664_
	);
	LUT3 #(
		.INIT('h10)
	) name10838 (
		_w16418_,
		_w16656_,
		_w16664_,
		_w16665_
	);
	LUT3 #(
		.INIT('h04)
	) name10839 (
		_w16410_,
		_w16408_,
		_w16585_,
		_w16666_
	);
	LUT3 #(
		.INIT('he0)
	) name10840 (
		_w16663_,
		_w16665_,
		_w16666_,
		_w16667_
	);
	LUT3 #(
		.INIT('ha9)
	) name10841 (
		\u1_L12_reg[3]/NET0131 ,
		_w16661_,
		_w16667_,
		_w16668_
	);
	LUT4 #(
		.INIT('h3400)
	) name10842 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16322_,
		_w16669_
	);
	LUT4 #(
		.INIT('hfd75)
	) name10843 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16670_
	);
	LUT4 #(
		.INIT('h0032)
	) name10844 (
		_w16322_,
		_w16342_,
		_w16670_,
		_w16669_,
		_w16671_
	);
	LUT4 #(
		.INIT('hd7fc)
	) name10845 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16672_
	);
	LUT4 #(
		.INIT('h8000)
	) name10846 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16322_,
		_w16673_
	);
	LUT4 #(
		.INIT('h0141)
	) name10847 (
		_w16317_,
		_w16319_,
		_w16321_,
		_w16322_,
		_w16674_
	);
	LUT3 #(
		.INIT('h10)
	) name10848 (
		_w16673_,
		_w16674_,
		_w16672_,
		_w16675_
	);
	LUT4 #(
		.INIT('h0040)
	) name10849 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16322_,
		_w16676_
	);
	LUT4 #(
		.INIT('h77ef)
	) name10850 (
		_w16317_,
		_w16318_,
		_w16319_,
		_w16321_,
		_w16677_
	);
	LUT3 #(
		.INIT('h31)
	) name10851 (
		_w16322_,
		_w16676_,
		_w16677_,
		_w16678_
	);
	LUT4 #(
		.INIT('hd800)
	) name10852 (
		_w16326_,
		_w16671_,
		_w16675_,
		_w16678_,
		_w16679_
	);
	LUT2 #(
		.INIT('h9)
	) name10853 (
		\u1_L12_reg[18]/P0001 ,
		_w16679_,
		_w16680_
	);
	LUT4 #(
		.INIT('hc963)
	) name10854 (
		decrypt_pad,
		\u1_R11_reg[3]/NET0131 ,
		\u1_uk_K_r11_reg[13]/NET0131 ,
		\u1_uk_K_r11_reg[18]/NET0131 ,
		_w16681_
	);
	LUT4 #(
		.INIT('hc693)
	) name10855 (
		decrypt_pad,
		\u1_R11_reg[1]/NET0131 ,
		\u1_uk_K_r11_reg[26]/NET0131 ,
		\u1_uk_K_r11_reg[46]/NET0131 ,
		_w16682_
	);
	LUT4 #(
		.INIT('hc963)
	) name10856 (
		decrypt_pad,
		\u1_R11_reg[5]/NET0131 ,
		\u1_uk_K_r11_reg[19]/NET0131 ,
		\u1_uk_K_r11_reg[24]/NET0131 ,
		_w16683_
	);
	LUT4 #(
		.INIT('hc693)
	) name10857 (
		decrypt_pad,
		\u1_R11_reg[2]/NET0131 ,
		\u1_uk_K_r11_reg[41]/NET0131 ,
		\u1_uk_K_r11_reg[4]/NET0131 ,
		_w16684_
	);
	LUT4 #(
		.INIT('hc963)
	) name10858 (
		decrypt_pad,
		\u1_R11_reg[32]/NET0131 ,
		\u1_uk_K_r11_reg[25]/NET0131 ,
		\u1_uk_K_r11_reg[5]/NET0131 ,
		_w16685_
	);
	LUT4 #(
		.INIT('hafa3)
	) name10859 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w16686_
	);
	LUT2 #(
		.INIT('h2)
	) name10860 (
		_w16681_,
		_w16686_,
		_w16687_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name10861 (
		_w16681_,
		_w16682_,
		_w16684_,
		_w16683_,
		_w16688_
	);
	LUT2 #(
		.INIT('h4)
	) name10862 (
		_w16688_,
		_w16685_,
		_w16689_
	);
	LUT2 #(
		.INIT('h2)
	) name10863 (
		_w16681_,
		_w16684_,
		_w16690_
	);
	LUT3 #(
		.INIT('hc4)
	) name10864 (
		_w16681_,
		_w16682_,
		_w16684_,
		_w16691_
	);
	LUT3 #(
		.INIT('h0e)
	) name10865 (
		_w16684_,
		_w16683_,
		_w16685_,
		_w16692_
	);
	LUT4 #(
		.INIT('hc963)
	) name10866 (
		decrypt_pad,
		\u1_R11_reg[4]/NET0131 ,
		\u1_uk_K_r11_reg[48]/NET0131 ,
		\u1_uk_K_r11_reg[53]/P0001 ,
		_w16693_
	);
	LUT3 #(
		.INIT('hb0)
	) name10867 (
		_w16691_,
		_w16692_,
		_w16693_,
		_w16694_
	);
	LUT3 #(
		.INIT('h10)
	) name10868 (
		_w16689_,
		_w16687_,
		_w16694_,
		_w16695_
	);
	LUT2 #(
		.INIT('h2)
	) name10869 (
		_w16681_,
		_w16685_,
		_w16696_
	);
	LUT3 #(
		.INIT('h08)
	) name10870 (
		_w16681_,
		_w16684_,
		_w16685_,
		_w16697_
	);
	LUT4 #(
		.INIT('h0080)
	) name10871 (
		_w16681_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w16698_
	);
	LUT4 #(
		.INIT('hff7c)
	) name10872 (
		_w16681_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w16699_
	);
	LUT2 #(
		.INIT('h2)
	) name10873 (
		_w16682_,
		_w16699_,
		_w16700_
	);
	LUT3 #(
		.INIT('h45)
	) name10874 (
		_w16681_,
		_w16684_,
		_w16685_,
		_w16701_
	);
	LUT4 #(
		.INIT('h2723)
	) name10875 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w16702_
	);
	LUT2 #(
		.INIT('h8)
	) name10876 (
		_w16701_,
		_w16702_,
		_w16703_
	);
	LUT2 #(
		.INIT('h8)
	) name10877 (
		_w16681_,
		_w16685_,
		_w16704_
	);
	LUT3 #(
		.INIT('h08)
	) name10878 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16705_
	);
	LUT2 #(
		.INIT('h8)
	) name10879 (
		_w16704_,
		_w16705_,
		_w16706_
	);
	LUT2 #(
		.INIT('h8)
	) name10880 (
		_w16683_,
		_w16685_,
		_w16707_
	);
	LUT3 #(
		.INIT('h0b)
	) name10881 (
		_w16681_,
		_w16682_,
		_w16684_,
		_w16708_
	);
	LUT3 #(
		.INIT('h15)
	) name10882 (
		_w16693_,
		_w16707_,
		_w16708_,
		_w16709_
	);
	LUT4 #(
		.INIT('h0100)
	) name10883 (
		_w16700_,
		_w16703_,
		_w16706_,
		_w16709_,
		_w16710_
	);
	LUT2 #(
		.INIT('h1)
	) name10884 (
		_w16682_,
		_w16683_,
		_w16711_
	);
	LUT4 #(
		.INIT('h7dbd)
	) name10885 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w16712_
	);
	LUT2 #(
		.INIT('h1)
	) name10886 (
		_w16681_,
		_w16712_,
		_w16713_
	);
	LUT2 #(
		.INIT('h8)
	) name10887 (
		_w16697_,
		_w16711_,
		_w16714_
	);
	LUT4 #(
		.INIT('h0200)
	) name10888 (
		_w16681_,
		_w16682_,
		_w16684_,
		_w16685_,
		_w16715_
	);
	LUT3 #(
		.INIT('h07)
	) name10889 (
		_w16697_,
		_w16711_,
		_w16715_,
		_w16716_
	);
	LUT2 #(
		.INIT('h4)
	) name10890 (
		_w16713_,
		_w16716_,
		_w16717_
	);
	LUT4 #(
		.INIT('ha955)
	) name10891 (
		\u1_L11_reg[31]/NET0131 ,
		_w16695_,
		_w16710_,
		_w16717_,
		_w16718_
	);
	LUT4 #(
		.INIT('hc963)
	) name10892 (
		decrypt_pad,
		\u1_R11_reg[24]/NET0131 ,
		\u1_uk_K_r11_reg[15]/NET0131 ,
		\u1_uk_K_r11_reg[52]/NET0131 ,
		_w16719_
	);
	LUT4 #(
		.INIT('hc693)
	) name10893 (
		decrypt_pad,
		\u1_R11_reg[23]/NET0131 ,
		\u1_uk_K_r11_reg[22]/NET0131 ,
		\u1_uk_K_r11_reg[44]/NET0131 ,
		_w16720_
	);
	LUT4 #(
		.INIT('hc693)
	) name10894 (
		decrypt_pad,
		\u1_R11_reg[21]/NET0131 ,
		\u1_uk_K_r11_reg[42]/NET0131 ,
		\u1_uk_K_r11_reg[9]/NET0131 ,
		_w16721_
	);
	LUT4 #(
		.INIT('hc693)
	) name10895 (
		decrypt_pad,
		\u1_R11_reg[20]/NET0131 ,
		\u1_uk_K_r11_reg[31]/NET0131 ,
		\u1_uk_K_r11_reg[49]/NET0131 ,
		_w16722_
	);
	LUT4 #(
		.INIT('hc963)
	) name10896 (
		decrypt_pad,
		\u1_R11_reg[22]/NET0131 ,
		\u1_uk_K_r11_reg[0]/NET0131 ,
		\u1_uk_K_r11_reg[9]/NET0131 ,
		_w16723_
	);
	LUT4 #(
		.INIT('hc963)
	) name10897 (
		decrypt_pad,
		\u1_R11_reg[25]/NET0131 ,
		\u1_uk_K_r11_reg[38]/NET0131 ,
		\u1_uk_K_r11_reg[43]/NET0131 ,
		_w16724_
	);
	LUT3 #(
		.INIT('hc4)
	) name10898 (
		_w16721_,
		_w16722_,
		_w16724_,
		_w16725_
	);
	LUT4 #(
		.INIT('h57db)
	) name10899 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16726_
	);
	LUT2 #(
		.INIT('h2)
	) name10900 (
		_w16720_,
		_w16726_,
		_w16727_
	);
	LUT4 #(
		.INIT('he020)
	) name10901 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16728_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name10902 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16729_
	);
	LUT3 #(
		.INIT('h01)
	) name10903 (
		_w16720_,
		_w16729_,
		_w16728_,
		_w16730_
	);
	LUT2 #(
		.INIT('h1)
	) name10904 (
		_w16723_,
		_w16720_,
		_w16731_
	);
	LUT4 #(
		.INIT('h0200)
	) name10905 (
		_w16722_,
		_w16723_,
		_w16720_,
		_w16724_,
		_w16732_
	);
	LUT2 #(
		.INIT('h4)
	) name10906 (
		_w16721_,
		_w16732_,
		_w16733_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10907 (
		_w16719_,
		_w16730_,
		_w16727_,
		_w16733_,
		_w16734_
	);
	LUT4 #(
		.INIT('h0028)
	) name10908 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16720_,
		_w16735_
	);
	LUT4 #(
		.INIT('h1000)
	) name10909 (
		_w16721_,
		_w16722_,
		_w16720_,
		_w16724_,
		_w16736_
	);
	LUT4 #(
		.INIT('h0008)
	) name10910 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16737_
	);
	LUT3 #(
		.INIT('h10)
	) name10911 (
		_w16722_,
		_w16723_,
		_w16720_,
		_w16738_
	);
	LUT3 #(
		.INIT('h01)
	) name10912 (
		_w16737_,
		_w16738_,
		_w16736_,
		_w16739_
	);
	LUT4 #(
		.INIT('haf8c)
	) name10913 (
		_w16721_,
		_w16723_,
		_w16720_,
		_w16724_,
		_w16740_
	);
	LUT3 #(
		.INIT('h8a)
	) name10914 (
		_w16722_,
		_w16723_,
		_w16720_,
		_w16741_
	);
	LUT4 #(
		.INIT('h4000)
	) name10915 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16742_
	);
	LUT3 #(
		.INIT('h0b)
	) name10916 (
		_w16740_,
		_w16741_,
		_w16742_,
		_w16743_
	);
	LUT4 #(
		.INIT('h00bf)
	) name10917 (
		_w16735_,
		_w16739_,
		_w16743_,
		_w16719_,
		_w16744_
	);
	LUT4 #(
		.INIT('heff7)
	) name10918 (
		_w16721_,
		_w16722_,
		_w16720_,
		_w16724_,
		_w16745_
	);
	LUT2 #(
		.INIT('h1)
	) name10919 (
		_w16723_,
		_w16745_,
		_w16746_
	);
	LUT4 #(
		.INIT('h0002)
	) name10920 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16747_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name10921 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16748_
	);
	LUT4 #(
		.INIT('h0001)
	) name10922 (
		_w16722_,
		_w16723_,
		_w16720_,
		_w16724_,
		_w16749_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name10923 (
		_w16721_,
		_w16720_,
		_w16748_,
		_w16749_,
		_w16750_
	);
	LUT2 #(
		.INIT('h4)
	) name10924 (
		_w16746_,
		_w16750_,
		_w16751_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name10925 (
		\u1_L11_reg[11]/NET0131 ,
		_w16744_,
		_w16734_,
		_w16751_,
		_w16752_
	);
	LUT4 #(
		.INIT('hc963)
	) name10926 (
		decrypt_pad,
		\u1_R11_reg[27]/NET0131 ,
		\u1_uk_K_r11_reg[35]/NET0131 ,
		\u1_uk_K_r11_reg[44]/NET0131 ,
		_w16753_
	);
	LUT4 #(
		.INIT('hc693)
	) name10927 (
		decrypt_pad,
		\u1_R11_reg[24]/NET0131 ,
		\u1_uk_K_r11_reg[15]/NET0131 ,
		\u1_uk_K_r11_reg[37]/NET0131 ,
		_w16754_
	);
	LUT4 #(
		.INIT('hc963)
	) name10928 (
		decrypt_pad,
		\u1_R11_reg[25]/NET0131 ,
		\u1_uk_K_r11_reg[45]/NET0131 ,
		\u1_uk_K_r11_reg[50]/NET0131 ,
		_w16755_
	);
	LUT4 #(
		.INIT('hc963)
	) name10929 (
		decrypt_pad,
		\u1_R11_reg[26]/NET0131 ,
		\u1_uk_K_r11_reg[2]/NET0131 ,
		\u1_uk_K_r11_reg[35]/NET0131 ,
		_w16756_
	);
	LUT4 #(
		.INIT('hc963)
	) name10930 (
		decrypt_pad,
		\u1_R11_reg[29]/NET0131 ,
		\u1_uk_K_r11_reg[14]/NET0131 ,
		\u1_uk_K_r11_reg[23]/NET0131 ,
		_w16757_
	);
	LUT4 #(
		.INIT('h2000)
	) name10931 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16758_
	);
	LUT4 #(
		.INIT('hd7f7)
	) name10932 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16759_
	);
	LUT2 #(
		.INIT('h2)
	) name10933 (
		_w16753_,
		_w16759_,
		_w16760_
	);
	LUT2 #(
		.INIT('h6)
	) name10934 (
		_w16754_,
		_w16755_,
		_w16761_
	);
	LUT4 #(
		.INIT('h3100)
	) name10935 (
		_w16756_,
		_w16753_,
		_w16755_,
		_w16757_,
		_w16762_
	);
	LUT2 #(
		.INIT('h8)
	) name10936 (
		_w16761_,
		_w16762_,
		_w16763_
	);
	LUT4 #(
		.INIT('h0001)
	) name10937 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16764_
	);
	LUT2 #(
		.INIT('h4)
	) name10938 (
		_w16754_,
		_w16757_,
		_w16765_
	);
	LUT4 #(
		.INIT('h0400)
	) name10939 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16766_
	);
	LUT4 #(
		.INIT('hc693)
	) name10940 (
		decrypt_pad,
		\u1_R11_reg[28]/NET0131 ,
		\u1_uk_K_r11_reg[0]/NET0131 ,
		\u1_uk_K_r11_reg[22]/NET0131 ,
		_w16767_
	);
	LUT3 #(
		.INIT('h04)
	) name10941 (
		_w16766_,
		_w16767_,
		_w16764_,
		_w16768_
	);
	LUT3 #(
		.INIT('h10)
	) name10942 (
		_w16760_,
		_w16763_,
		_w16768_,
		_w16769_
	);
	LUT2 #(
		.INIT('h6)
	) name10943 (
		_w16754_,
		_w16756_,
		_w16770_
	);
	LUT3 #(
		.INIT('hd0)
	) name10944 (
		_w16753_,
		_w16755_,
		_w16757_,
		_w16771_
	);
	LUT3 #(
		.INIT('h23)
	) name10945 (
		_w16770_,
		_w16767_,
		_w16771_,
		_w16772_
	);
	LUT4 #(
		.INIT('h0004)
	) name10946 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16773_
	);
	LUT3 #(
		.INIT('hca)
	) name10947 (
		_w16756_,
		_w16753_,
		_w16755_,
		_w16774_
	);
	LUT3 #(
		.INIT('h8a)
	) name10948 (
		_w16754_,
		_w16753_,
		_w16757_,
		_w16775_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name10949 (
		_w16753_,
		_w16773_,
		_w16774_,
		_w16775_,
		_w16776_
	);
	LUT2 #(
		.INIT('h8)
	) name10950 (
		_w16772_,
		_w16776_,
		_w16777_
	);
	LUT4 #(
		.INIT('h0900)
	) name10951 (
		_w16754_,
		_w16756_,
		_w16753_,
		_w16755_,
		_w16778_
	);
	LUT4 #(
		.INIT('hfbbf)
	) name10952 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16779_
	);
	LUT4 #(
		.INIT('hfbb4)
	) name10953 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16780_
	);
	LUT3 #(
		.INIT('h31)
	) name10954 (
		_w16753_,
		_w16778_,
		_w16780_,
		_w16781_
	);
	LUT4 #(
		.INIT('ha955)
	) name10955 (
		\u1_L11_reg[22]/NET0131 ,
		_w16769_,
		_w16777_,
		_w16781_,
		_w16782_
	);
	LUT4 #(
		.INIT('hc693)
	) name10956 (
		decrypt_pad,
		\u1_R11_reg[13]/NET0131 ,
		\u1_uk_K_r11_reg[13]/NET0131 ,
		\u1_uk_K_r11_reg[33]/NET0131 ,
		_w16783_
	);
	LUT4 #(
		.INIT('hc693)
	) name10957 (
		decrypt_pad,
		\u1_R11_reg[12]/NET0131 ,
		\u1_uk_K_r11_reg[19]/NET0131 ,
		\u1_uk_K_r11_reg[39]/NET0131 ,
		_w16784_
	);
	LUT4 #(
		.INIT('hc693)
	) name10958 (
		decrypt_pad,
		\u1_R11_reg[17]/NET0131 ,
		\u1_uk_K_r11_reg[3]/NET0131 ,
		\u1_uk_K_r11_reg[55]/NET0131 ,
		_w16785_
	);
	LUT4 #(
		.INIT('hc963)
	) name10959 (
		decrypt_pad,
		\u1_R11_reg[15]/NET0131 ,
		\u1_uk_K_r11_reg[10]/NET0131 ,
		\u1_uk_K_r11_reg[47]/NET0131 ,
		_w16786_
	);
	LUT4 #(
		.INIT('h2aa8)
	) name10960 (
		_w16786_,
		_w16784_,
		_w16783_,
		_w16785_,
		_w16787_
	);
	LUT4 #(
		.INIT('hc963)
	) name10961 (
		decrypt_pad,
		\u1_R11_reg[14]/NET0131 ,
		\u1_uk_K_r11_reg[34]/NET0131 ,
		\u1_uk_K_r11_reg[39]/NET0131 ,
		_w16788_
	);
	LUT3 #(
		.INIT('h08)
	) name10962 (
		_w16784_,
		_w16788_,
		_w16785_,
		_w16789_
	);
	LUT3 #(
		.INIT('h45)
	) name10963 (
		_w16786_,
		_w16783_,
		_w16785_,
		_w16790_
	);
	LUT3 #(
		.INIT('h45)
	) name10964 (
		_w16787_,
		_w16789_,
		_w16790_,
		_w16791_
	);
	LUT3 #(
		.INIT('h01)
	) name10965 (
		_w16784_,
		_w16788_,
		_w16785_,
		_w16792_
	);
	LUT4 #(
		.INIT('h0001)
	) name10966 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w16793_
	);
	LUT3 #(
		.INIT('h04)
	) name10967 (
		_w16784_,
		_w16783_,
		_w16785_,
		_w16794_
	);
	LUT4 #(
		.INIT('hffbe)
	) name10968 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w16795_
	);
	LUT4 #(
		.INIT('h0200)
	) name10969 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w16796_
	);
	LUT4 #(
		.INIT('hc963)
	) name10970 (
		decrypt_pad,
		\u1_R11_reg[16]/NET0131 ,
		\u1_uk_K_r11_reg[18]/NET0131 ,
		\u1_uk_K_r11_reg[55]/NET0131 ,
		_w16797_
	);
	LUT3 #(
		.INIT('h80)
	) name10971 (
		_w16786_,
		_w16783_,
		_w16788_,
		_w16798_
	);
	LUT4 #(
		.INIT('h2000)
	) name10972 (
		_w16786_,
		_w16784_,
		_w16783_,
		_w16788_,
		_w16799_
	);
	LUT4 #(
		.INIT('h0002)
	) name10973 (
		_w16795_,
		_w16797_,
		_w16799_,
		_w16796_,
		_w16800_
	);
	LUT2 #(
		.INIT('h4)
	) name10974 (
		_w16791_,
		_w16800_,
		_w16801_
	);
	LUT4 #(
		.INIT('h0001)
	) name10975 (
		_w16786_,
		_w16784_,
		_w16783_,
		_w16785_,
		_w16802_
	);
	LUT4 #(
		.INIT('h3ffe)
	) name10976 (
		_w16786_,
		_w16784_,
		_w16783_,
		_w16785_,
		_w16803_
	);
	LUT2 #(
		.INIT('h2)
	) name10977 (
		_w16788_,
		_w16803_,
		_w16804_
	);
	LUT2 #(
		.INIT('h2)
	) name10978 (
		_w16784_,
		_w16783_,
		_w16805_
	);
	LUT4 #(
		.INIT('h0014)
	) name10979 (
		_w16786_,
		_w16784_,
		_w16783_,
		_w16788_,
		_w16806_
	);
	LUT2 #(
		.INIT('h2)
	) name10980 (
		_w16797_,
		_w16806_,
		_w16807_
	);
	LUT4 #(
		.INIT('h0400)
	) name10981 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w16808_
	);
	LUT4 #(
		.INIT('h0080)
	) name10982 (
		_w16786_,
		_w16784_,
		_w16783_,
		_w16785_,
		_w16809_
	);
	LUT2 #(
		.INIT('h4)
	) name10983 (
		_w16784_,
		_w16785_,
		_w16810_
	);
	LUT4 #(
		.INIT('h0200)
	) name10984 (
		_w16786_,
		_w16784_,
		_w16783_,
		_w16785_,
		_w16811_
	);
	LUT3 #(
		.INIT('h01)
	) name10985 (
		_w16808_,
		_w16809_,
		_w16811_,
		_w16812_
	);
	LUT3 #(
		.INIT('h40)
	) name10986 (
		_w16804_,
		_w16807_,
		_w16812_,
		_w16813_
	);
	LUT4 #(
		.INIT('h0020)
	) name10987 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w16814_
	);
	LUT4 #(
		.INIT('heee4)
	) name10988 (
		_w16786_,
		_w16808_,
		_w16793_,
		_w16814_,
		_w16815_
	);
	LUT2 #(
		.INIT('h4)
	) name10989 (
		_w16788_,
		_w16809_,
		_w16816_
	);
	LUT2 #(
		.INIT('h1)
	) name10990 (
		_w16815_,
		_w16816_,
		_w16817_
	);
	LUT4 #(
		.INIT('ha955)
	) name10991 (
		\u1_L11_reg[20]/NET0131 ,
		_w16801_,
		_w16813_,
		_w16817_,
		_w16818_
	);
	LUT4 #(
		.INIT('h779a)
	) name10992 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16819_
	);
	LUT4 #(
		.INIT('h0e02)
	) name10993 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16820_
	);
	LUT4 #(
		.INIT('hf17d)
	) name10994 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16821_
	);
	LUT4 #(
		.INIT('h1000)
	) name10995 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16822_
	);
	LUT4 #(
		.INIT('h00e4)
	) name10996 (
		_w16720_,
		_w16821_,
		_w16819_,
		_w16822_,
		_w16823_
	);
	LUT2 #(
		.INIT('h1)
	) name10997 (
		_w16719_,
		_w16823_,
		_w16824_
	);
	LUT4 #(
		.INIT('hdd7d)
	) name10998 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16825_
	);
	LUT2 #(
		.INIT('h2)
	) name10999 (
		_w16720_,
		_w16825_,
		_w16826_
	);
	LUT3 #(
		.INIT('h48)
	) name11000 (
		_w16722_,
		_w16723_,
		_w16724_,
		_w16827_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name11001 (
		_w16721_,
		_w16723_,
		_w16720_,
		_w16724_,
		_w16828_
	);
	LUT3 #(
		.INIT('h01)
	) name11002 (
		_w16820_,
		_w16828_,
		_w16827_,
		_w16829_
	);
	LUT4 #(
		.INIT('h0004)
	) name11003 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16830_
	);
	LUT4 #(
		.INIT('h2000)
	) name11004 (
		_w16721_,
		_w16723_,
		_w16720_,
		_w16724_,
		_w16831_
	);
	LUT2 #(
		.INIT('h1)
	) name11005 (
		_w16830_,
		_w16831_,
		_w16832_
	);
	LUT4 #(
		.INIT('h5700)
	) name11006 (
		_w16719_,
		_w16826_,
		_w16829_,
		_w16832_,
		_w16833_
	);
	LUT3 #(
		.INIT('h9a)
	) name11007 (
		\u1_L11_reg[29]/NET0131 ,
		_w16824_,
		_w16833_,
		_w16834_
	);
	LUT4 #(
		.INIT('hc963)
	) name11008 (
		decrypt_pad,
		\u1_R11_reg[32]/NET0131 ,
		\u1_uk_K_r11_reg[42]/NET0131 ,
		\u1_uk_K_r11_reg[51]/NET0131 ,
		_w16835_
	);
	LUT4 #(
		.INIT('hc693)
	) name11009 (
		decrypt_pad,
		\u1_R11_reg[29]/NET0131 ,
		\u1_uk_K_r11_reg[1]/NET0131 ,
		\u1_uk_K_r11_reg[23]/NET0131 ,
		_w16836_
	);
	LUT4 #(
		.INIT('hc693)
	) name11010 (
		decrypt_pad,
		\u1_R11_reg[1]/NET0131 ,
		\u1_uk_K_r11_reg[45]/NET0131 ,
		\u1_uk_K_r11_reg[8]/NET0131 ,
		_w16837_
	);
	LUT4 #(
		.INIT('hc693)
	) name11011 (
		decrypt_pad,
		\u1_R11_reg[28]/NET0131 ,
		\u1_uk_K_r11_reg[29]/NET0131 ,
		\u1_uk_K_r11_reg[51]/NET0131 ,
		_w16838_
	);
	LUT4 #(
		.INIT('hc693)
	) name11012 (
		decrypt_pad,
		\u1_R11_reg[30]/NET0131 ,
		\u1_uk_K_r11_reg[2]/NET0131 ,
		\u1_uk_K_r11_reg[52]/NET0131 ,
		_w16839_
	);
	LUT4 #(
		.INIT('h0200)
	) name11013 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16840_
	);
	LUT4 #(
		.INIT('hc693)
	) name11014 (
		decrypt_pad,
		\u1_R11_reg[31]/NET0131 ,
		\u1_uk_K_r11_reg[14]/NET0131 ,
		\u1_uk_K_r11_reg[36]/NET0131 ,
		_w16841_
	);
	LUT2 #(
		.INIT('h4)
	) name11015 (
		_w16837_,
		_w16836_,
		_w16842_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name11016 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16843_
	);
	LUT3 #(
		.INIT('h02)
	) name11017 (
		_w16841_,
		_w16840_,
		_w16843_,
		_w16844_
	);
	LUT4 #(
		.INIT('h4000)
	) name11018 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16845_
	);
	LUT4 #(
		.INIT('h0009)
	) name11019 (
		_w16838_,
		_w16839_,
		_w16836_,
		_w16841_,
		_w16846_
	);
	LUT2 #(
		.INIT('h1)
	) name11020 (
		_w16845_,
		_w16846_,
		_w16847_
	);
	LUT3 #(
		.INIT('h8a)
	) name11021 (
		_w16835_,
		_w16844_,
		_w16847_,
		_w16848_
	);
	LUT3 #(
		.INIT('h10)
	) name11022 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16849_
	);
	LUT2 #(
		.INIT('h8)
	) name11023 (
		_w16837_,
		_w16836_,
		_w16850_
	);
	LUT3 #(
		.INIT('h07)
	) name11024 (
		_w16837_,
		_w16836_,
		_w16841_,
		_w16851_
	);
	LUT4 #(
		.INIT('h0020)
	) name11025 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16852_
	);
	LUT4 #(
		.INIT('hfb00)
	) name11026 (
		_w16838_,
		_w16837_,
		_w16836_,
		_w16841_,
		_w16853_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name11027 (
		_w16849_,
		_w16851_,
		_w16852_,
		_w16853_,
		_w16854_
	);
	LUT3 #(
		.INIT('h02)
	) name11028 (
		_w16838_,
		_w16839_,
		_w16841_,
		_w16855_
	);
	LUT4 #(
		.INIT('h8000)
	) name11029 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16856_
	);
	LUT3 #(
		.INIT('h01)
	) name11030 (
		_w16855_,
		_w16856_,
		_w16840_,
		_w16857_
	);
	LUT4 #(
		.INIT('h1000)
	) name11031 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16858_
	);
	LUT4 #(
		.INIT('h0040)
	) name11032 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16859_
	);
	LUT4 #(
		.INIT('hefb6)
	) name11033 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16860_
	);
	LUT4 #(
		.INIT('h3f15)
	) name11034 (
		_w16841_,
		_w16855_,
		_w16842_,
		_w16860_,
		_w16861_
	);
	LUT4 #(
		.INIT('hba00)
	) name11035 (
		_w16835_,
		_w16854_,
		_w16857_,
		_w16861_,
		_w16862_
	);
	LUT3 #(
		.INIT('h9a)
	) name11036 (
		\u1_L11_reg[5]/NET0131 ,
		_w16848_,
		_w16862_,
		_w16863_
	);
	LUT4 #(
		.INIT('h2000)
	) name11037 (
		_w16722_,
		_w16723_,
		_w16720_,
		_w16724_,
		_w16864_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11038 (
		_w16721_,
		_w16723_,
		_w16724_,
		_w16719_,
		_w16865_
	);
	LUT2 #(
		.INIT('h4)
	) name11039 (
		_w16864_,
		_w16865_,
		_w16866_
	);
	LUT3 #(
		.INIT('h51)
	) name11040 (
		_w16747_,
		_w16731_,
		_w16725_,
		_w16867_
	);
	LUT4 #(
		.INIT('hf070)
	) name11041 (
		_w16721_,
		_w16722_,
		_w16720_,
		_w16724_,
		_w16868_
	);
	LUT4 #(
		.INIT('hbcff)
	) name11042 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16869_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name11043 (
		_w16721_,
		_w16722_,
		_w16720_,
		_w16724_,
		_w16870_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name11044 (
		_w16822_,
		_w16868_,
		_w16869_,
		_w16870_,
		_w16871_
	);
	LUT3 #(
		.INIT('h01)
	) name11045 (
		_w16719_,
		_w16732_,
		_w16830_,
		_w16872_
	);
	LUT4 #(
		.INIT('h7077)
	) name11046 (
		_w16866_,
		_w16867_,
		_w16871_,
		_w16872_,
		_w16873_
	);
	LUT3 #(
		.INIT('h31)
	) name11047 (
		_w16721_,
		_w16722_,
		_w16724_,
		_w16874_
	);
	LUT4 #(
		.INIT('hd060)
	) name11048 (
		_w16721_,
		_w16722_,
		_w16720_,
		_w16724_,
		_w16875_
	);
	LUT4 #(
		.INIT('h070b)
	) name11049 (
		_w16721_,
		_w16722_,
		_w16720_,
		_w16724_,
		_w16876_
	);
	LUT4 #(
		.INIT('h3331)
	) name11050 (
		_w16723_,
		_w16749_,
		_w16876_,
		_w16875_,
		_w16877_
	);
	LUT3 #(
		.INIT('h65)
	) name11051 (
		\u1_L11_reg[4]/NET0131 ,
		_w16873_,
		_w16877_,
		_w16878_
	);
	LUT4 #(
		.INIT('hc693)
	) name11052 (
		decrypt_pad,
		\u1_R11_reg[6]/NET0131 ,
		\u1_uk_K_r11_reg[12]/NET0131 ,
		\u1_uk_K_r11_reg[32]/NET0131 ,
		_w16879_
	);
	LUT4 #(
		.INIT('hc693)
	) name11053 (
		decrypt_pad,
		\u1_R11_reg[9]/NET0131 ,
		\u1_uk_K_r11_reg[34]/NET0131 ,
		\u1_uk_K_r11_reg[54]/NET0131 ,
		_w16880_
	);
	LUT4 #(
		.INIT('hc963)
	) name11054 (
		decrypt_pad,
		\u1_R11_reg[5]/NET0131 ,
		\u1_uk_K_r11_reg[41]/NET0131 ,
		\u1_uk_K_r11_reg[46]/NET0131 ,
		_w16881_
	);
	LUT2 #(
		.INIT('h4)
	) name11055 (
		_w16880_,
		_w16881_,
		_w16882_
	);
	LUT4 #(
		.INIT('hc693)
	) name11056 (
		decrypt_pad,
		\u1_R11_reg[4]/NET0131 ,
		\u1_uk_K_r11_reg[10]/NET0131 ,
		\u1_uk_K_r11_reg[5]/NET0131 ,
		_w16883_
	);
	LUT2 #(
		.INIT('h2)
	) name11057 (
		_w16880_,
		_w16881_,
		_w16884_
	);
	LUT4 #(
		.INIT('h1012)
	) name11058 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16885_
	);
	LUT4 #(
		.INIT('hc963)
	) name11059 (
		decrypt_pad,
		\u1_R11_reg[7]/NET0131 ,
		\u1_uk_K_r11_reg[26]/NET0131 ,
		\u1_uk_K_r11_reg[6]/NET0131 ,
		_w16886_
	);
	LUT3 #(
		.INIT('h80)
	) name11060 (
		_w16886_,
		_w16879_,
		_w16883_,
		_w16887_
	);
	LUT4 #(
		.INIT('hc963)
	) name11061 (
		decrypt_pad,
		\u1_R11_reg[8]/NET0131 ,
		\u1_uk_K_r11_reg[17]/NET0131 ,
		\u1_uk_K_r11_reg[54]/NET0131 ,
		_w16888_
	);
	LUT4 #(
		.INIT('h0013)
	) name11062 (
		_w16884_,
		_w16885_,
		_w16887_,
		_w16888_,
		_w16889_
	);
	LUT2 #(
		.INIT('h2)
	) name11063 (
		_w16880_,
		_w16879_,
		_w16890_
	);
	LUT4 #(
		.INIT('h0004)
	) name11064 (
		_w16886_,
		_w16880_,
		_w16879_,
		_w16881_,
		_w16891_
	);
	LUT4 #(
		.INIT('h0080)
	) name11065 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16892_
	);
	LUT4 #(
		.INIT('h3bf5)
	) name11066 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16893_
	);
	LUT4 #(
		.INIT('h0302)
	) name11067 (
		_w16886_,
		_w16891_,
		_w16892_,
		_w16893_,
		_w16894_
	);
	LUT2 #(
		.INIT('h8)
	) name11068 (
		_w16889_,
		_w16894_,
		_w16895_
	);
	LUT2 #(
		.INIT('h8)
	) name11069 (
		_w16880_,
		_w16883_,
		_w16896_
	);
	LUT2 #(
		.INIT('h6)
	) name11070 (
		_w16880_,
		_w16883_,
		_w16897_
	);
	LUT4 #(
		.INIT('h0444)
	) name11071 (
		_w16886_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16898_
	);
	LUT2 #(
		.INIT('h4)
	) name11072 (
		_w16897_,
		_w16898_,
		_w16899_
	);
	LUT3 #(
		.INIT('h10)
	) name11073 (
		_w16880_,
		_w16879_,
		_w16883_,
		_w16900_
	);
	LUT4 #(
		.INIT('h0100)
	) name11074 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16901_
	);
	LUT4 #(
		.INIT('h2000)
	) name11075 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16902_
	);
	LUT4 #(
		.INIT('h0001)
	) name11076 (
		_w16886_,
		_w16880_,
		_w16881_,
		_w16883_,
		_w16903_
	);
	LUT4 #(
		.INIT('ha020)
	) name11077 (
		_w16886_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16904_
	);
	LUT4 #(
		.INIT('h0002)
	) name11078 (
		_w16888_,
		_w16902_,
		_w16903_,
		_w16904_,
		_w16905_
	);
	LUT3 #(
		.INIT('h10)
	) name11079 (
		_w16899_,
		_w16901_,
		_w16905_,
		_w16906_
	);
	LUT4 #(
		.INIT('h0004)
	) name11080 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16907_
	);
	LUT4 #(
		.INIT('hcffb)
	) name11081 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16908_
	);
	LUT2 #(
		.INIT('h9)
	) name11082 (
		_w16879_,
		_w16881_,
		_w16909_
	);
	LUT3 #(
		.INIT('h04)
	) name11083 (
		_w16886_,
		_w16880_,
		_w16883_,
		_w16910_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name11084 (
		_w16886_,
		_w16908_,
		_w16909_,
		_w16910_,
		_w16911_
	);
	LUT4 #(
		.INIT('ha955)
	) name11085 (
		\u1_L11_reg[2]/NET0131 ,
		_w16895_,
		_w16906_,
		_w16911_,
		_w16912_
	);
	LUT3 #(
		.INIT('h02)
	) name11086 (
		_w16786_,
		_w16794_,
		_w16796_,
		_w16913_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11087 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w16914_
	);
	LUT3 #(
		.INIT('h01)
	) name11088 (
		_w16786_,
		_w16808_,
		_w16914_,
		_w16915_
	);
	LUT4 #(
		.INIT('h6fff)
	) name11089 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w16916_
	);
	LUT4 #(
		.INIT('h02aa)
	) name11090 (
		_w16797_,
		_w16913_,
		_w16915_,
		_w16916_,
		_w16917_
	);
	LUT3 #(
		.INIT('h08)
	) name11091 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16918_
	);
	LUT4 #(
		.INIT('h0400)
	) name11092 (
		_w16786_,
		_w16784_,
		_w16788_,
		_w16785_,
		_w16919_
	);
	LUT3 #(
		.INIT('h01)
	) name11093 (
		_w16802_,
		_w16918_,
		_w16919_,
		_w16920_
	);
	LUT3 #(
		.INIT('h8a)
	) name11094 (
		_w16786_,
		_w16788_,
		_w16785_,
		_w16921_
	);
	LUT4 #(
		.INIT('h0200)
	) name11095 (
		_w16786_,
		_w16784_,
		_w16788_,
		_w16785_,
		_w16922_
	);
	LUT3 #(
		.INIT('h07)
	) name11096 (
		_w16805_,
		_w16921_,
		_w16922_,
		_w16923_
	);
	LUT4 #(
		.INIT('h1333)
	) name11097 (
		_w16795_,
		_w16797_,
		_w16920_,
		_w16923_,
		_w16924_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name11098 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w16925_
	);
	LUT2 #(
		.INIT('h1)
	) name11099 (
		_w16786_,
		_w16925_,
		_w16926_
	);
	LUT3 #(
		.INIT('h0b)
	) name11100 (
		_w16788_,
		_w16809_,
		_w16799_,
		_w16927_
	);
	LUT2 #(
		.INIT('h4)
	) name11101 (
		_w16926_,
		_w16927_,
		_w16928_
	);
	LUT4 #(
		.INIT('h5655)
	) name11102 (
		\u1_L11_reg[10]/NET0131 ,
		_w16924_,
		_w16917_,
		_w16928_,
		_w16929_
	);
	LUT3 #(
		.INIT('h54)
	) name11103 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16930_
	);
	LUT3 #(
		.INIT('ha2)
	) name11104 (
		_w16754_,
		_w16756_,
		_w16757_,
		_w16931_
	);
	LUT4 #(
		.INIT('h0189)
	) name11105 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16932_
	);
	LUT4 #(
		.INIT('h0816)
	) name11106 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16933_
	);
	LUT3 #(
		.INIT('h41)
	) name11107 (
		_w16753_,
		_w16755_,
		_w16757_,
		_w16934_
	);
	LUT3 #(
		.INIT('h53)
	) name11108 (
		_w16756_,
		_w16753_,
		_w16755_,
		_w16935_
	);
	LUT4 #(
		.INIT('h00f7)
	) name11109 (
		_w16754_,
		_w16756_,
		_w16753_,
		_w16767_,
		_w16936_
	);
	LUT4 #(
		.INIT('h0d00)
	) name11110 (
		_w16765_,
		_w16935_,
		_w16934_,
		_w16936_,
		_w16937_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name11111 (
		_w16754_,
		_w16753_,
		_w16755_,
		_w16757_,
		_w16938_
	);
	LUT2 #(
		.INIT('h4)
	) name11112 (
		_w16930_,
		_w16938_,
		_w16939_
	);
	LUT4 #(
		.INIT('h1248)
	) name11113 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w16940_
	);
	LUT4 #(
		.INIT('h00b0)
	) name11114 (
		_w16753_,
		_w16766_,
		_w16767_,
		_w16940_,
		_w16941_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name11115 (
		_w16933_,
		_w16937_,
		_w16939_,
		_w16941_,
		_w16942_
	);
	LUT2 #(
		.INIT('h6)
	) name11116 (
		\u1_L11_reg[12]/NET0131 ,
		_w16942_,
		_w16943_
	);
	LUT4 #(
		.INIT('h0008)
	) name11117 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16944_
	);
	LUT4 #(
		.INIT('hfea7)
	) name11118 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16945_
	);
	LUT4 #(
		.INIT('h4000)
	) name11119 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16946_
	);
	LUT4 #(
		.INIT('h9fff)
	) name11120 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16947_
	);
	LUT4 #(
		.INIT('h0155)
	) name11121 (
		_w16886_,
		_w16888_,
		_w16945_,
		_w16947_,
		_w16948_
	);
	LUT4 #(
		.INIT('he5fa)
	) name11122 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16949_
	);
	LUT2 #(
		.INIT('h2)
	) name11123 (
		_w16886_,
		_w16949_,
		_w16950_
	);
	LUT3 #(
		.INIT('h0e)
	) name11124 (
		_w16886_,
		_w16881_,
		_w16883_,
		_w16951_
	);
	LUT2 #(
		.INIT('h8)
	) name11125 (
		_w16890_,
		_w16951_,
		_w16952_
	);
	LUT3 #(
		.INIT('h0b)
	) name11126 (
		_w16882_,
		_w16887_,
		_w16888_,
		_w16953_
	);
	LUT3 #(
		.INIT('h10)
	) name11127 (
		_w16950_,
		_w16952_,
		_w16953_,
		_w16954_
	);
	LUT4 #(
		.INIT('h0010)
	) name11128 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16955_
	);
	LUT3 #(
		.INIT('h02)
	) name11129 (
		_w16888_,
		_w16902_,
		_w16955_,
		_w16956_
	);
	LUT2 #(
		.INIT('h1)
	) name11130 (
		_w16880_,
		_w16879_,
		_w16957_
	);
	LUT4 #(
		.INIT('h0501)
	) name11131 (
		_w16886_,
		_w16880_,
		_w16881_,
		_w16883_,
		_w16958_
	);
	LUT3 #(
		.INIT('h45)
	) name11132 (
		_w16946_,
		_w16957_,
		_w16958_,
		_w16959_
	);
	LUT4 #(
		.INIT('hfe76)
	) name11133 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w16960_
	);
	LUT4 #(
		.INIT('h0301)
	) name11134 (
		_w16886_,
		_w16891_,
		_w16892_,
		_w16960_,
		_w16961_
	);
	LUT3 #(
		.INIT('h80)
	) name11135 (
		_w16956_,
		_w16959_,
		_w16961_,
		_w16962_
	);
	LUT4 #(
		.INIT('h999a)
	) name11136 (
		\u1_L11_reg[13]/NET0131 ,
		_w16948_,
		_w16954_,
		_w16962_,
		_w16963_
	);
	LUT4 #(
		.INIT('h0002)
	) name11137 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16964_
	);
	LUT4 #(
		.INIT('h54bb)
	) name11138 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16965_
	);
	LUT4 #(
		.INIT('h5054)
	) name11139 (
		_w16835_,
		_w16841_,
		_w16964_,
		_w16965_,
		_w16966_
	);
	LUT2 #(
		.INIT('h4)
	) name11140 (
		_w16838_,
		_w16841_,
		_w16967_
	);
	LUT3 #(
		.INIT('h08)
	) name11141 (
		_w16837_,
		_w16839_,
		_w16836_,
		_w16968_
	);
	LUT2 #(
		.INIT('h4)
	) name11142 (
		_w16967_,
		_w16968_,
		_w16969_
	);
	LUT3 #(
		.INIT('h20)
	) name11143 (
		_w16838_,
		_w16839_,
		_w16836_,
		_w16970_
	);
	LUT2 #(
		.INIT('h4)
	) name11144 (
		_w16836_,
		_w16841_,
		_w16971_
	);
	LUT4 #(
		.INIT('h0100)
	) name11145 (
		_w16838_,
		_w16837_,
		_w16836_,
		_w16841_,
		_w16972_
	);
	LUT3 #(
		.INIT('h01)
	) name11146 (
		_w16858_,
		_w16972_,
		_w16970_,
		_w16973_
	);
	LUT4 #(
		.INIT('heb5e)
	) name11147 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16974_
	);
	LUT4 #(
		.INIT('h0004)
	) name11148 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16975_
	);
	LUT4 #(
		.INIT('hbffb)
	) name11149 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16976_
	);
	LUT4 #(
		.INIT('h0004)
	) name11150 (
		_w16835_,
		_w16838_,
		_w16836_,
		_w16841_,
		_w16977_
	);
	LUT4 #(
		.INIT('h00e4)
	) name11151 (
		_w16841_,
		_w16974_,
		_w16976_,
		_w16977_,
		_w16978_
	);
	LUT4 #(
		.INIT('h7500)
	) name11152 (
		_w16835_,
		_w16969_,
		_w16973_,
		_w16978_,
		_w16979_
	);
	LUT3 #(
		.INIT('h65)
	) name11153 (
		\u1_L11_reg[15]/P0001 ,
		_w16966_,
		_w16979_,
		_w16980_
	);
	LUT4 #(
		.INIT('h0201)
	) name11154 (
		_w16721_,
		_w16722_,
		_w16720_,
		_w16724_,
		_w16981_
	);
	LUT4 #(
		.INIT('hf700)
	) name11155 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16720_,
		_w16982_
	);
	LUT4 #(
		.INIT('h8000)
	) name11156 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16983_
	);
	LUT4 #(
		.INIT('h0045)
	) name11157 (
		_w16719_,
		_w16874_,
		_w16982_,
		_w16983_,
		_w16984_
	);
	LUT4 #(
		.INIT('h2010)
	) name11158 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16985_
	);
	LUT3 #(
		.INIT('h04)
	) name11159 (
		_w16736_,
		_w16719_,
		_w16985_,
		_w16986_
	);
	LUT4 #(
		.INIT('h010a)
	) name11160 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16724_,
		_w16987_
	);
	LUT4 #(
		.INIT('h0844)
	) name11161 (
		_w16721_,
		_w16722_,
		_w16723_,
		_w16720_,
		_w16988_
	);
	LUT2 #(
		.INIT('h1)
	) name11162 (
		_w16987_,
		_w16988_,
		_w16989_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name11163 (
		_w16981_,
		_w16984_,
		_w16986_,
		_w16989_,
		_w16990_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name11164 (
		_w16721_,
		_w16723_,
		_w16745_,
		_w16732_,
		_w16991_
	);
	LUT3 #(
		.INIT('h65)
	) name11165 (
		\u1_L11_reg[19]/P0001 ,
		_w16990_,
		_w16991_,
		_w16992_
	);
	LUT3 #(
		.INIT('h08)
	) name11166 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16993_
	);
	LUT2 #(
		.INIT('h4)
	) name11167 (
		_w16971_,
		_w16993_,
		_w16994_
	);
	LUT4 #(
		.INIT('h4555)
	) name11168 (
		_w16835_,
		_w16838_,
		_w16839_,
		_w16836_,
		_w16995_
	);
	LUT4 #(
		.INIT('h0040)
	) name11169 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16841_,
		_w16996_
	);
	LUT4 #(
		.INIT('h0010)
	) name11170 (
		_w16838_,
		_w16837_,
		_w16836_,
		_w16841_,
		_w16997_
	);
	LUT3 #(
		.INIT('h10)
	) name11171 (
		_w16996_,
		_w16997_,
		_w16995_,
		_w16998_
	);
	LUT4 #(
		.INIT('h0021)
	) name11172 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w16999_
	);
	LUT4 #(
		.INIT('hdd5f)
	) name11173 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w17000_
	);
	LUT3 #(
		.INIT('h31)
	) name11174 (
		_w16841_,
		_w16999_,
		_w17000_,
		_w17001_
	);
	LUT3 #(
		.INIT('h40)
	) name11175 (
		_w16994_,
		_w16998_,
		_w17001_,
		_w17002_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11176 (
		_w16838_,
		_w16839_,
		_w16836_,
		_w16841_,
		_w17003_
	);
	LUT4 #(
		.INIT('hbbf3)
	) name11177 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w17004_
	);
	LUT4 #(
		.INIT('h0080)
	) name11178 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w17005_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11179 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16841_,
		_w17006_
	);
	LUT4 #(
		.INIT('h7077)
	) name11180 (
		_w17003_,
		_w17004_,
		_w17005_,
		_w17006_,
		_w17007_
	);
	LUT4 #(
		.INIT('h2010)
	) name11181 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w17008_
	);
	LUT3 #(
		.INIT('h02)
	) name11182 (
		_w16835_,
		_w16975_,
		_w17008_,
		_w17009_
	);
	LUT2 #(
		.INIT('h4)
	) name11183 (
		_w17007_,
		_w17009_,
		_w17010_
	);
	LUT4 #(
		.INIT('h0100)
	) name11184 (
		_w16838_,
		_w16839_,
		_w16836_,
		_w16841_,
		_w17011_
	);
	LUT3 #(
		.INIT('h07)
	) name11185 (
		_w16850_,
		_w16855_,
		_w17011_,
		_w17012_
	);
	LUT4 #(
		.INIT('ha955)
	) name11186 (
		\u1_L11_reg[21]/NET0131 ,
		_w17002_,
		_w17010_,
		_w17012_,
		_w17013_
	);
	LUT4 #(
		.INIT('hccfd)
	) name11187 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17014_
	);
	LUT4 #(
		.INIT('h6fbf)
	) name11188 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17015_
	);
	LUT4 #(
		.INIT('h08aa)
	) name11189 (
		_w16786_,
		_w16797_,
		_w17014_,
		_w17015_,
		_w17016_
	);
	LUT4 #(
		.INIT('h220a)
	) name11190 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17017_
	);
	LUT4 #(
		.INIT('hfda8)
	) name11191 (
		_w16786_,
		_w16792_,
		_w16814_,
		_w17017_,
		_w17018_
	);
	LUT4 #(
		.INIT('h7bf7)
	) name11192 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17019_
	);
	LUT3 #(
		.INIT('h45)
	) name11193 (
		_w16797_,
		_w17018_,
		_w17019_,
		_w17020_
	);
	LUT4 #(
		.INIT('hb3fb)
	) name11194 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17021_
	);
	LUT4 #(
		.INIT('h0080)
	) name11195 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17022_
	);
	LUT4 #(
		.INIT('hef6f)
	) name11196 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17023_
	);
	LUT4 #(
		.INIT('h04cc)
	) name11197 (
		_w16786_,
		_w16797_,
		_w17021_,
		_w17023_,
		_w17024_
	);
	LUT2 #(
		.INIT('h1)
	) name11198 (
		_w16786_,
		_w16785_,
		_w17025_
	);
	LUT2 #(
		.INIT('h4)
	) name11199 (
		_w17023_,
		_w17025_,
		_w17026_
	);
	LUT2 #(
		.INIT('h1)
	) name11200 (
		_w17024_,
		_w17026_,
		_w17027_
	);
	LUT4 #(
		.INIT('h5655)
	) name11201 (
		\u1_L11_reg[1]/NET0131 ,
		_w17020_,
		_w17016_,
		_w17027_,
		_w17028_
	);
	LUT3 #(
		.INIT('h96)
	) name11202 (
		_w16682_,
		_w16683_,
		_w16685_,
		_w17029_
	);
	LUT4 #(
		.INIT('h1055)
	) name11203 (
		_w16681_,
		_w16682_,
		_w16684_,
		_w16685_,
		_w17030_
	);
	LUT2 #(
		.INIT('h8)
	) name11204 (
		_w17029_,
		_w17030_,
		_w17031_
	);
	LUT4 #(
		.INIT('h1000)
	) name11205 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w17032_
	);
	LUT4 #(
		.INIT('h0080)
	) name11206 (
		_w16681_,
		_w16682_,
		_w16683_,
		_w16685_,
		_w17033_
	);
	LUT4 #(
		.INIT('h0007)
	) name11207 (
		_w16704_,
		_w16705_,
		_w17032_,
		_w17033_,
		_w17034_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11208 (
		_w16693_,
		_w16714_,
		_w17031_,
		_w17034_,
		_w17035_
	);
	LUT4 #(
		.INIT('h5400)
	) name11209 (
		_w16681_,
		_w16682_,
		_w16684_,
		_w16685_,
		_w17036_
	);
	LUT3 #(
		.INIT('h7e)
	) name11210 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w17037_
	);
	LUT4 #(
		.INIT('h4500)
	) name11211 (
		_w16698_,
		_w16711_,
		_w17036_,
		_w17037_,
		_w17038_
	);
	LUT4 #(
		.INIT('h7def)
	) name11212 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w17039_
	);
	LUT2 #(
		.INIT('h1)
	) name11213 (
		_w16681_,
		_w17039_,
		_w17040_
	);
	LUT2 #(
		.INIT('h8)
	) name11214 (
		_w16684_,
		_w16693_,
		_w17041_
	);
	LUT4 #(
		.INIT('h0008)
	) name11215 (
		_w16681_,
		_w16682_,
		_w16683_,
		_w16685_,
		_w17042_
	);
	LUT3 #(
		.INIT('h45)
	) name11216 (
		_w16715_,
		_w17041_,
		_w17042_,
		_w17043_
	);
	LUT4 #(
		.INIT('h0e00)
	) name11217 (
		_w16693_,
		_w17038_,
		_w17040_,
		_w17043_,
		_w17044_
	);
	LUT3 #(
		.INIT('h9a)
	) name11218 (
		\u1_L11_reg[23]/NET0131 ,
		_w17035_,
		_w17044_,
		_w17045_
	);
	LUT4 #(
		.INIT('hc693)
	) name11219 (
		decrypt_pad,
		\u1_R11_reg[19]/NET0131 ,
		\u1_uk_K_r11_reg[21]/NET0131 ,
		\u1_uk_K_r11_reg[43]/NET0131 ,
		_w17046_
	);
	LUT4 #(
		.INIT('hc693)
	) name11220 (
		decrypt_pad,
		\u1_R11_reg[17]/NET0131 ,
		\u1_uk_K_r11_reg[16]/NET0131 ,
		\u1_uk_K_r11_reg[7]/NET0131 ,
		_w17047_
	);
	LUT4 #(
		.INIT('hc963)
	) name11221 (
		decrypt_pad,
		\u1_R11_reg[21]/NET0131 ,
		\u1_uk_K_r11_reg[28]/NET0131 ,
		\u1_uk_K_r11_reg[37]/NET0131 ,
		_w17048_
	);
	LUT4 #(
		.INIT('hc963)
	) name11222 (
		decrypt_pad,
		\u1_R11_reg[16]/NET0131 ,
		\u1_uk_K_r11_reg[16]/NET0131 ,
		\u1_uk_K_r11_reg[49]/NET0131 ,
		_w17049_
	);
	LUT4 #(
		.INIT('h00bf)
	) name11223 (
		_w17047_,
		_w17048_,
		_w17049_,
		_w17046_,
		_w17050_
	);
	LUT4 #(
		.INIT('hc963)
	) name11224 (
		decrypt_pad,
		\u1_R11_reg[18]/NET0131 ,
		\u1_uk_K_r11_reg[1]/NET0131 ,
		\u1_uk_K_r11_reg[38]/NET0131 ,
		_w17051_
	);
	LUT3 #(
		.INIT('h02)
	) name11225 (
		_w17047_,
		_w17051_,
		_w17049_,
		_w17052_
	);
	LUT2 #(
		.INIT('h2)
	) name11226 (
		_w17051_,
		_w17049_,
		_w17053_
	);
	LUT4 #(
		.INIT('h010d)
	) name11227 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17054_
	);
	LUT3 #(
		.INIT('h80)
	) name11228 (
		_w17047_,
		_w17048_,
		_w17049_,
		_w17055_
	);
	LUT4 #(
		.INIT('h7a00)
	) name11229 (
		_w17047_,
		_w17048_,
		_w17049_,
		_w17046_,
		_w17056_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name11230 (
		_w17050_,
		_w17052_,
		_w17054_,
		_w17056_,
		_w17057_
	);
	LUT4 #(
		.INIT('hd7df)
	) name11231 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17058_
	);
	LUT4 #(
		.INIT('hc963)
	) name11232 (
		decrypt_pad,
		\u1_R11_reg[20]/NET0131 ,
		\u1_uk_K_r11_reg[31]/NET0131 ,
		\u1_uk_K_r11_reg[36]/NET0131 ,
		_w17059_
	);
	LUT3 #(
		.INIT('hb0)
	) name11233 (
		_w17057_,
		_w17058_,
		_w17059_,
		_w17060_
	);
	LUT4 #(
		.INIT('hf7fb)
	) name11234 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17061_
	);
	LUT4 #(
		.INIT('hf7eb)
	) name11235 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17062_
	);
	LUT2 #(
		.INIT('h2)
	) name11236 (
		_w17046_,
		_w17062_,
		_w17063_
	);
	LUT3 #(
		.INIT('h20)
	) name11237 (
		_w17051_,
		_w17048_,
		_w17046_,
		_w17064_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name11238 (
		_w17051_,
		_w17048_,
		_w17049_,
		_w17046_,
		_w17065_
	);
	LUT3 #(
		.INIT('h02)
	) name11239 (
		_w17047_,
		_w17065_,
		_w17064_,
		_w17066_
	);
	LUT4 #(
		.INIT('h0015)
	) name11240 (
		_w17047_,
		_w17048_,
		_w17049_,
		_w17046_,
		_w17067_
	);
	LUT2 #(
		.INIT('h4)
	) name11241 (
		_w17053_,
		_w17067_,
		_w17068_
	);
	LUT4 #(
		.INIT('h2000)
	) name11242 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17069_
	);
	LUT4 #(
		.INIT('h0040)
	) name11243 (
		_w17047_,
		_w17051_,
		_w17049_,
		_w17046_,
		_w17070_
	);
	LUT2 #(
		.INIT('h1)
	) name11244 (
		_w17069_,
		_w17070_,
		_w17071_
	);
	LUT4 #(
		.INIT('hab00)
	) name11245 (
		_w17059_,
		_w17066_,
		_w17068_,
		_w17071_,
		_w17072_
	);
	LUT4 #(
		.INIT('h5655)
	) name11246 (
		\u1_L11_reg[25]/NET0131 ,
		_w17060_,
		_w17063_,
		_w17072_,
		_w17073_
	);
	LUT4 #(
		.INIT('ha040)
	) name11247 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w17074_
	);
	LUT4 #(
		.INIT('h3700)
	) name11248 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w17075_
	);
	LUT4 #(
		.INIT('h0002)
	) name11249 (
		_w16886_,
		_w16944_,
		_w17075_,
		_w17074_,
		_w17076_
	);
	LUT4 #(
		.INIT('hbff3)
	) name11250 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w17077_
	);
	LUT4 #(
		.INIT('h5515)
	) name11251 (
		_w16886_,
		_w16880_,
		_w16881_,
		_w16883_,
		_w17078_
	);
	LUT3 #(
		.INIT('h01)
	) name11252 (
		_w16880_,
		_w16879_,
		_w16883_,
		_w17079_
	);
	LUT4 #(
		.INIT('hfdee)
	) name11253 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w17080_
	);
	LUT3 #(
		.INIT('h80)
	) name11254 (
		_w17078_,
		_w17077_,
		_w17080_,
		_w17081_
	);
	LUT3 #(
		.INIT('ha8)
	) name11255 (
		_w16888_,
		_w17076_,
		_w17081_,
		_w17082_
	);
	LUT4 #(
		.INIT('h0551)
	) name11256 (
		_w16886_,
		_w16880_,
		_w16881_,
		_w16883_,
		_w17083_
	);
	LUT3 #(
		.INIT('h40)
	) name11257 (
		_w16900_,
		_w17077_,
		_w17083_,
		_w17084_
	);
	LUT4 #(
		.INIT('haa2a)
	) name11258 (
		_w16886_,
		_w16880_,
		_w16881_,
		_w16883_,
		_w17085_
	);
	LUT2 #(
		.INIT('h4)
	) name11259 (
		_w17079_,
		_w17085_,
		_w17086_
	);
	LUT4 #(
		.INIT('h4804)
	) name11260 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w17087_
	);
	LUT2 #(
		.INIT('h1)
	) name11261 (
		_w16888_,
		_w17087_,
		_w17088_
	);
	LUT3 #(
		.INIT('he0)
	) name11262 (
		_w17084_,
		_w17086_,
		_w17088_,
		_w17089_
	);
	LUT3 #(
		.INIT('ha9)
	) name11263 (
		\u1_L11_reg[28]/NET0131 ,
		_w17082_,
		_w17089_,
		_w17090_
	);
	LUT4 #(
		.INIT('hfd00)
	) name11264 (
		_w17047_,
		_w17051_,
		_w17049_,
		_w17046_,
		_w17091_
	);
	LUT4 #(
		.INIT('h3ffa)
	) name11265 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17092_
	);
	LUT2 #(
		.INIT('h8)
	) name11266 (
		_w17091_,
		_w17092_,
		_w17093_
	);
	LUT4 #(
		.INIT('h0100)
	) name11267 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17094_
	);
	LUT3 #(
		.INIT('h08)
	) name11268 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17095_
	);
	LUT4 #(
		.INIT('hf7a7)
	) name11269 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17096_
	);
	LUT4 #(
		.INIT('h0100)
	) name11270 (
		_w17046_,
		_w17069_,
		_w17094_,
		_w17096_,
		_w17097_
	);
	LUT4 #(
		.INIT('h4000)
	) name11271 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17098_
	);
	LUT4 #(
		.INIT('hbffd)
	) name11272 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17099_
	);
	LUT4 #(
		.INIT('h0155)
	) name11273 (
		_w17059_,
		_w17093_,
		_w17097_,
		_w17099_,
		_w17100_
	);
	LUT4 #(
		.INIT('hc52f)
	) name11274 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17101_
	);
	LUT2 #(
		.INIT('h2)
	) name11275 (
		_w17046_,
		_w17101_,
		_w17102_
	);
	LUT2 #(
		.INIT('h1)
	) name11276 (
		_w17051_,
		_w17046_,
		_w17103_
	);
	LUT3 #(
		.INIT('h08)
	) name11277 (
		_w17047_,
		_w17048_,
		_w17049_,
		_w17104_
	);
	LUT3 #(
		.INIT('hf6)
	) name11278 (
		_w17047_,
		_w17048_,
		_w17049_,
		_w17105_
	);
	LUT2 #(
		.INIT('h2)
	) name11279 (
		_w17103_,
		_w17105_,
		_w17106_
	);
	LUT2 #(
		.INIT('h9)
	) name11280 (
		_w17047_,
		_w17051_,
		_w17107_
	);
	LUT4 #(
		.INIT('h0600)
	) name11281 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17108_
	);
	LUT3 #(
		.INIT('ha2)
	) name11282 (
		_w17047_,
		_w17051_,
		_w17046_,
		_w17109_
	);
	LUT4 #(
		.INIT('hb000)
	) name11283 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17110_
	);
	LUT3 #(
		.INIT('h45)
	) name11284 (
		_w17108_,
		_w17109_,
		_w17110_,
		_w17111_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11285 (
		_w17059_,
		_w17102_,
		_w17106_,
		_w17111_,
		_w17112_
	);
	LUT4 #(
		.INIT('hfdfb)
	) name11286 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17113_
	);
	LUT4 #(
		.INIT('h0040)
	) name11287 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17114_
	);
	LUT4 #(
		.INIT('hffb7)
	) name11288 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17115_
	);
	LUT3 #(
		.INIT('hd8)
	) name11289 (
		_w17046_,
		_w17113_,
		_w17115_,
		_w17116_
	);
	LUT4 #(
		.INIT('h5655)
	) name11290 (
		\u1_L11_reg[14]/NET0131 ,
		_w17100_,
		_w17112_,
		_w17116_,
		_w17117_
	);
	LUT3 #(
		.INIT('h02)
	) name11291 (
		_w16786_,
		_w16808_,
		_w16796_,
		_w17118_
	);
	LUT4 #(
		.INIT('h0806)
	) name11292 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17119_
	);
	LUT4 #(
		.INIT('hefcc)
	) name11293 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17120_
	);
	LUT4 #(
		.INIT('h0504)
	) name11294 (
		_w16786_,
		_w16797_,
		_w17119_,
		_w17120_,
		_w17121_
	);
	LUT2 #(
		.INIT('h1)
	) name11295 (
		_w17118_,
		_w17121_,
		_w17122_
	);
	LUT4 #(
		.INIT('h0002)
	) name11296 (
		_w16786_,
		_w16784_,
		_w16783_,
		_w16785_,
		_w17123_
	);
	LUT4 #(
		.INIT('h0004)
	) name11297 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17124_
	);
	LUT4 #(
		.INIT('h0002)
	) name11298 (
		_w16797_,
		_w17022_,
		_w17123_,
		_w17124_,
		_w17125_
	);
	LUT4 #(
		.INIT('h54ff)
	) name11299 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16785_,
		_w17126_
	);
	LUT3 #(
		.INIT('h51)
	) name11300 (
		_w16786_,
		_w16784_,
		_w16788_,
		_w17127_
	);
	LUT4 #(
		.INIT('hcdff)
	) name11301 (
		_w16786_,
		_w16784_,
		_w16783_,
		_w16785_,
		_w17128_
	);
	LUT4 #(
		.INIT('hcf45)
	) name11302 (
		_w16788_,
		_w17126_,
		_w17127_,
		_w17128_,
		_w17129_
	);
	LUT2 #(
		.INIT('h2)
	) name11303 (
		_w16798_,
		_w16810_,
		_w17130_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11304 (
		_w16784_,
		_w16783_,
		_w16788_,
		_w16797_,
		_w17131_
	);
	LUT3 #(
		.INIT('h10)
	) name11305 (
		_w16808_,
		_w16809_,
		_w17131_,
		_w17132_
	);
	LUT4 #(
		.INIT('h7077)
	) name11306 (
		_w17125_,
		_w17129_,
		_w17130_,
		_w17132_,
		_w17133_
	);
	LUT3 #(
		.INIT('h56)
	) name11307 (
		\u1_L11_reg[26]/NET0131 ,
		_w17122_,
		_w17133_,
		_w17134_
	);
	LUT4 #(
		.INIT('h0400)
	) name11308 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17135_
	);
	LUT2 #(
		.INIT('h1)
	) name11309 (
		_w17046_,
		_w17135_,
		_w17136_
	);
	LUT3 #(
		.INIT('hd0)
	) name11310 (
		_w17048_,
		_w17049_,
		_w17046_,
		_w17137_
	);
	LUT3 #(
		.INIT('h54)
	) name11311 (
		_w17095_,
		_w17107_,
		_w17137_,
		_w17138_
	);
	LUT2 #(
		.INIT('h1)
	) name11312 (
		_w17136_,
		_w17138_,
		_w17139_
	);
	LUT4 #(
		.INIT('haffe)
	) name11313 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17140_
	);
	LUT4 #(
		.INIT('hfb00)
	) name11314 (
		_w17051_,
		_w17049_,
		_w17046_,
		_w17059_,
		_w17141_
	);
	LUT4 #(
		.INIT('hc400)
	) name11315 (
		_w17046_,
		_w17115_,
		_w17140_,
		_w17141_,
		_w17142_
	);
	LUT4 #(
		.INIT('h00b0)
	) name11316 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17143_
	);
	LUT2 #(
		.INIT('h2)
	) name11317 (
		_w17050_,
		_w17143_,
		_w17144_
	);
	LUT3 #(
		.INIT('h02)
	) name11318 (
		_w17046_,
		_w17055_,
		_w17094_,
		_w17145_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11319 (
		_w17047_,
		_w17051_,
		_w17049_,
		_w17059_,
		_w17146_
	);
	LUT2 #(
		.INIT('h8)
	) name11320 (
		_w17061_,
		_w17146_,
		_w17147_
	);
	LUT4 #(
		.INIT('h0155)
	) name11321 (
		_w17142_,
		_w17144_,
		_w17145_,
		_w17147_,
		_w17148_
	);
	LUT3 #(
		.INIT('h56)
	) name11322 (
		\u1_L11_reg[8]/NET0131 ,
		_w17139_,
		_w17148_,
		_w17149_
	);
	LUT4 #(
		.INIT('hbfd3)
	) name11323 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w17150_
	);
	LUT3 #(
		.INIT('h90)
	) name11324 (
		_w16838_,
		_w16837_,
		_w16836_,
		_w17151_
	);
	LUT3 #(
		.INIT('hb0)
	) name11325 (
		_w16838_,
		_w16839_,
		_w16841_,
		_w17152_
	);
	LUT4 #(
		.INIT('h00f1)
	) name11326 (
		_w16838_,
		_w16839_,
		_w16836_,
		_w16841_,
		_w17153_
	);
	LUT4 #(
		.INIT('h2700)
	) name11327 (
		_w17151_,
		_w17152_,
		_w17153_,
		_w17150_,
		_w17154_
	);
	LUT2 #(
		.INIT('h2)
	) name11328 (
		_w16835_,
		_w17154_,
		_w17155_
	);
	LUT4 #(
		.INIT('hef00)
	) name11329 (
		_w16837_,
		_w16839_,
		_w16836_,
		_w16841_,
		_w17156_
	);
	LUT4 #(
		.INIT('h2f33)
	) name11330 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w17157_
	);
	LUT2 #(
		.INIT('h8)
	) name11331 (
		_w17156_,
		_w17157_,
		_w17158_
	);
	LUT4 #(
		.INIT('h0080)
	) name11332 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16841_,
		_w17159_
	);
	LUT3 #(
		.INIT('h01)
	) name11333 (
		_w16859_,
		_w16997_,
		_w17159_,
		_w17160_
	);
	LUT3 #(
		.INIT('h45)
	) name11334 (
		_w16835_,
		_w17158_,
		_w17160_,
		_w17161_
	);
	LUT4 #(
		.INIT('heff7)
	) name11335 (
		_w16838_,
		_w16837_,
		_w16839_,
		_w16836_,
		_w17162_
	);
	LUT2 #(
		.INIT('h1)
	) name11336 (
		_w16841_,
		_w17162_,
		_w17163_
	);
	LUT4 #(
		.INIT('h0400)
	) name11337 (
		_w16837_,
		_w16839_,
		_w16836_,
		_w16841_,
		_w17164_
	);
	LUT3 #(
		.INIT('h07)
	) name11338 (
		_w16855_,
		_w16842_,
		_w17164_,
		_w17165_
	);
	LUT2 #(
		.INIT('h4)
	) name11339 (
		_w17163_,
		_w17165_,
		_w17166_
	);
	LUT4 #(
		.INIT('h5655)
	) name11340 (
		\u1_L11_reg[27]/NET0131 ,
		_w17155_,
		_w17161_,
		_w17166_,
		_w17167_
	);
	LUT3 #(
		.INIT('h40)
	) name11341 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w17168_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name11342 (
		_w16754_,
		_w16756_,
		_w16753_,
		_w16755_,
		_w17169_
	);
	LUT4 #(
		.INIT('hddd8)
	) name11343 (
		_w16753_,
		_w16766_,
		_w16758_,
		_w17168_,
		_w17170_
	);
	LUT4 #(
		.INIT('ha205)
	) name11344 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w17171_
	);
	LUT4 #(
		.INIT('h54a8)
	) name11345 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w17172_
	);
	LUT3 #(
		.INIT('h01)
	) name11346 (
		_w16753_,
		_w17171_,
		_w17172_,
		_w17173_
	);
	LUT3 #(
		.INIT('h8c)
	) name11347 (
		_w16756_,
		_w16755_,
		_w16757_,
		_w17174_
	);
	LUT2 #(
		.INIT('h2)
	) name11348 (
		_w16938_,
		_w17174_,
		_w17175_
	);
	LUT2 #(
		.INIT('h1)
	) name11349 (
		_w16753_,
		_w16755_,
		_w17176_
	);
	LUT3 #(
		.INIT('h08)
	) name11350 (
		_w16754_,
		_w16756_,
		_w16757_,
		_w17177_
	);
	LUT3 #(
		.INIT('h8a)
	) name11351 (
		_w16767_,
		_w17176_,
		_w17177_,
		_w17178_
	);
	LUT3 #(
		.INIT('h10)
	) name11352 (
		_w17175_,
		_w17173_,
		_w17178_,
		_w17179_
	);
	LUT4 #(
		.INIT('h5303)
	) name11353 (
		_w16756_,
		_w16753_,
		_w16755_,
		_w16757_,
		_w17180_
	);
	LUT2 #(
		.INIT('h2)
	) name11354 (
		_w16931_,
		_w17180_,
		_w17181_
	);
	LUT3 #(
		.INIT('h02)
	) name11355 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w17182_
	);
	LUT4 #(
		.INIT('h2202)
	) name11356 (
		_w16779_,
		_w16767_,
		_w16934_,
		_w17182_,
		_w17183_
	);
	LUT2 #(
		.INIT('h4)
	) name11357 (
		_w17181_,
		_w17183_,
		_w17184_
	);
	LUT4 #(
		.INIT('h6665)
	) name11358 (
		\u1_L11_reg[32]/NET0131 ,
		_w17170_,
		_w17179_,
		_w17184_,
		_w17185_
	);
	LUT4 #(
		.INIT('h0002)
	) name11359 (
		_w17059_,
		_w17069_,
		_w17104_,
		_w17135_,
		_w17186_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name11360 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17187_
	);
	LUT3 #(
		.INIT('h0e)
	) name11361 (
		_w17048_,
		_w17049_,
		_w17059_,
		_w17188_
	);
	LUT2 #(
		.INIT('h4)
	) name11362 (
		_w17187_,
		_w17188_,
		_w17189_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name11363 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17190_
	);
	LUT3 #(
		.INIT('h10)
	) name11364 (
		_w17046_,
		_w17098_,
		_w17190_,
		_w17191_
	);
	LUT3 #(
		.INIT('he0)
	) name11365 (
		_w17186_,
		_w17189_,
		_w17191_,
		_w17192_
	);
	LUT4 #(
		.INIT('h00df)
	) name11366 (
		_w17047_,
		_w17048_,
		_w17049_,
		_w17059_,
		_w17193_
	);
	LUT4 #(
		.INIT('hbf8b)
	) name11367 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17194_
	);
	LUT2 #(
		.INIT('h8)
	) name11368 (
		_w17193_,
		_w17194_,
		_w17195_
	);
	LUT4 #(
		.INIT('hcff5)
	) name11369 (
		_w17047_,
		_w17051_,
		_w17048_,
		_w17049_,
		_w17196_
	);
	LUT4 #(
		.INIT('h0200)
	) name11370 (
		_w17059_,
		_w17069_,
		_w17135_,
		_w17196_,
		_w17197_
	);
	LUT3 #(
		.INIT('h02)
	) name11371 (
		_w17046_,
		_w17094_,
		_w17114_,
		_w17198_
	);
	LUT3 #(
		.INIT('he0)
	) name11372 (
		_w17195_,
		_w17197_,
		_w17198_,
		_w17199_
	);
	LUT3 #(
		.INIT('ha9)
	) name11373 (
		\u1_L11_reg[3]/NET0131 ,
		_w17192_,
		_w17199_,
		_w17200_
	);
	LUT4 #(
		.INIT('hc963)
	) name11374 (
		decrypt_pad,
		\u1_R11_reg[11]/NET0131 ,
		\u1_uk_K_r11_reg[12]/NET0131 ,
		\u1_uk_K_r11_reg[17]/NET0131 ,
		_w17201_
	);
	LUT4 #(
		.INIT('hc963)
	) name11375 (
		decrypt_pad,
		\u1_R11_reg[12]/NET0131 ,
		\u1_uk_K_r11_reg[27]/P0001 ,
		\u1_uk_K_r11_reg[32]/NET0131 ,
		_w17202_
	);
	LUT4 #(
		.INIT('hc693)
	) name11376 (
		decrypt_pad,
		\u1_R11_reg[13]/NET0131 ,
		\u1_uk_K_r11_reg[20]/NET0131 ,
		\u1_uk_K_r11_reg[40]/NET0131 ,
		_w17203_
	);
	LUT4 #(
		.INIT('hc963)
	) name11377 (
		decrypt_pad,
		\u1_R11_reg[9]/NET0131 ,
		\u1_uk_K_r11_reg[3]/NET0131 ,
		\u1_uk_K_r11_reg[40]/NET0131 ,
		_w17204_
	);
	LUT4 #(
		.INIT('hc963)
	) name11378 (
		decrypt_pad,
		\u1_R11_reg[10]/NET0131 ,
		\u1_uk_K_r11_reg[11]/NET0131 ,
		\u1_uk_K_r11_reg[48]/NET0131 ,
		_w17205_
	);
	LUT4 #(
		.INIT('hc693)
	) name11379 (
		decrypt_pad,
		\u1_R11_reg[8]/NET0131 ,
		\u1_uk_K_r11_reg[11]/NET0131 ,
		\u1_uk_K_r11_reg[6]/NET0131 ,
		_w17206_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name11380 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17207_
	);
	LUT4 #(
		.INIT('h95b5)
	) name11381 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17208_
	);
	LUT2 #(
		.INIT('h1)
	) name11382 (
		_w17203_,
		_w17206_,
		_w17209_
	);
	LUT4 #(
		.INIT('h0001)
	) name11383 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17210_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name11384 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17211_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11385 (
		_w17202_,
		_w17201_,
		_w17208_,
		_w17211_,
		_w17212_
	);
	LUT2 #(
		.INIT('h6)
	) name11386 (
		_w17204_,
		_w17205_,
		_w17213_
	);
	LUT2 #(
		.INIT('h8)
	) name11387 (
		_w17203_,
		_w17206_,
		_w17214_
	);
	LUT3 #(
		.INIT('h46)
	) name11388 (
		_w17203_,
		_w17206_,
		_w17201_,
		_w17215_
	);
	LUT2 #(
		.INIT('h1)
	) name11389 (
		_w17213_,
		_w17215_,
		_w17216_
	);
	LUT3 #(
		.INIT('h40)
	) name11390 (
		_w17206_,
		_w17204_,
		_w17201_,
		_w17217_
	);
	LUT4 #(
		.INIT('h0660)
	) name11391 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17218_
	);
	LUT3 #(
		.INIT('h45)
	) name11392 (
		_w17202_,
		_w17217_,
		_w17218_,
		_w17219_
	);
	LUT3 #(
		.INIT('h80)
	) name11393 (
		_w17204_,
		_w17205_,
		_w17202_,
		_w17220_
	);
	LUT2 #(
		.INIT('h8)
	) name11394 (
		_w17209_,
		_w17220_,
		_w17221_
	);
	LUT3 #(
		.INIT('h0b)
	) name11395 (
		_w17203_,
		_w17204_,
		_w17201_,
		_w17222_
	);
	LUT3 #(
		.INIT('h51)
	) name11396 (
		_w17206_,
		_w17204_,
		_w17205_,
		_w17223_
	);
	LUT3 #(
		.INIT('hd0)
	) name11397 (
		_w17203_,
		_w17204_,
		_w17202_,
		_w17224_
	);
	LUT3 #(
		.INIT('h40)
	) name11398 (
		_w17223_,
		_w17222_,
		_w17224_,
		_w17225_
	);
	LUT4 #(
		.INIT('h1011)
	) name11399 (
		_w17221_,
		_w17225_,
		_w17216_,
		_w17219_,
		_w17226_
	);
	LUT3 #(
		.INIT('h65)
	) name11400 (
		\u1_L11_reg[6]/NET0131 ,
		_w17212_,
		_w17226_,
		_w17227_
	);
	LUT3 #(
		.INIT('h48)
	) name11401 (
		_w16754_,
		_w16755_,
		_w16757_,
		_w17228_
	);
	LUT4 #(
		.INIT('h4080)
	) name11402 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w17229_
	);
	LUT3 #(
		.INIT('h21)
	) name11403 (
		_w16754_,
		_w16756_,
		_w16757_,
		_w17230_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name11404 (
		_w16754_,
		_w16753_,
		_w16755_,
		_w16757_,
		_w17231_
	);
	LUT4 #(
		.INIT('h5455)
	) name11405 (
		_w16767_,
		_w17230_,
		_w17229_,
		_w17231_,
		_w17232_
	);
	LUT4 #(
		.INIT('h2210)
	) name11406 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w17233_
	);
	LUT2 #(
		.INIT('h2)
	) name11407 (
		_w16753_,
		_w17233_,
		_w17234_
	);
	LUT3 #(
		.INIT('h04)
	) name11408 (
		_w16932_,
		_w17169_,
		_w17228_,
		_w17235_
	);
	LUT4 #(
		.INIT('h4880)
	) name11409 (
		_w16754_,
		_w16756_,
		_w16755_,
		_w16757_,
		_w17236_
	);
	LUT2 #(
		.INIT('h2)
	) name11410 (
		_w16767_,
		_w17236_,
		_w17237_
	);
	LUT4 #(
		.INIT('h0155)
	) name11411 (
		_w17232_,
		_w17234_,
		_w17235_,
		_w17237_,
		_w17238_
	);
	LUT2 #(
		.INIT('h4)
	) name11412 (
		_w16753_,
		_w17236_,
		_w17239_
	);
	LUT2 #(
		.INIT('h4)
	) name11413 (
		_w16753_,
		_w16767_,
		_w17240_
	);
	LUT4 #(
		.INIT('h00dc)
	) name11414 (
		_w16753_,
		_w16773_,
		_w17233_,
		_w17240_,
		_w17241_
	);
	LUT2 #(
		.INIT('h1)
	) name11415 (
		_w17239_,
		_w17241_,
		_w17242_
	);
	LUT3 #(
		.INIT('h65)
	) name11416 (
		\u1_L11_reg[7]/NET0131 ,
		_w17238_,
		_w17242_,
		_w17243_
	);
	LUT4 #(
		.INIT('h8448)
	) name11417 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w17244_
	);
	LUT3 #(
		.INIT('h19)
	) name11418 (
		_w16682_,
		_w16683_,
		_w16685_,
		_w17245_
	);
	LUT3 #(
		.INIT('h10)
	) name11419 (
		_w16684_,
		_w16683_,
		_w16685_,
		_w17246_
	);
	LUT4 #(
		.INIT('h0200)
	) name11420 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w17247_
	);
	LUT4 #(
		.INIT('h0007)
	) name11421 (
		_w16690_,
		_w17245_,
		_w17244_,
		_w17247_,
		_w17248_
	);
	LUT3 #(
		.INIT('h28)
	) name11422 (
		_w16681_,
		_w16682_,
		_w16683_,
		_w17249_
	);
	LUT4 #(
		.INIT('h0141)
	) name11423 (
		_w16681_,
		_w16682_,
		_w16683_,
		_w16685_,
		_w17250_
	);
	LUT4 #(
		.INIT('h9ffb)
	) name11424 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w17251_
	);
	LUT4 #(
		.INIT('h4500)
	) name11425 (
		_w17250_,
		_w17246_,
		_w17249_,
		_w17251_,
		_w17252_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name11426 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w17253_
	);
	LUT2 #(
		.INIT('h1)
	) name11427 (
		_w16681_,
		_w17253_,
		_w17254_
	);
	LUT4 #(
		.INIT('h0e04)
	) name11428 (
		_w16693_,
		_w17252_,
		_w17254_,
		_w17248_,
		_w17255_
	);
	LUT2 #(
		.INIT('h9)
	) name11429 (
		\u1_L11_reg[9]/NET0131 ,
		_w17255_,
		_w17256_
	);
	LUT3 #(
		.INIT('h80)
	) name11430 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17257_
	);
	LUT4 #(
		.INIT('h6979)
	) name11431 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17201_,
		_w17258_
	);
	LUT2 #(
		.INIT('h1)
	) name11432 (
		_w17205_,
		_w17258_,
		_w17259_
	);
	LUT4 #(
		.INIT('h0014)
	) name11433 (
		_w17203_,
		_w17206_,
		_w17205_,
		_w17201_,
		_w17260_
	);
	LUT4 #(
		.INIT('h2000)
	) name11434 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17261_
	);
	LUT3 #(
		.INIT('h02)
	) name11435 (
		_w17202_,
		_w17260_,
		_w17261_,
		_w17262_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name11436 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17263_
	);
	LUT2 #(
		.INIT('h1)
	) name11437 (
		_w17201_,
		_w17263_,
		_w17264_
	);
	LUT4 #(
		.INIT('h6800)
	) name11438 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17201_,
		_w17265_
	);
	LUT3 #(
		.INIT('h01)
	) name11439 (
		_w17202_,
		_w17210_,
		_w17265_,
		_w17266_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name11440 (
		_w17259_,
		_w17262_,
		_w17264_,
		_w17266_,
		_w17267_
	);
	LUT4 #(
		.INIT('h4100)
	) name11441 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17268_
	);
	LUT2 #(
		.INIT('h8)
	) name11442 (
		_w17206_,
		_w17205_,
		_w17269_
	);
	LUT4 #(
		.INIT('h00df)
	) name11443 (
		_w17206_,
		_w17204_,
		_w17205_,
		_w17201_,
		_w17270_
	);
	LUT3 #(
		.INIT('h0d)
	) name11444 (
		_w17201_,
		_w17268_,
		_w17270_,
		_w17271_
	);
	LUT3 #(
		.INIT('h56)
	) name11445 (
		\u1_L11_reg[16]/NET0131 ,
		_w17267_,
		_w17271_,
		_w17272_
	);
	LUT4 #(
		.INIT('h6660)
	) name11446 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17273_
	);
	LUT4 #(
		.INIT('h0009)
	) name11447 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17274_
	);
	LUT4 #(
		.INIT('h551b)
	) name11448 (
		_w17202_,
		_w17207_,
		_w17273_,
		_w17274_,
		_w17275_
	);
	LUT4 #(
		.INIT('h1df2)
	) name11449 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17276_
	);
	LUT2 #(
		.INIT('h2)
	) name11450 (
		_w17202_,
		_w17276_,
		_w17277_
	);
	LUT4 #(
		.INIT('h0020)
	) name11451 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17278_
	);
	LUT4 #(
		.INIT('h0004)
	) name11452 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17279_
	);
	LUT3 #(
		.INIT('h02)
	) name11453 (
		_w17201_,
		_w17278_,
		_w17279_,
		_w17280_
	);
	LUT4 #(
		.INIT('he0ee)
	) name11454 (
		_w17201_,
		_w17275_,
		_w17277_,
		_w17280_,
		_w17281_
	);
	LUT2 #(
		.INIT('h2)
	) name11455 (
		_w17205_,
		_w17201_,
		_w17282_
	);
	LUT2 #(
		.INIT('h8)
	) name11456 (
		_w17257_,
		_w17282_,
		_w17283_
	);
	LUT4 #(
		.INIT('h0400)
	) name11457 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17284_
	);
	LUT3 #(
		.INIT('hed)
	) name11458 (
		_w17203_,
		_w17206_,
		_w17205_,
		_w17285_
	);
	LUT3 #(
		.INIT('h10)
	) name11459 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17286_
	);
	LUT4 #(
		.INIT('he2cd)
	) name11460 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17287_
	);
	LUT4 #(
		.INIT('h5054)
	) name11461 (
		_w17202_,
		_w17201_,
		_w17284_,
		_w17287_,
		_w17288_
	);
	LUT2 #(
		.INIT('h1)
	) name11462 (
		_w17283_,
		_w17288_,
		_w17289_
	);
	LUT3 #(
		.INIT('h65)
	) name11463 (
		\u1_L11_reg[24]/NET0131 ,
		_w17281_,
		_w17289_,
		_w17290_
	);
	LUT3 #(
		.INIT('h20)
	) name11464 (
		_w17201_,
		_w17279_,
		_w17285_,
		_w17291_
	);
	LUT3 #(
		.INIT('h07)
	) name11465 (
		_w17206_,
		_w17205_,
		_w17201_,
		_w17292_
	);
	LUT2 #(
		.INIT('h4)
	) name11466 (
		_w17286_,
		_w17292_,
		_w17293_
	);
	LUT3 #(
		.INIT('ha8)
	) name11467 (
		_w17202_,
		_w17291_,
		_w17293_,
		_w17294_
	);
	LUT4 #(
		.INIT('hdd02)
	) name11468 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17295_
	);
	LUT4 #(
		.INIT('hf450)
	) name11469 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17201_,
		_w17296_
	);
	LUT2 #(
		.INIT('h1)
	) name11470 (
		_w17295_,
		_w17296_,
		_w17297_
	);
	LUT4 #(
		.INIT('h73af)
	) name11471 (
		_w17203_,
		_w17206_,
		_w17204_,
		_w17205_,
		_w17298_
	);
	LUT3 #(
		.INIT('h51)
	) name11472 (
		_w17202_,
		_w17201_,
		_w17298_,
		_w17299_
	);
	LUT2 #(
		.INIT('h4)
	) name11473 (
		_w17297_,
		_w17299_,
		_w17300_
	);
	LUT3 #(
		.INIT('h20)
	) name11474 (
		_w17203_,
		_w17204_,
		_w17201_,
		_w17301_
	);
	LUT2 #(
		.INIT('h8)
	) name11475 (
		_w17269_,
		_w17301_,
		_w17302_
	);
	LUT4 #(
		.INIT('h0040)
	) name11476 (
		_w17203_,
		_w17204_,
		_w17205_,
		_w17201_,
		_w17303_
	);
	LUT3 #(
		.INIT('h0d)
	) name11477 (
		_w17220_,
		_w17214_,
		_w17303_,
		_w17304_
	);
	LUT2 #(
		.INIT('h4)
	) name11478 (
		_w17302_,
		_w17304_,
		_w17305_
	);
	LUT4 #(
		.INIT('h56aa)
	) name11479 (
		\u1_L11_reg[30]/NET0131 ,
		_w17294_,
		_w17300_,
		_w17305_,
		_w17306_
	);
	LUT4 #(
		.INIT('hbefe)
	) name11480 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w17307_
	);
	LUT3 #(
		.INIT('h53)
	) name11481 (
		_w16886_,
		_w16879_,
		_w16881_,
		_w17308_
	);
	LUT4 #(
		.INIT('h0043)
	) name11482 (
		_w16886_,
		_w16879_,
		_w16881_,
		_w16883_,
		_w17309_
	);
	LUT4 #(
		.INIT('h0d00)
	) name11483 (
		_w16896_,
		_w17308_,
		_w17309_,
		_w17307_,
		_w17310_
	);
	LUT4 #(
		.INIT('h2028)
	) name11484 (
		_w16886_,
		_w16880_,
		_w16881_,
		_w16883_,
		_w17311_
	);
	LUT3 #(
		.INIT('hd8)
	) name11485 (
		_w16880_,
		_w16879_,
		_w16881_,
		_w17312_
	);
	LUT2 #(
		.INIT('h4)
	) name11486 (
		_w16886_,
		_w16883_,
		_w17313_
	);
	LUT4 #(
		.INIT('h1011)
	) name11487 (
		_w16907_,
		_w17311_,
		_w17312_,
		_w17313_,
		_w17314_
	);
	LUT3 #(
		.INIT('h80)
	) name11488 (
		_w16880_,
		_w16879_,
		_w16883_,
		_w17315_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name11489 (
		_w16886_,
		_w16955_,
		_w17078_,
		_w17315_,
		_w17316_
	);
	LUT4 #(
		.INIT('h0d08)
	) name11490 (
		_w16888_,
		_w17314_,
		_w17316_,
		_w17310_,
		_w17317_
	);
	LUT2 #(
		.INIT('h9)
	) name11491 (
		\u1_L11_reg[18]/P0001 ,
		_w17317_,
		_w17318_
	);
	LUT4 #(
		.INIT('hc963)
	) name11492 (
		decrypt_pad,
		\u1_R10_reg[28]/NET0131 ,
		\u1_uk_K_r10_reg[36]/NET0131 ,
		\u1_uk_K_r10_reg[45]/P0001 ,
		_w17319_
	);
	LUT4 #(
		.INIT('hc963)
	) name11493 (
		decrypt_pad,
		\u1_R10_reg[26]/NET0131 ,
		\u1_uk_K_r10_reg[16]/NET0131 ,
		\u1_uk_K_r10_reg[21]/NET0131 ,
		_w17320_
	);
	LUT4 #(
		.INIT('hc963)
	) name11494 (
		decrypt_pad,
		\u1_R10_reg[25]/NET0131 ,
		\u1_uk_K_r10_reg[0]/NET0131 ,
		\u1_uk_K_r10_reg[36]/NET0131 ,
		_w17321_
	);
	LUT4 #(
		.INIT('hc963)
	) name11495 (
		decrypt_pad,
		\u1_R10_reg[29]/NET0131 ,
		\u1_uk_K_r10_reg[28]/NET0131 ,
		\u1_uk_K_r10_reg[9]/NET0131 ,
		_w17322_
	);
	LUT3 #(
		.INIT('hea)
	) name11496 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17323_
	);
	LUT4 #(
		.INIT('hc693)
	) name11497 (
		decrypt_pad,
		\u1_R10_reg[24]/NET0131 ,
		\u1_uk_K_r10_reg[1]/NET0131 ,
		\u1_uk_K_r10_reg[51]/NET0131 ,
		_w17324_
	);
	LUT4 #(
		.INIT('hc693)
	) name11498 (
		decrypt_pad,
		\u1_R10_reg[27]/NET0131 ,
		\u1_uk_K_r10_reg[30]/NET0131 ,
		\u1_uk_K_r10_reg[49]/NET0131 ,
		_w17325_
	);
	LUT3 #(
		.INIT('h70)
	) name11499 (
		_w17320_,
		_w17321_,
		_w17325_,
		_w17326_
	);
	LUT4 #(
		.INIT('h7000)
	) name11500 (
		_w17320_,
		_w17321_,
		_w17324_,
		_w17325_,
		_w17327_
	);
	LUT2 #(
		.INIT('h8)
	) name11501 (
		_w17323_,
		_w17327_,
		_w17328_
	);
	LUT4 #(
		.INIT('h1000)
	) name11502 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17329_
	);
	LUT4 #(
		.INIT('hef3f)
	) name11503 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17330_
	);
	LUT2 #(
		.INIT('h2)
	) name11504 (
		_w17322_,
		_w17324_,
		_w17331_
	);
	LUT4 #(
		.INIT('h0020)
	) name11505 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17332_
	);
	LUT4 #(
		.INIT('hffde)
	) name11506 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17333_
	);
	LUT3 #(
		.INIT('he0)
	) name11507 (
		_w17325_,
		_w17330_,
		_w17333_,
		_w17334_
	);
	LUT3 #(
		.INIT('h8a)
	) name11508 (
		_w17319_,
		_w17328_,
		_w17334_,
		_w17335_
	);
	LUT4 #(
		.INIT('h0072)
	) name11509 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17325_,
		_w17336_
	);
	LUT4 #(
		.INIT('h10f0)
	) name11510 (
		_w17320_,
		_w17321_,
		_w17324_,
		_w17325_,
		_w17337_
	);
	LUT2 #(
		.INIT('h4)
	) name11511 (
		_w17336_,
		_w17337_,
		_w17338_
	);
	LUT4 #(
		.INIT('h0002)
	) name11512 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17339_
	);
	LUT2 #(
		.INIT('h6)
	) name11513 (
		_w17320_,
		_w17324_,
		_w17340_
	);
	LUT3 #(
		.INIT('h8c)
	) name11514 (
		_w17321_,
		_w17322_,
		_w17325_,
		_w17341_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name11515 (
		_w17339_,
		_w17325_,
		_w17340_,
		_w17341_,
		_w17342_
	);
	LUT4 #(
		.INIT('h0008)
	) name11516 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17343_
	);
	LUT4 #(
		.INIT('hfcd7)
	) name11517 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17344_
	);
	LUT4 #(
		.INIT('h0084)
	) name11518 (
		_w17320_,
		_w17321_,
		_w17324_,
		_w17325_,
		_w17345_
	);
	LUT4 #(
		.INIT('h0100)
	) name11519 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17325_,
		_w17346_
	);
	LUT4 #(
		.INIT('h0031)
	) name11520 (
		_w17325_,
		_w17345_,
		_w17344_,
		_w17346_,
		_w17347_
	);
	LUT4 #(
		.INIT('hba00)
	) name11521 (
		_w17319_,
		_w17338_,
		_w17342_,
		_w17347_,
		_w17348_
	);
	LUT3 #(
		.INIT('h65)
	) name11522 (
		\u1_L10_reg[22]/NET0131 ,
		_w17335_,
		_w17348_,
		_w17349_
	);
	LUT4 #(
		.INIT('hc963)
	) name11523 (
		decrypt_pad,
		\u1_R10_reg[3]/NET0131 ,
		\u1_uk_K_r10_reg[27]/NET0131 ,
		\u1_uk_K_r10_reg[4]/NET0131 ,
		_w17350_
	);
	LUT4 #(
		.INIT('hc693)
	) name11524 (
		decrypt_pad,
		\u1_R10_reg[1]/NET0131 ,
		\u1_uk_K_r10_reg[12]/NET0131 ,
		\u1_uk_K_r10_reg[3]/NET0131 ,
		_w17351_
	);
	LUT4 #(
		.INIT('hc963)
	) name11525 (
		decrypt_pad,
		\u1_R10_reg[32]/NET0131 ,
		\u1_uk_K_r10_reg[39]/NET0131 ,
		\u1_uk_K_r10_reg[48]/NET0131 ,
		_w17352_
	);
	LUT4 #(
		.INIT('hc693)
	) name11526 (
		decrypt_pad,
		\u1_R10_reg[5]/NET0131 ,
		\u1_uk_K_r10_reg[10]/NET0131 ,
		\u1_uk_K_r10_reg[33]/NET0131 ,
		_w17353_
	);
	LUT4 #(
		.INIT('hc963)
	) name11527 (
		decrypt_pad,
		\u1_R10_reg[2]/NET0131 ,
		\u1_uk_K_r10_reg[18]/NET0131 ,
		\u1_uk_K_r10_reg[27]/NET0131 ,
		_w17354_
	);
	LUT4 #(
		.INIT('h4000)
	) name11528 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17355_
	);
	LUT2 #(
		.INIT('h8)
	) name11529 (
		_w17350_,
		_w17355_,
		_w17356_
	);
	LUT4 #(
		.INIT('hc693)
	) name11530 (
		decrypt_pad,
		\u1_R10_reg[4]/NET0131 ,
		\u1_uk_K_r10_reg[39]/NET0131 ,
		\u1_uk_K_r10_reg[5]/NET0131 ,
		_w17357_
	);
	LUT4 #(
		.INIT('h0080)
	) name11531 (
		_w17353_,
		_w17354_,
		_w17350_,
		_w17352_,
		_w17358_
	);
	LUT3 #(
		.INIT('h13)
	) name11532 (
		_w17351_,
		_w17357_,
		_w17358_,
		_w17359_
	);
	LUT2 #(
		.INIT('h9)
	) name11533 (
		_w17354_,
		_w17352_,
		_w17360_
	);
	LUT4 #(
		.INIT('h010d)
	) name11534 (
		_w17353_,
		_w17351_,
		_w17350_,
		_w17352_,
		_w17361_
	);
	LUT4 #(
		.INIT('h5dbb)
	) name11535 (
		_w17353_,
		_w17351_,
		_w17350_,
		_w17352_,
		_w17362_
	);
	LUT4 #(
		.INIT('h6f2a)
	) name11536 (
		_w17354_,
		_w17352_,
		_w17361_,
		_w17362_,
		_w17363_
	);
	LUT4 #(
		.INIT('h4e11)
	) name11537 (
		_w17353_,
		_w17354_,
		_w17350_,
		_w17352_,
		_w17364_
	);
	LUT2 #(
		.INIT('h2)
	) name11538 (
		_w17350_,
		_w17352_,
		_w17365_
	);
	LUT4 #(
		.INIT('h0060)
	) name11539 (
		_w17353_,
		_w17354_,
		_w17350_,
		_w17352_,
		_w17366_
	);
	LUT4 #(
		.INIT('h0c08)
	) name11540 (
		_w17351_,
		_w17357_,
		_w17366_,
		_w17364_,
		_w17367_
	);
	LUT4 #(
		.INIT('h00bf)
	) name11541 (
		_w17356_,
		_w17359_,
		_w17363_,
		_w17367_,
		_w17368_
	);
	LUT4 #(
		.INIT('h8000)
	) name11542 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17369_
	);
	LUT3 #(
		.INIT('h04)
	) name11543 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17370_
	);
	LUT4 #(
		.INIT('h0020)
	) name11544 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17371_
	);
	LUT3 #(
		.INIT('h80)
	) name11545 (
		_w17351_,
		_w17352_,
		_w17357_,
		_w17372_
	);
	LUT4 #(
		.INIT('h0001)
	) name11546 (
		_w17371_,
		_w17369_,
		_w17372_,
		_w17370_,
		_w17373_
	);
	LUT3 #(
		.INIT('h10)
	) name11547 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17374_
	);
	LUT4 #(
		.INIT('h1000)
	) name11548 (
		_w17351_,
		_w17354_,
		_w17350_,
		_w17352_,
		_w17375_
	);
	LUT3 #(
		.INIT('h07)
	) name11549 (
		_w17365_,
		_w17374_,
		_w17375_,
		_w17376_
	);
	LUT3 #(
		.INIT('he0)
	) name11550 (
		_w17350_,
		_w17373_,
		_w17376_,
		_w17377_
	);
	LUT3 #(
		.INIT('h65)
	) name11551 (
		\u1_L10_reg[31]/NET0131 ,
		_w17368_,
		_w17377_,
		_w17378_
	);
	LUT4 #(
		.INIT('hc963)
	) name11552 (
		decrypt_pad,
		\u1_R10_reg[24]/NET0131 ,
		\u1_uk_K_r10_reg[29]/NET0131 ,
		\u1_uk_K_r10_reg[38]/NET0131 ,
		_w17379_
	);
	LUT4 #(
		.INIT('hc963)
	) name11553 (
		decrypt_pad,
		\u1_R10_reg[22]/NET0131 ,
		\u1_uk_K_r10_reg[14]/NET0131 ,
		\u1_uk_K_r10_reg[50]/NET0131 ,
		_w17380_
	);
	LUT4 #(
		.INIT('hc963)
	) name11554 (
		decrypt_pad,
		\u1_R10_reg[21]/NET0131 ,
		\u1_uk_K_r10_reg[23]/NET0131 ,
		\u1_uk_K_r10_reg[28]/NET0131 ,
		_w17381_
	);
	LUT4 #(
		.INIT('hc693)
	) name11555 (
		decrypt_pad,
		\u1_R10_reg[20]/NET0131 ,
		\u1_uk_K_r10_reg[44]/NET0131 ,
		\u1_uk_K_r10_reg[8]/NET0131 ,
		_w17382_
	);
	LUT4 #(
		.INIT('hc693)
	) name11556 (
		decrypt_pad,
		\u1_R10_reg[25]/NET0131 ,
		\u1_uk_K_r10_reg[29]/NET0131 ,
		\u1_uk_K_r10_reg[52]/NET0131 ,
		_w17383_
	);
	LUT4 #(
		.INIT('he020)
	) name11557 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17384_
	);
	LUT4 #(
		.INIT('hc963)
	) name11558 (
		decrypt_pad,
		\u1_R10_reg[23]/NET0131 ,
		\u1_uk_K_r10_reg[31]/NET0131 ,
		\u1_uk_K_r10_reg[8]/NET0131 ,
		_w17385_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name11559 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17386_
	);
	LUT3 #(
		.INIT('h01)
	) name11560 (
		_w17385_,
		_w17386_,
		_w17384_,
		_w17387_
	);
	LUT2 #(
		.INIT('h2)
	) name11561 (
		_w17382_,
		_w17383_,
		_w17388_
	);
	LUT2 #(
		.INIT('h1)
	) name11562 (
		_w17381_,
		_w17380_,
		_w17389_
	);
	LUT4 #(
		.INIT('h0004)
	) name11563 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17390_
	);
	LUT4 #(
		.INIT('h57db)
	) name11564 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17391_
	);
	LUT2 #(
		.INIT('h1)
	) name11565 (
		_w17380_,
		_w17385_,
		_w17392_
	);
	LUT4 #(
		.INIT('h0200)
	) name11566 (
		_w17382_,
		_w17380_,
		_w17385_,
		_w17383_,
		_w17393_
	);
	LUT2 #(
		.INIT('h4)
	) name11567 (
		_w17381_,
		_w17393_,
		_w17394_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name11568 (
		_w17381_,
		_w17385_,
		_w17391_,
		_w17393_,
		_w17395_
	);
	LUT3 #(
		.INIT('h8a)
	) name11569 (
		_w17379_,
		_w17387_,
		_w17395_,
		_w17396_
	);
	LUT4 #(
		.INIT('h0010)
	) name11570 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17397_
	);
	LUT3 #(
		.INIT('hac)
	) name11571 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17398_
	);
	LUT4 #(
		.INIT('h5300)
	) name11572 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17385_,
		_w17399_
	);
	LUT2 #(
		.INIT('h4)
	) name11573 (
		_w17397_,
		_w17399_,
		_w17400_
	);
	LUT4 #(
		.INIT('h0028)
	) name11574 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17385_,
		_w17401_
	);
	LUT3 #(
		.INIT('hdc)
	) name11575 (
		_w17381_,
		_w17380_,
		_w17385_,
		_w17402_
	);
	LUT4 #(
		.INIT('h4000)
	) name11576 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17403_
	);
	LUT4 #(
		.INIT('h0051)
	) name11577 (
		_w17401_,
		_w17388_,
		_w17402_,
		_w17403_,
		_w17404_
	);
	LUT3 #(
		.INIT('h45)
	) name11578 (
		_w17379_,
		_w17400_,
		_w17404_,
		_w17405_
	);
	LUT3 #(
		.INIT('h40)
	) name11579 (
		_w17382_,
		_w17385_,
		_w17383_,
		_w17406_
	);
	LUT2 #(
		.INIT('h2)
	) name11580 (
		_w17382_,
		_w17385_,
		_w17407_
	);
	LUT3 #(
		.INIT('h02)
	) name11581 (
		_w17381_,
		_w17380_,
		_w17383_,
		_w17408_
	);
	LUT4 #(
		.INIT('h0777)
	) name11582 (
		_w17389_,
		_w17406_,
		_w17407_,
		_w17408_,
		_w17409_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name11583 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17410_
	);
	LUT4 #(
		.INIT('hb030)
	) name11584 (
		_w17382_,
		_w17380_,
		_w17385_,
		_w17383_,
		_w17411_
	);
	LUT3 #(
		.INIT('h01)
	) name11585 (
		_w17381_,
		_w17382_,
		_w17383_,
		_w17412_
	);
	LUT4 #(
		.INIT('h45cf)
	) name11586 (
		_w17392_,
		_w17410_,
		_w17411_,
		_w17412_,
		_w17413_
	);
	LUT2 #(
		.INIT('h8)
	) name11587 (
		_w17409_,
		_w17413_,
		_w17414_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name11588 (
		\u1_L10_reg[11]/NET0131 ,
		_w17405_,
		_w17396_,
		_w17414_,
		_w17415_
	);
	LUT4 #(
		.INIT('hc693)
	) name11589 (
		decrypt_pad,
		\u1_R10_reg[13]/NET0131 ,
		\u1_uk_K_r10_reg[24]/NET0131 ,
		\u1_uk_K_r10_reg[47]/NET0131 ,
		_w17416_
	);
	LUT4 #(
		.INIT('hc963)
	) name11590 (
		decrypt_pad,
		\u1_R10_reg[12]/NET0131 ,
		\u1_uk_K_r10_reg[53]/NET0131 ,
		\u1_uk_K_r10_reg[5]/NET0131 ,
		_w17417_
	);
	LUT4 #(
		.INIT('hc963)
	) name11591 (
		decrypt_pad,
		\u1_R10_reg[17]/NET0131 ,
		\u1_uk_K_r10_reg[12]/NET0131 ,
		\u1_uk_K_r10_reg[46]/NET0131 ,
		_w17418_
	);
	LUT4 #(
		.INIT('hc963)
	) name11592 (
		decrypt_pad,
		\u1_R10_reg[15]/NET0131 ,
		\u1_uk_K_r10_reg[24]/NET0131 ,
		\u1_uk_K_r10_reg[33]/NET0131 ,
		_w17419_
	);
	LUT3 #(
		.INIT('h01)
	) name11593 (
		_w17417_,
		_w17416_,
		_w17418_,
		_w17420_
	);
	LUT4 #(
		.INIT('h2aa8)
	) name11594 (
		_w17419_,
		_w17417_,
		_w17416_,
		_w17418_,
		_w17421_
	);
	LUT4 #(
		.INIT('hc693)
	) name11595 (
		decrypt_pad,
		\u1_R10_reg[14]/NET0131 ,
		\u1_uk_K_r10_reg[25]/NET0131 ,
		\u1_uk_K_r10_reg[48]/NET0131 ,
		_w17422_
	);
	LUT3 #(
		.INIT('h08)
	) name11596 (
		_w17417_,
		_w17422_,
		_w17418_,
		_w17423_
	);
	LUT3 #(
		.INIT('h45)
	) name11597 (
		_w17419_,
		_w17416_,
		_w17418_,
		_w17424_
	);
	LUT3 #(
		.INIT('h45)
	) name11598 (
		_w17421_,
		_w17423_,
		_w17424_,
		_w17425_
	);
	LUT4 #(
		.INIT('h0001)
	) name11599 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17426_
	);
	LUT3 #(
		.INIT('h04)
	) name11600 (
		_w17417_,
		_w17416_,
		_w17418_,
		_w17427_
	);
	LUT4 #(
		.INIT('hffbe)
	) name11601 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17428_
	);
	LUT3 #(
		.INIT('h80)
	) name11602 (
		_w17419_,
		_w17416_,
		_w17422_,
		_w17429_
	);
	LUT4 #(
		.INIT('h2000)
	) name11603 (
		_w17419_,
		_w17417_,
		_w17416_,
		_w17422_,
		_w17430_
	);
	LUT4 #(
		.INIT('hc963)
	) name11604 (
		decrypt_pad,
		\u1_R10_reg[16]/NET0131 ,
		\u1_uk_K_r10_reg[32]/NET0131 ,
		\u1_uk_K_r10_reg[41]/P0001 ,
		_w17431_
	);
	LUT2 #(
		.INIT('h2)
	) name11605 (
		_w17417_,
		_w17416_,
		_w17432_
	);
	LUT4 #(
		.INIT('h0200)
	) name11606 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17433_
	);
	LUT4 #(
		.INIT('h0002)
	) name11607 (
		_w17428_,
		_w17431_,
		_w17430_,
		_w17433_,
		_w17434_
	);
	LUT2 #(
		.INIT('h4)
	) name11608 (
		_w17425_,
		_w17434_,
		_w17435_
	);
	LUT2 #(
		.INIT('h4)
	) name11609 (
		_w17417_,
		_w17418_,
		_w17436_
	);
	LUT4 #(
		.INIT('h0200)
	) name11610 (
		_w17419_,
		_w17417_,
		_w17416_,
		_w17418_,
		_w17437_
	);
	LUT2 #(
		.INIT('h2)
	) name11611 (
		_w17431_,
		_w17437_,
		_w17438_
	);
	LUT4 #(
		.INIT('h0400)
	) name11612 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17439_
	);
	LUT4 #(
		.INIT('h0080)
	) name11613 (
		_w17419_,
		_w17417_,
		_w17416_,
		_w17418_,
		_w17440_
	);
	LUT4 #(
		.INIT('h8000)
	) name11614 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17441_
	);
	LUT3 #(
		.INIT('h01)
	) name11615 (
		_w17439_,
		_w17440_,
		_w17441_,
		_w17442_
	);
	LUT2 #(
		.INIT('h9)
	) name11616 (
		_w17417_,
		_w17416_,
		_w17443_
	);
	LUT4 #(
		.INIT('h0014)
	) name11617 (
		_w17419_,
		_w17417_,
		_w17416_,
		_w17422_,
		_w17444_
	);
	LUT2 #(
		.INIT('h4)
	) name11618 (
		_w17419_,
		_w17422_,
		_w17445_
	);
	LUT3 #(
		.INIT('h13)
	) name11619 (
		_w17420_,
		_w17444_,
		_w17445_,
		_w17446_
	);
	LUT3 #(
		.INIT('h80)
	) name11620 (
		_w17438_,
		_w17442_,
		_w17446_,
		_w17447_
	);
	LUT4 #(
		.INIT('h0020)
	) name11621 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17448_
	);
	LUT4 #(
		.INIT('heee4)
	) name11622 (
		_w17419_,
		_w17439_,
		_w17448_,
		_w17426_,
		_w17449_
	);
	LUT2 #(
		.INIT('h4)
	) name11623 (
		_w17422_,
		_w17440_,
		_w17450_
	);
	LUT2 #(
		.INIT('h1)
	) name11624 (
		_w17449_,
		_w17450_,
		_w17451_
	);
	LUT4 #(
		.INIT('ha955)
	) name11625 (
		\u1_L10_reg[20]/NET0131 ,
		_w17435_,
		_w17447_,
		_w17451_,
		_w17452_
	);
	LUT4 #(
		.INIT('h6fff)
	) name11626 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17453_
	);
	LUT3 #(
		.INIT('h02)
	) name11627 (
		_w17419_,
		_w17427_,
		_w17433_,
		_w17454_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11628 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17455_
	);
	LUT3 #(
		.INIT('h01)
	) name11629 (
		_w17419_,
		_w17439_,
		_w17455_,
		_w17456_
	);
	LUT4 #(
		.INIT('h222a)
	) name11630 (
		_w17431_,
		_w17453_,
		_w17454_,
		_w17456_,
		_w17457_
	);
	LUT3 #(
		.INIT('h8a)
	) name11631 (
		_w17419_,
		_w17422_,
		_w17418_,
		_w17458_
	);
	LUT3 #(
		.INIT('h2a)
	) name11632 (
		_w17428_,
		_w17432_,
		_w17458_,
		_w17459_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name11633 (
		_w17419_,
		_w17417_,
		_w17416_,
		_w17418_,
		_w17460_
	);
	LUT4 #(
		.INIT('hf5ee)
	) name11634 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17461_
	);
	LUT4 #(
		.INIT('hfca8)
	) name11635 (
		_w17419_,
		_w17422_,
		_w17460_,
		_w17461_,
		_w17462_
	);
	LUT3 #(
		.INIT('h15)
	) name11636 (
		_w17431_,
		_w17459_,
		_w17462_,
		_w17463_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name11637 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17464_
	);
	LUT2 #(
		.INIT('h1)
	) name11638 (
		_w17419_,
		_w17464_,
		_w17465_
	);
	LUT3 #(
		.INIT('h0b)
	) name11639 (
		_w17422_,
		_w17440_,
		_w17430_,
		_w17466_
	);
	LUT2 #(
		.INIT('h4)
	) name11640 (
		_w17465_,
		_w17466_,
		_w17467_
	);
	LUT4 #(
		.INIT('h5655)
	) name11641 (
		\u1_L10_reg[10]/NET0131 ,
		_w17463_,
		_w17457_,
		_w17467_,
		_w17468_
	);
	LUT4 #(
		.INIT('h0006)
	) name11642 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17469_
	);
	LUT3 #(
		.INIT('h47)
	) name11643 (
		_w17320_,
		_w17321_,
		_w17325_,
		_w17470_
	);
	LUT4 #(
		.INIT('h0051)
	) name11644 (
		_w17319_,
		_w17331_,
		_w17470_,
		_w17469_,
		_w17471_
	);
	LUT3 #(
		.INIT('h10)
	) name11645 (
		_w17320_,
		_w17322_,
		_w17324_,
		_w17472_
	);
	LUT4 #(
		.INIT('h2100)
	) name11646 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17473_
	);
	LUT2 #(
		.INIT('h6)
	) name11647 (
		_w17321_,
		_w17322_,
		_w17474_
	);
	LUT4 #(
		.INIT('h143c)
	) name11648 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17475_
	);
	LUT3 #(
		.INIT('h32)
	) name11649 (
		_w17325_,
		_w17473_,
		_w17475_,
		_w17476_
	);
	LUT2 #(
		.INIT('h8)
	) name11650 (
		_w17471_,
		_w17476_,
		_w17477_
	);
	LUT2 #(
		.INIT('h4)
	) name11651 (
		_w17325_,
		_w17332_,
		_w17478_
	);
	LUT3 #(
		.INIT('h02)
	) name11652 (
		_w17319_,
		_w17329_,
		_w17343_,
		_w17479_
	);
	LUT4 #(
		.INIT('h0240)
	) name11653 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17480_
	);
	LUT4 #(
		.INIT('h33fe)
	) name11654 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17481_
	);
	LUT3 #(
		.INIT('h31)
	) name11655 (
		_w17325_,
		_w17480_,
		_w17481_,
		_w17482_
	);
	LUT3 #(
		.INIT('h40)
	) name11656 (
		_w17478_,
		_w17479_,
		_w17482_,
		_w17483_
	);
	LUT3 #(
		.INIT('ha9)
	) name11657 (
		\u1_L10_reg[12]/NET0131 ,
		_w17477_,
		_w17483_,
		_w17484_
	);
	LUT4 #(
		.INIT('hc693)
	) name11658 (
		decrypt_pad,
		\u1_R10_reg[20]/NET0131 ,
		\u1_uk_K_r10_reg[22]/NET0131 ,
		\u1_uk_K_r10_reg[45]/P0001 ,
		_w17485_
	);
	LUT4 #(
		.INIT('hc963)
	) name11659 (
		decrypt_pad,
		\u1_R10_reg[19]/NET0131 ,
		\u1_uk_K_r10_reg[2]/NET0131 ,
		\u1_uk_K_r10_reg[7]/NET0131 ,
		_w17486_
	);
	LUT4 #(
		.INIT('hc963)
	) name11660 (
		decrypt_pad,
		\u1_R10_reg[17]/NET0131 ,
		\u1_uk_K_r10_reg[21]/NET0131 ,
		\u1_uk_K_r10_reg[2]/NET0131 ,
		_w17487_
	);
	LUT4 #(
		.INIT('hc963)
	) name11661 (
		decrypt_pad,
		\u1_R10_reg[16]/NET0131 ,
		\u1_uk_K_r10_reg[30]/NET0131 ,
		\u1_uk_K_r10_reg[35]/NET0131 ,
		_w17488_
	);
	LUT4 #(
		.INIT('hc693)
	) name11662 (
		decrypt_pad,
		\u1_R10_reg[21]/NET0131 ,
		\u1_uk_K_r10_reg[23]/NET0131 ,
		\u1_uk_K_r10_reg[42]/NET0131 ,
		_w17489_
	);
	LUT2 #(
		.INIT('h2)
	) name11663 (
		_w17488_,
		_w17489_,
		_w17490_
	);
	LUT4 #(
		.INIT('hc963)
	) name11664 (
		decrypt_pad,
		\u1_R10_reg[18]/NET0131 ,
		\u1_uk_K_r10_reg[15]/NET0131 ,
		\u1_uk_K_r10_reg[51]/NET0131 ,
		_w17491_
	);
	LUT4 #(
		.INIT('h938f)
	) name11665 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17492_
	);
	LUT2 #(
		.INIT('h2)
	) name11666 (
		_w17486_,
		_w17492_,
		_w17493_
	);
	LUT3 #(
		.INIT('hbe)
	) name11667 (
		_w17488_,
		_w17489_,
		_w17487_,
		_w17494_
	);
	LUT2 #(
		.INIT('h1)
	) name11668 (
		_w17491_,
		_w17486_,
		_w17495_
	);
	LUT2 #(
		.INIT('h4)
	) name11669 (
		_w17494_,
		_w17495_,
		_w17496_
	);
	LUT3 #(
		.INIT('h80)
	) name11670 (
		_w17488_,
		_w17489_,
		_w17487_,
		_w17497_
	);
	LUT2 #(
		.INIT('h2)
	) name11671 (
		_w17491_,
		_w17486_,
		_w17498_
	);
	LUT4 #(
		.INIT('h0400)
	) name11672 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17499_
	);
	LUT4 #(
		.INIT('h0008)
	) name11673 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17500_
	);
	LUT4 #(
		.INIT('hfbb7)
	) name11674 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17501_
	);
	LUT3 #(
		.INIT('h70)
	) name11675 (
		_w17497_,
		_w17498_,
		_w17501_,
		_w17502_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11676 (
		_w17485_,
		_w17493_,
		_w17496_,
		_w17502_,
		_w17503_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11677 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17486_,
		_w17504_
	);
	LUT4 #(
		.INIT('heefc)
	) name11678 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17505_
	);
	LUT2 #(
		.INIT('h8)
	) name11679 (
		_w17504_,
		_w17505_,
		_w17506_
	);
	LUT3 #(
		.INIT('h04)
	) name11680 (
		_w17488_,
		_w17489_,
		_w17487_,
		_w17507_
	);
	LUT4 #(
		.INIT('h00df)
	) name11681 (
		_w17491_,
		_w17489_,
		_w17487_,
		_w17486_,
		_w17508_
	);
	LUT4 #(
		.INIT('h0004)
	) name11682 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17509_
	);
	LUT4 #(
		.INIT('h4000)
	) name11683 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17510_
	);
	LUT4 #(
		.INIT('hbffb)
	) name11684 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17511_
	);
	LUT3 #(
		.INIT('h40)
	) name11685 (
		_w17507_,
		_w17508_,
		_w17511_,
		_w17512_
	);
	LUT4 #(
		.INIT('h0080)
	) name11686 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17513_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name11687 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17514_
	);
	LUT4 #(
		.INIT('h001f)
	) name11688 (
		_w17506_,
		_w17512_,
		_w17514_,
		_w17485_,
		_w17515_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name11689 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17516_
	);
	LUT4 #(
		.INIT('h0020)
	) name11690 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17517_
	);
	LUT4 #(
		.INIT('hfddf)
	) name11691 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17518_
	);
	LUT3 #(
		.INIT('hd8)
	) name11692 (
		_w17486_,
		_w17516_,
		_w17518_,
		_w17519_
	);
	LUT4 #(
		.INIT('h5655)
	) name11693 (
		\u1_L10_reg[14]/NET0131 ,
		_w17515_,
		_w17503_,
		_w17519_,
		_w17520_
	);
	LUT4 #(
		.INIT('hddea)
	) name11694 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17521_
	);
	LUT2 #(
		.INIT('h9)
	) name11695 (
		_w17353_,
		_w17351_,
		_w17522_
	);
	LUT4 #(
		.INIT('h9000)
	) name11696 (
		_w17353_,
		_w17351_,
		_w17350_,
		_w17352_,
		_w17523_
	);
	LUT4 #(
		.INIT('hbfdf)
	) name11697 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17524_
	);
	LUT4 #(
		.INIT('h3200)
	) name11698 (
		_w17350_,
		_w17523_,
		_w17521_,
		_w17524_,
		_w17525_
	);
	LUT2 #(
		.INIT('h8)
	) name11699 (
		_w17351_,
		_w17366_,
		_w17526_
	);
	LUT4 #(
		.INIT('h0200)
	) name11700 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17527_
	);
	LUT4 #(
		.INIT('hfd03)
	) name11701 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17528_
	);
	LUT4 #(
		.INIT('h8480)
	) name11702 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17529_
	);
	LUT4 #(
		.INIT('h0c01)
	) name11703 (
		_w17351_,
		_w17354_,
		_w17350_,
		_w17352_,
		_w17530_
	);
	LUT4 #(
		.INIT('h0031)
	) name11704 (
		_w17350_,
		_w17529_,
		_w17528_,
		_w17530_,
		_w17531_
	);
	LUT4 #(
		.INIT('h3120)
	) name11705 (
		_w17357_,
		_w17526_,
		_w17531_,
		_w17525_,
		_w17532_
	);
	LUT2 #(
		.INIT('h9)
	) name11706 (
		\u1_L10_reg[17]/NET0131 ,
		_w17532_,
		_w17533_
	);
	LUT4 #(
		.INIT('hc693)
	) name11707 (
		decrypt_pad,
		\u1_R10_reg[30]/NET0131 ,
		\u1_uk_K_r10_reg[43]/NET0131 ,
		\u1_uk_K_r10_reg[7]/NET0131 ,
		_w17534_
	);
	LUT4 #(
		.INIT('hc963)
	) name11708 (
		decrypt_pad,
		\u1_R10_reg[1]/NET0131 ,
		\u1_uk_K_r10_reg[22]/NET0131 ,
		\u1_uk_K_r10_reg[31]/NET0131 ,
		_w17535_
	);
	LUT4 #(
		.INIT('hc693)
	) name11709 (
		decrypt_pad,
		\u1_R10_reg[28]/NET0131 ,
		\u1_uk_K_r10_reg[15]/NET0131 ,
		\u1_uk_K_r10_reg[38]/NET0131 ,
		_w17536_
	);
	LUT4 #(
		.INIT('hc963)
	) name11710 (
		decrypt_pad,
		\u1_R10_reg[29]/NET0131 ,
		\u1_uk_K_r10_reg[37]/NET0131 ,
		\u1_uk_K_r10_reg[42]/NET0131 ,
		_w17537_
	);
	LUT4 #(
		.INIT('hf100)
	) name11711 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17538_
	);
	LUT4 #(
		.INIT('h0ef3)
	) name11712 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17539_
	);
	LUT4 #(
		.INIT('hc693)
	) name11713 (
		decrypt_pad,
		\u1_R10_reg[31]/P0001 ,
		\u1_uk_K_r10_reg[0]/NET0131 ,
		\u1_uk_K_r10_reg[50]/NET0131 ,
		_w17540_
	);
	LUT4 #(
		.INIT('h0010)
	) name11714 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17541_
	);
	LUT4 #(
		.INIT('hc963)
	) name11715 (
		decrypt_pad,
		\u1_R10_reg[32]/NET0131 ,
		\u1_uk_K_r10_reg[1]/NET0131 ,
		\u1_uk_K_r10_reg[37]/NET0131 ,
		_w17542_
	);
	LUT4 #(
		.INIT('h00f4)
	) name11716 (
		_w17539_,
		_w17540_,
		_w17541_,
		_w17542_,
		_w17543_
	);
	LUT4 #(
		.INIT('h0200)
	) name11717 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17544_
	);
	LUT4 #(
		.INIT('h0001)
	) name11718 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17545_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name11719 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17546_
	);
	LUT2 #(
		.INIT('h2)
	) name11720 (
		_w17534_,
		_w17537_,
		_w17547_
	);
	LUT4 #(
		.INIT('hf95e)
	) name11721 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17548_
	);
	LUT2 #(
		.INIT('h1)
	) name11722 (
		_w17540_,
		_w17548_,
		_w17549_
	);
	LUT3 #(
		.INIT('h40)
	) name11723 (
		_w17534_,
		_w17536_,
		_w17537_,
		_w17550_
	);
	LUT2 #(
		.INIT('h4)
	) name11724 (
		_w17536_,
		_w17540_,
		_w17551_
	);
	LUT3 #(
		.INIT('h08)
	) name11725 (
		_w17534_,
		_w17535_,
		_w17537_,
		_w17552_
	);
	LUT3 #(
		.INIT('h45)
	) name11726 (
		_w17550_,
		_w17551_,
		_w17552_,
		_w17553_
	);
	LUT4 #(
		.INIT('h0100)
	) name11727 (
		_w17535_,
		_w17536_,
		_w17537_,
		_w17540_,
		_w17554_
	);
	LUT2 #(
		.INIT('h1)
	) name11728 (
		_w17554_,
		_w17544_,
		_w17555_
	);
	LUT4 #(
		.INIT('h0004)
	) name11729 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17556_
	);
	LUT4 #(
		.INIT('h0800)
	) name11730 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17557_
	);
	LUT4 #(
		.INIT('hf7fb)
	) name11731 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17558_
	);
	LUT4 #(
		.INIT('h0002)
	) name11732 (
		_w17536_,
		_w17537_,
		_w17540_,
		_w17542_,
		_w17559_
	);
	LUT3 #(
		.INIT('h0d)
	) name11733 (
		_w17540_,
		_w17558_,
		_w17559_,
		_w17560_
	);
	LUT4 #(
		.INIT('hd500)
	) name11734 (
		_w17542_,
		_w17553_,
		_w17555_,
		_w17560_,
		_w17561_
	);
	LUT4 #(
		.INIT('h5655)
	) name11735 (
		\u1_L10_reg[15]/P0001 ,
		_w17543_,
		_w17549_,
		_w17561_,
		_w17562_
	);
	LUT4 #(
		.INIT('hccfd)
	) name11736 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17563_
	);
	LUT4 #(
		.INIT('h6fbf)
	) name11737 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17564_
	);
	LUT4 #(
		.INIT('h08aa)
	) name11738 (
		_w17419_,
		_w17431_,
		_w17563_,
		_w17564_,
		_w17565_
	);
	LUT3 #(
		.INIT('h01)
	) name11739 (
		_w17417_,
		_w17422_,
		_w17418_,
		_w17566_
	);
	LUT4 #(
		.INIT('h220a)
	) name11740 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17567_
	);
	LUT4 #(
		.INIT('hfda8)
	) name11741 (
		_w17419_,
		_w17448_,
		_w17566_,
		_w17567_,
		_w17568_
	);
	LUT4 #(
		.INIT('h7bf7)
	) name11742 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17569_
	);
	LUT3 #(
		.INIT('h45)
	) name11743 (
		_w17431_,
		_w17568_,
		_w17569_,
		_w17570_
	);
	LUT4 #(
		.INIT('hb3fb)
	) name11744 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17571_
	);
	LUT4 #(
		.INIT('h1090)
	) name11745 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17572_
	);
	LUT4 #(
		.INIT('hcc04)
	) name11746 (
		_w17419_,
		_w17431_,
		_w17571_,
		_w17572_,
		_w17573_
	);
	LUT3 #(
		.INIT('h04)
	) name11747 (
		_w17419_,
		_w17422_,
		_w17418_,
		_w17574_
	);
	LUT2 #(
		.INIT('h8)
	) name11748 (
		_w17443_,
		_w17574_,
		_w17575_
	);
	LUT2 #(
		.INIT('h1)
	) name11749 (
		_w17573_,
		_w17575_,
		_w17576_
	);
	LUT4 #(
		.INIT('h5655)
	) name11750 (
		\u1_L10_reg[1]/NET0131 ,
		_w17570_,
		_w17565_,
		_w17576_,
		_w17577_
	);
	LUT4 #(
		.INIT('h0020)
	) name11751 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17578_
	);
	LUT2 #(
		.INIT('h8)
	) name11752 (
		_w17535_,
		_w17536_,
		_w17579_
	);
	LUT3 #(
		.INIT('hba)
	) name11753 (
		_w17534_,
		_w17537_,
		_w17540_,
		_w17580_
	);
	LUT4 #(
		.INIT('h00df)
	) name11754 (
		_w17534_,
		_w17536_,
		_w17537_,
		_w17542_,
		_w17581_
	);
	LUT4 #(
		.INIT('h0d00)
	) name11755 (
		_w17579_,
		_w17580_,
		_w17578_,
		_w17581_,
		_w17582_
	);
	LUT4 #(
		.INIT('hcf5f)
	) name11756 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17583_
	);
	LUT2 #(
		.INIT('h2)
	) name11757 (
		_w17540_,
		_w17583_,
		_w17584_
	);
	LUT4 #(
		.INIT('h0008)
	) name11758 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17540_,
		_w17585_
	);
	LUT4 #(
		.INIT('h0010)
	) name11759 (
		_w17535_,
		_w17536_,
		_w17537_,
		_w17540_,
		_w17586_
	);
	LUT3 #(
		.INIT('h01)
	) name11760 (
		_w17545_,
		_w17586_,
		_w17585_,
		_w17587_
	);
	LUT3 #(
		.INIT('h40)
	) name11761 (
		_w17584_,
		_w17587_,
		_w17582_,
		_w17588_
	);
	LUT4 #(
		.INIT('h1090)
	) name11762 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17589_
	);
	LUT3 #(
		.INIT('h80)
	) name11763 (
		_w17534_,
		_w17536_,
		_w17537_,
		_w17590_
	);
	LUT4 #(
		.INIT('hf3bb)
	) name11764 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17591_
	);
	LUT4 #(
		.INIT('he4ee)
	) name11765 (
		_w17540_,
		_w17589_,
		_w17590_,
		_w17591_,
		_w17592_
	);
	LUT4 #(
		.INIT('h2002)
	) name11766 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17593_
	);
	LUT3 #(
		.INIT('h02)
	) name11767 (
		_w17542_,
		_w17556_,
		_w17593_,
		_w17594_
	);
	LUT2 #(
		.INIT('h4)
	) name11768 (
		_w17592_,
		_w17594_,
		_w17595_
	);
	LUT4 #(
		.INIT('h0100)
	) name11769 (
		_w17534_,
		_w17536_,
		_w17537_,
		_w17540_,
		_w17596_
	);
	LUT3 #(
		.INIT('h04)
	) name11770 (
		_w17534_,
		_w17537_,
		_w17540_,
		_w17597_
	);
	LUT3 #(
		.INIT('h13)
	) name11771 (
		_w17579_,
		_w17596_,
		_w17597_,
		_w17598_
	);
	LUT4 #(
		.INIT('ha955)
	) name11772 (
		\u1_L10_reg[21]/NET0131 ,
		_w17588_,
		_w17595_,
		_w17598_,
		_w17599_
	);
	LUT4 #(
		.INIT('h3dc8)
	) name11773 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17600_
	);
	LUT4 #(
		.INIT('hee3f)
	) name11774 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17601_
	);
	LUT4 #(
		.INIT('ha7ff)
	) name11775 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17602_
	);
	LUT4 #(
		.INIT('hd800)
	) name11776 (
		_w17486_,
		_w17600_,
		_w17601_,
		_w17602_,
		_w17603_
	);
	LUT2 #(
		.INIT('h2)
	) name11777 (
		_w17485_,
		_w17603_,
		_w17604_
	);
	LUT4 #(
		.INIT('hddf3)
	) name11778 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17605_
	);
	LUT2 #(
		.INIT('h1)
	) name11779 (
		_w17486_,
		_w17605_,
		_w17606_
	);
	LUT4 #(
		.INIT('h1000)
	) name11780 (
		_w17491_,
		_w17489_,
		_w17487_,
		_w17486_,
		_w17607_
	);
	LUT4 #(
		.INIT('h0001)
	) name11781 (
		_w17491_,
		_w17488_,
		_w17487_,
		_w17486_,
		_w17608_
	);
	LUT4 #(
		.INIT('h2000)
	) name11782 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17609_
	);
	LUT3 #(
		.INIT('h01)
	) name11783 (
		_w17608_,
		_w17609_,
		_w17607_,
		_w17610_
	);
	LUT4 #(
		.INIT('hf7ed)
	) name11784 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17611_
	);
	LUT4 #(
		.INIT('h0008)
	) name11785 (
		_w17491_,
		_w17488_,
		_w17487_,
		_w17486_,
		_w17612_
	);
	LUT4 #(
		.INIT('h0031)
	) name11786 (
		_w17486_,
		_w17510_,
		_w17611_,
		_w17612_,
		_w17613_
	);
	LUT4 #(
		.INIT('hba00)
	) name11787 (
		_w17485_,
		_w17606_,
		_w17610_,
		_w17613_,
		_w17614_
	);
	LUT3 #(
		.INIT('h65)
	) name11788 (
		\u1_L10_reg[25]/NET0131 ,
		_w17604_,
		_w17614_,
		_w17615_
	);
	LUT4 #(
		.INIT('hc963)
	) name11789 (
		decrypt_pad,
		\u1_R10_reg[6]/NET0131 ,
		\u1_uk_K_r10_reg[46]/NET0131 ,
		\u1_uk_K_r10_reg[55]/NET0131 ,
		_w17616_
	);
	LUT4 #(
		.INIT('hc963)
	) name11790 (
		decrypt_pad,
		\u1_R10_reg[4]/NET0131 ,
		\u1_uk_K_r10_reg[19]/NET0131 ,
		\u1_uk_K_r10_reg[53]/NET0131 ,
		_w17617_
	);
	LUT4 #(
		.INIT('hc963)
	) name11791 (
		decrypt_pad,
		\u1_R10_reg[9]/NET0131 ,
		\u1_uk_K_r10_reg[11]/NET0131 ,
		\u1_uk_K_r10_reg[20]/NET0131 ,
		_w17618_
	);
	LUT4 #(
		.INIT('hc693)
	) name11792 (
		decrypt_pad,
		\u1_R10_reg[5]/NET0131 ,
		\u1_uk_K_r10_reg[32]/NET0131 ,
		\u1_uk_K_r10_reg[55]/NET0131 ,
		_w17619_
	);
	LUT4 #(
		.INIT('h1000)
	) name11793 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17620_
	);
	LUT4 #(
		.INIT('hc693)
	) name11794 (
		decrypt_pad,
		\u1_R10_reg[7]/NET0131 ,
		\u1_uk_K_r10_reg[17]/NET0131 ,
		\u1_uk_K_r10_reg[40]/NET0131 ,
		_w17621_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name11795 (
		_w17621_,
		_w17617_,
		_w17618_,
		_w17619_,
		_w17622_
	);
	LUT3 #(
		.INIT('h45)
	) name11796 (
		_w17621_,
		_w17619_,
		_w17616_,
		_w17623_
	);
	LUT2 #(
		.INIT('h4)
	) name11797 (
		_w17621_,
		_w17617_,
		_w17624_
	);
	LUT4 #(
		.INIT('habaa)
	) name11798 (
		_w17621_,
		_w17617_,
		_w17619_,
		_w17616_,
		_w17625_
	);
	LUT4 #(
		.INIT('hbfae)
	) name11799 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17626_
	);
	LUT2 #(
		.INIT('h8)
	) name11800 (
		_w17617_,
		_w17616_,
		_w17627_
	);
	LUT4 #(
		.INIT('h2000)
	) name11801 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17628_
	);
	LUT4 #(
		.INIT('h9fae)
	) name11802 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17629_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name11803 (
		_w17620_,
		_w17622_,
		_w17625_,
		_w17629_,
		_w17630_
	);
	LUT4 #(
		.INIT('h0400)
	) name11804 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17631_
	);
	LUT4 #(
		.INIT('hc693)
	) name11805 (
		decrypt_pad,
		\u1_R10_reg[8]/NET0131 ,
		\u1_uk_K_r10_reg[40]/NET0131 ,
		\u1_uk_K_r10_reg[6]/NET0131 ,
		_w17632_
	);
	LUT2 #(
		.INIT('h2)
	) name11806 (
		_w17617_,
		_w17616_,
		_w17633_
	);
	LUT3 #(
		.INIT('h51)
	) name11807 (
		_w17621_,
		_w17618_,
		_w17619_,
		_w17634_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11808 (
		_w17632_,
		_w17633_,
		_w17634_,
		_w17631_,
		_w17635_
	);
	LUT4 #(
		.INIT('h5b59)
	) name11809 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17636_
	);
	LUT4 #(
		.INIT('h7077)
	) name11810 (
		_w17621_,
		_w17626_,
		_w17625_,
		_w17636_,
		_w17637_
	);
	LUT2 #(
		.INIT('h6)
	) name11811 (
		_w17617_,
		_w17618_,
		_w17638_
	);
	LUT4 #(
		.INIT('h0900)
	) name11812 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17639_
	);
	LUT3 #(
		.INIT('h01)
	) name11813 (
		_w17632_,
		_w17628_,
		_w17639_,
		_w17640_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name11814 (
		_w17630_,
		_w17635_,
		_w17637_,
		_w17640_,
		_w17641_
	);
	LUT2 #(
		.INIT('h6)
	) name11815 (
		\u1_L10_reg[28]/NET0131 ,
		_w17641_,
		_w17642_
	);
	LUT4 #(
		.INIT('h779a)
	) name11816 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17643_
	);
	LUT4 #(
		.INIT('h0e02)
	) name11817 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17644_
	);
	LUT4 #(
		.INIT('hf17d)
	) name11818 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17645_
	);
	LUT4 #(
		.INIT('h1000)
	) name11819 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17646_
	);
	LUT4 #(
		.INIT('h00e4)
	) name11820 (
		_w17385_,
		_w17645_,
		_w17643_,
		_w17646_,
		_w17647_
	);
	LUT2 #(
		.INIT('h1)
	) name11821 (
		_w17379_,
		_w17647_,
		_w17648_
	);
	LUT4 #(
		.INIT('hdd7d)
	) name11822 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17649_
	);
	LUT2 #(
		.INIT('h2)
	) name11823 (
		_w17385_,
		_w17649_,
		_w17650_
	);
	LUT3 #(
		.INIT('h48)
	) name11824 (
		_w17382_,
		_w17380_,
		_w17383_,
		_w17651_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name11825 (
		_w17381_,
		_w17380_,
		_w17385_,
		_w17383_,
		_w17652_
	);
	LUT3 #(
		.INIT('h01)
	) name11826 (
		_w17652_,
		_w17644_,
		_w17651_,
		_w17653_
	);
	LUT4 #(
		.INIT('h2000)
	) name11827 (
		_w17381_,
		_w17380_,
		_w17385_,
		_w17383_,
		_w17654_
	);
	LUT2 #(
		.INIT('h1)
	) name11828 (
		_w17390_,
		_w17654_,
		_w17655_
	);
	LUT4 #(
		.INIT('h5700)
	) name11829 (
		_w17379_,
		_w17650_,
		_w17653_,
		_w17655_,
		_w17656_
	);
	LUT3 #(
		.INIT('h9a)
	) name11830 (
		\u1_L10_reg[29]/NET0131 ,
		_w17648_,
		_w17656_,
		_w17657_
	);
	LUT4 #(
		.INIT('h0001)
	) name11831 (
		_w17621_,
		_w17617_,
		_w17618_,
		_w17619_,
		_w17658_
	);
	LUT4 #(
		.INIT('h0080)
	) name11832 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17659_
	);
	LUT3 #(
		.INIT('h02)
	) name11833 (
		_w17632_,
		_w17659_,
		_w17658_,
		_w17660_
	);
	LUT4 #(
		.INIT('h1500)
	) name11834 (
		_w17621_,
		_w17617_,
		_w17619_,
		_w17616_,
		_w17661_
	);
	LUT4 #(
		.INIT('h0002)
	) name11835 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17662_
	);
	LUT4 #(
		.INIT('h80a0)
	) name11836 (
		_w17621_,
		_w17617_,
		_w17619_,
		_w17616_,
		_w17663_
	);
	LUT4 #(
		.INIT('h0203)
	) name11837 (
		_w17638_,
		_w17662_,
		_w17663_,
		_w17661_,
		_w17664_
	);
	LUT4 #(
		.INIT('h0034)
	) name11838 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17665_
	);
	LUT4 #(
		.INIT('h0800)
	) name11839 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17666_
	);
	LUT4 #(
		.INIT('h0105)
	) name11840 (
		_w17632_,
		_w17621_,
		_w17665_,
		_w17666_,
		_w17667_
	);
	LUT4 #(
		.INIT('h51f3)
	) name11841 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17668_
	);
	LUT4 #(
		.INIT('h5515)
	) name11842 (
		_w17621_,
		_w17617_,
		_w17618_,
		_w17619_,
		_w17669_
	);
	LUT2 #(
		.INIT('h2)
	) name11843 (
		_w17618_,
		_w17616_,
		_w17670_
	);
	LUT4 #(
		.INIT('h0004)
	) name11844 (
		_w17621_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17671_
	);
	LUT4 #(
		.INIT('h4000)
	) name11845 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17672_
	);
	LUT4 #(
		.INIT('h000b)
	) name11846 (
		_w17668_,
		_w17669_,
		_w17671_,
		_w17672_,
		_w17673_
	);
	LUT4 #(
		.INIT('h0777)
	) name11847 (
		_w17660_,
		_w17664_,
		_w17667_,
		_w17673_,
		_w17674_
	);
	LUT3 #(
		.INIT('h10)
	) name11848 (
		_w17618_,
		_w17619_,
		_w17616_,
		_w17675_
	);
	LUT4 #(
		.INIT('h0100)
	) name11849 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17676_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name11850 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17677_
	);
	LUT4 #(
		.INIT('h4404)
	) name11851 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17678_
	);
	LUT4 #(
		.INIT('h31f5)
	) name11852 (
		_w17621_,
		_w17623_,
		_w17677_,
		_w17678_,
		_w17679_
	);
	LUT3 #(
		.INIT('h65)
	) name11853 (
		\u1_L10_reg[2]/NET0131 ,
		_w17674_,
		_w17679_,
		_w17680_
	);
	LUT3 #(
		.INIT('he0)
	) name11854 (
		_w17380_,
		_w17385_,
		_w17383_,
		_w17681_
	);
	LUT4 #(
		.INIT('h0002)
	) name11855 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17682_
	);
	LUT4 #(
		.INIT('h002a)
	) name11856 (
		_w17379_,
		_w17398_,
		_w17681_,
		_w17682_,
		_w17683_
	);
	LUT4 #(
		.INIT('hbc77)
	) name11857 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17684_
	);
	LUT4 #(
		.INIT('h0100)
	) name11858 (
		_w17379_,
		_w17390_,
		_w17393_,
		_w17684_,
		_w17685_
	);
	LUT3 #(
		.INIT('hde)
	) name11859 (
		_w17381_,
		_w17382_,
		_w17383_,
		_w17686_
	);
	LUT4 #(
		.INIT('h2090)
	) name11860 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17687_
	);
	LUT2 #(
		.INIT('h2)
	) name11861 (
		_w17385_,
		_w17687_,
		_w17688_
	);
	LUT3 #(
		.INIT('he0)
	) name11862 (
		_w17683_,
		_w17685_,
		_w17688_,
		_w17689_
	);
	LUT4 #(
		.INIT('hfcf4)
	) name11863 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17690_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11864 (
		_w17379_,
		_w17398_,
		_w17681_,
		_w17690_,
		_w17691_
	);
	LUT4 #(
		.INIT('hefdd)
	) name11865 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17692_
	);
	LUT4 #(
		.INIT('h0100)
	) name11866 (
		_w17379_,
		_w17390_,
		_w17393_,
		_w17692_,
		_w17693_
	);
	LUT4 #(
		.INIT('h8040)
	) name11867 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17694_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name11868 (
		_w17382_,
		_w17380_,
		_w17385_,
		_w17383_,
		_w17695_
	);
	LUT2 #(
		.INIT('h4)
	) name11869 (
		_w17694_,
		_w17695_,
		_w17696_
	);
	LUT3 #(
		.INIT('he0)
	) name11870 (
		_w17691_,
		_w17693_,
		_w17696_,
		_w17697_
	);
	LUT3 #(
		.INIT('ha9)
	) name11871 (
		\u1_L10_reg[4]/NET0131 ,
		_w17689_,
		_w17697_,
		_w17698_
	);
	LUT3 #(
		.INIT('h02)
	) name11872 (
		_w17419_,
		_w17439_,
		_w17433_,
		_w17699_
	);
	LUT4 #(
		.INIT('h0806)
	) name11873 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17700_
	);
	LUT4 #(
		.INIT('hefcc)
	) name11874 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17701_
	);
	LUT4 #(
		.INIT('h0504)
	) name11875 (
		_w17419_,
		_w17431_,
		_w17700_,
		_w17701_,
		_w17702_
	);
	LUT2 #(
		.INIT('h1)
	) name11876 (
		_w17699_,
		_w17702_,
		_w17703_
	);
	LUT4 #(
		.INIT('h0084)
	) name11877 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17704_
	);
	LUT4 #(
		.INIT('h0002)
	) name11878 (
		_w17419_,
		_w17417_,
		_w17416_,
		_w17418_,
		_w17705_
	);
	LUT3 #(
		.INIT('h02)
	) name11879 (
		_w17431_,
		_w17705_,
		_w17704_,
		_w17706_
	);
	LUT4 #(
		.INIT('hcdff)
	) name11880 (
		_w17419_,
		_w17417_,
		_w17416_,
		_w17418_,
		_w17707_
	);
	LUT4 #(
		.INIT('h54ff)
	) name11881 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17418_,
		_w17708_
	);
	LUT3 #(
		.INIT('h51)
	) name11882 (
		_w17419_,
		_w17417_,
		_w17422_,
		_w17709_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name11883 (
		_w17422_,
		_w17707_,
		_w17708_,
		_w17709_,
		_w17710_
	);
	LUT2 #(
		.INIT('h2)
	) name11884 (
		_w17429_,
		_w17436_,
		_w17711_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11885 (
		_w17417_,
		_w17416_,
		_w17422_,
		_w17431_,
		_w17712_
	);
	LUT3 #(
		.INIT('h10)
	) name11886 (
		_w17439_,
		_w17440_,
		_w17712_,
		_w17713_
	);
	LUT4 #(
		.INIT('h7077)
	) name11887 (
		_w17706_,
		_w17710_,
		_w17711_,
		_w17713_,
		_w17714_
	);
	LUT3 #(
		.INIT('h56)
	) name11888 (
		\u1_L10_reg[26]/NET0131 ,
		_w17703_,
		_w17714_,
		_w17715_
	);
	LUT4 #(
		.INIT('h3b19)
	) name11889 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17716_
	);
	LUT4 #(
		.INIT('h8000)
	) name11890 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17717_
	);
	LUT4 #(
		.INIT('h0e04)
	) name11891 (
		_w17385_,
		_w17686_,
		_w17717_,
		_w17716_,
		_w17718_
	);
	LUT2 #(
		.INIT('h1)
	) name11892 (
		_w17379_,
		_w17718_,
		_w17719_
	);
	LUT4 #(
		.INIT('ha4f5)
	) name11893 (
		_w17382_,
		_w17380_,
		_w17385_,
		_w17383_,
		_w17720_
	);
	LUT2 #(
		.INIT('h1)
	) name11894 (
		_w17381_,
		_w17720_,
		_w17721_
	);
	LUT4 #(
		.INIT('h2010)
	) name11895 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17383_,
		_w17722_
	);
	LUT4 #(
		.INIT('h0800)
	) name11896 (
		_w17381_,
		_w17382_,
		_w17380_,
		_w17385_,
		_w17723_
	);
	LUT3 #(
		.INIT('h01)
	) name11897 (
		_w17408_,
		_w17722_,
		_w17723_,
		_w17724_
	);
	LUT3 #(
		.INIT('h8a)
	) name11898 (
		_w17379_,
		_w17721_,
		_w17724_,
		_w17725_
	);
	LUT2 #(
		.INIT('h2)
	) name11899 (
		_w17409_,
		_w17394_,
		_w17726_
	);
	LUT4 #(
		.INIT('h5655)
	) name11900 (
		\u1_L10_reg[19]/P0001 ,
		_w17725_,
		_w17719_,
		_w17726_,
		_w17727_
	);
	LUT3 #(
		.INIT('h96)
	) name11901 (
		_w17353_,
		_w17351_,
		_w17352_,
		_w17728_
	);
	LUT3 #(
		.INIT('hb0)
	) name11902 (
		_w17353_,
		_w17354_,
		_w17352_,
		_w17729_
	);
	LUT4 #(
		.INIT('h040f)
	) name11903 (
		_w17353_,
		_w17354_,
		_w17350_,
		_w17352_,
		_w17730_
	);
	LUT2 #(
		.INIT('h8)
	) name11904 (
		_w17728_,
		_w17730_,
		_w17731_
	);
	LUT4 #(
		.INIT('hc080)
	) name11905 (
		_w17353_,
		_w17351_,
		_w17350_,
		_w17352_,
		_w17732_
	);
	LUT2 #(
		.INIT('h4)
	) name11906 (
		_w17729_,
		_w17732_,
		_w17733_
	);
	LUT3 #(
		.INIT('h07)
	) name11907 (
		_w17365_,
		_w17374_,
		_w17527_,
		_w17734_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11908 (
		_w17357_,
		_w17731_,
		_w17733_,
		_w17734_,
		_w17735_
	);
	LUT4 #(
		.INIT('h13ff)
	) name11909 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17736_
	);
	LUT4 #(
		.INIT('h0400)
	) name11910 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17737_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name11911 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17738_
	);
	LUT4 #(
		.INIT('hf400)
	) name11912 (
		_w17369_,
		_w17357_,
		_w17736_,
		_w17738_,
		_w17739_
	);
	LUT3 #(
		.INIT('h0b)
	) name11913 (
		_w17353_,
		_w17351_,
		_w17352_,
		_w17740_
	);
	LUT4 #(
		.INIT('h1030)
	) name11914 (
		_w17351_,
		_w17354_,
		_w17350_,
		_w17352_,
		_w17741_
	);
	LUT2 #(
		.INIT('h4)
	) name11915 (
		_w17740_,
		_w17741_,
		_w17742_
	);
	LUT3 #(
		.INIT('h81)
	) name11916 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17743_
	);
	LUT4 #(
		.INIT('h0040)
	) name11917 (
		_w17353_,
		_w17351_,
		_w17350_,
		_w17352_,
		_w17744_
	);
	LUT4 #(
		.INIT('h5554)
	) name11918 (
		_w17357_,
		_w17358_,
		_w17744_,
		_w17743_,
		_w17745_
	);
	LUT4 #(
		.INIT('h0302)
	) name11919 (
		_w17350_,
		_w17742_,
		_w17745_,
		_w17739_,
		_w17746_
	);
	LUT3 #(
		.INIT('h9a)
	) name11920 (
		\u1_L10_reg[23]/NET0131 ,
		_w17735_,
		_w17746_,
		_w17747_
	);
	LUT4 #(
		.INIT('hc3fa)
	) name11921 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17748_
	);
	LUT4 #(
		.INIT('h0040)
	) name11922 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17749_
	);
	LUT4 #(
		.INIT('h1000)
	) name11923 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17750_
	);
	LUT4 #(
		.INIT('hedbf)
	) name11924 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17751_
	);
	LUT4 #(
		.INIT('h0455)
	) name11925 (
		_w17540_,
		_w17542_,
		_w17748_,
		_w17751_,
		_w17752_
	);
	LUT3 #(
		.INIT('hb0)
	) name11926 (
		_w17535_,
		_w17536_,
		_w17540_,
		_w17753_
	);
	LUT4 #(
		.INIT('hf79b)
	) name11927 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w17754_
	);
	LUT4 #(
		.INIT('h80cc)
	) name11928 (
		_w17538_,
		_w17542_,
		_w17753_,
		_w17754_,
		_w17755_
	);
	LUT4 #(
		.INIT('haf8d)
	) name11929 (
		_w17535_,
		_w17536_,
		_w17540_,
		_w17542_,
		_w17756_
	);
	LUT2 #(
		.INIT('h2)
	) name11930 (
		_w17547_,
		_w17756_,
		_w17757_
	);
	LUT4 #(
		.INIT('hdf00)
	) name11931 (
		_w17534_,
		_w17536_,
		_w17537_,
		_w17540_,
		_w17758_
	);
	LUT3 #(
		.INIT('h63)
	) name11932 (
		_w17534_,
		_w17535_,
		_w17537_,
		_w17759_
	);
	LUT4 #(
		.INIT('h0080)
	) name11933 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17540_,
		_w17760_
	);
	LUT4 #(
		.INIT('h0111)
	) name11934 (
		_w17586_,
		_w17760_,
		_w17758_,
		_w17759_,
		_w17761_
	);
	LUT4 #(
		.INIT('h0032)
	) name11935 (
		_w17542_,
		_w17757_,
		_w17761_,
		_w17755_,
		_w17762_
	);
	LUT3 #(
		.INIT('h65)
	) name11936 (
		\u1_L10_reg[27]/NET0131 ,
		_w17752_,
		_w17762_,
		_w17763_
	);
	LUT2 #(
		.INIT('h9)
	) name11937 (
		_w17322_,
		_w17324_,
		_w17764_
	);
	LUT4 #(
		.INIT('hd003)
	) name11938 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17765_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name11939 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17766_
	);
	LUT3 #(
		.INIT('h01)
	) name11940 (
		_w17325_,
		_w17766_,
		_w17765_,
		_w17767_
	);
	LUT4 #(
		.INIT('h0800)
	) name11941 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17768_
	);
	LUT4 #(
		.INIT('hb5bc)
	) name11942 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17769_
	);
	LUT3 #(
		.INIT('h31)
	) name11943 (
		_w17325_,
		_w17768_,
		_w17769_,
		_w17770_
	);
	LUT3 #(
		.INIT('h8a)
	) name11944 (
		_w17319_,
		_w17767_,
		_w17770_,
		_w17771_
	);
	LUT3 #(
		.INIT('h40)
	) name11945 (
		_w17321_,
		_w17322_,
		_w17324_,
		_w17772_
	);
	LUT4 #(
		.INIT('hab89)
	) name11946 (
		_w17325_,
		_w17472_,
		_w17474_,
		_w17772_,
		_w17773_
	);
	LUT4 #(
		.INIT('h7bd7)
	) name11947 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17774_
	);
	LUT4 #(
		.INIT('h00c8)
	) name11948 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17325_,
		_w17775_
	);
	LUT4 #(
		.INIT('h135f)
	) name11949 (
		_w17325_,
		_w17340_,
		_w17332_,
		_w17775_,
		_w17776_
	);
	LUT4 #(
		.INIT('hba00)
	) name11950 (
		_w17319_,
		_w17773_,
		_w17774_,
		_w17776_,
		_w17777_
	);
	LUT3 #(
		.INIT('h65)
	) name11951 (
		\u1_L10_reg[32]/NET0131 ,
		_w17771_,
		_w17777_,
		_w17778_
	);
	LUT4 #(
		.INIT('hc963)
	) name11952 (
		decrypt_pad,
		\u1_R10_reg[11]/NET0131 ,
		\u1_uk_K_r10_reg[26]/NET0131 ,
		\u1_uk_K_r10_reg[3]/NET0131 ,
		_w17779_
	);
	LUT4 #(
		.INIT('hc693)
	) name11953 (
		decrypt_pad,
		\u1_R10_reg[12]/NET0131 ,
		\u1_uk_K_r10_reg[18]/NET0131 ,
		\u1_uk_K_r10_reg[41]/P0001 ,
		_w17780_
	);
	LUT4 #(
		.INIT('hc963)
	) name11954 (
		decrypt_pad,
		\u1_R10_reg[13]/NET0131 ,
		\u1_uk_K_r10_reg[54]/NET0131 ,
		\u1_uk_K_r10_reg[6]/NET0131 ,
		_w17781_
	);
	LUT4 #(
		.INIT('hc963)
	) name11955 (
		decrypt_pad,
		\u1_R10_reg[9]/NET0131 ,
		\u1_uk_K_r10_reg[17]/NET0131 ,
		\u1_uk_K_r10_reg[26]/NET0131 ,
		_w17782_
	);
	LUT4 #(
		.INIT('hc963)
	) name11956 (
		decrypt_pad,
		\u1_R10_reg[10]/NET0131 ,
		\u1_uk_K_r10_reg[25]/NET0131 ,
		\u1_uk_K_r10_reg[34]/NET0131 ,
		_w17783_
	);
	LUT4 #(
		.INIT('hc963)
	) name11957 (
		decrypt_pad,
		\u1_R10_reg[8]/NET0131 ,
		\u1_uk_K_r10_reg[20]/NET0131 ,
		\u1_uk_K_r10_reg[54]/NET0131 ,
		_w17784_
	);
	LUT4 #(
		.INIT('h95b5)
	) name11958 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17785_
	);
	LUT2 #(
		.INIT('h1)
	) name11959 (
		_w17781_,
		_w17784_,
		_w17786_
	);
	LUT4 #(
		.INIT('h0001)
	) name11960 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17787_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name11961 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17788_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11962 (
		_w17780_,
		_w17779_,
		_w17785_,
		_w17788_,
		_w17789_
	);
	LUT2 #(
		.INIT('h6)
	) name11963 (
		_w17782_,
		_w17783_,
		_w17790_
	);
	LUT2 #(
		.INIT('h8)
	) name11964 (
		_w17781_,
		_w17784_,
		_w17791_
	);
	LUT2 #(
		.INIT('h8)
	) name11965 (
		_w17781_,
		_w17779_,
		_w17792_
	);
	LUT3 #(
		.INIT('h46)
	) name11966 (
		_w17781_,
		_w17784_,
		_w17779_,
		_w17793_
	);
	LUT2 #(
		.INIT('h1)
	) name11967 (
		_w17790_,
		_w17793_,
		_w17794_
	);
	LUT4 #(
		.INIT('h6660)
	) name11968 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17795_
	);
	LUT4 #(
		.INIT('h353f)
	) name11969 (
		_w17781_,
		_w17782_,
		_w17783_,
		_w17779_,
		_w17796_
	);
	LUT3 #(
		.INIT('h15)
	) name11970 (
		_w17780_,
		_w17795_,
		_w17796_,
		_w17797_
	);
	LUT3 #(
		.INIT('h80)
	) name11971 (
		_w17782_,
		_w17783_,
		_w17780_,
		_w17798_
	);
	LUT3 #(
		.INIT('h51)
	) name11972 (
		_w17784_,
		_w17782_,
		_w17783_,
		_w17799_
	);
	LUT2 #(
		.INIT('h9)
	) name11973 (
		_w17781_,
		_w17782_,
		_w17800_
	);
	LUT4 #(
		.INIT('h0090)
	) name11974 (
		_w17781_,
		_w17782_,
		_w17780_,
		_w17779_,
		_w17801_
	);
	LUT4 #(
		.INIT('h7077)
	) name11975 (
		_w17786_,
		_w17798_,
		_w17799_,
		_w17801_,
		_w17802_
	);
	LUT4 #(
		.INIT('h4500)
	) name11976 (
		_w17789_,
		_w17794_,
		_w17797_,
		_w17802_,
		_w17803_
	);
	LUT2 #(
		.INIT('h9)
	) name11977 (
		\u1_L10_reg[6]/NET0131 ,
		_w17803_,
		_w17804_
	);
	LUT4 #(
		.INIT('hf126)
	) name11978 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17805_
	);
	LUT4 #(
		.INIT('h2880)
	) name11979 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17806_
	);
	LUT4 #(
		.INIT('h5004)
	) name11980 (
		_w17320_,
		_w17321_,
		_w17322_,
		_w17324_,
		_w17807_
	);
	LUT4 #(
		.INIT('h1302)
	) name11981 (
		_w17325_,
		_w17806_,
		_w17807_,
		_w17805_,
		_w17808_
	);
	LUT2 #(
		.INIT('h2)
	) name11982 (
		_w17319_,
		_w17808_,
		_w17809_
	);
	LUT2 #(
		.INIT('h4)
	) name11983 (
		_w17325_,
		_w17806_,
		_w17810_
	);
	LUT2 #(
		.INIT('h2)
	) name11984 (
		_w17319_,
		_w17325_,
		_w17811_
	);
	LUT3 #(
		.INIT('h4c)
	) name11985 (
		_w17321_,
		_w17322_,
		_w17324_,
		_w17812_
	);
	LUT4 #(
		.INIT('h8a00)
	) name11986 (
		_w17320_,
		_w17322_,
		_w17324_,
		_w17325_,
		_w17813_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name11987 (
		_w17326_,
		_w17764_,
		_w17812_,
		_w17813_,
		_w17814_
	);
	LUT3 #(
		.INIT('h45)
	) name11988 (
		_w17339_,
		_w17325_,
		_w17807_,
		_w17815_
	);
	LUT4 #(
		.INIT('h0133)
	) name11989 (
		_w17319_,
		_w17811_,
		_w17814_,
		_w17815_,
		_w17816_
	);
	LUT4 #(
		.INIT('h5556)
	) name11990 (
		\u1_L10_reg[7]/NET0131 ,
		_w17810_,
		_w17816_,
		_w17809_,
		_w17817_
	);
	LUT3 #(
		.INIT('h02)
	) name11991 (
		_w17486_,
		_w17509_,
		_w17497_,
		_w17818_
	);
	LUT4 #(
		.INIT('h3010)
	) name11992 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17819_
	);
	LUT4 #(
		.INIT('h00f7)
	) name11993 (
		_w17488_,
		_w17489_,
		_w17487_,
		_w17486_,
		_w17820_
	);
	LUT2 #(
		.INIT('h4)
	) name11994 (
		_w17819_,
		_w17820_,
		_w17821_
	);
	LUT4 #(
		.INIT('he6fd)
	) name11995 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17822_
	);
	LUT4 #(
		.INIT('h0155)
	) name11996 (
		_w17485_,
		_w17818_,
		_w17821_,
		_w17822_,
		_w17823_
	);
	LUT4 #(
		.INIT('h0001)
	) name11997 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17824_
	);
	LUT4 #(
		.INIT('hff3e)
	) name11998 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17825_
	);
	LUT3 #(
		.INIT('h04)
	) name11999 (
		_w17491_,
		_w17488_,
		_w17486_,
		_w17826_
	);
	LUT4 #(
		.INIT('h00c4)
	) name12000 (
		_w17486_,
		_w17518_,
		_w17825_,
		_w17826_,
		_w17827_
	);
	LUT4 #(
		.INIT('he5df)
	) name12001 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17828_
	);
	LUT4 #(
		.INIT('haf23)
	) name12002 (
		_w17489_,
		_w17486_,
		_w17612_,
		_w17828_,
		_w17829_
	);
	LUT3 #(
		.INIT('hd0)
	) name12003 (
		_w17485_,
		_w17827_,
		_w17829_,
		_w17830_
	);
	LUT3 #(
		.INIT('h65)
	) name12004 (
		\u1_L10_reg[8]/NET0131 ,
		_w17823_,
		_w17830_,
		_w17831_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name12005 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17832_
	);
	LUT4 #(
		.INIT('hebed)
	) name12006 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17833_
	);
	LUT4 #(
		.INIT('h0313)
	) name12007 (
		_w17632_,
		_w17621_,
		_w17832_,
		_w17833_,
		_w17834_
	);
	LUT3 #(
		.INIT('h06)
	) name12008 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17835_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name12009 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17836_
	);
	LUT3 #(
		.INIT('h02)
	) name12010 (
		_w17621_,
		_w17836_,
		_w17835_,
		_w17837_
	);
	LUT3 #(
		.INIT('h8a)
	) name12011 (
		_w17621_,
		_w17618_,
		_w17619_,
		_w17838_
	);
	LUT3 #(
		.INIT('h32)
	) name12012 (
		_w17621_,
		_w17617_,
		_w17619_,
		_w17839_
	);
	LUT4 #(
		.INIT('h135f)
	) name12013 (
		_w17627_,
		_w17670_,
		_w17838_,
		_w17839_,
		_w17840_
	);
	LUT3 #(
		.INIT('h45)
	) name12014 (
		_w17632_,
		_w17837_,
		_w17840_,
		_w17841_
	);
	LUT3 #(
		.INIT('h01)
	) name12015 (
		_w17618_,
		_w17619_,
		_w17616_,
		_w17842_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12016 (
		_w17621_,
		_w17617_,
		_w17618_,
		_w17616_,
		_w17843_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12017 (
		_w17675_,
		_w17669_,
		_w17842_,
		_w17843_,
		_w17844_
	);
	LUT4 #(
		.INIT('hdf6f)
	) name12018 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17845_
	);
	LUT3 #(
		.INIT('h10)
	) name12019 (
		_w17671_,
		_w17672_,
		_w17845_,
		_w17846_
	);
	LUT3 #(
		.INIT('h8a)
	) name12020 (
		_w17632_,
		_w17844_,
		_w17846_,
		_w17847_
	);
	LUT4 #(
		.INIT('haaa9)
	) name12021 (
		\u1_L10_reg[13]/NET0131 ,
		_w17841_,
		_w17834_,
		_w17847_,
		_w17848_
	);
	LUT3 #(
		.INIT('h10)
	) name12022 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17849_
	);
	LUT3 #(
		.INIT('h28)
	) name12023 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17850_
	);
	LUT4 #(
		.INIT('h6979)
	) name12024 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17779_,
		_w17851_
	);
	LUT3 #(
		.INIT('h07)
	) name12025 (
		_w17784_,
		_w17783_,
		_w17779_,
		_w17852_
	);
	LUT4 #(
		.INIT('h0014)
	) name12026 (
		_w17781_,
		_w17784_,
		_w17783_,
		_w17779_,
		_w17853_
	);
	LUT4 #(
		.INIT('h2000)
	) name12027 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17854_
	);
	LUT4 #(
		.INIT('h000e)
	) name12028 (
		_w17783_,
		_w17851_,
		_w17853_,
		_w17854_,
		_w17855_
	);
	LUT4 #(
		.INIT('h6800)
	) name12029 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17779_,
		_w17856_
	);
	LUT4 #(
		.INIT('h00ab)
	) name12030 (
		_w17781_,
		_w17784_,
		_w17783_,
		_w17779_,
		_w17857_
	);
	LUT4 #(
		.INIT('h0045)
	) name12031 (
		_w17787_,
		_w17850_,
		_w17857_,
		_w17856_,
		_w17858_
	);
	LUT4 #(
		.INIT('h4100)
	) name12032 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17859_
	);
	LUT3 #(
		.INIT('h20)
	) name12033 (
		_w17784_,
		_w17782_,
		_w17783_,
		_w17860_
	);
	LUT4 #(
		.INIT('h00df)
	) name12034 (
		_w17784_,
		_w17782_,
		_w17783_,
		_w17779_,
		_w17861_
	);
	LUT3 #(
		.INIT('h0d)
	) name12035 (
		_w17779_,
		_w17859_,
		_w17861_,
		_w17862_
	);
	LUT4 #(
		.INIT('h00d8)
	) name12036 (
		_w17780_,
		_w17855_,
		_w17858_,
		_w17862_,
		_w17863_
	);
	LUT2 #(
		.INIT('h9)
	) name12037 (
		\u1_L10_reg[16]/NET0131 ,
		_w17863_,
		_w17864_
	);
	LUT3 #(
		.INIT('h02)
	) name12038 (
		_w17781_,
		_w17784_,
		_w17783_,
		_w17865_
	);
	LUT3 #(
		.INIT('hed)
	) name12039 (
		_w17781_,
		_w17784_,
		_w17783_,
		_w17866_
	);
	LUT4 #(
		.INIT('he2cd)
	) name12040 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17867_
	);
	LUT4 #(
		.INIT('h0400)
	) name12041 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17868_
	);
	LUT4 #(
		.INIT('h0009)
	) name12042 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17869_
	);
	LUT4 #(
		.INIT('h9db6)
	) name12043 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17870_
	);
	LUT4 #(
		.INIT('h3210)
	) name12044 (
		_w17779_,
		_w17868_,
		_w17870_,
		_w17867_,
		_w17871_
	);
	LUT2 #(
		.INIT('h1)
	) name12045 (
		_w17780_,
		_w17871_,
		_w17872_
	);
	LUT4 #(
		.INIT('h1d00)
	) name12046 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17873_
	);
	LUT3 #(
		.INIT('hd0)
	) name12047 (
		_w17782_,
		_w17783_,
		_w17779_,
		_w17874_
	);
	LUT3 #(
		.INIT('h10)
	) name12048 (
		_w17865_,
		_w17873_,
		_w17874_,
		_w17875_
	);
	LUT3 #(
		.INIT('h01)
	) name12049 (
		_w17779_,
		_w17795_,
		_w17869_,
		_w17876_
	);
	LUT2 #(
		.INIT('h2)
	) name12050 (
		_w17783_,
		_w17779_,
		_w17877_
	);
	LUT3 #(
		.INIT('h80)
	) name12051 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17878_
	);
	LUT4 #(
		.INIT('h0600)
	) name12052 (
		_w17781_,
		_w17784_,
		_w17783_,
		_w17779_,
		_w17879_
	);
	LUT4 #(
		.INIT('h153f)
	) name12053 (
		_w17800_,
		_w17877_,
		_w17878_,
		_w17879_,
		_w17880_
	);
	LUT4 #(
		.INIT('h5700)
	) name12054 (
		_w17780_,
		_w17875_,
		_w17876_,
		_w17880_,
		_w17881_
	);
	LUT3 #(
		.INIT('h65)
	) name12055 (
		\u1_L10_reg[24]/NET0131 ,
		_w17872_,
		_w17881_,
		_w17882_
	);
	LUT2 #(
		.INIT('h4)
	) name12056 (
		_w17849_,
		_w17852_,
		_w17883_
	);
	LUT4 #(
		.INIT('h0004)
	) name12057 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17884_
	);
	LUT3 #(
		.INIT('h08)
	) name12058 (
		_w17779_,
		_w17866_,
		_w17884_,
		_w17885_
	);
	LUT3 #(
		.INIT('ha8)
	) name12059 (
		_w17780_,
		_w17883_,
		_w17885_,
		_w17886_
	);
	LUT4 #(
		.INIT('h73af)
	) name12060 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17887_
	);
	LUT2 #(
		.INIT('h2)
	) name12061 (
		_w17779_,
		_w17887_,
		_w17888_
	);
	LUT2 #(
		.INIT('h1)
	) name12062 (
		_w17780_,
		_w17869_,
		_w17889_
	);
	LUT4 #(
		.INIT('h0200)
	) name12063 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17783_,
		_w17890_
	);
	LUT3 #(
		.INIT('hac)
	) name12064 (
		_w17781_,
		_w17784_,
		_w17782_,
		_w17891_
	);
	LUT3 #(
		.INIT('h13)
	) name12065 (
		_w17852_,
		_w17890_,
		_w17891_,
		_w17892_
	);
	LUT3 #(
		.INIT('h40)
	) name12066 (
		_w17888_,
		_w17889_,
		_w17892_,
		_w17893_
	);
	LUT2 #(
		.INIT('h2)
	) name12067 (
		_w17798_,
		_w17791_,
		_w17894_
	);
	LUT4 #(
		.INIT('h0040)
	) name12068 (
		_w17781_,
		_w17782_,
		_w17783_,
		_w17779_,
		_w17895_
	);
	LUT3 #(
		.INIT('h07)
	) name12069 (
		_w17792_,
		_w17860_,
		_w17895_,
		_w17896_
	);
	LUT2 #(
		.INIT('h4)
	) name12070 (
		_w17894_,
		_w17896_,
		_w17897_
	);
	LUT4 #(
		.INIT('h56aa)
	) name12071 (
		\u1_L10_reg[30]/NET0131 ,
		_w17886_,
		_w17893_,
		_w17897_,
		_w17898_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name12072 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17899_
	);
	LUT2 #(
		.INIT('h2)
	) name12073 (
		_w17486_,
		_w17899_,
		_w17900_
	);
	LUT4 #(
		.INIT('h0040)
	) name12074 (
		_w17488_,
		_w17489_,
		_w17487_,
		_w17486_,
		_w17901_
	);
	LUT4 #(
		.INIT('h0004)
	) name12075 (
		_w17510_,
		_w17485_,
		_w17500_,
		_w17901_,
		_w17902_
	);
	LUT4 #(
		.INIT('he3ef)
	) name12076 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17903_
	);
	LUT2 #(
		.INIT('h2)
	) name12077 (
		_w17486_,
		_w17903_,
		_w17904_
	);
	LUT4 #(
		.INIT('h5010)
	) name12078 (
		_w17491_,
		_w17488_,
		_w17489_,
		_w17487_,
		_w17905_
	);
	LUT3 #(
		.INIT('hd0)
	) name12079 (
		_w17491_,
		_w17487_,
		_w17486_,
		_w17906_
	);
	LUT4 #(
		.INIT('h5554)
	) name12080 (
		_w17485_,
		_w17490_,
		_w17906_,
		_w17905_,
		_w17907_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12081 (
		_w17900_,
		_w17902_,
		_w17904_,
		_w17907_,
		_w17908_
	);
	LUT3 #(
		.INIT('h02)
	) name12082 (
		_w17486_,
		_w17509_,
		_w17517_,
		_w17909_
	);
	LUT4 #(
		.INIT('h0001)
	) name12083 (
		_w17486_,
		_w17513_,
		_w17499_,
		_w17824_,
		_w17910_
	);
	LUT2 #(
		.INIT('h1)
	) name12084 (
		_w17909_,
		_w17910_,
		_w17911_
	);
	LUT3 #(
		.INIT('h56)
	) name12085 (
		\u1_L10_reg[3]/NET0131 ,
		_w17908_,
		_w17911_,
		_w17912_
	);
	LUT4 #(
		.INIT('h9060)
	) name12086 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17913_
	);
	LUT4 #(
		.INIT('h002a)
	) name12087 (
		_w17357_,
		_w17522_,
		_w17741_,
		_w17737_,
		_w17914_
	);
	LUT4 #(
		.INIT('he0f0)
	) name12088 (
		_w17353_,
		_w17354_,
		_w17350_,
		_w17352_,
		_w17915_
	);
	LUT2 #(
		.INIT('h4)
	) name12089 (
		_w17522_,
		_w17915_,
		_w17916_
	);
	LUT4 #(
		.INIT('h2010)
	) name12090 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17917_
	);
	LUT4 #(
		.INIT('h0109)
	) name12091 (
		_w17353_,
		_w17351_,
		_w17350_,
		_w17352_,
		_w17918_
	);
	LUT4 #(
		.INIT('h0800)
	) name12092 (
		_w17353_,
		_w17351_,
		_w17354_,
		_w17352_,
		_w17919_
	);
	LUT4 #(
		.INIT('h0001)
	) name12093 (
		_w17357_,
		_w17918_,
		_w17919_,
		_w17917_,
		_w17920_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12094 (
		_w17913_,
		_w17914_,
		_w17916_,
		_w17920_,
		_w17921_
	);
	LUT3 #(
		.INIT('h08)
	) name12095 (
		_w17353_,
		_w17351_,
		_w17350_,
		_w17922_
	);
	LUT2 #(
		.INIT('h4)
	) name12096 (
		_w17360_,
		_w17922_,
		_w17923_
	);
	LUT3 #(
		.INIT('h56)
	) name12097 (
		\u1_L10_reg[9]/NET0131 ,
		_w17921_,
		_w17923_,
		_w17924_
	);
	LUT4 #(
		.INIT('hd7fc)
	) name12098 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17925_
	);
	LUT4 #(
		.INIT('h8000)
	) name12099 (
		_w17621_,
		_w17617_,
		_w17618_,
		_w17619_,
		_w17926_
	);
	LUT4 #(
		.INIT('h1003)
	) name12100 (
		_w17621_,
		_w17617_,
		_w17619_,
		_w17616_,
		_w17927_
	);
	LUT4 #(
		.INIT('h5455)
	) name12101 (
		_w17632_,
		_w17926_,
		_w17927_,
		_w17925_,
		_w17928_
	);
	LUT4 #(
		.INIT('h0a20)
	) name12102 (
		_w17621_,
		_w17617_,
		_w17618_,
		_w17619_,
		_w17929_
	);
	LUT3 #(
		.INIT('he4)
	) name12103 (
		_w17618_,
		_w17619_,
		_w17616_,
		_w17930_
	);
	LUT4 #(
		.INIT('h0031)
	) name12104 (
		_w17624_,
		_w17676_,
		_w17930_,
		_w17929_,
		_w17931_
	);
	LUT4 #(
		.INIT('h1000)
	) name12105 (
		_w17621_,
		_w17617_,
		_w17618_,
		_w17619_,
		_w17932_
	);
	LUT4 #(
		.INIT('h77ef)
	) name12106 (
		_w17617_,
		_w17618_,
		_w17619_,
		_w17616_,
		_w17933_
	);
	LUT3 #(
		.INIT('h31)
	) name12107 (
		_w17621_,
		_w17932_,
		_w17933_,
		_w17934_
	);
	LUT4 #(
		.INIT('h0d00)
	) name12108 (
		_w17632_,
		_w17931_,
		_w17928_,
		_w17934_,
		_w17935_
	);
	LUT2 #(
		.INIT('h9)
	) name12109 (
		\u1_L10_reg[18]/P0001 ,
		_w17935_,
		_w17936_
	);
	LUT4 #(
		.INIT('hc963)
	) name12110 (
		decrypt_pad,
		\u1_R9_reg[4]/NET0131 ,
		\u1_uk_K_r9_reg[19]/NET0131 ,
		\u1_uk_K_r9_reg[25]/NET0131 ,
		_w17937_
	);
	LUT4 #(
		.INIT('hc963)
	) name12111 (
		decrypt_pad,
		\u1_R9_reg[3]/NET0131 ,
		\u1_uk_K_r9_reg[41]/NET0131 ,
		\u1_uk_K_r9_reg[47]/NET0131 ,
		_w17938_
	);
	LUT4 #(
		.INIT('hc963)
	) name12112 (
		decrypt_pad,
		\u1_R9_reg[5]/NET0131 ,
		\u1_uk_K_r9_reg[47]/NET0131 ,
		\u1_uk_K_r9_reg[53]/NET0131 ,
		_w17939_
	);
	LUT4 #(
		.INIT('hc963)
	) name12113 (
		decrypt_pad,
		\u1_R9_reg[1]/NET0131 ,
		\u1_uk_K_r9_reg[17]/NET0131 ,
		\u1_uk_K_r9_reg[55]/NET0131 ,
		_w17940_
	);
	LUT2 #(
		.INIT('h2)
	) name12114 (
		_w17939_,
		_w17940_,
		_w17941_
	);
	LUT4 #(
		.INIT('hc693)
	) name12115 (
		decrypt_pad,
		\u1_R9_reg[2]/NET0131 ,
		\u1_uk_K_r9_reg[13]/NET0131 ,
		\u1_uk_K_r9_reg[32]/NET0131 ,
		_w17942_
	);
	LUT4 #(
		.INIT('hc693)
	) name12116 (
		decrypt_pad,
		\u1_R9_reg[32]/NET0131 ,
		\u1_uk_K_r9_reg[34]/NET0131 ,
		\u1_uk_K_r9_reg[53]/NET0131 ,
		_w17943_
	);
	LUT4 #(
		.INIT('hfd0d)
	) name12117 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w17944_
	);
	LUT2 #(
		.INIT('h2)
	) name12118 (
		_w17938_,
		_w17944_,
		_w17945_
	);
	LUT2 #(
		.INIT('h9)
	) name12119 (
		_w17942_,
		_w17943_,
		_w17946_
	);
	LUT4 #(
		.INIT('h0026)
	) name12120 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w17947_
	);
	LUT2 #(
		.INIT('h4)
	) name12121 (
		_w17938_,
		_w17940_,
		_w17948_
	);
	LUT3 #(
		.INIT('h40)
	) name12122 (
		_w17938_,
		_w17943_,
		_w17940_,
		_w17949_
	);
	LUT2 #(
		.INIT('h4)
	) name12123 (
		_w17943_,
		_w17939_,
		_w17950_
	);
	LUT2 #(
		.INIT('h2)
	) name12124 (
		_w17938_,
		_w17942_,
		_w17951_
	);
	LUT3 #(
		.INIT('hd0)
	) name12125 (
		_w17938_,
		_w17942_,
		_w17940_,
		_w17952_
	);
	LUT4 #(
		.INIT('h0051)
	) name12126 (
		_w17949_,
		_w17950_,
		_w17952_,
		_w17947_,
		_w17953_
	);
	LUT3 #(
		.INIT('h8a)
	) name12127 (
		_w17937_,
		_w17945_,
		_w17953_,
		_w17954_
	);
	LUT2 #(
		.INIT('h6)
	) name12128 (
		_w17943_,
		_w17939_,
		_w17955_
	);
	LUT3 #(
		.INIT('h01)
	) name12129 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17956_
	);
	LUT4 #(
		.INIT('hf77c)
	) name12130 (
		_w17938_,
		_w17942_,
		_w17943_,
		_w17939_,
		_w17957_
	);
	LUT2 #(
		.INIT('h4)
	) name12131 (
		_w17957_,
		_w17940_,
		_w17958_
	);
	LUT3 #(
		.INIT('h40)
	) name12132 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17959_
	);
	LUT2 #(
		.INIT('h4)
	) name12133 (
		_w17948_,
		_w17959_,
		_w17960_
	);
	LUT2 #(
		.INIT('h2)
	) name12134 (
		_w17942_,
		_w17940_,
		_w17961_
	);
	LUT3 #(
		.INIT('hc4)
	) name12135 (
		_w17942_,
		_w17943_,
		_w17940_,
		_w17962_
	);
	LUT3 #(
		.INIT('h51)
	) name12136 (
		_w17938_,
		_w17942_,
		_w17943_,
		_w17963_
	);
	LUT3 #(
		.INIT('h10)
	) name12137 (
		_w17941_,
		_w17962_,
		_w17963_,
		_w17964_
	);
	LUT4 #(
		.INIT('h00fe)
	) name12138 (
		_w17958_,
		_w17960_,
		_w17964_,
		_w17937_,
		_w17965_
	);
	LUT4 #(
		.INIT('h7adf)
	) name12139 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w17966_
	);
	LUT2 #(
		.INIT('h1)
	) name12140 (
		_w17938_,
		_w17966_,
		_w17967_
	);
	LUT3 #(
		.INIT('h02)
	) name12141 (
		_w17938_,
		_w17943_,
		_w17939_,
		_w17968_
	);
	LUT4 #(
		.INIT('h0020)
	) name12142 (
		_w17938_,
		_w17942_,
		_w17943_,
		_w17940_,
		_w17969_
	);
	LUT3 #(
		.INIT('h07)
	) name12143 (
		_w17961_,
		_w17968_,
		_w17969_,
		_w17970_
	);
	LUT2 #(
		.INIT('h4)
	) name12144 (
		_w17967_,
		_w17970_,
		_w17971_
	);
	LUT4 #(
		.INIT('h5655)
	) name12145 (
		\u1_L9_reg[31]/NET0131 ,
		_w17965_,
		_w17954_,
		_w17971_,
		_w17972_
	);
	LUT4 #(
		.INIT('hc963)
	) name12146 (
		decrypt_pad,
		\u1_R9_reg[24]/NET0131 ,
		\u1_uk_K_r9_reg[43]/NET0131 ,
		\u1_uk_K_r9_reg[51]/NET0131 ,
		_w17973_
	);
	LUT4 #(
		.INIT('hc963)
	) name12147 (
		decrypt_pad,
		\u1_R9_reg[23]/NET0131 ,
		\u1_uk_K_r9_reg[45]/NET0131 ,
		\u1_uk_K_r9_reg[49]/NET0131 ,
		_w17974_
	);
	LUT4 #(
		.INIT('hc963)
	) name12148 (
		decrypt_pad,
		\u1_R9_reg[22]/NET0131 ,
		\u1_uk_K_r9_reg[28]/NET0131 ,
		\u1_uk_K_r9_reg[36]/NET0131 ,
		_w17975_
	);
	LUT4 #(
		.INIT('hc963)
	) name12149 (
		decrypt_pad,
		\u1_R9_reg[20]/NET0131 ,
		\u1_uk_K_r9_reg[22]/NET0131 ,
		\u1_uk_K_r9_reg[30]/NET0131 ,
		_w17976_
	);
	LUT4 #(
		.INIT('hc693)
	) name12150 (
		decrypt_pad,
		\u1_R9_reg[21]/NET0131 ,
		\u1_uk_K_r9_reg[14]/NET0131 ,
		\u1_uk_K_r9_reg[37]/NET0131 ,
		_w17977_
	);
	LUT4 #(
		.INIT('h4555)
	) name12151 (
		_w17974_,
		_w17976_,
		_w17977_,
		_w17975_,
		_w17978_
	);
	LUT4 #(
		.INIT('h1862)
	) name12152 (
		_w17974_,
		_w17976_,
		_w17977_,
		_w17975_,
		_w17979_
	);
	LUT4 #(
		.INIT('hc693)
	) name12153 (
		decrypt_pad,
		\u1_R9_reg[25]/NET0131 ,
		\u1_uk_K_r9_reg[15]/NET0131 ,
		\u1_uk_K_r9_reg[7]/NET0131 ,
		_w17980_
	);
	LUT4 #(
		.INIT('h0004)
	) name12154 (
		_w17974_,
		_w17976_,
		_w17980_,
		_w17975_,
		_w17981_
	);
	LUT4 #(
		.INIT('h0800)
	) name12155 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w17982_
	);
	LUT4 #(
		.INIT('h0020)
	) name12156 (
		_w17974_,
		_w17976_,
		_w17980_,
		_w17977_,
		_w17983_
	);
	LUT4 #(
		.INIT('h0020)
	) name12157 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w17984_
	);
	LUT4 #(
		.INIT('h0001)
	) name12158 (
		_w17983_,
		_w17981_,
		_w17982_,
		_w17984_,
		_w17985_
	);
	LUT3 #(
		.INIT('h45)
	) name12159 (
		_w17973_,
		_w17979_,
		_w17985_,
		_w17986_
	);
	LUT4 #(
		.INIT('h0002)
	) name12160 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w17987_
	);
	LUT4 #(
		.INIT('h2f7d)
	) name12161 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w17988_
	);
	LUT2 #(
		.INIT('h2)
	) name12162 (
		_w17974_,
		_w17988_,
		_w17989_
	);
	LUT4 #(
		.INIT('h00b7)
	) name12163 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w17990_
	);
	LUT3 #(
		.INIT('h80)
	) name12164 (
		_w17976_,
		_w17980_,
		_w17975_,
		_w17991_
	);
	LUT3 #(
		.INIT('h02)
	) name12165 (
		_w17978_,
		_w17991_,
		_w17990_,
		_w17992_
	);
	LUT3 #(
		.INIT('hde)
	) name12166 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17993_
	);
	LUT4 #(
		.INIT('h0004)
	) name12167 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w17994_
	);
	LUT4 #(
		.INIT('h77eb)
	) name12168 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w17995_
	);
	LUT4 #(
		.INIT('hfe54)
	) name12169 (
		_w17974_,
		_w17975_,
		_w17993_,
		_w17995_,
		_w17996_
	);
	LUT4 #(
		.INIT('h5700)
	) name12170 (
		_w17973_,
		_w17989_,
		_w17992_,
		_w17996_,
		_w17997_
	);
	LUT3 #(
		.INIT('h9a)
	) name12171 (
		\u1_L9_reg[11]/NET0131 ,
		_w17986_,
		_w17997_,
		_w17998_
	);
	LUT4 #(
		.INIT('hc693)
	) name12172 (
		decrypt_pad,
		\u1_R9_reg[28]/NET0131 ,
		\u1_uk_K_r9_reg[31]/P0001 ,
		\u1_uk_K_r9_reg[50]/NET0131 ,
		_w17999_
	);
	LUT4 #(
		.INIT('hc963)
	) name12173 (
		decrypt_pad,
		\u1_R9_reg[26]/NET0131 ,
		\u1_uk_K_r9_reg[30]/NET0131 ,
		\u1_uk_K_r9_reg[7]/NET0131 ,
		_w18000_
	);
	LUT4 #(
		.INIT('hc963)
	) name12174 (
		decrypt_pad,
		\u1_R9_reg[25]/NET0131 ,
		\u1_uk_K_r9_reg[14]/NET0131 ,
		\u1_uk_K_r9_reg[22]/NET0131 ,
		_w18001_
	);
	LUT4 #(
		.INIT('hc963)
	) name12175 (
		decrypt_pad,
		\u1_R9_reg[29]/NET0131 ,
		\u1_uk_K_r9_reg[42]/NET0131 ,
		\u1_uk_K_r9_reg[50]/NET0131 ,
		_w18002_
	);
	LUT3 #(
		.INIT('hea)
	) name12176 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18003_
	);
	LUT4 #(
		.INIT('hc963)
	) name12177 (
		decrypt_pad,
		\u1_R9_reg[24]/NET0131 ,
		\u1_uk_K_r9_reg[38]/NET0131 ,
		\u1_uk_K_r9_reg[42]/NET0131 ,
		_w18004_
	);
	LUT4 #(
		.INIT('hc693)
	) name12178 (
		decrypt_pad,
		\u1_R9_reg[27]/NET0131 ,
		\u1_uk_K_r9_reg[16]/NET0131 ,
		\u1_uk_K_r9_reg[8]/NET0131 ,
		_w18005_
	);
	LUT3 #(
		.INIT('h70)
	) name12179 (
		_w18000_,
		_w18001_,
		_w18005_,
		_w18006_
	);
	LUT4 #(
		.INIT('h7000)
	) name12180 (
		_w18000_,
		_w18001_,
		_w18004_,
		_w18005_,
		_w18007_
	);
	LUT2 #(
		.INIT('h8)
	) name12181 (
		_w18003_,
		_w18007_,
		_w18008_
	);
	LUT4 #(
		.INIT('h1000)
	) name12182 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18009_
	);
	LUT4 #(
		.INIT('hef3f)
	) name12183 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18010_
	);
	LUT2 #(
		.INIT('h2)
	) name12184 (
		_w18002_,
		_w18004_,
		_w18011_
	);
	LUT4 #(
		.INIT('h0020)
	) name12185 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18012_
	);
	LUT4 #(
		.INIT('hffde)
	) name12186 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18013_
	);
	LUT3 #(
		.INIT('he0)
	) name12187 (
		_w18005_,
		_w18010_,
		_w18013_,
		_w18014_
	);
	LUT3 #(
		.INIT('h8a)
	) name12188 (
		_w17999_,
		_w18008_,
		_w18014_,
		_w18015_
	);
	LUT4 #(
		.INIT('h0072)
	) name12189 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18005_,
		_w18016_
	);
	LUT4 #(
		.INIT('h10f0)
	) name12190 (
		_w18000_,
		_w18001_,
		_w18004_,
		_w18005_,
		_w18017_
	);
	LUT2 #(
		.INIT('h4)
	) name12191 (
		_w18016_,
		_w18017_,
		_w18018_
	);
	LUT4 #(
		.INIT('h0002)
	) name12192 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18019_
	);
	LUT2 #(
		.INIT('h6)
	) name12193 (
		_w18000_,
		_w18004_,
		_w18020_
	);
	LUT3 #(
		.INIT('h8c)
	) name12194 (
		_w18001_,
		_w18002_,
		_w18005_,
		_w18021_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name12195 (
		_w18019_,
		_w18005_,
		_w18020_,
		_w18021_,
		_w18022_
	);
	LUT4 #(
		.INIT('h0008)
	) name12196 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18023_
	);
	LUT4 #(
		.INIT('hfcd7)
	) name12197 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18024_
	);
	LUT4 #(
		.INIT('h0084)
	) name12198 (
		_w18000_,
		_w18001_,
		_w18004_,
		_w18005_,
		_w18025_
	);
	LUT4 #(
		.INIT('h0100)
	) name12199 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18005_,
		_w18026_
	);
	LUT4 #(
		.INIT('h0031)
	) name12200 (
		_w18005_,
		_w18025_,
		_w18024_,
		_w18026_,
		_w18027_
	);
	LUT4 #(
		.INIT('hba00)
	) name12201 (
		_w17999_,
		_w18018_,
		_w18022_,
		_w18027_,
		_w18028_
	);
	LUT3 #(
		.INIT('h65)
	) name12202 (
		\u1_L9_reg[22]/NET0131 ,
		_w18015_,
		_w18028_,
		_w18029_
	);
	LUT4 #(
		.INIT('hc693)
	) name12203 (
		decrypt_pad,
		\u1_R9_reg[13]/NET0131 ,
		\u1_uk_K_r9_reg[10]/NET0131 ,
		\u1_uk_K_r9_reg[4]/NET0131 ,
		_w18030_
	);
	LUT4 #(
		.INIT('hc963)
	) name12204 (
		decrypt_pad,
		\u1_R9_reg[15]/NET0131 ,
		\u1_uk_K_r9_reg[13]/NET0131 ,
		\u1_uk_K_r9_reg[19]/NET0131 ,
		_w18031_
	);
	LUT4 #(
		.INIT('hc963)
	) name12205 (
		decrypt_pad,
		\u1_R9_reg[12]/NET0131 ,
		\u1_uk_K_r9_reg[10]/NET0131 ,
		\u1_uk_K_r9_reg[48]/NET0131 ,
		_w18032_
	);
	LUT4 #(
		.INIT('hc693)
	) name12206 (
		decrypt_pad,
		\u1_R9_reg[14]/NET0131 ,
		\u1_uk_K_r9_reg[11]/NET0131 ,
		\u1_uk_K_r9_reg[5]/NET0131 ,
		_w18033_
	);
	LUT4 #(
		.INIT('h4000)
	) name12207 (
		_w18032_,
		_w18030_,
		_w18031_,
		_w18033_,
		_w18034_
	);
	LUT4 #(
		.INIT('hc693)
	) name12208 (
		decrypt_pad,
		\u1_R9_reg[16]/NET0131 ,
		\u1_uk_K_r9_reg[27]/P0001 ,
		\u1_uk_K_r9_reg[46]/NET0131 ,
		_w18035_
	);
	LUT2 #(
		.INIT('h1)
	) name12209 (
		_w18034_,
		_w18035_,
		_w18036_
	);
	LUT4 #(
		.INIT('hc963)
	) name12210 (
		decrypt_pad,
		\u1_R9_reg[17]/NET0131 ,
		\u1_uk_K_r9_reg[26]/NET0131 ,
		\u1_uk_K_r9_reg[32]/NET0131 ,
		_w18037_
	);
	LUT4 #(
		.INIT('h8000)
	) name12211 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18031_,
		_w18038_
	);
	LUT4 #(
		.INIT('h0008)
	) name12212 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18039_
	);
	LUT2 #(
		.INIT('h4)
	) name12213 (
		_w18030_,
		_w18031_,
		_w18040_
	);
	LUT4 #(
		.INIT('h0100)
	) name12214 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18031_,
		_w18041_
	);
	LUT3 #(
		.INIT('h01)
	) name12215 (
		_w18039_,
		_w18041_,
		_w18038_,
		_w18042_
	);
	LUT2 #(
		.INIT('h2)
	) name12216 (
		_w18032_,
		_w18037_,
		_w18043_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name12217 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18044_
	);
	LUT2 #(
		.INIT('h4)
	) name12218 (
		_w18032_,
		_w18030_,
		_w18045_
	);
	LUT2 #(
		.INIT('h4)
	) name12219 (
		_w18037_,
		_w18033_,
		_w18046_
	);
	LUT4 #(
		.INIT('h1000)
	) name12220 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18047_
	);
	LUT4 #(
		.INIT('heffe)
	) name12221 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18048_
	);
	LUT3 #(
		.INIT('he0)
	) name12222 (
		_w18031_,
		_w18044_,
		_w18048_,
		_w18049_
	);
	LUT3 #(
		.INIT('h80)
	) name12223 (
		_w18036_,
		_w18042_,
		_w18049_,
		_w18050_
	);
	LUT2 #(
		.INIT('h1)
	) name12224 (
		_w18030_,
		_w18031_,
		_w18051_
	);
	LUT4 #(
		.INIT('h0001)
	) name12225 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18031_,
		_w18052_
	);
	LUT4 #(
		.INIT('h7f7e)
	) name12226 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18031_,
		_w18053_
	);
	LUT2 #(
		.INIT('h2)
	) name12227 (
		_w18033_,
		_w18053_,
		_w18054_
	);
	LUT2 #(
		.INIT('h9)
	) name12228 (
		_w18032_,
		_w18030_,
		_w18055_
	);
	LUT4 #(
		.INIT('h0006)
	) name12229 (
		_w18032_,
		_w18030_,
		_w18031_,
		_w18033_,
		_w18056_
	);
	LUT4 #(
		.INIT('h2000)
	) name12230 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18031_,
		_w18057_
	);
	LUT4 #(
		.INIT('h0040)
	) name12231 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18058_
	);
	LUT2 #(
		.INIT('h4)
	) name12232 (
		_w18032_,
		_w18037_,
		_w18059_
	);
	LUT4 #(
		.INIT('h0400)
	) name12233 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18031_,
		_w18060_
	);
	LUT4 #(
		.INIT('h0004)
	) name12234 (
		_w18057_,
		_w18035_,
		_w18058_,
		_w18060_,
		_w18061_
	);
	LUT3 #(
		.INIT('h10)
	) name12235 (
		_w18056_,
		_w18054_,
		_w18061_,
		_w18062_
	);
	LUT3 #(
		.INIT('hde)
	) name12236 (
		_w18032_,
		_w18037_,
		_w18033_,
		_w18063_
	);
	LUT2 #(
		.INIT('h2)
	) name12237 (
		_w18040_,
		_w18063_,
		_w18064_
	);
	LUT3 #(
		.INIT('h02)
	) name12238 (
		_w18037_,
		_w18031_,
		_w18033_,
		_w18065_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name12239 (
		_w18057_,
		_w18033_,
		_w18045_,
		_w18065_,
		_w18066_
	);
	LUT2 #(
		.INIT('h4)
	) name12240 (
		_w18064_,
		_w18066_,
		_w18067_
	);
	LUT4 #(
		.INIT('ha955)
	) name12241 (
		\u1_L9_reg[20]/NET0131 ,
		_w18050_,
		_w18062_,
		_w18067_,
		_w18068_
	);
	LUT4 #(
		.INIT('hc963)
	) name12242 (
		decrypt_pad,
		\u1_R9_reg[6]/NET0131 ,
		\u1_uk_K_r9_reg[3]/NET0131 ,
		\u1_uk_K_r9_reg[41]/NET0131 ,
		_w18069_
	);
	LUT4 #(
		.INIT('hc963)
	) name12243 (
		decrypt_pad,
		\u1_R9_reg[9]/NET0131 ,
		\u1_uk_K_r9_reg[25]/NET0131 ,
		\u1_uk_K_r9_reg[6]/NET0131 ,
		_w18070_
	);
	LUT4 #(
		.INIT('hc963)
	) name12244 (
		decrypt_pad,
		\u1_R9_reg[5]/NET0131 ,
		\u1_uk_K_r9_reg[12]/NET0131 ,
		\u1_uk_K_r9_reg[18]/NET0131 ,
		_w18071_
	);
	LUT4 #(
		.INIT('hc963)
	) name12245 (
		decrypt_pad,
		\u1_R9_reg[4]/NET0131 ,
		\u1_uk_K_r9_reg[33]/NET0131 ,
		\u1_uk_K_r9_reg[39]/NET0131 ,
		_w18072_
	);
	LUT4 #(
		.INIT('h0310)
	) name12246 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18073_
	);
	LUT4 #(
		.INIT('hc693)
	) name12247 (
		decrypt_pad,
		\u1_R9_reg[7]/NET0131 ,
		\u1_uk_K_r9_reg[3]/NET0131 ,
		\u1_uk_K_r9_reg[54]/NET0131 ,
		_w18074_
	);
	LUT4 #(
		.INIT('h0010)
	) name12248 (
		_w18074_,
		_w18072_,
		_w18070_,
		_w18071_,
		_w18075_
	);
	LUT4 #(
		.INIT('hc963)
	) name12249 (
		decrypt_pad,
		\u1_R9_reg[8]/NET0131 ,
		\u1_uk_K_r9_reg[20]/NET0131 ,
		\u1_uk_K_r9_reg[26]/NET0131 ,
		_w18076_
	);
	LUT3 #(
		.INIT('h01)
	) name12250 (
		_w18075_,
		_w18073_,
		_w18076_,
		_w18077_
	);
	LUT2 #(
		.INIT('h4)
	) name12251 (
		_w18069_,
		_w18070_,
		_w18078_
	);
	LUT4 #(
		.INIT('h0010)
	) name12252 (
		_w18074_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18079_
	);
	LUT4 #(
		.INIT('h4000)
	) name12253 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18080_
	);
	LUT2 #(
		.INIT('h8)
	) name12254 (
		_w18072_,
		_w18069_,
		_w18081_
	);
	LUT3 #(
		.INIT('h51)
	) name12255 (
		_w18074_,
		_w18070_,
		_w18071_,
		_w18082_
	);
	LUT3 #(
		.INIT('ha6)
	) name12256 (
		_w18074_,
		_w18070_,
		_w18071_,
		_w18083_
	);
	LUT4 #(
		.INIT('h1101)
	) name12257 (
		_w18079_,
		_w18080_,
		_w18081_,
		_w18083_,
		_w18084_
	);
	LUT2 #(
		.INIT('h8)
	) name12258 (
		_w18077_,
		_w18084_,
		_w18085_
	);
	LUT2 #(
		.INIT('h4)
	) name12259 (
		_w18072_,
		_w18069_,
		_w18086_
	);
	LUT2 #(
		.INIT('h8)
	) name12260 (
		_w18074_,
		_w18071_,
		_w18087_
	);
	LUT4 #(
		.INIT('h0002)
	) name12261 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18088_
	);
	LUT3 #(
		.INIT('h54)
	) name12262 (
		_w18086_,
		_w18087_,
		_w18088_,
		_w18089_
	);
	LUT2 #(
		.INIT('h8)
	) name12263 (
		_w18072_,
		_w18070_,
		_w18090_
	);
	LUT2 #(
		.INIT('h6)
	) name12264 (
		_w18072_,
		_w18070_,
		_w18091_
	);
	LUT4 #(
		.INIT('h1050)
	) name12265 (
		_w18074_,
		_w18072_,
		_w18069_,
		_w18071_,
		_w18092_
	);
	LUT2 #(
		.INIT('h4)
	) name12266 (
		_w18091_,
		_w18092_,
		_w18093_
	);
	LUT2 #(
		.INIT('h2)
	) name12267 (
		_w18072_,
		_w18069_,
		_w18094_
	);
	LUT4 #(
		.INIT('h2000)
	) name12268 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18095_
	);
	LUT4 #(
		.INIT('h0001)
	) name12269 (
		_w18074_,
		_w18072_,
		_w18070_,
		_w18071_,
		_w18096_
	);
	LUT3 #(
		.INIT('h02)
	) name12270 (
		_w18076_,
		_w18095_,
		_w18096_,
		_w18097_
	);
	LUT3 #(
		.INIT('h10)
	) name12271 (
		_w18093_,
		_w18089_,
		_w18097_,
		_w18098_
	);
	LUT4 #(
		.INIT('h0004)
	) name12272 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18099_
	);
	LUT4 #(
		.INIT('hddfb)
	) name12273 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18100_
	);
	LUT3 #(
		.INIT('hba)
	) name12274 (
		_w18074_,
		_w18069_,
		_w18071_,
		_w18101_
	);
	LUT4 #(
		.INIT('h5010)
	) name12275 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18102_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name12276 (
		_w18074_,
		_w18100_,
		_w18101_,
		_w18102_,
		_w18103_
	);
	LUT4 #(
		.INIT('ha955)
	) name12277 (
		\u1_L9_reg[2]/NET0131 ,
		_w18085_,
		_w18098_,
		_w18103_,
		_w18104_
	);
	LUT4 #(
		.INIT('hdf27)
	) name12278 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18105_
	);
	LUT4 #(
		.INIT('h6d7c)
	) name12279 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18106_
	);
	LUT4 #(
		.INIT('h0400)
	) name12280 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18107_
	);
	LUT4 #(
		.INIT('h00d8)
	) name12281 (
		_w17974_,
		_w18106_,
		_w18105_,
		_w18107_,
		_w18108_
	);
	LUT2 #(
		.INIT('h1)
	) name12282 (
		_w17973_,
		_w18108_,
		_w18109_
	);
	LUT4 #(
		.INIT('h9faf)
	) name12283 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18110_
	);
	LUT2 #(
		.INIT('h2)
	) name12284 (
		_w17974_,
		_w18110_,
		_w18111_
	);
	LUT4 #(
		.INIT('h66fe)
	) name12285 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18112_
	);
	LUT2 #(
		.INIT('h1)
	) name12286 (
		_w17974_,
		_w18112_,
		_w18113_
	);
	LUT4 #(
		.INIT('hfefb)
	) name12287 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18114_
	);
	LUT3 #(
		.INIT('h10)
	) name12288 (
		_w17981_,
		_w17982_,
		_w18114_,
		_w18115_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name12289 (
		_w17973_,
		_w18111_,
		_w18113_,
		_w18115_,
		_w18116_
	);
	LUT4 #(
		.INIT('h0080)
	) name12290 (
		_w17974_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18117_
	);
	LUT2 #(
		.INIT('h1)
	) name12291 (
		_w17987_,
		_w18117_,
		_w18118_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name12292 (
		\u1_L9_reg[29]/NET0131 ,
		_w18116_,
		_w18109_,
		_w18118_,
		_w18119_
	);
	LUT4 #(
		.INIT('hd79b)
	) name12293 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18120_
	);
	LUT4 #(
		.INIT('h6100)
	) name12294 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18121_
	);
	LUT4 #(
		.INIT('hcc04)
	) name12295 (
		_w17973_,
		_w17974_,
		_w18120_,
		_w18121_,
		_w18122_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12296 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18123_
	);
	LUT4 #(
		.INIT('h7dee)
	) name12297 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18124_
	);
	LUT4 #(
		.INIT('h0233)
	) name12298 (
		_w17973_,
		_w17974_,
		_w18123_,
		_w18124_,
		_w18125_
	);
	LUT4 #(
		.INIT('heb67)
	) name12299 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18126_
	);
	LUT4 #(
		.INIT('h5051)
	) name12300 (
		_w17973_,
		_w17974_,
		_w17987_,
		_w18126_,
		_w18127_
	);
	LUT4 #(
		.INIT('h0080)
	) name12301 (
		_w17974_,
		_w17976_,
		_w17980_,
		_w17975_,
		_w18128_
	);
	LUT4 #(
		.INIT('h3fef)
	) name12302 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18129_
	);
	LUT3 #(
		.INIT('h8a)
	) name12303 (
		_w17973_,
		_w18128_,
		_w18129_,
		_w18130_
	);
	LUT4 #(
		.INIT('h0001)
	) name12304 (
		_w18122_,
		_w18127_,
		_w18125_,
		_w18130_,
		_w18131_
	);
	LUT2 #(
		.INIT('h9)
	) name12305 (
		\u1_L9_reg[4]/NET0131 ,
		_w18131_,
		_w18132_
	);
	LUT4 #(
		.INIT('hc963)
	) name12306 (
		decrypt_pad,
		\u1_R9_reg[32]/NET0131 ,
		\u1_uk_K_r9_reg[15]/NET0131 ,
		\u1_uk_K_r9_reg[23]/NET0131 ,
		_w18133_
	);
	LUT4 #(
		.INIT('hc693)
	) name12307 (
		decrypt_pad,
		\u1_R9_reg[31]/NET0131 ,
		\u1_uk_K_r9_reg[45]/NET0131 ,
		\u1_uk_K_r9_reg[9]/NET0131 ,
		_w18134_
	);
	LUT4 #(
		.INIT('hc693)
	) name12308 (
		decrypt_pad,
		\u1_R9_reg[29]/NET0131 ,
		\u1_uk_K_r9_reg[28]/NET0131 ,
		\u1_uk_K_r9_reg[51]/NET0131 ,
		_w18135_
	);
	LUT4 #(
		.INIT('hc963)
	) name12309 (
		decrypt_pad,
		\u1_R9_reg[1]/NET0131 ,
		\u1_uk_K_r9_reg[36]/NET0131 ,
		\u1_uk_K_r9_reg[44]/NET0131 ,
		_w18136_
	);
	LUT4 #(
		.INIT('hc963)
	) name12310 (
		decrypt_pad,
		\u1_R9_reg[30]/NET0131 ,
		\u1_uk_K_r9_reg[21]/NET0131 ,
		\u1_uk_K_r9_reg[29]/NET0131 ,
		_w18137_
	);
	LUT4 #(
		.INIT('hc693)
	) name12311 (
		decrypt_pad,
		\u1_R9_reg[28]/NET0131 ,
		\u1_uk_K_r9_reg[1]/NET0131 ,
		\u1_uk_K_r9_reg[52]/NET0131 ,
		_w18138_
	);
	LUT3 #(
		.INIT('h08)
	) name12312 (
		_w18138_,
		_w18136_,
		_w18137_,
		_w18139_
	);
	LUT4 #(
		.INIT('hf359)
	) name12313 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18140_
	);
	LUT3 #(
		.INIT('h01)
	) name12314 (
		_w18138_,
		_w18135_,
		_w18137_,
		_w18141_
	);
	LUT4 #(
		.INIT('h4000)
	) name12315 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18142_
	);
	LUT4 #(
		.INIT('h008d)
	) name12316 (
		_w18134_,
		_w18140_,
		_w18141_,
		_w18142_,
		_w18143_
	);
	LUT2 #(
		.INIT('h2)
	) name12317 (
		_w18133_,
		_w18143_,
		_w18144_
	);
	LUT2 #(
		.INIT('h1)
	) name12318 (
		_w18137_,
		_w18134_,
		_w18145_
	);
	LUT4 #(
		.INIT('h7d70)
	) name12319 (
		_w18135_,
		_w18136_,
		_w18137_,
		_w18134_,
		_w18146_
	);
	LUT2 #(
		.INIT('h2)
	) name12320 (
		_w18138_,
		_w18146_,
		_w18147_
	);
	LUT4 #(
		.INIT('h0200)
	) name12321 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18148_
	);
	LUT4 #(
		.INIT('hef00)
	) name12322 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18134_,
		_w18149_
	);
	LUT3 #(
		.INIT('h10)
	) name12323 (
		_w18138_,
		_w18136_,
		_w18137_,
		_w18150_
	);
	LUT3 #(
		.INIT('h07)
	) name12324 (
		_w18135_,
		_w18136_,
		_w18134_,
		_w18151_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12325 (
		_w18148_,
		_w18149_,
		_w18150_,
		_w18151_,
		_w18152_
	);
	LUT3 #(
		.INIT('h0e)
	) name12326 (
		_w18147_,
		_w18152_,
		_w18133_,
		_w18153_
	);
	LUT4 #(
		.INIT('h0400)
	) name12327 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18154_
	);
	LUT4 #(
		.INIT('hfbdf)
	) name12328 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18155_
	);
	LUT4 #(
		.INIT('h1000)
	) name12329 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18156_
	);
	LUT4 #(
		.INIT('h0001)
	) name12330 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18157_
	);
	LUT4 #(
		.INIT('hebde)
	) name12331 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18158_
	);
	LUT2 #(
		.INIT('h2)
	) name12332 (
		_w18134_,
		_w18158_,
		_w18159_
	);
	LUT3 #(
		.INIT('h20)
	) name12333 (
		_w18138_,
		_w18135_,
		_w18133_,
		_w18160_
	);
	LUT3 #(
		.INIT('h08)
	) name12334 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18161_
	);
	LUT4 #(
		.INIT('hcedf)
	) name12335 (
		_w18137_,
		_w18134_,
		_w18160_,
		_w18161_,
		_w18162_
	);
	LUT2 #(
		.INIT('h4)
	) name12336 (
		_w18159_,
		_w18162_,
		_w18163_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name12337 (
		\u1_L9_reg[5]/NET0131 ,
		_w18153_,
		_w18144_,
		_w18163_,
		_w18164_
	);
	LUT4 #(
		.INIT('h8400)
	) name12338 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18165_
	);
	LUT4 #(
		.INIT('hefe7)
	) name12339 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18166_
	);
	LUT2 #(
		.INIT('h2)
	) name12340 (
		_w18031_,
		_w18166_,
		_w18167_
	);
	LUT3 #(
		.INIT('h31)
	) name12341 (
		_w18030_,
		_w18031_,
		_w18033_,
		_w18168_
	);
	LUT4 #(
		.INIT('h153f)
	) name12342 (
		_w18043_,
		_w18045_,
		_w18065_,
		_w18168_,
		_w18169_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name12343 (
		_w18035_,
		_w18167_,
		_w18165_,
		_w18169_,
		_w18170_
	);
	LUT3 #(
		.INIT('h08)
	) name12344 (
		_w18037_,
		_w18031_,
		_w18033_,
		_w18171_
	);
	LUT4 #(
		.INIT('h0040)
	) name12345 (
		_w18032_,
		_w18037_,
		_w18031_,
		_w18033_,
		_w18172_
	);
	LUT3 #(
		.INIT('ha2)
	) name12346 (
		_w18032_,
		_w18037_,
		_w18033_,
		_w18173_
	);
	LUT4 #(
		.INIT('h0013)
	) name12347 (
		_w18040_,
		_w18052_,
		_w18173_,
		_w18172_,
		_w18174_
	);
	LUT4 #(
		.INIT('hff31)
	) name12348 (
		_w18037_,
		_w18030_,
		_w18031_,
		_w18033_,
		_w18175_
	);
	LUT3 #(
		.INIT('hc4)
	) name12349 (
		_w18032_,
		_w18048_,
		_w18175_,
		_w18176_
	);
	LUT3 #(
		.INIT('h15)
	) name12350 (
		_w18035_,
		_w18174_,
		_w18176_,
		_w18177_
	);
	LUT4 #(
		.INIT('h7bfe)
	) name12351 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18178_
	);
	LUT2 #(
		.INIT('h1)
	) name12352 (
		_w18031_,
		_w18178_,
		_w18179_
	);
	LUT3 #(
		.INIT('h0d)
	) name12353 (
		_w18057_,
		_w18033_,
		_w18034_,
		_w18180_
	);
	LUT2 #(
		.INIT('h4)
	) name12354 (
		_w18179_,
		_w18180_,
		_w18181_
	);
	LUT4 #(
		.INIT('h5655)
	) name12355 (
		\u1_L9_reg[10]/NET0131 ,
		_w18177_,
		_w18170_,
		_w18181_,
		_w18182_
	);
	LUT4 #(
		.INIT('h0006)
	) name12356 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18183_
	);
	LUT3 #(
		.INIT('h47)
	) name12357 (
		_w18000_,
		_w18001_,
		_w18005_,
		_w18184_
	);
	LUT4 #(
		.INIT('h0051)
	) name12358 (
		_w17999_,
		_w18011_,
		_w18184_,
		_w18183_,
		_w18185_
	);
	LUT3 #(
		.INIT('h10)
	) name12359 (
		_w18000_,
		_w18002_,
		_w18004_,
		_w18186_
	);
	LUT4 #(
		.INIT('h2100)
	) name12360 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18187_
	);
	LUT2 #(
		.INIT('h6)
	) name12361 (
		_w18001_,
		_w18002_,
		_w18188_
	);
	LUT4 #(
		.INIT('h143c)
	) name12362 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18189_
	);
	LUT3 #(
		.INIT('h32)
	) name12363 (
		_w18005_,
		_w18187_,
		_w18189_,
		_w18190_
	);
	LUT2 #(
		.INIT('h8)
	) name12364 (
		_w18185_,
		_w18190_,
		_w18191_
	);
	LUT2 #(
		.INIT('h4)
	) name12365 (
		_w18005_,
		_w18012_,
		_w18192_
	);
	LUT3 #(
		.INIT('h02)
	) name12366 (
		_w17999_,
		_w18009_,
		_w18023_,
		_w18193_
	);
	LUT4 #(
		.INIT('h0240)
	) name12367 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18194_
	);
	LUT4 #(
		.INIT('h33fe)
	) name12368 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18195_
	);
	LUT3 #(
		.INIT('h31)
	) name12369 (
		_w18005_,
		_w18194_,
		_w18195_,
		_w18196_
	);
	LUT3 #(
		.INIT('h40)
	) name12370 (
		_w18192_,
		_w18193_,
		_w18196_,
		_w18197_
	);
	LUT3 #(
		.INIT('ha9)
	) name12371 (
		\u1_L9_reg[12]/NET0131 ,
		_w18191_,
		_w18197_,
		_w18198_
	);
	LUT4 #(
		.INIT('haaa2)
	) name12372 (
		_w18074_,
		_w18072_,
		_w18070_,
		_w18071_,
		_w18199_
	);
	LUT4 #(
		.INIT('hfd50)
	) name12373 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18200_
	);
	LUT2 #(
		.INIT('h2)
	) name12374 (
		_w18199_,
		_w18200_,
		_w18201_
	);
	LUT3 #(
		.INIT('h32)
	) name12375 (
		_w18074_,
		_w18072_,
		_w18071_,
		_w18202_
	);
	LUT2 #(
		.INIT('h8)
	) name12376 (
		_w18078_,
		_w18202_,
		_w18203_
	);
	LUT3 #(
		.INIT('h8a)
	) name12377 (
		_w18074_,
		_w18070_,
		_w18071_,
		_w18204_
	);
	LUT3 #(
		.INIT('h13)
	) name12378 (
		_w18081_,
		_w18076_,
		_w18204_,
		_w18205_
	);
	LUT3 #(
		.INIT('h10)
	) name12379 (
		_w18201_,
		_w18203_,
		_w18205_,
		_w18206_
	);
	LUT4 #(
		.INIT('h00ac)
	) name12380 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18207_
	);
	LUT3 #(
		.INIT('h40)
	) name12381 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18208_
	);
	LUT3 #(
		.INIT('h01)
	) name12382 (
		_w18069_,
		_w18070_,
		_w18071_,
		_w18209_
	);
	LUT4 #(
		.INIT('heee4)
	) name12383 (
		_w18074_,
		_w18207_,
		_w18209_,
		_w18208_,
		_w18210_
	);
	LUT4 #(
		.INIT('h0800)
	) name12384 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18211_
	);
	LUT4 #(
		.INIT('hd7ff)
	) name12385 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18212_
	);
	LUT4 #(
		.INIT('h0100)
	) name12386 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18213_
	);
	LUT4 #(
		.INIT('h0010)
	) name12387 (
		_w18079_,
		_w18080_,
		_w18076_,
		_w18213_,
		_w18214_
	);
	LUT3 #(
		.INIT('h40)
	) name12388 (
		_w18210_,
		_w18212_,
		_w18214_,
		_w18215_
	);
	LUT4 #(
		.INIT('h0040)
	) name12389 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18216_
	);
	LUT4 #(
		.INIT('hfabd)
	) name12390 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18217_
	);
	LUT4 #(
		.INIT('h0515)
	) name12391 (
		_w18074_,
		_w18076_,
		_w18212_,
		_w18217_,
		_w18218_
	);
	LUT4 #(
		.INIT('haa56)
	) name12392 (
		\u1_L9_reg[13]/NET0131 ,
		_w18206_,
		_w18215_,
		_w18218_,
		_w18219_
	);
	LUT4 #(
		.INIT('hc963)
	) name12393 (
		decrypt_pad,
		\u1_R9_reg[20]/NET0131 ,
		\u1_uk_K_r9_reg[0]/P0001 ,
		\u1_uk_K_r9_reg[8]/NET0131 ,
		_w18220_
	);
	LUT4 #(
		.INIT('hc963)
	) name12394 (
		decrypt_pad,
		\u1_R9_reg[19]/NET0131 ,
		\u1_uk_K_r9_reg[16]/NET0131 ,
		\u1_uk_K_r9_reg[52]/NET0131 ,
		_w18221_
	);
	LUT4 #(
		.INIT('hc693)
	) name12395 (
		decrypt_pad,
		\u1_R9_reg[16]/NET0131 ,
		\u1_uk_K_r9_reg[21]/NET0131 ,
		\u1_uk_K_r9_reg[44]/NET0131 ,
		_w18222_
	);
	LUT4 #(
		.INIT('hc963)
	) name12396 (
		decrypt_pad,
		\u1_R9_reg[21]/NET0131 ,
		\u1_uk_K_r9_reg[1]/NET0131 ,
		\u1_uk_K_r9_reg[9]/NET0131 ,
		_w18223_
	);
	LUT4 #(
		.INIT('hc963)
	) name12397 (
		decrypt_pad,
		\u1_R9_reg[17]/NET0131 ,
		\u1_uk_K_r9_reg[35]/NET0131 ,
		\u1_uk_K_r9_reg[43]/NET0131 ,
		_w18224_
	);
	LUT4 #(
		.INIT('hc963)
	) name12398 (
		decrypt_pad,
		\u1_R9_reg[18]/NET0131 ,
		\u1_uk_K_r9_reg[29]/NET0131 ,
		\u1_uk_K_r9_reg[37]/NET0131 ,
		_w18225_
	);
	LUT4 #(
		.INIT('h87b3)
	) name12399 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18226_
	);
	LUT2 #(
		.INIT('h2)
	) name12400 (
		_w18221_,
		_w18226_,
		_w18227_
	);
	LUT2 #(
		.INIT('h1)
	) name12401 (
		_w18225_,
		_w18221_,
		_w18228_
	);
	LUT3 #(
		.INIT('hde)
	) name12402 (
		_w18223_,
		_w18222_,
		_w18224_,
		_w18229_
	);
	LUT2 #(
		.INIT('h2)
	) name12403 (
		_w18228_,
		_w18229_,
		_w18230_
	);
	LUT3 #(
		.INIT('h80)
	) name12404 (
		_w18223_,
		_w18222_,
		_w18224_,
		_w18231_
	);
	LUT2 #(
		.INIT('h2)
	) name12405 (
		_w18225_,
		_w18221_,
		_w18232_
	);
	LUT4 #(
		.INIT('h0020)
	) name12406 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18233_
	);
	LUT4 #(
		.INIT('hef9f)
	) name12407 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18234_
	);
	LUT3 #(
		.INIT('h70)
	) name12408 (
		_w18231_,
		_w18232_,
		_w18234_,
		_w18235_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name12409 (
		_w18220_,
		_w18230_,
		_w18227_,
		_w18235_,
		_w18236_
	);
	LUT3 #(
		.INIT('h74)
	) name12410 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18237_
	);
	LUT4 #(
		.INIT('h0180)
	) name12411 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18238_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12412 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18221_,
		_w18239_
	);
	LUT4 #(
		.INIT('hfafc)
	) name12413 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18240_
	);
	LUT2 #(
		.INIT('h8)
	) name12414 (
		_w18239_,
		_w18240_,
		_w18241_
	);
	LUT4 #(
		.INIT('h4000)
	) name12415 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18242_
	);
	LUT4 #(
		.INIT('h0010)
	) name12416 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18243_
	);
	LUT4 #(
		.INIT('hddf3)
	) name12417 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18244_
	);
	LUT4 #(
		.INIT('h0100)
	) name12418 (
		_w18221_,
		_w18243_,
		_w18242_,
		_w18244_,
		_w18245_
	);
	LUT4 #(
		.INIT('h00ab)
	) name12419 (
		_w18238_,
		_w18241_,
		_w18245_,
		_w18220_,
		_w18246_
	);
	LUT4 #(
		.INIT('h0008)
	) name12420 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18247_
	);
	LUT4 #(
		.INIT('h0208)
	) name12421 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18248_
	);
	LUT4 #(
		.INIT('heffd)
	) name12422 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18249_
	);
	LUT3 #(
		.INIT('hb1)
	) name12423 (
		_w18221_,
		_w18248_,
		_w18249_,
		_w18250_
	);
	LUT4 #(
		.INIT('h5655)
	) name12424 (
		\u1_L9_reg[14]/NET0131 ,
		_w18246_,
		_w18236_,
		_w18250_,
		_w18251_
	);
	LUT4 #(
		.INIT('h7773)
	) name12425 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18252_
	);
	LUT4 #(
		.INIT('h6763)
	) name12426 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18253_
	);
	LUT4 #(
		.INIT('h0002)
	) name12427 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18254_
	);
	LUT4 #(
		.INIT('h3302)
	) name12428 (
		_w18134_,
		_w18133_,
		_w18253_,
		_w18254_,
		_w18255_
	);
	LUT4 #(
		.INIT('hd9be)
	) name12429 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18256_
	);
	LUT2 #(
		.INIT('h1)
	) name12430 (
		_w18134_,
		_w18256_,
		_w18257_
	);
	LUT3 #(
		.INIT('h08)
	) name12431 (
		_w18138_,
		_w18135_,
		_w18137_,
		_w18258_
	);
	LUT4 #(
		.INIT('h0040)
	) name12432 (
		_w18135_,
		_w18136_,
		_w18137_,
		_w18134_,
		_w18259_
	);
	LUT3 #(
		.INIT('h01)
	) name12433 (
		_w18154_,
		_w18258_,
		_w18259_,
		_w18260_
	);
	LUT4 #(
		.INIT('h2000)
	) name12434 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18261_
	);
	LUT4 #(
		.INIT('h0100)
	) name12435 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18134_,
		_w18262_
	);
	LUT2 #(
		.INIT('h1)
	) name12436 (
		_w18261_,
		_w18262_,
		_w18263_
	);
	LUT4 #(
		.INIT('hbfef)
	) name12437 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18264_
	);
	LUT4 #(
		.INIT('h0002)
	) name12438 (
		_w18138_,
		_w18135_,
		_w18134_,
		_w18133_,
		_w18265_
	);
	LUT3 #(
		.INIT('h0d)
	) name12439 (
		_w18134_,
		_w18264_,
		_w18265_,
		_w18266_
	);
	LUT4 #(
		.INIT('hd500)
	) name12440 (
		_w18133_,
		_w18260_,
		_w18263_,
		_w18266_,
		_w18267_
	);
	LUT4 #(
		.INIT('h5655)
	) name12441 (
		\u1_L9_reg[15]/P0001 ,
		_w18255_,
		_w18257_,
		_w18267_,
		_w18268_
	);
	LUT4 #(
		.INIT('h2100)
	) name12442 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18269_
	);
	LUT2 #(
		.INIT('h1)
	) name12443 (
		_w18031_,
		_w18269_,
		_w18270_
	);
	LUT4 #(
		.INIT('hf3f1)
	) name12444 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18271_
	);
	LUT2 #(
		.INIT('h2)
	) name12445 (
		_w18035_,
		_w18271_,
		_w18272_
	);
	LUT3 #(
		.INIT('h02)
	) name12446 (
		_w18031_,
		_w18047_,
		_w18165_,
		_w18273_
	);
	LUT3 #(
		.INIT('h45)
	) name12447 (
		_w18270_,
		_w18272_,
		_w18273_,
		_w18274_
	);
	LUT4 #(
		.INIT('h2500)
	) name12448 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18275_
	);
	LUT4 #(
		.INIT('h080c)
	) name12449 (
		_w18037_,
		_w18030_,
		_w18031_,
		_w18033_,
		_w18276_
	);
	LUT4 #(
		.INIT('h080a)
	) name12450 (
		_w18035_,
		_w18173_,
		_w18275_,
		_w18276_,
		_w18277_
	);
	LUT3 #(
		.INIT('h08)
	) name12451 (
		_w18037_,
		_w18030_,
		_w18033_,
		_w18278_
	);
	LUT3 #(
		.INIT('h8a)
	) name12452 (
		_w18032_,
		_w18030_,
		_w18031_,
		_w18279_
	);
	LUT3 #(
		.INIT('h10)
	) name12453 (
		_w18046_,
		_w18278_,
		_w18279_,
		_w18280_
	);
	LUT4 #(
		.INIT('hfdee)
	) name12454 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18281_
	);
	LUT4 #(
		.INIT('h0301)
	) name12455 (
		_w18031_,
		_w18035_,
		_w18058_,
		_w18281_,
		_w18282_
	);
	LUT3 #(
		.INIT('h45)
	) name12456 (
		_w18277_,
		_w18280_,
		_w18282_,
		_w18283_
	);
	LUT3 #(
		.INIT('h56)
	) name12457 (
		\u1_L9_reg[1]/NET0131 ,
		_w18274_,
		_w18283_,
		_w18284_
	);
	LUT4 #(
		.INIT('hfb9f)
	) name12458 (
		_w17974_,
		_w17976_,
		_w17980_,
		_w17977_,
		_w18285_
	);
	LUT2 #(
		.INIT('h1)
	) name12459 (
		_w17975_,
		_w18285_,
		_w18286_
	);
	LUT4 #(
		.INIT('h1001)
	) name12460 (
		_w17974_,
		_w17976_,
		_w17980_,
		_w17977_,
		_w18287_
	);
	LUT4 #(
		.INIT('h45e5)
	) name12461 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18288_
	);
	LUT4 #(
		.INIT('h8000)
	) name12462 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18289_
	);
	LUT4 #(
		.INIT('h0051)
	) name12463 (
		_w17973_,
		_w17974_,
		_w18288_,
		_w18289_,
		_w18290_
	);
	LUT3 #(
		.INIT('h04)
	) name12464 (
		_w17974_,
		_w17976_,
		_w17977_,
		_w18291_
	);
	LUT4 #(
		.INIT('haa8a)
	) name12465 (
		_w17973_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18292_
	);
	LUT3 #(
		.INIT('h10)
	) name12466 (
		_w17994_,
		_w18291_,
		_w18292_,
		_w18293_
	);
	LUT4 #(
		.INIT('h4100)
	) name12467 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18294_
	);
	LUT4 #(
		.INIT('hfb5b)
	) name12468 (
		_w17976_,
		_w17980_,
		_w17977_,
		_w17975_,
		_w18295_
	);
	LUT3 #(
		.INIT('h31)
	) name12469 (
		_w17974_,
		_w18294_,
		_w18295_,
		_w18296_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name12470 (
		_w18287_,
		_w18290_,
		_w18293_,
		_w18296_,
		_w18297_
	);
	LUT3 #(
		.INIT('h56)
	) name12471 (
		\u1_L9_reg[19]/NET0131 ,
		_w18286_,
		_w18297_,
		_w18298_
	);
	LUT4 #(
		.INIT('h378f)
	) name12472 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18299_
	);
	LUT2 #(
		.INIT('h2)
	) name12473 (
		_w18134_,
		_w18299_,
		_w18300_
	);
	LUT4 #(
		.INIT('hd5f5)
	) name12474 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18301_
	);
	LUT3 #(
		.INIT('h0b)
	) name12475 (
		_w18136_,
		_w18137_,
		_w18134_,
		_w18302_
	);
	LUT4 #(
		.INIT('hf6ef)
	) name12476 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18303_
	);
	LUT3 #(
		.INIT('hb0)
	) name12477 (
		_w18301_,
		_w18302_,
		_w18303_,
		_w18304_
	);
	LUT3 #(
		.INIT('h8a)
	) name12478 (
		_w18133_,
		_w18300_,
		_w18304_,
		_w18305_
	);
	LUT4 #(
		.INIT('hb9ff)
	) name12479 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18306_
	);
	LUT4 #(
		.INIT('h0040)
	) name12480 (
		_w18138_,
		_w18136_,
		_w18137_,
		_w18134_,
		_w18307_
	);
	LUT4 #(
		.INIT('h0004)
	) name12481 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18134_,
		_w18308_
	);
	LUT3 #(
		.INIT('h10)
	) name12482 (
		_w18307_,
		_w18308_,
		_w18306_,
		_w18309_
	);
	LUT2 #(
		.INIT('h4)
	) name12483 (
		_w18135_,
		_w18134_,
		_w18310_
	);
	LUT3 #(
		.INIT('h31)
	) name12484 (
		_w18139_,
		_w18157_,
		_w18310_,
		_w18311_
	);
	LUT3 #(
		.INIT('h15)
	) name12485 (
		_w18133_,
		_w18309_,
		_w18311_,
		_w18312_
	);
	LUT4 #(
		.INIT('hd5f7)
	) name12486 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18313_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name12487 (
		_w18134_,
		_w18133_,
		_w18141_,
		_w18313_,
		_w18314_
	);
	LUT3 #(
		.INIT('h80)
	) name12488 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18315_
	);
	LUT2 #(
		.INIT('h8)
	) name12489 (
		_w18145_,
		_w18315_,
		_w18316_
	);
	LUT2 #(
		.INIT('h1)
	) name12490 (
		_w18314_,
		_w18316_,
		_w18317_
	);
	LUT4 #(
		.INIT('h5655)
	) name12491 (
		\u1_L9_reg[21]/NET0131 ,
		_w18305_,
		_w18312_,
		_w18317_,
		_w18318_
	);
	LUT4 #(
		.INIT('h337f)
	) name12492 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w18319_
	);
	LUT2 #(
		.INIT('h1)
	) name12493 (
		_w17938_,
		_w18319_,
		_w18320_
	);
	LUT3 #(
		.INIT('h23)
	) name12494 (
		_w17938_,
		_w17939_,
		_w17940_,
		_w18321_
	);
	LUT3 #(
		.INIT('h35)
	) name12495 (
		_w17942_,
		_w17943_,
		_w17940_,
		_w18322_
	);
	LUT2 #(
		.INIT('h8)
	) name12496 (
		_w18321_,
		_w18322_,
		_w18323_
	);
	LUT3 #(
		.INIT('h80)
	) name12497 (
		_w17942_,
		_w17939_,
		_w17940_,
		_w18324_
	);
	LUT4 #(
		.INIT('h0800)
	) name12498 (
		_w17938_,
		_w17942_,
		_w17943_,
		_w17939_,
		_w18325_
	);
	LUT3 #(
		.INIT('h01)
	) name12499 (
		_w17937_,
		_w18325_,
		_w18324_,
		_w18326_
	);
	LUT3 #(
		.INIT('h10)
	) name12500 (
		_w18320_,
		_w18323_,
		_w18326_,
		_w18327_
	);
	LUT2 #(
		.INIT('h8)
	) name12501 (
		_w17938_,
		_w17940_,
		_w18328_
	);
	LUT4 #(
		.INIT('ha800)
	) name12502 (
		_w17938_,
		_w17942_,
		_w17939_,
		_w17940_,
		_w18329_
	);
	LUT2 #(
		.INIT('h8)
	) name12503 (
		_w17955_,
		_w18329_,
		_w18330_
	);
	LUT4 #(
		.INIT('h0040)
	) name12504 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w18331_
	);
	LUT4 #(
		.INIT('h004c)
	) name12505 (
		_w17961_,
		_w17937_,
		_w17968_,
		_w18331_,
		_w18332_
	);
	LUT2 #(
		.INIT('h4)
	) name12506 (
		_w18330_,
		_w18332_,
		_w18333_
	);
	LUT3 #(
		.INIT('h69)
	) name12507 (
		_w17943_,
		_w17939_,
		_w17940_,
		_w18334_
	);
	LUT4 #(
		.INIT('h3b00)
	) name12508 (
		_w17942_,
		_w17943_,
		_w17940_,
		_w17937_,
		_w18335_
	);
	LUT4 #(
		.INIT('h7bef)
	) name12509 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w18336_
	);
	LUT4 #(
		.INIT('h1055)
	) name12510 (
		_w17938_,
		_w18334_,
		_w18335_,
		_w18336_,
		_w18337_
	);
	LUT3 #(
		.INIT('h13)
	) name12511 (
		_w17956_,
		_w17969_,
		_w18328_,
		_w18338_
	);
	LUT2 #(
		.INIT('h4)
	) name12512 (
		_w18337_,
		_w18338_,
		_w18339_
	);
	LUT4 #(
		.INIT('h56aa)
	) name12513 (
		\u1_L9_reg[23]/NET0131 ,
		_w18327_,
		_w18333_,
		_w18339_,
		_w18340_
	);
	LUT4 #(
		.INIT('h3de0)
	) name12514 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18341_
	);
	LUT4 #(
		.INIT('hfa3f)
	) name12515 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18342_
	);
	LUT4 #(
		.INIT('h6400)
	) name12516 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18343_
	);
	LUT4 #(
		.INIT('h00d8)
	) name12517 (
		_w18221_,
		_w18341_,
		_w18342_,
		_w18343_,
		_w18344_
	);
	LUT2 #(
		.INIT('h2)
	) name12518 (
		_w18220_,
		_w18344_,
		_w18345_
	);
	LUT4 #(
		.INIT('hdff9)
	) name12519 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18346_
	);
	LUT2 #(
		.INIT('h2)
	) name12520 (
		_w18221_,
		_w18346_,
		_w18347_
	);
	LUT2 #(
		.INIT('h4)
	) name12521 (
		_w18223_,
		_w18221_,
		_w18348_
	);
	LUT4 #(
		.INIT('hf5cf)
	) name12522 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18349_
	);
	LUT3 #(
		.INIT('hb0)
	) name12523 (
		_w18223_,
		_w18224_,
		_w18221_,
		_w18350_
	);
	LUT4 #(
		.INIT('h5501)
	) name12524 (
		_w18225_,
		_w18222_,
		_w18224_,
		_w18221_,
		_w18351_
	);
	LUT4 #(
		.INIT('he0ee)
	) name12525 (
		_w18348_,
		_w18349_,
		_w18350_,
		_w18351_,
		_w18352_
	);
	LUT4 #(
		.INIT('h0008)
	) name12526 (
		_w18225_,
		_w18222_,
		_w18224_,
		_w18221_,
		_w18353_
	);
	LUT2 #(
		.INIT('h1)
	) name12527 (
		_w18242_,
		_w18353_,
		_w18354_
	);
	LUT4 #(
		.INIT('h0e00)
	) name12528 (
		_w18220_,
		_w18352_,
		_w18347_,
		_w18354_,
		_w18355_
	);
	LUT3 #(
		.INIT('h65)
	) name12529 (
		\u1_L9_reg[25]/NET0131 ,
		_w18345_,
		_w18355_,
		_w18356_
	);
	LUT4 #(
		.INIT('h0092)
	) name12530 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18357_
	);
	LUT3 #(
		.INIT('h8c)
	) name12531 (
		_w18032_,
		_w18037_,
		_w18033_,
		_w18358_
	);
	LUT2 #(
		.INIT('h1)
	) name12532 (
		_w18030_,
		_w18035_,
		_w18359_
	);
	LUT4 #(
		.INIT('h5150)
	) name12533 (
		_w18031_,
		_w18358_,
		_w18357_,
		_w18359_,
		_w18360_
	);
	LUT4 #(
		.INIT('h2010)
	) name12534 (
		_w18032_,
		_w18037_,
		_w18030_,
		_w18033_,
		_w18361_
	);
	LUT4 #(
		.INIT('h0f01)
	) name12535 (
		_w18032_,
		_w18030_,
		_w18031_,
		_w18033_,
		_w18362_
	);
	LUT2 #(
		.INIT('h8)
	) name12536 (
		_w18358_,
		_w18362_,
		_w18363_
	);
	LUT3 #(
		.INIT('h40)
	) name12537 (
		_w18032_,
		_w18037_,
		_w18033_,
		_w18364_
	);
	LUT4 #(
		.INIT('h2022)
	) name12538 (
		_w18035_,
		_w18041_,
		_w18051_,
		_w18364_,
		_w18365_
	);
	LUT3 #(
		.INIT('h10)
	) name12539 (
		_w18363_,
		_w18361_,
		_w18365_,
		_w18366_
	);
	LUT3 #(
		.INIT('h80)
	) name12540 (
		_w18030_,
		_w18031_,
		_w18033_,
		_w18367_
	);
	LUT2 #(
		.INIT('h4)
	) name12541 (
		_w18059_,
		_w18367_,
		_w18368_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12542 (
		_w18032_,
		_w18030_,
		_w18033_,
		_w18035_,
		_w18369_
	);
	LUT3 #(
		.INIT('h10)
	) name12543 (
		_w18057_,
		_w18058_,
		_w18369_,
		_w18370_
	);
	LUT2 #(
		.INIT('h4)
	) name12544 (
		_w18368_,
		_w18370_,
		_w18371_
	);
	LUT2 #(
		.INIT('h4)
	) name12545 (
		_w18055_,
		_w18171_,
		_w18372_
	);
	LUT4 #(
		.INIT('h000e)
	) name12546 (
		_w18366_,
		_w18371_,
		_w18372_,
		_w18360_,
		_w18373_
	);
	LUT2 #(
		.INIT('h9)
	) name12547 (
		\u1_L9_reg[26]/NET0131 ,
		_w18373_,
		_w18374_
	);
	LUT4 #(
		.INIT('haefe)
	) name12548 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18375_
	);
	LUT3 #(
		.INIT('h04)
	) name12549 (
		_w18072_,
		_w18069_,
		_w18071_,
		_w18376_
	);
	LUT4 #(
		.INIT('h5545)
	) name12550 (
		_w18074_,
		_w18072_,
		_w18069_,
		_w18071_,
		_w18377_
	);
	LUT4 #(
		.INIT('h55ad)
	) name12551 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18378_
	);
	LUT4 #(
		.INIT('h7277)
	) name12552 (
		_w18074_,
		_w18375_,
		_w18376_,
		_w18378_,
		_w18379_
	);
	LUT4 #(
		.INIT('h0084)
	) name12553 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18380_
	);
	LUT3 #(
		.INIT('h01)
	) name12554 (
		_w18076_,
		_w18211_,
		_w18380_,
		_w18381_
	);
	LUT4 #(
		.INIT('ha400)
	) name12555 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18382_
	);
	LUT4 #(
		.INIT('ha6fe)
	) name12556 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18383_
	);
	LUT4 #(
		.INIT('h31f5)
	) name12557 (
		_w18199_,
		_w18377_,
		_w18382_,
		_w18383_,
		_w18384_
	);
	LUT4 #(
		.INIT('h00d0)
	) name12558 (
		_w18094_,
		_w18082_,
		_w18076_,
		_w18216_,
		_w18385_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12559 (
		_w18379_,
		_w18381_,
		_w18384_,
		_w18385_,
		_w18386_
	);
	LUT2 #(
		.INIT('h6)
	) name12560 (
		\u1_L9_reg[28]/NET0131 ,
		_w18386_,
		_w18387_
	);
	LUT4 #(
		.INIT('hff3e)
	) name12561 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18388_
	);
	LUT3 #(
		.INIT('h04)
	) name12562 (
		_w18225_,
		_w18222_,
		_w18221_,
		_w18389_
	);
	LUT4 #(
		.INIT('h0031)
	) name12563 (
		_w18221_,
		_w18248_,
		_w18388_,
		_w18389_,
		_w18390_
	);
	LUT2 #(
		.INIT('h2)
	) name12564 (
		_w18220_,
		_w18390_,
		_w18391_
	);
	LUT3 #(
		.INIT('h02)
	) name12565 (
		_w18221_,
		_w18243_,
		_w18231_,
		_w18392_
	);
	LUT4 #(
		.INIT('h0c04)
	) name12566 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18393_
	);
	LUT4 #(
		.INIT('h00f7)
	) name12567 (
		_w18223_,
		_w18222_,
		_w18224_,
		_w18221_,
		_w18394_
	);
	LUT2 #(
		.INIT('h4)
	) name12568 (
		_w18393_,
		_w18394_,
		_w18395_
	);
	LUT4 #(
		.INIT('hdafd)
	) name12569 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18396_
	);
	LUT4 #(
		.INIT('h0155)
	) name12570 (
		_w18220_,
		_w18392_,
		_w18395_,
		_w18396_,
		_w18397_
	);
	LUT4 #(
		.INIT('hd9f7)
	) name12571 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18398_
	);
	LUT4 #(
		.INIT('haf23)
	) name12572 (
		_w18223_,
		_w18221_,
		_w18353_,
		_w18398_,
		_w18399_
	);
	LUT4 #(
		.INIT('h5655)
	) name12573 (
		\u1_L9_reg[8]/NET0131 ,
		_w18397_,
		_w18391_,
		_w18399_,
		_w18400_
	);
	LUT4 #(
		.INIT('hb7a6)
	) name12574 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18401_
	);
	LUT2 #(
		.INIT('h1)
	) name12575 (
		_w18134_,
		_w18401_,
		_w18402_
	);
	LUT3 #(
		.INIT('hd0)
	) name12576 (
		_w18138_,
		_w18136_,
		_w18134_,
		_w18403_
	);
	LUT4 #(
		.INIT('hbdcf)
	) name12577 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18404_
	);
	LUT3 #(
		.INIT('hb0)
	) name12578 (
		_w18252_,
		_w18403_,
		_w18404_,
		_w18405_
	);
	LUT3 #(
		.INIT('h8a)
	) name12579 (
		_w18133_,
		_w18402_,
		_w18405_,
		_w18406_
	);
	LUT4 #(
		.INIT('hfd00)
	) name12580 (
		_w18135_,
		_w18136_,
		_w18137_,
		_w18134_,
		_w18407_
	);
	LUT4 #(
		.INIT('h0bcf)
	) name12581 (
		_w18138_,
		_w18135_,
		_w18136_,
		_w18137_,
		_w18408_
	);
	LUT2 #(
		.INIT('h8)
	) name12582 (
		_w18407_,
		_w18408_,
		_w18409_
	);
	LUT4 #(
		.INIT('h0080)
	) name12583 (
		_w18138_,
		_w18136_,
		_w18137_,
		_w18134_,
		_w18410_
	);
	LUT3 #(
		.INIT('h01)
	) name12584 (
		_w18156_,
		_w18308_,
		_w18410_,
		_w18411_
	);
	LUT3 #(
		.INIT('h45)
	) name12585 (
		_w18133_,
		_w18409_,
		_w18411_,
		_w18412_
	);
	LUT2 #(
		.INIT('h1)
	) name12586 (
		_w18134_,
		_w18155_,
		_w18413_
	);
	LUT4 #(
		.INIT('h1000)
	) name12587 (
		_w18135_,
		_w18136_,
		_w18137_,
		_w18134_,
		_w18414_
	);
	LUT3 #(
		.INIT('h07)
	) name12588 (
		_w18145_,
		_w18161_,
		_w18414_,
		_w18415_
	);
	LUT2 #(
		.INIT('h4)
	) name12589 (
		_w18413_,
		_w18415_,
		_w18416_
	);
	LUT4 #(
		.INIT('h5655)
	) name12590 (
		\u1_L9_reg[27]/NET0131 ,
		_w18406_,
		_w18412_,
		_w18416_,
		_w18417_
	);
	LUT3 #(
		.INIT('h02)
	) name12591 (
		_w18221_,
		_w18243_,
		_w18247_,
		_w18418_
	);
	LUT4 #(
		.INIT('h1001)
	) name12592 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18419_
	);
	LUT3 #(
		.INIT('h0e)
	) name12593 (
		_w18228_,
		_w18394_,
		_w18419_,
		_w18420_
	);
	LUT2 #(
		.INIT('h1)
	) name12594 (
		_w18418_,
		_w18420_,
		_w18421_
	);
	LUT3 #(
		.INIT('h04)
	) name12595 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18422_
	);
	LUT4 #(
		.INIT('hbf00)
	) name12596 (
		_w18223_,
		_w18222_,
		_w18224_,
		_w18221_,
		_w18423_
	);
	LUT4 #(
		.INIT('h7077)
	) name12597 (
		_w18237_,
		_w18394_,
		_w18422_,
		_w18423_,
		_w18424_
	);
	LUT4 #(
		.INIT('h008a)
	) name12598 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18425_
	);
	LUT2 #(
		.INIT('h1)
	) name12599 (
		_w18220_,
		_w18425_,
		_w18426_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name12600 (
		_w18225_,
		_w18223_,
		_w18222_,
		_w18224_,
		_w18427_
	);
	LUT2 #(
		.INIT('h2)
	) name12601 (
		_w18221_,
		_w18427_,
		_w18428_
	);
	LUT4 #(
		.INIT('h0020)
	) name12602 (
		_w18223_,
		_w18222_,
		_w18224_,
		_w18221_,
		_w18429_
	);
	LUT4 #(
		.INIT('h0004)
	) name12603 (
		_w18242_,
		_w18220_,
		_w18233_,
		_w18429_,
		_w18430_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12604 (
		_w18424_,
		_w18426_,
		_w18428_,
		_w18430_,
		_w18431_
	);
	LUT3 #(
		.INIT('h56)
	) name12605 (
		\u1_L9_reg[3]/NET0131 ,
		_w18421_,
		_w18431_,
		_w18432_
	);
	LUT4 #(
		.INIT('hc963)
	) name12606 (
		decrypt_pad,
		\u1_R9_reg[11]/NET0131 ,
		\u1_uk_K_r9_reg[40]/NET0131 ,
		\u1_uk_K_r9_reg[46]/NET0131 ,
		_w18433_
	);
	LUT4 #(
		.INIT('hc693)
	) name12607 (
		decrypt_pad,
		\u1_R9_reg[12]/NET0131 ,
		\u1_uk_K_r9_reg[4]/NET0131 ,
		\u1_uk_K_r9_reg[55]/NET0131 ,
		_w18434_
	);
	LUT4 #(
		.INIT('hc693)
	) name12608 (
		decrypt_pad,
		\u1_R9_reg[10]/NET0131 ,
		\u1_uk_K_r9_reg[20]/NET0131 ,
		\u1_uk_K_r9_reg[39]/NET0131 ,
		_w18435_
	);
	LUT4 #(
		.INIT('hc963)
	) name12609 (
		decrypt_pad,
		\u1_R9_reg[8]/NET0131 ,
		\u1_uk_K_r9_reg[34]/NET0131 ,
		\u1_uk_K_r9_reg[40]/NET0131 ,
		_w18436_
	);
	LUT4 #(
		.INIT('hc963)
	) name12610 (
		decrypt_pad,
		\u1_R9_reg[13]/NET0131 ,
		\u1_uk_K_r9_reg[11]/NET0131 ,
		\u1_uk_K_r9_reg[17]/NET0131 ,
		_w18437_
	);
	LUT4 #(
		.INIT('hc693)
	) name12611 (
		decrypt_pad,
		\u1_R9_reg[9]/NET0131 ,
		\u1_uk_K_r9_reg[12]/NET0131 ,
		\u1_uk_K_r9_reg[6]/NET0131 ,
		_w18438_
	);
	LUT4 #(
		.INIT('h93d3)
	) name12612 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18439_
	);
	LUT4 #(
		.INIT('h0001)
	) name12613 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18440_
	);
	LUT4 #(
		.INIT('hf3fe)
	) name12614 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18441_
	);
	LUT4 #(
		.INIT('h08cc)
	) name12615 (
		_w18434_,
		_w18433_,
		_w18439_,
		_w18441_,
		_w18442_
	);
	LUT2 #(
		.INIT('h8)
	) name12616 (
		_w18437_,
		_w18433_,
		_w18443_
	);
	LUT3 #(
		.INIT('h80)
	) name12617 (
		_w18437_,
		_w18438_,
		_w18433_,
		_w18444_
	);
	LUT2 #(
		.INIT('h9)
	) name12618 (
		_w18436_,
		_w18437_,
		_w18445_
	);
	LUT2 #(
		.INIT('h1)
	) name12619 (
		_w18438_,
		_w18435_,
		_w18446_
	);
	LUT2 #(
		.INIT('h6)
	) name12620 (
		_w18438_,
		_w18435_,
		_w18447_
	);
	LUT4 #(
		.INIT('h0660)
	) name12621 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18448_
	);
	LUT2 #(
		.INIT('h4)
	) name12622 (
		_w18444_,
		_w18448_,
		_w18449_
	);
	LUT3 #(
		.INIT('h26)
	) name12623 (
		_w18436_,
		_w18437_,
		_w18433_,
		_w18450_
	);
	LUT3 #(
		.INIT('h54)
	) name12624 (
		_w18434_,
		_w18450_,
		_w18447_,
		_w18451_
	);
	LUT2 #(
		.INIT('h1)
	) name12625 (
		_w18436_,
		_w18437_,
		_w18452_
	);
	LUT3 #(
		.INIT('h80)
	) name12626 (
		_w18438_,
		_w18435_,
		_w18434_,
		_w18453_
	);
	LUT4 #(
		.INIT('h5d0d)
	) name12627 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18454_
	);
	LUT4 #(
		.INIT('h00b0)
	) name12628 (
		_w18437_,
		_w18438_,
		_w18434_,
		_w18433_,
		_w18455_
	);
	LUT4 #(
		.INIT('h7077)
	) name12629 (
		_w18452_,
		_w18453_,
		_w18454_,
		_w18455_,
		_w18456_
	);
	LUT4 #(
		.INIT('h4500)
	) name12630 (
		_w18442_,
		_w18449_,
		_w18451_,
		_w18456_,
		_w18457_
	);
	LUT2 #(
		.INIT('h9)
	) name12631 (
		\u1_L9_reg[6]/NET0131 ,
		_w18457_,
		_w18458_
	);
	LUT4 #(
		.INIT('h8228)
	) name12632 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w18459_
	);
	LUT3 #(
		.INIT('h43)
	) name12633 (
		_w17943_,
		_w17939_,
		_w17940_,
		_w18460_
	);
	LUT4 #(
		.INIT('h0400)
	) name12634 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w18461_
	);
	LUT4 #(
		.INIT('h002a)
	) name12635 (
		_w17937_,
		_w17951_,
		_w18460_,
		_w18461_,
		_w18462_
	);
	LUT4 #(
		.INIT('h1005)
	) name12636 (
		_w17938_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w18463_
	);
	LUT2 #(
		.INIT('h1)
	) name12637 (
		_w17937_,
		_w18463_,
		_w18464_
	);
	LUT4 #(
		.INIT('h41c3)
	) name12638 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w18465_
	);
	LUT4 #(
		.INIT('h4082)
	) name12639 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w18466_
	);
	LUT3 #(
		.INIT('h04)
	) name12640 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w18467_
	);
	LUT3 #(
		.INIT('h28)
	) name12641 (
		_w17938_,
		_w17939_,
		_w17940_,
		_w18468_
	);
	LUT3 #(
		.INIT('h45)
	) name12642 (
		_w18466_,
		_w18467_,
		_w18468_,
		_w18469_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name12643 (
		_w18459_,
		_w18462_,
		_w18464_,
		_w18469_,
		_w18470_
	);
	LUT3 #(
		.INIT('h40)
	) name12644 (
		_w17938_,
		_w17939_,
		_w17940_,
		_w18471_
	);
	LUT2 #(
		.INIT('h4)
	) name12645 (
		_w17946_,
		_w18471_,
		_w18472_
	);
	LUT3 #(
		.INIT('h56)
	) name12646 (
		\u1_L9_reg[9]/NET0131 ,
		_w18470_,
		_w18472_,
		_w18473_
	);
	LUT2 #(
		.INIT('h9)
	) name12647 (
		_w18002_,
		_w18004_,
		_w18474_
	);
	LUT4 #(
		.INIT('hd003)
	) name12648 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18475_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name12649 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18476_
	);
	LUT3 #(
		.INIT('h01)
	) name12650 (
		_w18005_,
		_w18476_,
		_w18475_,
		_w18477_
	);
	LUT4 #(
		.INIT('h0800)
	) name12651 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18478_
	);
	LUT4 #(
		.INIT('hb5bc)
	) name12652 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18479_
	);
	LUT3 #(
		.INIT('h31)
	) name12653 (
		_w18005_,
		_w18478_,
		_w18479_,
		_w18480_
	);
	LUT3 #(
		.INIT('h8a)
	) name12654 (
		_w17999_,
		_w18477_,
		_w18480_,
		_w18481_
	);
	LUT3 #(
		.INIT('h40)
	) name12655 (
		_w18001_,
		_w18002_,
		_w18004_,
		_w18482_
	);
	LUT4 #(
		.INIT('hab89)
	) name12656 (
		_w18005_,
		_w18186_,
		_w18188_,
		_w18482_,
		_w18483_
	);
	LUT4 #(
		.INIT('h7bd7)
	) name12657 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18484_
	);
	LUT4 #(
		.INIT('h00c8)
	) name12658 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18005_,
		_w18485_
	);
	LUT4 #(
		.INIT('h135f)
	) name12659 (
		_w18005_,
		_w18020_,
		_w18012_,
		_w18485_,
		_w18486_
	);
	LUT4 #(
		.INIT('hba00)
	) name12660 (
		_w17999_,
		_w18483_,
		_w18484_,
		_w18486_,
		_w18487_
	);
	LUT3 #(
		.INIT('h65)
	) name12661 (
		\u1_L9_reg[32]/NET0131 ,
		_w18481_,
		_w18487_,
		_w18488_
	);
	LUT4 #(
		.INIT('hf126)
	) name12662 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18489_
	);
	LUT4 #(
		.INIT('h2880)
	) name12663 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18490_
	);
	LUT4 #(
		.INIT('h5004)
	) name12664 (
		_w18000_,
		_w18001_,
		_w18002_,
		_w18004_,
		_w18491_
	);
	LUT4 #(
		.INIT('h1302)
	) name12665 (
		_w18005_,
		_w18490_,
		_w18491_,
		_w18489_,
		_w18492_
	);
	LUT2 #(
		.INIT('h2)
	) name12666 (
		_w17999_,
		_w18492_,
		_w18493_
	);
	LUT2 #(
		.INIT('h4)
	) name12667 (
		_w18005_,
		_w18490_,
		_w18494_
	);
	LUT2 #(
		.INIT('h2)
	) name12668 (
		_w17999_,
		_w18005_,
		_w18495_
	);
	LUT3 #(
		.INIT('h4c)
	) name12669 (
		_w18001_,
		_w18002_,
		_w18004_,
		_w18496_
	);
	LUT4 #(
		.INIT('h8a00)
	) name12670 (
		_w18000_,
		_w18002_,
		_w18004_,
		_w18005_,
		_w18497_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name12671 (
		_w18006_,
		_w18474_,
		_w18496_,
		_w18497_,
		_w18498_
	);
	LUT3 #(
		.INIT('h45)
	) name12672 (
		_w18019_,
		_w18005_,
		_w18491_,
		_w18499_
	);
	LUT4 #(
		.INIT('h0133)
	) name12673 (
		_w17999_,
		_w18495_,
		_w18498_,
		_w18499_,
		_w18500_
	);
	LUT4 #(
		.INIT('h5556)
	) name12674 (
		\u1_L9_reg[7]/NET0131 ,
		_w18494_,
		_w18500_,
		_w18493_,
		_w18501_
	);
	LUT3 #(
		.INIT('h10)
	) name12675 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18502_
	);
	LUT2 #(
		.INIT('h8)
	) name12676 (
		_w18436_,
		_w18437_,
		_w18503_
	);
	LUT3 #(
		.INIT('h80)
	) name12677 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18504_
	);
	LUT4 #(
		.INIT('h6979)
	) name12678 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18433_,
		_w18505_
	);
	LUT2 #(
		.INIT('h1)
	) name12679 (
		_w18435_,
		_w18505_,
		_w18506_
	);
	LUT4 #(
		.INIT('h4000)
	) name12680 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18507_
	);
	LUT4 #(
		.INIT('h0100)
	) name12681 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18508_
	);
	LUT3 #(
		.INIT('h12)
	) name12682 (
		_w18436_,
		_w18437_,
		_w18435_,
		_w18509_
	);
	LUT4 #(
		.INIT('h020f)
	) name12683 (
		_w18433_,
		_w18508_,
		_w18507_,
		_w18509_,
		_w18510_
	);
	LUT3 #(
		.INIT('h8a)
	) name12684 (
		_w18434_,
		_w18506_,
		_w18510_,
		_w18511_
	);
	LUT4 #(
		.INIT('h7b6a)
	) name12685 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18512_
	);
	LUT4 #(
		.INIT('h6800)
	) name12686 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18433_,
		_w18513_
	);
	LUT4 #(
		.INIT('h00f2)
	) name12687 (
		_w18433_,
		_w18440_,
		_w18512_,
		_w18513_,
		_w18514_
	);
	LUT3 #(
		.INIT('h20)
	) name12688 (
		_w18436_,
		_w18438_,
		_w18435_,
		_w18515_
	);
	LUT4 #(
		.INIT('h00df)
	) name12689 (
		_w18436_,
		_w18438_,
		_w18435_,
		_w18433_,
		_w18516_
	);
	LUT4 #(
		.INIT('h2000)
	) name12690 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18517_
	);
	LUT4 #(
		.INIT('h3331)
	) name12691 (
		_w18433_,
		_w18516_,
		_w18508_,
		_w18517_,
		_w18518_
	);
	LUT3 #(
		.INIT('h0e)
	) name12692 (
		_w18434_,
		_w18514_,
		_w18518_,
		_w18519_
	);
	LUT3 #(
		.INIT('h65)
	) name12693 (
		\u1_L9_reg[16]/NET0131 ,
		_w18511_,
		_w18519_,
		_w18520_
	);
	LUT4 #(
		.INIT('h0a20)
	) name12694 (
		_w18074_,
		_w18072_,
		_w18070_,
		_w18071_,
		_w18521_
	);
	LUT3 #(
		.INIT('hb8)
	) name12695 (
		_w18069_,
		_w18070_,
		_w18071_,
		_w18522_
	);
	LUT2 #(
		.INIT('h4)
	) name12696 (
		_w18074_,
		_w18072_,
		_w18523_
	);
	LUT4 #(
		.INIT('h1011)
	) name12697 (
		_w18099_,
		_w18521_,
		_w18522_,
		_w18523_,
		_w18524_
	);
	LUT4 #(
		.INIT('h1003)
	) name12698 (
		_w18074_,
		_w18072_,
		_w18069_,
		_w18071_,
		_w18525_
	);
	LUT3 #(
		.INIT('h53)
	) name12699 (
		_w18074_,
		_w18069_,
		_w18071_,
		_w18526_
	);
	LUT4 #(
		.INIT('hf7fc)
	) name12700 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18527_
	);
	LUT4 #(
		.INIT('h0d00)
	) name12701 (
		_w18090_,
		_w18526_,
		_w18525_,
		_w18527_,
		_w18528_
	);
	LUT4 #(
		.INIT('h1000)
	) name12702 (
		_w18074_,
		_w18072_,
		_w18070_,
		_w18071_,
		_w18529_
	);
	LUT4 #(
		.INIT('h7e7f)
	) name12703 (
		_w18072_,
		_w18069_,
		_w18070_,
		_w18071_,
		_w18530_
	);
	LUT3 #(
		.INIT('h31)
	) name12704 (
		_w18074_,
		_w18529_,
		_w18530_,
		_w18531_
	);
	LUT4 #(
		.INIT('he400)
	) name12705 (
		_w18076_,
		_w18528_,
		_w18524_,
		_w18531_,
		_w18532_
	);
	LUT2 #(
		.INIT('h9)
	) name12706 (
		\u1_L9_reg[18]/P0001 ,
		_w18532_,
		_w18533_
	);
	LUT4 #(
		.INIT('h0009)
	) name12707 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18534_
	);
	LUT4 #(
		.INIT('h99d6)
	) name12708 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18535_
	);
	LUT3 #(
		.INIT('h32)
	) name12709 (
		_w18434_,
		_w18433_,
		_w18535_,
		_w18536_
	);
	LUT4 #(
		.INIT('h0042)
	) name12710 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18537_
	);
	LUT4 #(
		.INIT('heb00)
	) name12711 (
		_w18436_,
		_w18437_,
		_w18435_,
		_w18433_,
		_w18538_
	);
	LUT4 #(
		.INIT('he5ef)
	) name12712 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18539_
	);
	LUT4 #(
		.INIT('h3222)
	) name12713 (
		_w18434_,
		_w18537_,
		_w18538_,
		_w18539_,
		_w18540_
	);
	LUT2 #(
		.INIT('h1)
	) name12714 (
		_w18536_,
		_w18540_,
		_w18541_
	);
	LUT2 #(
		.INIT('h2)
	) name12715 (
		_w18435_,
		_w18433_,
		_w18542_
	);
	LUT2 #(
		.INIT('h8)
	) name12716 (
		_w18504_,
		_w18542_,
		_w18543_
	);
	LUT4 #(
		.INIT('h1bf4)
	) name12717 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18544_
	);
	LUT2 #(
		.INIT('h2)
	) name12718 (
		_w18433_,
		_w18544_,
		_w18545_
	);
	LUT3 #(
		.INIT('h0e)
	) name12719 (
		_w18438_,
		_w18435_,
		_w18433_,
		_w18546_
	);
	LUT4 #(
		.INIT('h153f)
	) name12720 (
		_w18445_,
		_w18450_,
		_w18446_,
		_w18546_,
		_w18547_
	);
	LUT4 #(
		.INIT('h1311)
	) name12721 (
		_w18434_,
		_w18543_,
		_w18545_,
		_w18547_,
		_w18548_
	);
	LUT3 #(
		.INIT('h65)
	) name12722 (
		\u1_L9_reg[24]/NET0131 ,
		_w18541_,
		_w18548_,
		_w18549_
	);
	LUT4 #(
		.INIT('h0002)
	) name12723 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18550_
	);
	LUT3 #(
		.INIT('h07)
	) name12724 (
		_w18436_,
		_w18435_,
		_w18433_,
		_w18551_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name12725 (
		_w18502_,
		_w18538_,
		_w18550_,
		_w18551_,
		_w18552_
	);
	LUT4 #(
		.INIT('h008a)
	) name12726 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18553_
	);
	LUT4 #(
		.INIT('h00bf)
	) name12727 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18433_,
		_w18554_
	);
	LUT4 #(
		.INIT('h8a00)
	) name12728 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18555_
	);
	LUT4 #(
		.INIT('hfb00)
	) name12729 (
		_w18437_,
		_w18438_,
		_w18435_,
		_w18433_,
		_w18556_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12730 (
		_w18553_,
		_w18554_,
		_w18555_,
		_w18556_,
		_w18557_
	);
	LUT4 #(
		.INIT('h0400)
	) name12731 (
		_w18436_,
		_w18437_,
		_w18438_,
		_w18435_,
		_w18558_
	);
	LUT3 #(
		.INIT('h01)
	) name12732 (
		_w18434_,
		_w18534_,
		_w18558_,
		_w18559_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name12733 (
		_w18434_,
		_w18552_,
		_w18557_,
		_w18559_,
		_w18560_
	);
	LUT2 #(
		.INIT('h8)
	) name12734 (
		_w18443_,
		_w18515_,
		_w18561_
	);
	LUT4 #(
		.INIT('h0040)
	) name12735 (
		_w18437_,
		_w18438_,
		_w18435_,
		_w18433_,
		_w18562_
	);
	LUT3 #(
		.INIT('h0d)
	) name12736 (
		_w18453_,
		_w18503_,
		_w18562_,
		_w18563_
	);
	LUT2 #(
		.INIT('h4)
	) name12737 (
		_w18561_,
		_w18563_,
		_w18564_
	);
	LUT3 #(
		.INIT('h9a)
	) name12738 (
		\u1_L9_reg[30]/NET0131 ,
		_w18560_,
		_w18564_,
		_w18565_
	);
	LUT4 #(
		.INIT('hc693)
	) name12739 (
		decrypt_pad,
		\u1_R8_reg[28]/NET0131 ,
		\u1_uk_K_r8_reg[44]/NET0131 ,
		\u1_uk_K_r8_reg[9]/NET0131 ,
		_w18566_
	);
	LUT4 #(
		.INIT('hc963)
	) name12740 (
		decrypt_pad,
		\u1_R8_reg[27]/NET0131 ,
		\u1_uk_K_r8_reg[22]/NET0131 ,
		\u1_uk_K_r8_reg[2]/NET0131 ,
		_w18567_
	);
	LUT4 #(
		.INIT('hc693)
	) name12741 (
		decrypt_pad,
		\u1_R8_reg[24]/NET0131 ,
		\u1_uk_K_r8_reg[28]/NET0131 ,
		\u1_uk_K_r8_reg[52]/NET0131 ,
		_w18568_
	);
	LUT2 #(
		.INIT('h8)
	) name12742 (
		_w18567_,
		_w18568_,
		_w18569_
	);
	LUT4 #(
		.INIT('hc963)
	) name12743 (
		decrypt_pad,
		\u1_R8_reg[26]/NET0131 ,
		\u1_uk_K_r8_reg[44]/NET0131 ,
		\u1_uk_K_r8_reg[52]/NET0131 ,
		_w18570_
	);
	LUT4 #(
		.INIT('hc963)
	) name12744 (
		decrypt_pad,
		\u1_R8_reg[25]/NET0131 ,
		\u1_uk_K_r8_reg[28]/NET0131 ,
		\u1_uk_K_r8_reg[8]/NET0131 ,
		_w18571_
	);
	LUT4 #(
		.INIT('hc963)
	) name12745 (
		decrypt_pad,
		\u1_R8_reg[29]/NET0131 ,
		\u1_uk_K_r8_reg[1]/NET0131 ,
		\u1_uk_K_r8_reg[36]/NET0131 ,
		_w18572_
	);
	LUT3 #(
		.INIT('h9d)
	) name12746 (
		_w18570_,
		_w18571_,
		_w18572_,
		_w18573_
	);
	LUT2 #(
		.INIT('h2)
	) name12747 (
		_w18569_,
		_w18573_,
		_w18574_
	);
	LUT4 #(
		.INIT('he3ff)
	) name12748 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18575_
	);
	LUT4 #(
		.INIT('h0200)
	) name12749 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18576_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name12750 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18577_
	);
	LUT3 #(
		.INIT('he0)
	) name12751 (
		_w18567_,
		_w18575_,
		_w18577_,
		_w18578_
	);
	LUT3 #(
		.INIT('h8a)
	) name12752 (
		_w18566_,
		_w18574_,
		_w18578_,
		_w18579_
	);
	LUT4 #(
		.INIT('h0002)
	) name12753 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18580_
	);
	LUT4 #(
		.INIT('h5a2d)
	) name12754 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18581_
	);
	LUT4 #(
		.INIT('h0200)
	) name12755 (
		_w18567_,
		_w18570_,
		_w18571_,
		_w18568_,
		_w18582_
	);
	LUT4 #(
		.INIT('h8400)
	) name12756 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18583_
	);
	LUT4 #(
		.INIT('h000e)
	) name12757 (
		_w18567_,
		_w18581_,
		_w18582_,
		_w18583_,
		_w18584_
	);
	LUT4 #(
		.INIT('h1545)
	) name12758 (
		_w18567_,
		_w18570_,
		_w18571_,
		_w18568_,
		_w18585_
	);
	LUT4 #(
		.INIT('h0008)
	) name12759 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18586_
	);
	LUT4 #(
		.INIT('hffc6)
	) name12760 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18587_
	);
	LUT4 #(
		.INIT('h3133)
	) name12761 (
		_w18567_,
		_w18585_,
		_w18576_,
		_w18587_,
		_w18588_
	);
	LUT3 #(
		.INIT('h0e)
	) name12762 (
		_w18584_,
		_w18566_,
		_w18588_,
		_w18589_
	);
	LUT3 #(
		.INIT('h65)
	) name12763 (
		\u1_L8_reg[22]/NET0131 ,
		_w18579_,
		_w18589_,
		_w18590_
	);
	LUT4 #(
		.INIT('hc963)
	) name12764 (
		decrypt_pad,
		\u1_R8_reg[24]/NET0131 ,
		\u1_uk_K_r8_reg[2]/NET0131 ,
		\u1_uk_K_r8_reg[37]/P0001 ,
		_w18591_
	);
	LUT4 #(
		.INIT('hc963)
	) name12765 (
		decrypt_pad,
		\u1_R8_reg[23]/NET0131 ,
		\u1_uk_K_r8_reg[0]/NET0131 ,
		\u1_uk_K_r8_reg[35]/NET0131 ,
		_w18592_
	);
	LUT4 #(
		.INIT('hc693)
	) name12766 (
		decrypt_pad,
		\u1_R8_reg[21]/NET0131 ,
		\u1_uk_K_r8_reg[0]/NET0131 ,
		\u1_uk_K_r8_reg[51]/NET0131 ,
		_w18593_
	);
	LUT4 #(
		.INIT('hc693)
	) name12767 (
		decrypt_pad,
		\u1_R8_reg[20]/NET0131 ,
		\u1_uk_K_r8_reg[16]/NET0131 ,
		\u1_uk_K_r8_reg[36]/NET0131 ,
		_w18594_
	);
	LUT4 #(
		.INIT('hc693)
	) name12768 (
		decrypt_pad,
		\u1_R8_reg[22]/NET0131 ,
		\u1_uk_K_r8_reg[22]/NET0131 ,
		\u1_uk_K_r8_reg[42]/NET0131 ,
		_w18595_
	);
	LUT4 #(
		.INIT('h4555)
	) name12769 (
		_w18592_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18596_
	);
	LUT4 #(
		.INIT('h4155)
	) name12770 (
		_w18592_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18597_
	);
	LUT4 #(
		.INIT('hc693)
	) name12771 (
		decrypt_pad,
		\u1_R8_reg[25]/NET0131 ,
		\u1_uk_K_r8_reg[1]/NET0131 ,
		\u1_uk_K_r8_reg[21]/NET0131 ,
		_w18598_
	);
	LUT4 #(
		.INIT('haaa2)
	) name12772 (
		_w18592_,
		_w18598_,
		_w18594_,
		_w18593_,
		_w18599_
	);
	LUT3 #(
		.INIT('he6)
	) name12773 (
		_w18594_,
		_w18595_,
		_w18593_,
		_w18600_
	);
	LUT3 #(
		.INIT('h13)
	) name12774 (
		_w18599_,
		_w18597_,
		_w18600_,
		_w18601_
	);
	LUT4 #(
		.INIT('h0080)
	) name12775 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18602_
	);
	LUT2 #(
		.INIT('h4)
	) name12776 (
		_w18598_,
		_w18594_,
		_w18603_
	);
	LUT3 #(
		.INIT('hce)
	) name12777 (
		_w18592_,
		_w18595_,
		_w18593_,
		_w18604_
	);
	LUT3 #(
		.INIT('h31)
	) name12778 (
		_w18603_,
		_w18602_,
		_w18604_,
		_w18605_
	);
	LUT3 #(
		.INIT('h45)
	) name12779 (
		_w18591_,
		_w18601_,
		_w18605_,
		_w18606_
	);
	LUT4 #(
		.INIT('h0004)
	) name12780 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18607_
	);
	LUT4 #(
		.INIT('h47fb)
	) name12781 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18608_
	);
	LUT2 #(
		.INIT('h2)
	) name12782 (
		_w18592_,
		_w18608_,
		_w18609_
	);
	LUT4 #(
		.INIT('h0040)
	) name12783 (
		_w18592_,
		_w18598_,
		_w18594_,
		_w18595_,
		_w18610_
	);
	LUT2 #(
		.INIT('h4)
	) name12784 (
		_w18593_,
		_w18610_,
		_w18611_
	);
	LUT4 #(
		.INIT('h7270)
	) name12785 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18612_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name12786 (
		_w18593_,
		_w18610_,
		_w18596_,
		_w18612_,
		_w18613_
	);
	LUT3 #(
		.INIT('h8a)
	) name12787 (
		_w18591_,
		_w18609_,
		_w18613_,
		_w18614_
	);
	LUT4 #(
		.INIT('h4555)
	) name12788 (
		_w18592_,
		_w18598_,
		_w18594_,
		_w18593_,
		_w18615_
	);
	LUT3 #(
		.INIT('h01)
	) name12789 (
		_w18595_,
		_w18615_,
		_w18599_,
		_w18616_
	);
	LUT4 #(
		.INIT('h0100)
	) name12790 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18617_
	);
	LUT4 #(
		.INIT('h7e7f)
	) name12791 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18618_
	);
	LUT3 #(
		.INIT('h01)
	) name12792 (
		_w18598_,
		_w18594_,
		_w18593_,
		_w18619_
	);
	LUT4 #(
		.INIT('he4f5)
	) name12793 (
		_w18592_,
		_w18595_,
		_w18618_,
		_w18619_,
		_w18620_
	);
	LUT2 #(
		.INIT('h4)
	) name12794 (
		_w18616_,
		_w18620_,
		_w18621_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name12795 (
		\u1_L8_reg[11]/NET0131 ,
		_w18614_,
		_w18606_,
		_w18621_,
		_w18622_
	);
	LUT4 #(
		.INIT('hc693)
	) name12796 (
		decrypt_pad,
		\u1_R8_reg[16]/NET0131 ,
		\u1_uk_K_r8_reg[13]/P0001 ,
		\u1_uk_K_r8_reg[3]/NET0131 ,
		_w18623_
	);
	LUT4 #(
		.INIT('hc963)
	) name12797 (
		decrypt_pad,
		\u1_R8_reg[15]/NET0131 ,
		\u1_uk_K_r8_reg[27]/NET0131 ,
		\u1_uk_K_r8_reg[5]/NET0131 ,
		_w18624_
	);
	LUT4 #(
		.INIT('hc693)
	) name12798 (
		decrypt_pad,
		\u1_R8_reg[17]/NET0131 ,
		\u1_uk_K_r8_reg[18]/NET0131 ,
		\u1_uk_K_r8_reg[40]/NET0131 ,
		_w18625_
	);
	LUT4 #(
		.INIT('hc963)
	) name12799 (
		decrypt_pad,
		\u1_R8_reg[13]/NET0131 ,
		\u1_uk_K_r8_reg[18]/NET0131 ,
		\u1_uk_K_r8_reg[53]/NET0131 ,
		_w18626_
	);
	LUT4 #(
		.INIT('hc963)
	) name12800 (
		decrypt_pad,
		\u1_R8_reg[14]/NET0131 ,
		\u1_uk_K_r8_reg[19]/NET0131 ,
		\u1_uk_K_r8_reg[54]/NET0131 ,
		_w18627_
	);
	LUT4 #(
		.INIT('hc963)
	) name12801 (
		decrypt_pad,
		\u1_R8_reg[12]/NET0131 ,
		\u1_uk_K_r8_reg[24]/NET0131 ,
		\u1_uk_K_r8_reg[34]/NET0131 ,
		_w18628_
	);
	LUT4 #(
		.INIT('hbf15)
	) name12802 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18629_
	);
	LUT2 #(
		.INIT('h1)
	) name12803 (
		_w18624_,
		_w18629_,
		_w18630_
	);
	LUT2 #(
		.INIT('h8)
	) name12804 (
		_w18626_,
		_w18624_,
		_w18631_
	);
	LUT4 #(
		.INIT('h8000)
	) name12805 (
		_w18625_,
		_w18628_,
		_w18626_,
		_w18624_,
		_w18632_
	);
	LUT4 #(
		.INIT('h1000)
	) name12806 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18633_
	);
	LUT2 #(
		.INIT('h8)
	) name12807 (
		_w18627_,
		_w18624_,
		_w18634_
	);
	LUT4 #(
		.INIT('h4000)
	) name12808 (
		_w18628_,
		_w18627_,
		_w18626_,
		_w18624_,
		_w18635_
	);
	LUT3 #(
		.INIT('h01)
	) name12809 (
		_w18633_,
		_w18635_,
		_w18632_,
		_w18636_
	);
	LUT3 #(
		.INIT('h02)
	) name12810 (
		_w18628_,
		_w18627_,
		_w18626_,
		_w18637_
	);
	LUT4 #(
		.INIT('h0008)
	) name12811 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18638_
	);
	LUT3 #(
		.INIT('h01)
	) name12812 (
		_w18625_,
		_w18628_,
		_w18626_,
		_w18639_
	);
	LUT2 #(
		.INIT('h2)
	) name12813 (
		_w18627_,
		_w18624_,
		_w18640_
	);
	LUT3 #(
		.INIT('h31)
	) name12814 (
		_w18639_,
		_w18638_,
		_w18640_,
		_w18641_
	);
	LUT4 #(
		.INIT('h4555)
	) name12815 (
		_w18623_,
		_w18630_,
		_w18636_,
		_w18641_,
		_w18642_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name12816 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18643_
	);
	LUT4 #(
		.INIT('h00de)
	) name12817 (
		_w18628_,
		_w18627_,
		_w18626_,
		_w18624_,
		_w18644_
	);
	LUT4 #(
		.INIT('h0200)
	) name12818 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18645_
	);
	LUT4 #(
		.INIT('h7dff)
	) name12819 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18646_
	);
	LUT4 #(
		.INIT('h4000)
	) name12820 (
		_w18625_,
		_w18628_,
		_w18626_,
		_w18624_,
		_w18647_
	);
	LUT4 #(
		.INIT('hbdff)
	) name12821 (
		_w18625_,
		_w18628_,
		_w18626_,
		_w18624_,
		_w18648_
	);
	LUT4 #(
		.INIT('h8a00)
	) name12822 (
		_w18646_,
		_w18643_,
		_w18644_,
		_w18648_,
		_w18649_
	);
	LUT4 #(
		.INIT('hffbe)
	) name12823 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18650_
	);
	LUT2 #(
		.INIT('h2)
	) name12824 (
		_w18624_,
		_w18650_,
		_w18651_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name12825 (
		_w18627_,
		_w18645_,
		_w18624_,
		_w18647_,
		_w18652_
	);
	LUT4 #(
		.INIT('h0d00)
	) name12826 (
		_w18623_,
		_w18649_,
		_w18651_,
		_w18652_,
		_w18653_
	);
	LUT3 #(
		.INIT('h65)
	) name12827 (
		\u1_L8_reg[20]/NET0131 ,
		_w18642_,
		_w18653_,
		_w18654_
	);
	LUT4 #(
		.INIT('hc963)
	) name12828 (
		decrypt_pad,
		\u1_R8_reg[31]/P0001 ,
		\u1_uk_K_r8_reg[23]/NET0131 ,
		\u1_uk_K_r8_reg[31]/NET0131 ,
		_w18655_
	);
	LUT4 #(
		.INIT('hc693)
	) name12829 (
		decrypt_pad,
		\u1_R8_reg[28]/NET0131 ,
		\u1_uk_K_r8_reg[42]/NET0131 ,
		\u1_uk_K_r8_reg[7]/NET0131 ,
		_w18656_
	);
	LUT4 #(
		.INIT('hc693)
	) name12830 (
		decrypt_pad,
		\u1_R8_reg[30]/NET0131 ,
		\u1_uk_K_r8_reg[15]/NET0131 ,
		\u1_uk_K_r8_reg[35]/NET0131 ,
		_w18657_
	);
	LUT2 #(
		.INIT('h2)
	) name12831 (
		_w18656_,
		_w18657_,
		_w18658_
	);
	LUT4 #(
		.INIT('hc693)
	) name12832 (
		decrypt_pad,
		\u1_R8_reg[1]/NET0131 ,
		\u1_uk_K_r8_reg[30]/NET0131 ,
		\u1_uk_K_r8_reg[50]/NET0131 ,
		_w18659_
	);
	LUT4 #(
		.INIT('hc693)
	) name12833 (
		decrypt_pad,
		\u1_R8_reg[29]/NET0131 ,
		\u1_uk_K_r8_reg[14]/NET0131 ,
		\u1_uk_K_r8_reg[38]/NET0131 ,
		_w18660_
	);
	LUT2 #(
		.INIT('h4)
	) name12834 (
		_w18659_,
		_w18660_,
		_w18661_
	);
	LUT4 #(
		.INIT('hc963)
	) name12835 (
		decrypt_pad,
		\u1_R8_reg[32]/NET0131 ,
		\u1_uk_K_r8_reg[29]/NET0131 ,
		\u1_uk_K_r8_reg[9]/NET0131 ,
		_w18662_
	);
	LUT4 #(
		.INIT('h0020)
	) name12836 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18663_
	);
	LUT4 #(
		.INIT('h1000)
	) name12837 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18664_
	);
	LUT2 #(
		.INIT('h1)
	) name12838 (
		_w18660_,
		_w18657_,
		_w18665_
	);
	LUT4 #(
		.INIT('heff7)
	) name12839 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18666_
	);
	LUT4 #(
		.INIT('h0400)
	) name12840 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18667_
	);
	LUT3 #(
		.INIT('h01)
	) name12841 (
		_w18656_,
		_w18660_,
		_w18657_,
		_w18668_
	);
	LUT4 #(
		.INIT('h0001)
	) name12842 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18669_
	);
	LUT4 #(
		.INIT('hebf6)
	) name12843 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18670_
	);
	LUT4 #(
		.INIT('hd700)
	) name12844 (
		_w18662_,
		_w18658_,
		_w18661_,
		_w18670_,
		_w18671_
	);
	LUT2 #(
		.INIT('h2)
	) name12845 (
		_w18655_,
		_w18671_,
		_w18672_
	);
	LUT4 #(
		.INIT('h0200)
	) name12846 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18673_
	);
	LUT4 #(
		.INIT('haa8a)
	) name12847 (
		_w18655_,
		_w18656_,
		_w18659_,
		_w18660_,
		_w18674_
	);
	LUT3 #(
		.INIT('h10)
	) name12848 (
		_w18656_,
		_w18659_,
		_w18657_,
		_w18675_
	);
	LUT3 #(
		.INIT('h15)
	) name12849 (
		_w18655_,
		_w18659_,
		_w18660_,
		_w18676_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12850 (
		_w18673_,
		_w18674_,
		_w18675_,
		_w18676_,
		_w18677_
	);
	LUT4 #(
		.INIT('h8000)
	) name12851 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18678_
	);
	LUT3 #(
		.INIT('h04)
	) name12852 (
		_w18655_,
		_w18656_,
		_w18657_,
		_w18679_
	);
	LUT3 #(
		.INIT('h01)
	) name12853 (
		_w18663_,
		_w18679_,
		_w18678_,
		_w18680_
	);
	LUT3 #(
		.INIT('h45)
	) name12854 (
		_w18662_,
		_w18677_,
		_w18680_,
		_w18681_
	);
	LUT2 #(
		.INIT('h4)
	) name12855 (
		_w18655_,
		_w18663_,
		_w18682_
	);
	LUT4 #(
		.INIT('h4000)
	) name12856 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18683_
	);
	LUT4 #(
		.INIT('hb5fa)
	) name12857 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18684_
	);
	LUT4 #(
		.INIT('h00a2)
	) name12858 (
		_w18662_,
		_w18655_,
		_w18683_,
		_w18684_,
		_w18685_
	);
	LUT2 #(
		.INIT('h1)
	) name12859 (
		_w18682_,
		_w18685_,
		_w18686_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name12860 (
		\u1_L8_reg[5]/NET0131 ,
		_w18681_,
		_w18672_,
		_w18686_,
		_w18687_
	);
	LUT4 #(
		.INIT('hdcfe)
	) name12861 (
		_w18625_,
		_w18628_,
		_w18626_,
		_w18624_,
		_w18688_
	);
	LUT2 #(
		.INIT('h1)
	) name12862 (
		_w18634_,
		_w18688_,
		_w18689_
	);
	LUT3 #(
		.INIT('hf2)
	) name12863 (
		_w18625_,
		_w18627_,
		_w18626_,
		_w18690_
	);
	LUT2 #(
		.INIT('h8)
	) name12864 (
		_w18628_,
		_w18624_,
		_w18691_
	);
	LUT4 #(
		.INIT('h0008)
	) name12865 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18624_,
		_w18692_
	);
	LUT4 #(
		.INIT('he3ff)
	) name12866 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18693_
	);
	LUT4 #(
		.INIT('h2300)
	) name12867 (
		_w18690_,
		_w18692_,
		_w18691_,
		_w18693_,
		_w18694_
	);
	LUT3 #(
		.INIT('h45)
	) name12868 (
		_w18623_,
		_w18689_,
		_w18694_,
		_w18695_
	);
	LUT4 #(
		.INIT('hb1bb)
	) name12869 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18696_
	);
	LUT4 #(
		.INIT('h00df)
	) name12870 (
		_w18628_,
		_w18627_,
		_w18626_,
		_w18624_,
		_w18697_
	);
	LUT2 #(
		.INIT('h4)
	) name12871 (
		_w18696_,
		_w18697_,
		_w18698_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name12872 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18699_
	);
	LUT4 #(
		.INIT('h1d00)
	) name12873 (
		_w18625_,
		_w18628_,
		_w18626_,
		_w18624_,
		_w18700_
	);
	LUT3 #(
		.INIT('h2a)
	) name12874 (
		_w18699_,
		_w18690_,
		_w18700_,
		_w18701_
	);
	LUT3 #(
		.INIT('h8a)
	) name12875 (
		_w18623_,
		_w18698_,
		_w18701_,
		_w18702_
	);
	LUT4 #(
		.INIT('h7fde)
	) name12876 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18703_
	);
	LUT2 #(
		.INIT('h1)
	) name12877 (
		_w18624_,
		_w18703_,
		_w18704_
	);
	LUT3 #(
		.INIT('h0b)
	) name12878 (
		_w18627_,
		_w18647_,
		_w18635_,
		_w18705_
	);
	LUT2 #(
		.INIT('h4)
	) name12879 (
		_w18704_,
		_w18705_,
		_w18706_
	);
	LUT4 #(
		.INIT('h5655)
	) name12880 (
		\u1_L8_reg[10]/NET0131 ,
		_w18702_,
		_w18695_,
		_w18706_,
		_w18707_
	);
	LUT4 #(
		.INIT('h2000)
	) name12881 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18708_
	);
	LUT4 #(
		.INIT('h0006)
	) name12882 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18709_
	);
	LUT4 #(
		.INIT('h0800)
	) name12883 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18710_
	);
	LUT4 #(
		.INIT('h0001)
	) name12884 (
		_w18566_,
		_w18709_,
		_w18708_,
		_w18710_,
		_w18711_
	);
	LUT3 #(
		.INIT('h04)
	) name12885 (
		_w18570_,
		_w18568_,
		_w18572_,
		_w18712_
	);
	LUT4 #(
		.INIT('h5545)
	) name12886 (
		_w18567_,
		_w18570_,
		_w18568_,
		_w18572_,
		_w18713_
	);
	LUT2 #(
		.INIT('h6)
	) name12887 (
		_w18568_,
		_w18572_,
		_w18714_
	);
	LUT4 #(
		.INIT('h0310)
	) name12888 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18715_
	);
	LUT2 #(
		.INIT('h6)
	) name12889 (
		_w18571_,
		_w18572_,
		_w18716_
	);
	LUT4 #(
		.INIT('h134c)
	) name12890 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18717_
	);
	LUT4 #(
		.INIT('h1f0a)
	) name12891 (
		_w18567_,
		_w18712_,
		_w18715_,
		_w18717_,
		_w18718_
	);
	LUT2 #(
		.INIT('h8)
	) name12892 (
		_w18711_,
		_w18718_,
		_w18719_
	);
	LUT4 #(
		.INIT('h1400)
	) name12893 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18720_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name12894 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w18721_
	);
	LUT2 #(
		.INIT('h2)
	) name12895 (
		_w18567_,
		_w18721_,
		_w18722_
	);
	LUT4 #(
		.INIT('h0c04)
	) name12896 (
		_w18567_,
		_w18570_,
		_w18571_,
		_w18568_,
		_w18723_
	);
	LUT4 #(
		.INIT('h0222)
	) name12897 (
		_w18566_,
		_w18586_,
		_w18714_,
		_w18723_,
		_w18724_
	);
	LUT3 #(
		.INIT('h10)
	) name12898 (
		_w18722_,
		_w18720_,
		_w18724_,
		_w18725_
	);
	LUT3 #(
		.INIT('ha9)
	) name12899 (
		\u1_L8_reg[12]/NET0131 ,
		_w18719_,
		_w18725_,
		_w18726_
	);
	LUT4 #(
		.INIT('hc963)
	) name12900 (
		decrypt_pad,
		\u1_R8_reg[19]/NET0131 ,
		\u1_uk_K_r8_reg[30]/NET0131 ,
		\u1_uk_K_r8_reg[38]/NET0131 ,
		_w18727_
	);
	LUT4 #(
		.INIT('hc963)
	) name12901 (
		decrypt_pad,
		\u1_R8_reg[21]/NET0131 ,
		\u1_uk_K_r8_reg[15]/NET0131 ,
		\u1_uk_K_r8_reg[50]/NET0131 ,
		_w18728_
	);
	LUT4 #(
		.INIT('hc693)
	) name12902 (
		decrypt_pad,
		\u1_R8_reg[17]/NET0131 ,
		\u1_uk_K_r8_reg[29]/NET0131 ,
		\u1_uk_K_r8_reg[49]/NET0131 ,
		_w18729_
	);
	LUT4 #(
		.INIT('hc963)
	) name12903 (
		decrypt_pad,
		\u1_R8_reg[16]/NET0131 ,
		\u1_uk_K_r8_reg[31]/NET0131 ,
		\u1_uk_K_r8_reg[7]/NET0131 ,
		_w18730_
	);
	LUT4 #(
		.INIT('hc693)
	) name12904 (
		decrypt_pad,
		\u1_R8_reg[18]/NET0131 ,
		\u1_uk_K_r8_reg[23]/NET0131 ,
		\u1_uk_K_r8_reg[43]/NET0131 ,
		_w18731_
	);
	LUT2 #(
		.INIT('h6)
	) name12905 (
		_w18728_,
		_w18729_,
		_w18732_
	);
	LUT4 #(
		.INIT('hcb79)
	) name12906 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18733_
	);
	LUT3 #(
		.INIT('h04)
	) name12907 (
		_w18730_,
		_w18729_,
		_w18731_,
		_w18734_
	);
	LUT4 #(
		.INIT('h76ae)
	) name12908 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18735_
	);
	LUT4 #(
		.INIT('h0810)
	) name12909 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18736_
	);
	LUT4 #(
		.INIT('h00b8)
	) name12910 (
		_w18735_,
		_w18727_,
		_w18733_,
		_w18736_,
		_w18737_
	);
	LUT4 #(
		.INIT('hc963)
	) name12911 (
		decrypt_pad,
		\u1_R8_reg[20]/NET0131 ,
		\u1_uk_K_r8_reg[14]/NET0131 ,
		\u1_uk_K_r8_reg[49]/NET0131 ,
		_w18738_
	);
	LUT2 #(
		.INIT('h1)
	) name12912 (
		_w18737_,
		_w18738_,
		_w18739_
	);
	LUT2 #(
		.INIT('h2)
	) name12913 (
		_w18731_,
		_w18727_,
		_w18740_
	);
	LUT3 #(
		.INIT('h80)
	) name12914 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18741_
	);
	LUT2 #(
		.INIT('h8)
	) name12915 (
		_w18740_,
		_w18741_,
		_w18742_
	);
	LUT3 #(
		.INIT('h01)
	) name12916 (
		_w18730_,
		_w18731_,
		_w18727_,
		_w18743_
	);
	LUT4 #(
		.INIT('h0200)
	) name12917 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18744_
	);
	LUT3 #(
		.INIT('h0b)
	) name12918 (
		_w18732_,
		_w18743_,
		_w18744_,
		_w18745_
	);
	LUT4 #(
		.INIT('h0028)
	) name12919 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18746_
	);
	LUT3 #(
		.INIT('h90)
	) name12920 (
		_w18730_,
		_w18728_,
		_w18731_,
		_w18747_
	);
	LUT3 #(
		.INIT('he0)
	) name12921 (
		_w18728_,
		_w18729_,
		_w18727_,
		_w18748_
	);
	LUT4 #(
		.INIT('h3233)
	) name12922 (
		_w18734_,
		_w18746_,
		_w18747_,
		_w18748_,
		_w18749_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name12923 (
		_w18738_,
		_w18742_,
		_w18745_,
		_w18749_,
		_w18750_
	);
	LUT4 #(
		.INIT('h0020)
	) name12924 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18751_
	);
	LUT4 #(
		.INIT('hfedf)
	) name12925 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18752_
	);
	LUT4 #(
		.INIT('h0400)
	) name12926 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18753_
	);
	LUT4 #(
		.INIT('hebff)
	) name12927 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18754_
	);
	LUT3 #(
		.INIT('hd8)
	) name12928 (
		_w18727_,
		_w18752_,
		_w18754_,
		_w18755_
	);
	LUT4 #(
		.INIT('h5655)
	) name12929 (
		\u1_L8_reg[14]/NET0131 ,
		_w18739_,
		_w18750_,
		_w18755_,
		_w18756_
	);
	LUT4 #(
		.INIT('h5b4b)
	) name12930 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18757_
	);
	LUT4 #(
		.INIT('h0002)
	) name12931 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18758_
	);
	LUT4 #(
		.INIT('h5504)
	) name12932 (
		_w18662_,
		_w18655_,
		_w18757_,
		_w18758_,
		_w18759_
	);
	LUT4 #(
		.INIT('h0004)
	) name12933 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18760_
	);
	LUT3 #(
		.INIT('h02)
	) name12934 (
		_w18655_,
		_w18683_,
		_w18760_,
		_w18761_
	);
	LUT4 #(
		.INIT('h0040)
	) name12935 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18762_
	);
	LUT4 #(
		.INIT('h0c04)
	) name12936 (
		_w18662_,
		_w18656_,
		_w18660_,
		_w18657_,
		_w18763_
	);
	LUT4 #(
		.INIT('h0001)
	) name12937 (
		_w18655_,
		_w18664_,
		_w18762_,
		_w18763_,
		_w18764_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name12938 (
		_w18655_,
		_w18656_,
		_w18659_,
		_w18657_,
		_w18765_
	);
	LUT3 #(
		.INIT('h0e)
	) name12939 (
		_w18655_,
		_w18659_,
		_w18660_,
		_w18766_
	);
	LUT4 #(
		.INIT('h0800)
	) name12940 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18767_
	);
	LUT4 #(
		.INIT('he75f)
	) name12941 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18768_
	);
	LUT4 #(
		.INIT('h20aa)
	) name12942 (
		_w18662_,
		_w18765_,
		_w18766_,
		_w18768_,
		_w18769_
	);
	LUT4 #(
		.INIT('h00dc)
	) name12943 (
		_w18669_,
		_w18761_,
		_w18764_,
		_w18769_,
		_w18770_
	);
	LUT3 #(
		.INIT('h65)
	) name12944 (
		\u1_L8_reg[15]/P0001 ,
		_w18759_,
		_w18770_,
		_w18771_
	);
	LUT4 #(
		.INIT('h4010)
	) name12945 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18772_
	);
	LUT2 #(
		.INIT('h1)
	) name12946 (
		_w18624_,
		_w18772_,
		_w18773_
	);
	LUT4 #(
		.INIT('hff51)
	) name12947 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18774_
	);
	LUT2 #(
		.INIT('h2)
	) name12948 (
		_w18623_,
		_w18774_,
		_w18775_
	);
	LUT3 #(
		.INIT('h20)
	) name12949 (
		_w18624_,
		_w18633_,
		_w18699_,
		_w18776_
	);
	LUT3 #(
		.INIT('h45)
	) name12950 (
		_w18773_,
		_w18775_,
		_w18776_,
		_w18777_
	);
	LUT4 #(
		.INIT('hfebe)
	) name12951 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18778_
	);
	LUT2 #(
		.INIT('h2)
	) name12952 (
		_w18624_,
		_w18778_,
		_w18779_
	);
	LUT3 #(
		.INIT('h4c)
	) name12953 (
		_w18625_,
		_w18628_,
		_w18626_,
		_w18780_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12954 (
		_w18625_,
		_w18627_,
		_w18626_,
		_w18624_,
		_w18781_
	);
	LUT4 #(
		.INIT('h0444)
	) name12955 (
		_w18623_,
		_w18646_,
		_w18780_,
		_w18781_,
		_w18782_
	);
	LUT3 #(
		.INIT('h2b)
	) name12956 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18783_
	);
	LUT4 #(
		.INIT('hbf94)
	) name12957 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18624_,
		_w18784_
	);
	LUT4 #(
		.INIT('haa8a)
	) name12958 (
		_w18623_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18785_
	);
	LUT3 #(
		.INIT('hd0)
	) name12959 (
		_w18626_,
		_w18784_,
		_w18785_,
		_w18786_
	);
	LUT3 #(
		.INIT('h0b)
	) name12960 (
		_w18779_,
		_w18782_,
		_w18786_,
		_w18787_
	);
	LUT3 #(
		.INIT('h56)
	) name12961 (
		\u1_L8_reg[1]/NET0131 ,
		_w18777_,
		_w18787_,
		_w18788_
	);
	LUT4 #(
		.INIT('hc693)
	) name12962 (
		decrypt_pad,
		\u1_R8_reg[5]/NET0131 ,
		\u1_uk_K_r8_reg[39]/NET0131 ,
		\u1_uk_K_r8_reg[4]/NET0131 ,
		_w18789_
	);
	LUT4 #(
		.INIT('hc693)
	) name12963 (
		decrypt_pad,
		\u1_R8_reg[2]/NET0131 ,
		\u1_uk_K_r8_reg[24]/NET0131 ,
		\u1_uk_K_r8_reg[46]/NET0131 ,
		_w18790_
	);
	LUT4 #(
		.INIT('hc693)
	) name12964 (
		decrypt_pad,
		\u1_R8_reg[1]/NET0131 ,
		\u1_uk_K_r8_reg[41]/NET0131 ,
		\u1_uk_K_r8_reg[6]/NET0131 ,
		_w18791_
	);
	LUT4 #(
		.INIT('hc963)
	) name12965 (
		decrypt_pad,
		\u1_R8_reg[32]/NET0131 ,
		\u1_uk_K_r8_reg[10]/NET0131 ,
		\u1_uk_K_r8_reg[20]/NET0131 ,
		_w18792_
	);
	LUT4 #(
		.INIT('h0208)
	) name12966 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w18793_
	);
	LUT4 #(
		.INIT('hc693)
	) name12967 (
		decrypt_pad,
		\u1_R8_reg[3]/NET0131 ,
		\u1_uk_K_r8_reg[33]/NET0131 ,
		\u1_uk_K_r8_reg[55]/NET0131 ,
		_w18794_
	);
	LUT4 #(
		.INIT('h6f00)
	) name12968 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18794_,
		_w18795_
	);
	LUT3 #(
		.INIT('h41)
	) name12969 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18796_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name12970 (
		_w18789_,
		_w18792_,
		_w18794_,
		_w18790_,
		_w18797_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12971 (
		_w18793_,
		_w18795_,
		_w18796_,
		_w18797_,
		_w18798_
	);
	LUT4 #(
		.INIT('h2400)
	) name12972 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w18799_
	);
	LUT4 #(
		.INIT('hc693)
	) name12973 (
		decrypt_pad,
		\u1_R8_reg[4]/NET0131 ,
		\u1_uk_K_r8_reg[11]/NET0131 ,
		\u1_uk_K_r8_reg[33]/NET0131 ,
		_w18800_
	);
	LUT2 #(
		.INIT('h1)
	) name12974 (
		_w18799_,
		_w18800_,
		_w18801_
	);
	LUT4 #(
		.INIT('h0040)
	) name12975 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w18802_
	);
	LUT4 #(
		.INIT('hf0b5)
	) name12976 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w18803_
	);
	LUT2 #(
		.INIT('h2)
	) name12977 (
		_w18794_,
		_w18803_,
		_w18804_
	);
	LUT4 #(
		.INIT('h0c01)
	) name12978 (
		_w18791_,
		_w18792_,
		_w18794_,
		_w18790_,
		_w18805_
	);
	LUT3 #(
		.INIT('h20)
	) name12979 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18806_
	);
	LUT4 #(
		.INIT('h0020)
	) name12980 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w18807_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12981 (
		_w18791_,
		_w18789_,
		_w18790_,
		_w18800_,
		_w18808_
	);
	LUT3 #(
		.INIT('h10)
	) name12982 (
		_w18807_,
		_w18805_,
		_w18808_,
		_w18809_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12983 (
		_w18798_,
		_w18801_,
		_w18804_,
		_w18809_,
		_w18810_
	);
	LUT2 #(
		.INIT('h6)
	) name12984 (
		\u1_L8_reg[17]/NET0131 ,
		_w18810_,
		_w18811_
	);
	LUT4 #(
		.INIT('h5551)
	) name12985 (
		_w18655_,
		_w18656_,
		_w18659_,
		_w18657_,
		_w18812_
	);
	LUT4 #(
		.INIT('he040)
	) name12986 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18813_
	);
	LUT4 #(
		.INIT('haaa2)
	) name12987 (
		_w18655_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18814_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name12988 (
		_w18767_,
		_w18812_,
		_w18813_,
		_w18814_,
		_w18815_
	);
	LUT4 #(
		.INIT('h2100)
	) name12989 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18816_
	);
	LUT3 #(
		.INIT('h02)
	) name12990 (
		_w18662_,
		_w18760_,
		_w18816_,
		_w18817_
	);
	LUT2 #(
		.INIT('h4)
	) name12991 (
		_w18815_,
		_w18817_,
		_w18818_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name12992 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18819_
	);
	LUT4 #(
		.INIT('h0040)
	) name12993 (
		_w18655_,
		_w18656_,
		_w18659_,
		_w18657_,
		_w18820_
	);
	LUT4 #(
		.INIT('h0888)
	) name12994 (
		_w18655_,
		_w18656_,
		_w18659_,
		_w18660_,
		_w18821_
	);
	LUT4 #(
		.INIT('h2300)
	) name12995 (
		_w18665_,
		_w18820_,
		_w18821_,
		_w18819_,
		_w18822_
	);
	LUT4 #(
		.INIT('hccef)
	) name12996 (
		_w18655_,
		_w18656_,
		_w18659_,
		_w18660_,
		_w18823_
	);
	LUT2 #(
		.INIT('h2)
	) name12997 (
		_w18657_,
		_w18823_,
		_w18824_
	);
	LUT4 #(
		.INIT('h0080)
	) name12998 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w18825_
	);
	LUT4 #(
		.INIT('h0100)
	) name12999 (
		_w18655_,
		_w18656_,
		_w18659_,
		_w18660_,
		_w18826_
	);
	LUT3 #(
		.INIT('h01)
	) name13000 (
		_w18662_,
		_w18826_,
		_w18825_,
		_w18827_
	);
	LUT3 #(
		.INIT('h40)
	) name13001 (
		_w18824_,
		_w18827_,
		_w18822_,
		_w18828_
	);
	LUT4 #(
		.INIT('h0002)
	) name13002 (
		_w18655_,
		_w18656_,
		_w18660_,
		_w18657_,
		_w18829_
	);
	LUT3 #(
		.INIT('h0b)
	) name13003 (
		_w18655_,
		_w18825_,
		_w18829_,
		_w18830_
	);
	LUT4 #(
		.INIT('ha955)
	) name13004 (
		\u1_L8_reg[21]/NET0131 ,
		_w18818_,
		_w18828_,
		_w18830_,
		_w18831_
	);
	LUT3 #(
		.INIT('h08)
	) name13005 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18832_
	);
	LUT4 #(
		.INIT('h00f7)
	) name13006 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18727_,
		_w18833_
	);
	LUT4 #(
		.INIT('h7a00)
	) name13007 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18727_,
		_w18834_
	);
	LUT4 #(
		.INIT('heefc)
	) name13008 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18835_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name13009 (
		_w18734_,
		_w18833_,
		_w18834_,
		_w18835_,
		_w18836_
	);
	LUT3 #(
		.INIT('h40)
	) name13010 (
		_w18728_,
		_w18729_,
		_w18731_,
		_w18837_
	);
	LUT4 #(
		.INIT('h2000)
	) name13011 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18838_
	);
	LUT4 #(
		.INIT('hf700)
	) name13012 (
		_w18728_,
		_w18729_,
		_w18731_,
		_w18738_,
		_w18839_
	);
	LUT2 #(
		.INIT('h4)
	) name13013 (
		_w18838_,
		_w18839_,
		_w18840_
	);
	LUT3 #(
		.INIT('hb0)
	) name13014 (
		_w18728_,
		_w18729_,
		_w18727_,
		_w18841_
	);
	LUT3 #(
		.INIT('h0e)
	) name13015 (
		_w18730_,
		_w18729_,
		_w18727_,
		_w18842_
	);
	LUT4 #(
		.INIT('h0f01)
	) name13016 (
		_w18730_,
		_w18729_,
		_w18731_,
		_w18727_,
		_w18843_
	);
	LUT2 #(
		.INIT('h4)
	) name13017 (
		_w18841_,
		_w18843_,
		_w18844_
	);
	LUT4 #(
		.INIT('h5702)
	) name13018 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18845_
	);
	LUT3 #(
		.INIT('h40)
	) name13019 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18846_
	);
	LUT4 #(
		.INIT('h4000)
	) name13020 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18847_
	);
	LUT4 #(
		.INIT('h0111)
	) name13021 (
		_w18738_,
		_w18847_,
		_w18842_,
		_w18845_,
		_w18848_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name13022 (
		_w18836_,
		_w18840_,
		_w18844_,
		_w18848_,
		_w18849_
	);
	LUT4 #(
		.INIT('hdeff)
	) name13023 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18850_
	);
	LUT4 #(
		.INIT('hdefb)
	) name13024 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18851_
	);
	LUT4 #(
		.INIT('h0020)
	) name13025 (
		_w18730_,
		_w18729_,
		_w18731_,
		_w18727_,
		_w18852_
	);
	LUT4 #(
		.INIT('h0080)
	) name13026 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w18853_
	);
	LUT4 #(
		.INIT('h0301)
	) name13027 (
		_w18727_,
		_w18852_,
		_w18853_,
		_w18851_,
		_w18854_
	);
	LUT3 #(
		.INIT('h65)
	) name13028 (
		\u1_L8_reg[25]/NET0131 ,
		_w18849_,
		_w18854_,
		_w18855_
	);
	LUT4 #(
		.INIT('h6100)
	) name13029 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18856_
	);
	LUT4 #(
		.INIT('hdfce)
	) name13030 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18857_
	);
	LUT4 #(
		.INIT('h7f7d)
	) name13031 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18858_
	);
	LUT4 #(
		.INIT('ha820)
	) name13032 (
		_w18623_,
		_w18624_,
		_w18858_,
		_w18857_,
		_w18859_
	);
	LUT2 #(
		.INIT('h2)
	) name13033 (
		_w18631_,
		_w18783_,
		_w18860_
	);
	LUT3 #(
		.INIT('h01)
	) name13034 (
		_w18623_,
		_w18645_,
		_w18637_,
		_w18861_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name13035 (
		_w18856_,
		_w18859_,
		_w18860_,
		_w18861_,
		_w18862_
	);
	LUT4 #(
		.INIT('h0904)
	) name13036 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18863_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13037 (
		_w18625_,
		_w18628_,
		_w18627_,
		_w18626_,
		_w18864_
	);
	LUT4 #(
		.INIT('h0032)
	) name13038 (
		_w18623_,
		_w18624_,
		_w18864_,
		_w18863_,
		_w18865_
	);
	LUT3 #(
		.INIT('h04)
	) name13039 (
		_w18645_,
		_w18624_,
		_w18638_,
		_w18866_
	);
	LUT2 #(
		.INIT('h1)
	) name13040 (
		_w18865_,
		_w18866_,
		_w18867_
	);
	LUT3 #(
		.INIT('h56)
	) name13041 (
		\u1_L8_reg[26]/NET0131 ,
		_w18862_,
		_w18867_,
		_w18868_
	);
	LUT4 #(
		.INIT('h67ba)
	) name13042 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18869_
	);
	LUT4 #(
		.INIT('hb4f7)
	) name13043 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18870_
	);
	LUT4 #(
		.INIT('h0020)
	) name13044 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18871_
	);
	LUT4 #(
		.INIT('h00e4)
	) name13045 (
		_w18592_,
		_w18870_,
		_w18869_,
		_w18871_,
		_w18872_
	);
	LUT2 #(
		.INIT('h1)
	) name13046 (
		_w18591_,
		_w18872_,
		_w18873_
	);
	LUT4 #(
		.INIT('h9cff)
	) name13047 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18874_
	);
	LUT2 #(
		.INIT('h2)
	) name13048 (
		_w18592_,
		_w18874_,
		_w18875_
	);
	LUT4 #(
		.INIT('h6f6e)
	) name13049 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18876_
	);
	LUT2 #(
		.INIT('h1)
	) name13050 (
		_w18592_,
		_w18876_,
		_w18877_
	);
	LUT4 #(
		.INIT('h0012)
	) name13051 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18878_
	);
	LUT4 #(
		.INIT('h0010)
	) name13052 (
		_w18592_,
		_w18598_,
		_w18594_,
		_w18595_,
		_w18879_
	);
	LUT3 #(
		.INIT('h01)
	) name13053 (
		_w18602_,
		_w18878_,
		_w18879_,
		_w18880_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name13054 (
		_w18591_,
		_w18875_,
		_w18877_,
		_w18880_,
		_w18881_
	);
	LUT4 #(
		.INIT('h0800)
	) name13055 (
		_w18592_,
		_w18598_,
		_w18595_,
		_w18593_,
		_w18882_
	);
	LUT2 #(
		.INIT('h1)
	) name13056 (
		_w18607_,
		_w18882_,
		_w18883_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name13057 (
		\u1_L8_reg[29]/NET0131 ,
		_w18881_,
		_w18873_,
		_w18883_,
		_w18884_
	);
	LUT4 #(
		.INIT('hc693)
	) name13058 (
		decrypt_pad,
		\u1_R8_reg[8]/NET0131 ,
		\u1_uk_K_r8_reg[12]/NET0131 ,
		\u1_uk_K_r8_reg[34]/NET0131 ,
		_w18885_
	);
	LUT4 #(
		.INIT('hc963)
	) name13059 (
		decrypt_pad,
		\u1_R8_reg[7]/NET0131 ,
		\u1_uk_K_r8_reg[11]/NET0131 ,
		\u1_uk_K_r8_reg[46]/NET0131 ,
		_w18886_
	);
	LUT4 #(
		.INIT('hc963)
	) name13060 (
		decrypt_pad,
		\u1_R8_reg[5]/NET0131 ,
		\u1_uk_K_r8_reg[26]/NET0131 ,
		\u1_uk_K_r8_reg[4]/NET0131 ,
		_w18887_
	);
	LUT4 #(
		.INIT('hc693)
	) name13061 (
		decrypt_pad,
		\u1_R8_reg[4]/NET0131 ,
		\u1_uk_K_r8_reg[25]/NET0131 ,
		\u1_uk_K_r8_reg[47]/NET0131 ,
		_w18888_
	);
	LUT4 #(
		.INIT('hc693)
	) name13062 (
		decrypt_pad,
		\u1_R8_reg[9]/NET0131 ,
		\u1_uk_K_r8_reg[17]/NET0131 ,
		\u1_uk_K_r8_reg[39]/NET0131 ,
		_w18889_
	);
	LUT4 #(
		.INIT('hc963)
	) name13063 (
		decrypt_pad,
		\u1_R8_reg[6]/NET0131 ,
		\u1_uk_K_r8_reg[17]/NET0131 ,
		\u1_uk_K_r8_reg[27]/NET0131 ,
		_w18890_
	);
	LUT3 #(
		.INIT('h5d)
	) name13064 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18891_
	);
	LUT4 #(
		.INIT('h59fb)
	) name13065 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18892_
	);
	LUT2 #(
		.INIT('h1)
	) name13066 (
		_w18886_,
		_w18892_,
		_w18893_
	);
	LUT4 #(
		.INIT('h0034)
	) name13067 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18894_
	);
	LUT4 #(
		.INIT('h0800)
	) name13068 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18895_
	);
	LUT2 #(
		.INIT('h2)
	) name13069 (
		_w18889_,
		_w18890_,
		_w18896_
	);
	LUT4 #(
		.INIT('h0004)
	) name13070 (
		_w18886_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18897_
	);
	LUT4 #(
		.INIT('h4000)
	) name13071 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18898_
	);
	LUT4 #(
		.INIT('h0007)
	) name13072 (
		_w18886_,
		_w18895_,
		_w18897_,
		_w18898_,
		_w18899_
	);
	LUT4 #(
		.INIT('h5455)
	) name13073 (
		_w18885_,
		_w18893_,
		_w18894_,
		_w18899_,
		_w18900_
	);
	LUT4 #(
		.INIT('h0002)
	) name13074 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18901_
	);
	LUT4 #(
		.INIT('h0001)
	) name13075 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18887_,
		_w18902_
	);
	LUT4 #(
		.INIT('h80a0)
	) name13076 (
		_w18886_,
		_w18888_,
		_w18887_,
		_w18890_,
		_w18903_
	);
	LUT3 #(
		.INIT('h01)
	) name13077 (
		_w18902_,
		_w18903_,
		_w18901_,
		_w18904_
	);
	LUT4 #(
		.INIT('h0080)
	) name13078 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18905_
	);
	LUT4 #(
		.INIT('h4500)
	) name13079 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18890_,
		_w18906_
	);
	LUT3 #(
		.INIT('h13)
	) name13080 (
		_w18891_,
		_w18905_,
		_w18906_,
		_w18907_
	);
	LUT4 #(
		.INIT('h4004)
	) name13081 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18908_
	);
	LUT3 #(
		.INIT('h10)
	) name13082 (
		_w18889_,
		_w18887_,
		_w18890_,
		_w18909_
	);
	LUT4 #(
		.INIT('h0100)
	) name13083 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18910_
	);
	LUT3 #(
		.INIT('h08)
	) name13084 (
		_w18888_,
		_w18887_,
		_w18890_,
		_w18911_
	);
	LUT4 #(
		.INIT('heee4)
	) name13085 (
		_w18886_,
		_w18908_,
		_w18911_,
		_w18910_,
		_w18912_
	);
	LUT4 #(
		.INIT('h00d5)
	) name13086 (
		_w18885_,
		_w18904_,
		_w18907_,
		_w18912_,
		_w18913_
	);
	LUT3 #(
		.INIT('h65)
	) name13087 (
		\u1_L8_reg[2]/NET0131 ,
		_w18900_,
		_w18913_,
		_w18914_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name13088 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18915_
	);
	LUT2 #(
		.INIT('h2)
	) name13089 (
		_w18886_,
		_w18915_,
		_w18916_
	);
	LUT4 #(
		.INIT('hbfae)
	) name13090 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18917_
	);
	LUT2 #(
		.INIT('h1)
	) name13091 (
		_w18886_,
		_w18917_,
		_w18918_
	);
	LUT2 #(
		.INIT('h8)
	) name13092 (
		_w18886_,
		_w18888_,
		_w18919_
	);
	LUT4 #(
		.INIT('h7737)
	) name13093 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18887_,
		_w18920_
	);
	LUT4 #(
		.INIT('h0400)
	) name13094 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18921_
	);
	LUT3 #(
		.INIT('h0e)
	) name13095 (
		_w18890_,
		_w18920_,
		_w18921_,
		_w18922_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name13096 (
		_w18885_,
		_w18918_,
		_w18916_,
		_w18922_,
		_w18923_
	);
	LUT4 #(
		.INIT('hdaff)
	) name13097 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18924_
	);
	LUT2 #(
		.INIT('h1)
	) name13098 (
		_w18886_,
		_w18924_,
		_w18925_
	);
	LUT3 #(
		.INIT('h02)
	) name13099 (
		_w18888_,
		_w18889_,
		_w18890_,
		_w18926_
	);
	LUT4 #(
		.INIT('h1145)
	) name13100 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18887_,
		_w18927_
	);
	LUT4 #(
		.INIT('h7077)
	) name13101 (
		_w18886_,
		_w18917_,
		_w18926_,
		_w18927_,
		_w18928_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name13102 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18929_
	);
	LUT4 #(
		.INIT('h2322)
	) name13103 (
		_w18885_,
		_w18925_,
		_w18928_,
		_w18929_,
		_w18930_
	);
	LUT3 #(
		.INIT('h65)
	) name13104 (
		\u1_L8_reg[28]/NET0131 ,
		_w18923_,
		_w18930_,
		_w18931_
	);
	LUT4 #(
		.INIT('hb97d)
	) name13105 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18932_
	);
	LUT2 #(
		.INIT('h2)
	) name13106 (
		_w18592_,
		_w18932_,
		_w18933_
	);
	LUT3 #(
		.INIT('h01)
	) name13107 (
		_w18591_,
		_w18607_,
		_w18610_,
		_w18934_
	);
	LUT3 #(
		.INIT('h80)
	) name13108 (
		_w18598_,
		_w18595_,
		_w18593_,
		_w18935_
	);
	LUT4 #(
		.INIT('h0080)
	) name13109 (
		_w18592_,
		_w18598_,
		_w18594_,
		_w18595_,
		_w18936_
	);
	LUT4 #(
		.INIT('h0002)
	) name13110 (
		_w18591_,
		_w18617_,
		_w18936_,
		_w18935_,
		_w18937_
	);
	LUT3 #(
		.INIT('h0b)
	) name13111 (
		_w18933_,
		_w18934_,
		_w18937_,
		_w18938_
	);
	LUT4 #(
		.INIT('heedf)
	) name13112 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18939_
	);
	LUT3 #(
		.INIT('h01)
	) name13113 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18940_
	);
	LUT4 #(
		.INIT('hf8fc)
	) name13114 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18941_
	);
	LUT4 #(
		.INIT('h3210)
	) name13115 (
		_w18591_,
		_w18940_,
		_w18939_,
		_w18941_,
		_w18942_
	);
	LUT4 #(
		.INIT('h1545)
	) name13116 (
		_w18592_,
		_w18598_,
		_w18594_,
		_w18593_,
		_w18943_
	);
	LUT4 #(
		.INIT('h82a8)
	) name13117 (
		_w18592_,
		_w18598_,
		_w18594_,
		_w18593_,
		_w18944_
	);
	LUT3 #(
		.INIT('h02)
	) name13118 (
		_w18595_,
		_w18944_,
		_w18943_,
		_w18945_
	);
	LUT3 #(
		.INIT('h0e)
	) name13119 (
		_w18592_,
		_w18942_,
		_w18945_,
		_w18946_
	);
	LUT3 #(
		.INIT('h65)
	) name13120 (
		\u1_L8_reg[4]/NET0131 ,
		_w18938_,
		_w18946_,
		_w18947_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name13121 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18948_
	);
	LUT4 #(
		.INIT('hcb6d)
	) name13122 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18949_
	);
	LUT2 #(
		.INIT('h1)
	) name13123 (
		_w18886_,
		_w18949_,
		_w18950_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name13124 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18951_
	);
	LUT4 #(
		.INIT('haa82)
	) name13125 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18887_,
		_w18952_
	);
	LUT2 #(
		.INIT('h4)
	) name13126 (
		_w18951_,
		_w18952_,
		_w18953_
	);
	LUT3 #(
		.INIT('hb0)
	) name13127 (
		_w18889_,
		_w18887_,
		_w18890_,
		_w18954_
	);
	LUT2 #(
		.INIT('h8)
	) name13128 (
		_w18919_,
		_w18954_,
		_w18955_
	);
	LUT3 #(
		.INIT('h32)
	) name13129 (
		_w18886_,
		_w18888_,
		_w18887_,
		_w18956_
	);
	LUT3 #(
		.INIT('h15)
	) name13130 (
		_w18885_,
		_w18896_,
		_w18956_,
		_w18957_
	);
	LUT4 #(
		.INIT('h0100)
	) name13131 (
		_w18955_,
		_w18950_,
		_w18953_,
		_w18957_,
		_w18958_
	);
	LUT3 #(
		.INIT('h01)
	) name13132 (
		_w18889_,
		_w18887_,
		_w18890_,
		_w18959_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name13133 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18890_,
		_w18960_
	);
	LUT4 #(
		.INIT('h5515)
	) name13134 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18887_,
		_w18961_
	);
	LUT4 #(
		.INIT('h8acf)
	) name13135 (
		_w18909_,
		_w18959_,
		_w18960_,
		_w18961_,
		_w18962_
	);
	LUT4 #(
		.INIT('h0010)
	) name13136 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w18963_
	);
	LUT4 #(
		.INIT('h0002)
	) name13137 (
		_w18885_,
		_w18897_,
		_w18898_,
		_w18963_,
		_w18964_
	);
	LUT3 #(
		.INIT('h20)
	) name13138 (
		_w18948_,
		_w18962_,
		_w18964_,
		_w18965_
	);
	LUT3 #(
		.INIT('h56)
	) name13139 (
		\u1_L8_reg[13]/NET0131 ,
		_w18958_,
		_w18965_,
		_w18966_
	);
	LUT4 #(
		.INIT('h0401)
	) name13140 (
		_w18592_,
		_w18598_,
		_w18594_,
		_w18593_,
		_w18967_
	);
	LUT4 #(
		.INIT('h2e33)
	) name13141 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18968_
	);
	LUT4 #(
		.INIT('h8000)
	) name13142 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18969_
	);
	LUT4 #(
		.INIT('h0051)
	) name13143 (
		_w18591_,
		_w18592_,
		_w18968_,
		_w18969_,
		_w18970_
	);
	LUT4 #(
		.INIT('h0800)
	) name13144 (
		_w18592_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18971_
	);
	LUT4 #(
		.INIT('h2000)
	) name13145 (
		_w18598_,
		_w18594_,
		_w18595_,
		_w18593_,
		_w18972_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name13146 (
		_w18591_,
		_w18598_,
		_w18595_,
		_w18593_,
		_w18973_
	);
	LUT3 #(
		.INIT('h10)
	) name13147 (
		_w18972_,
		_w18971_,
		_w18973_,
		_w18974_
	);
	LUT4 #(
		.INIT('h0058)
	) name13148 (
		_w18592_,
		_w18598_,
		_w18594_,
		_w18593_,
		_w18975_
	);
	LUT2 #(
		.INIT('h1)
	) name13149 (
		_w18878_,
		_w18975_,
		_w18976_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name13150 (
		_w18967_,
		_w18970_,
		_w18974_,
		_w18976_,
		_w18977_
	);
	LUT2 #(
		.INIT('h1)
	) name13151 (
		_w18611_,
		_w18616_,
		_w18978_
	);
	LUT3 #(
		.INIT('h65)
	) name13152 (
		\u1_L8_reg[19]/P0001 ,
		_w18977_,
		_w18978_,
		_w18979_
	);
	LUT4 #(
		.INIT('he9f9)
	) name13153 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w18980_
	);
	LUT4 #(
		.INIT('h8000)
	) name13154 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w18981_
	);
	LUT4 #(
		.INIT('h5504)
	) name13155 (
		_w18794_,
		_w18800_,
		_w18980_,
		_w18981_,
		_w18982_
	);
	LUT4 #(
		.INIT('h0800)
	) name13156 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18794_,
		_w18983_
	);
	LUT3 #(
		.INIT('h02)
	) name13157 (
		_w18800_,
		_w18802_,
		_w18983_,
		_w18984_
	);
	LUT2 #(
		.INIT('h8)
	) name13158 (
		_w18794_,
		_w18790_,
		_w18985_
	);
	LUT3 #(
		.INIT('h10)
	) name13159 (
		_w18789_,
		_w18792_,
		_w18790_,
		_w18986_
	);
	LUT2 #(
		.INIT('h4)
	) name13160 (
		_w18791_,
		_w18794_,
		_w18987_
	);
	LUT4 #(
		.INIT('h0777)
	) name13161 (
		_w18806_,
		_w18985_,
		_w18986_,
		_w18987_,
		_w18988_
	);
	LUT4 #(
		.INIT('h2000)
	) name13162 (
		_w18789_,
		_w18792_,
		_w18794_,
		_w18790_,
		_w18989_
	);
	LUT4 #(
		.INIT('h0200)
	) name13163 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18794_,
		_w18990_
	);
	LUT3 #(
		.INIT('h01)
	) name13164 (
		_w18800_,
		_w18990_,
		_w18989_,
		_w18991_
	);
	LUT3 #(
		.INIT('h81)
	) name13165 (
		_w18791_,
		_w18789_,
		_w18790_,
		_w18992_
	);
	LUT3 #(
		.INIT('h15)
	) name13166 (
		_w18791_,
		_w18789_,
		_w18790_,
		_w18993_
	);
	LUT2 #(
		.INIT('h2)
	) name13167 (
		_w18792_,
		_w18794_,
		_w18994_
	);
	LUT3 #(
		.INIT('h45)
	) name13168 (
		_w18992_,
		_w18993_,
		_w18994_,
		_w18995_
	);
	LUT4 #(
		.INIT('h0777)
	) name13169 (
		_w18984_,
		_w18988_,
		_w18991_,
		_w18995_,
		_w18996_
	);
	LUT4 #(
		.INIT('haddb)
	) name13170 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18794_,
		_w18997_
	);
	LUT2 #(
		.INIT('h1)
	) name13171 (
		_w18790_,
		_w18997_,
		_w18998_
	);
	LUT4 #(
		.INIT('haaa9)
	) name13172 (
		\u1_L8_reg[23]/NET0131 ,
		_w18982_,
		_w18996_,
		_w18998_,
		_w18999_
	);
	LUT4 #(
		.INIT('h8090)
	) name13173 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w19000_
	);
	LUT3 #(
		.INIT('h60)
	) name13174 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w19001_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name13175 (
		_w18655_,
		_w18668_,
		_w19000_,
		_w19001_,
		_w19002_
	);
	LUT4 #(
		.INIT('hbdf3)
	) name13176 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w19003_
	);
	LUT3 #(
		.INIT('h8a)
	) name13177 (
		_w18662_,
		_w19002_,
		_w19003_,
		_w19004_
	);
	LUT4 #(
		.INIT('hdc0c)
	) name13178 (
		_w18656_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w19005_
	);
	LUT4 #(
		.INIT('haa8a)
	) name13179 (
		_w18655_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w19006_
	);
	LUT4 #(
		.INIT('h4544)
	) name13180 (
		_w18662_,
		_w18667_,
		_w19005_,
		_w19006_,
		_w19007_
	);
	LUT2 #(
		.INIT('h1)
	) name13181 (
		_w18655_,
		_w18666_,
		_w19008_
	);
	LUT4 #(
		.INIT('h4000)
	) name13182 (
		_w18655_,
		_w18656_,
		_w18659_,
		_w18657_,
		_w19009_
	);
	LUT3 #(
		.INIT('h54)
	) name13183 (
		_w18662_,
		_w18826_,
		_w19009_,
		_w19010_
	);
	LUT4 #(
		.INIT('h0200)
	) name13184 (
		_w18655_,
		_w18659_,
		_w18660_,
		_w18657_,
		_w19011_
	);
	LUT3 #(
		.INIT('h0b)
	) name13185 (
		_w18655_,
		_w18663_,
		_w19011_,
		_w19012_
	);
	LUT4 #(
		.INIT('h0100)
	) name13186 (
		_w19007_,
		_w19008_,
		_w19010_,
		_w19012_,
		_w19013_
	);
	LUT3 #(
		.INIT('h65)
	) name13187 (
		\u1_L8_reg[27]/NET0131 ,
		_w19004_,
		_w19013_,
		_w19014_
	);
	LUT4 #(
		.INIT('h8048)
	) name13188 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w19015_
	);
	LUT4 #(
		.INIT('hcfaf)
	) name13189 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w19016_
	);
	LUT2 #(
		.INIT('h2)
	) name13190 (
		_w18567_,
		_w19016_,
		_w19017_
	);
	LUT3 #(
		.INIT('h51)
	) name13191 (
		_w18576_,
		_w18713_,
		_w18716_,
		_w19018_
	);
	LUT4 #(
		.INIT('h5455)
	) name13192 (
		_w18566_,
		_w19015_,
		_w19017_,
		_w19018_,
		_w19019_
	);
	LUT4 #(
		.INIT('h1001)
	) name13193 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w19020_
	);
	LUT4 #(
		.INIT('hcee2)
	) name13194 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w19021_
	);
	LUT3 #(
		.INIT('h01)
	) name13195 (
		_w18567_,
		_w19021_,
		_w19020_,
		_w19022_
	);
	LUT4 #(
		.INIT('hbbfc)
	) name13196 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w19023_
	);
	LUT3 #(
		.INIT('h08)
	) name13197 (
		_w18570_,
		_w18568_,
		_w18572_,
		_w19024_
	);
	LUT4 #(
		.INIT('h11f5)
	) name13198 (
		_w18567_,
		_w18571_,
		_w19023_,
		_w19024_,
		_w19025_
	);
	LUT4 #(
		.INIT('h4151)
	) name13199 (
		_w18567_,
		_w18570_,
		_w18568_,
		_w18572_,
		_w19026_
	);
	LUT4 #(
		.INIT('h00e4)
	) name13200 (
		_w18567_,
		_w18571_,
		_w18576_,
		_w19026_,
		_w19027_
	);
	LUT4 #(
		.INIT('h0075)
	) name13201 (
		_w18566_,
		_w19022_,
		_w19025_,
		_w19027_,
		_w19028_
	);
	LUT3 #(
		.INIT('h65)
	) name13202 (
		\u1_L8_reg[32]/NET0131 ,
		_w19019_,
		_w19028_,
		_w19029_
	);
	LUT4 #(
		.INIT('hc693)
	) name13203 (
		decrypt_pad,
		\u1_R8_reg[11]/NET0131 ,
		\u1_uk_K_r8_reg[32]/NET0131 ,
		\u1_uk_K_r8_reg[54]/NET0131 ,
		_w19030_
	);
	LUT4 #(
		.INIT('hc963)
	) name13204 (
		decrypt_pad,
		\u1_R8_reg[13]/NET0131 ,
		\u1_uk_K_r8_reg[25]/NET0131 ,
		\u1_uk_K_r8_reg[3]/NET0131 ,
		_w19031_
	);
	LUT4 #(
		.INIT('hc963)
	) name13205 (
		decrypt_pad,
		\u1_R8_reg[9]/NET0131 ,
		\u1_uk_K_r8_reg[20]/NET0131 ,
		\u1_uk_K_r8_reg[55]/NET0131 ,
		_w19032_
	);
	LUT4 #(
		.INIT('hc963)
	) name13206 (
		decrypt_pad,
		\u1_R8_reg[10]/NET0131 ,
		\u1_uk_K_r8_reg[53]/NET0131 ,
		\u1_uk_K_r8_reg[6]/NET0131 ,
		_w19033_
	);
	LUT4 #(
		.INIT('hc693)
	) name13207 (
		decrypt_pad,
		\u1_R8_reg[8]/NET0131 ,
		\u1_uk_K_r8_reg[26]/NET0131 ,
		\u1_uk_K_r8_reg[48]/NET0131 ,
		_w19034_
	);
	LUT2 #(
		.INIT('h2)
	) name13208 (
		_w19031_,
		_w19034_,
		_w19035_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name13209 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19036_
	);
	LUT4 #(
		.INIT('h9b55)
	) name13210 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19037_
	);
	LUT4 #(
		.INIT('hc963)
	) name13211 (
		decrypt_pad,
		\u1_R8_reg[12]/NET0131 ,
		\u1_uk_K_r8_reg[12]/NET0131 ,
		\u1_uk_K_r8_reg[47]/NET0131 ,
		_w19038_
	);
	LUT4 #(
		.INIT('h0001)
	) name13212 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19039_
	);
	LUT4 #(
		.INIT('hff5e)
	) name13213 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19040_
	);
	LUT4 #(
		.INIT('h20aa)
	) name13214 (
		_w19030_,
		_w19037_,
		_w19038_,
		_w19040_,
		_w19041_
	);
	LUT3 #(
		.INIT('h45)
	) name13215 (
		_w19030_,
		_w19031_,
		_w19032_,
		_w19042_
	);
	LUT4 #(
		.INIT('h30bb)
	) name13216 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19043_
	);
	LUT4 #(
		.INIT('h1000)
	) name13217 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19044_
	);
	LUT4 #(
		.INIT('h00a2)
	) name13218 (
		_w19038_,
		_w19042_,
		_w19043_,
		_w19044_,
		_w19045_
	);
	LUT2 #(
		.INIT('h4)
	) name13219 (
		_w19031_,
		_w19034_,
		_w19046_
	);
	LUT4 #(
		.INIT('hffcb)
	) name13220 (
		_w19030_,
		_w19031_,
		_w19034_,
		_w19032_,
		_w19047_
	);
	LUT2 #(
		.INIT('h1)
	) name13221 (
		_w19033_,
		_w19047_,
		_w19048_
	);
	LUT4 #(
		.INIT('h2000)
	) name13222 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19049_
	);
	LUT2 #(
		.INIT('h4)
	) name13223 (
		_w19030_,
		_w19049_,
		_w19050_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name13224 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19051_
	);
	LUT4 #(
		.INIT('h0990)
	) name13225 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19052_
	);
	LUT4 #(
		.INIT('h4000)
	) name13226 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19053_
	);
	LUT4 #(
		.INIT('h0200)
	) name13227 (
		_w19030_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19054_
	);
	LUT4 #(
		.INIT('h0001)
	) name13228 (
		_w19038_,
		_w19053_,
		_w19052_,
		_w19054_,
		_w19055_
	);
	LUT4 #(
		.INIT('h5455)
	) name13229 (
		_w19045_,
		_w19050_,
		_w19048_,
		_w19055_,
		_w19056_
	);
	LUT3 #(
		.INIT('h56)
	) name13230 (
		\u1_L8_reg[6]/NET0131 ,
		_w19041_,
		_w19056_,
		_w19057_
	);
	LUT4 #(
		.INIT('hf7f6)
	) name13231 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w19058_
	);
	LUT3 #(
		.INIT('h02)
	) name13232 (
		_w18730_,
		_w18731_,
		_w18727_,
		_w19059_
	);
	LUT4 #(
		.INIT('h00c4)
	) name13233 (
		_w18727_,
		_w18754_,
		_w19058_,
		_w19059_,
		_w19060_
	);
	LUT2 #(
		.INIT('h2)
	) name13234 (
		_w18738_,
		_w19060_,
		_w19061_
	);
	LUT4 #(
		.INIT('h4044)
	) name13235 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w19062_
	);
	LUT4 #(
		.INIT('h0002)
	) name13236 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w19063_
	);
	LUT4 #(
		.INIT('hfe54)
	) name13237 (
		_w18727_,
		_w18832_,
		_w19062_,
		_w19063_,
		_w19064_
	);
	LUT4 #(
		.INIT('h8000)
	) name13238 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18727_,
		_w19065_
	);
	LUT3 #(
		.INIT('h04)
	) name13239 (
		_w18734_,
		_w18850_,
		_w19065_,
		_w19066_
	);
	LUT3 #(
		.INIT('h45)
	) name13240 (
		_w18738_,
		_w19064_,
		_w19066_,
		_w19067_
	);
	LUT2 #(
		.INIT('h1)
	) name13241 (
		_w18727_,
		_w18744_,
		_w19068_
	);
	LUT2 #(
		.INIT('h9)
	) name13242 (
		_w18729_,
		_w18731_,
		_w19069_
	);
	LUT3 #(
		.INIT('hb0)
	) name13243 (
		_w18730_,
		_w18728_,
		_w18727_,
		_w19070_
	);
	LUT3 #(
		.INIT('h54)
	) name13244 (
		_w18837_,
		_w19069_,
		_w19070_,
		_w19071_
	);
	LUT2 #(
		.INIT('h1)
	) name13245 (
		_w19068_,
		_w19071_,
		_w19072_
	);
	LUT4 #(
		.INIT('h5556)
	) name13246 (
		\u1_L8_reg[8]/NET0131 ,
		_w19067_,
		_w19072_,
		_w19061_,
		_w19073_
	);
	LUT2 #(
		.INIT('h2)
	) name13247 (
		_w18567_,
		_w18566_,
		_w19074_
	);
	LUT4 #(
		.INIT('h877a)
	) name13248 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w19075_
	);
	LUT2 #(
		.INIT('h2)
	) name13249 (
		_w19074_,
		_w19075_,
		_w19076_
	);
	LUT4 #(
		.INIT('h5004)
	) name13250 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w19077_
	);
	LUT4 #(
		.INIT('hd77f)
	) name13251 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w19078_
	);
	LUT2 #(
		.INIT('h4)
	) name13252 (
		_w18567_,
		_w18566_,
		_w19079_
	);
	LUT2 #(
		.INIT('h9)
	) name13253 (
		_w18567_,
		_w18566_,
		_w19080_
	);
	LUT3 #(
		.INIT('h20)
	) name13254 (
		_w19078_,
		_w19077_,
		_w19080_,
		_w19081_
	);
	LUT3 #(
		.INIT('h09)
	) name13255 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w19082_
	);
	LUT4 #(
		.INIT('h0ce0)
	) name13256 (
		_w18570_,
		_w18571_,
		_w18568_,
		_w18572_,
		_w19083_
	);
	LUT4 #(
		.INIT('h0008)
	) name13257 (
		_w19078_,
		_w19079_,
		_w19083_,
		_w19082_,
		_w19084_
	);
	LUT4 #(
		.INIT('h00ab)
	) name13258 (
		_w18580_,
		_w19076_,
		_w19081_,
		_w19084_,
		_w19085_
	);
	LUT2 #(
		.INIT('h6)
	) name13259 (
		\u1_L8_reg[7]/NET0131 ,
		_w19085_,
		_w19086_
	);
	LUT3 #(
		.INIT('h02)
	) name13260 (
		_w19030_,
		_w19033_,
		_w19032_,
		_w19087_
	);
	LUT4 #(
		.INIT('h3310)
	) name13261 (
		_w19030_,
		_w19035_,
		_w19051_,
		_w19087_,
		_w19088_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name13262 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19089_
	);
	LUT3 #(
		.INIT('hc4)
	) name13263 (
		_w19030_,
		_w19038_,
		_w19089_,
		_w19090_
	);
	LUT3 #(
		.INIT('h10)
	) name13264 (
		_w19048_,
		_w19088_,
		_w19090_,
		_w19091_
	);
	LUT4 #(
		.INIT('ha8a2)
	) name13265 (
		_w19030_,
		_w19031_,
		_w19034_,
		_w19033_,
		_w19092_
	);
	LUT3 #(
		.INIT('h10)
	) name13266 (
		_w19031_,
		_w19034_,
		_w19032_,
		_w19093_
	);
	LUT4 #(
		.INIT('hee3f)
	) name13267 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19094_
	);
	LUT2 #(
		.INIT('h8)
	) name13268 (
		_w19092_,
		_w19094_,
		_w19095_
	);
	LUT4 #(
		.INIT('h0009)
	) name13269 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19096_
	);
	LUT3 #(
		.INIT('h04)
	) name13270 (
		_w19030_,
		_w19036_,
		_w19096_,
		_w19097_
	);
	LUT4 #(
		.INIT('h0040)
	) name13271 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19098_
	);
	LUT2 #(
		.INIT('h1)
	) name13272 (
		_w19038_,
		_w19098_,
		_w19099_
	);
	LUT3 #(
		.INIT('he0)
	) name13273 (
		_w19095_,
		_w19097_,
		_w19099_,
		_w19100_
	);
	LUT2 #(
		.INIT('h4)
	) name13274 (
		_w19030_,
		_w19033_,
		_w19101_
	);
	LUT2 #(
		.INIT('h8)
	) name13275 (
		_w19031_,
		_w19034_,
		_w19102_
	);
	LUT3 #(
		.INIT('h80)
	) name13276 (
		_w19031_,
		_w19034_,
		_w19032_,
		_w19103_
	);
	LUT2 #(
		.INIT('h8)
	) name13277 (
		_w19101_,
		_w19103_,
		_w19104_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name13278 (
		_w19031_,
		_w19034_,
		_w19054_,
		_w19087_,
		_w19105_
	);
	LUT2 #(
		.INIT('h4)
	) name13279 (
		_w19104_,
		_w19105_,
		_w19106_
	);
	LUT4 #(
		.INIT('ha955)
	) name13280 (
		\u1_L8_reg[24]/NET0131 ,
		_w19091_,
		_w19100_,
		_w19106_,
		_w19107_
	);
	LUT3 #(
		.INIT('h15)
	) name13281 (
		_w19030_,
		_w19034_,
		_w19033_,
		_w19108_
	);
	LUT3 #(
		.INIT('h23)
	) name13282 (
		_w19093_,
		_w19092_,
		_w19108_,
		_w19109_
	);
	LUT4 #(
		.INIT('h7000)
	) name13283 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19110_
	);
	LUT4 #(
		.INIT('h002a)
	) name13284 (
		_w19038_,
		_w19046_,
		_w19087_,
		_w19110_,
		_w19111_
	);
	LUT2 #(
		.INIT('h4)
	) name13285 (
		_w19109_,
		_w19111_,
		_w19112_
	);
	LUT4 #(
		.INIT('h7a3f)
	) name13286 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19113_
	);
	LUT2 #(
		.INIT('h2)
	) name13287 (
		_w19030_,
		_w19113_,
		_w19114_
	);
	LUT3 #(
		.INIT('h72)
	) name13288 (
		_w19034_,
		_w19033_,
		_w19032_,
		_w19115_
	);
	LUT2 #(
		.INIT('h8)
	) name13289 (
		_w19042_,
		_w19115_,
		_w19116_
	);
	LUT4 #(
		.INIT('h0020)
	) name13290 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w19117_
	);
	LUT3 #(
		.INIT('h01)
	) name13291 (
		_w19038_,
		_w19096_,
		_w19117_,
		_w19118_
	);
	LUT3 #(
		.INIT('h10)
	) name13292 (
		_w19114_,
		_w19116_,
		_w19118_,
		_w19119_
	);
	LUT3 #(
		.INIT('h08)
	) name13293 (
		_w19030_,
		_w19033_,
		_w19032_,
		_w19120_
	);
	LUT4 #(
		.INIT('h1000)
	) name13294 (
		_w19030_,
		_w19031_,
		_w19033_,
		_w19032_,
		_w19121_
	);
	LUT3 #(
		.INIT('h07)
	) name13295 (
		_w19102_,
		_w19120_,
		_w19121_,
		_w19122_
	);
	LUT4 #(
		.INIT('h56aa)
	) name13296 (
		\u1_L8_reg[30]/NET0131 ,
		_w19112_,
		_w19119_,
		_w19122_,
		_w19123_
	);
	LUT4 #(
		.INIT('h0002)
	) name13297 (
		_w18738_,
		_w18744_,
		_w18853_,
		_w18846_,
		_w19124_
	);
	LUT4 #(
		.INIT('h0d00)
	) name13298 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w19125_
	);
	LUT4 #(
		.INIT('h22e6)
	) name13299 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w19126_
	);
	LUT3 #(
		.INIT('h10)
	) name13300 (
		_w18738_,
		_w19125_,
		_w19126_,
		_w19127_
	);
	LUT4 #(
		.INIT('hf7fe)
	) name13301 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w19128_
	);
	LUT3 #(
		.INIT('h10)
	) name13302 (
		_w18727_,
		_w18751_,
		_w19128_,
		_w19129_
	);
	LUT3 #(
		.INIT('he0)
	) name13303 (
		_w19124_,
		_w19127_,
		_w19129_,
		_w19130_
	);
	LUT4 #(
		.INIT('h1098)
	) name13304 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w19131_
	);
	LUT4 #(
		.INIT('h0002)
	) name13305 (
		_w18738_,
		_w18744_,
		_w18853_,
		_w19131_,
		_w19132_
	);
	LUT4 #(
		.INIT('h2064)
	) name13306 (
		_w18730_,
		_w18728_,
		_w18729_,
		_w18731_,
		_w19133_
	);
	LUT3 #(
		.INIT('h01)
	) name13307 (
		_w18738_,
		_w19125_,
		_w19133_,
		_w19134_
	);
	LUT3 #(
		.INIT('h02)
	) name13308 (
		_w18727_,
		_w18753_,
		_w19063_,
		_w19135_
	);
	LUT3 #(
		.INIT('he0)
	) name13309 (
		_w19132_,
		_w19134_,
		_w19135_,
		_w19136_
	);
	LUT3 #(
		.INIT('ha9)
	) name13310 (
		\u1_L8_reg[3]/NET0131 ,
		_w19130_,
		_w19136_,
		_w19137_
	);
	LUT4 #(
		.INIT('h9600)
	) name13311 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w19138_
	);
	LUT3 #(
		.INIT('h19)
	) name13312 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w19139_
	);
	LUT2 #(
		.INIT('h2)
	) name13313 (
		_w18794_,
		_w18790_,
		_w19140_
	);
	LUT4 #(
		.INIT('h0015)
	) name13314 (
		_w18807_,
		_w19139_,
		_w19140_,
		_w19138_,
		_w19141_
	);
	LUT2 #(
		.INIT('h2)
	) name13315 (
		_w18800_,
		_w19141_,
		_w19142_
	);
	LUT4 #(
		.INIT('h0019)
	) name13316 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18794_,
		_w19143_
	);
	LUT3 #(
		.INIT('h08)
	) name13317 (
		_w18791_,
		_w18792_,
		_w18790_,
		_w19144_
	);
	LUT4 #(
		.INIT('h0080)
	) name13318 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w19145_
	);
	LUT2 #(
		.INIT('h1)
	) name13319 (
		_w19143_,
		_w19145_,
		_w19146_
	);
	LUT4 #(
		.INIT('h4100)
	) name13320 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w19147_
	);
	LUT3 #(
		.INIT('h60)
	) name13321 (
		_w18791_,
		_w18789_,
		_w18794_,
		_w19148_
	);
	LUT3 #(
		.INIT('h45)
	) name13322 (
		_w19147_,
		_w19144_,
		_w19148_,
		_w19149_
	);
	LUT4 #(
		.INIT('hf77f)
	) name13323 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w19150_
	);
	LUT2 #(
		.INIT('h1)
	) name13324 (
		_w18794_,
		_w19150_,
		_w19151_
	);
	LUT4 #(
		.INIT('h00ea)
	) name13325 (
		_w18800_,
		_w19146_,
		_w19149_,
		_w19151_,
		_w19152_
	);
	LUT3 #(
		.INIT('h65)
	) name13326 (
		\u1_L8_reg[9]/NET0131 ,
		_w19142_,
		_w19152_,
		_w19153_
	);
	LUT4 #(
		.INIT('h0a20)
	) name13327 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18887_,
		_w19154_
	);
	LUT4 #(
		.INIT('hfd75)
	) name13328 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w19155_
	);
	LUT4 #(
		.INIT('h0032)
	) name13329 (
		_w18886_,
		_w18910_,
		_w19155_,
		_w19154_,
		_w19156_
	);
	LUT4 #(
		.INIT('h8000)
	) name13330 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18887_,
		_w19157_
	);
	LUT4 #(
		.INIT('hdffc)
	) name13331 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w19158_
	);
	LUT4 #(
		.INIT('h1003)
	) name13332 (
		_w18886_,
		_w18888_,
		_w18887_,
		_w18890_,
		_w19159_
	);
	LUT4 #(
		.INIT('h0100)
	) name13333 (
		_w18895_,
		_w19157_,
		_w19159_,
		_w19158_,
		_w19160_
	);
	LUT4 #(
		.INIT('h1000)
	) name13334 (
		_w18886_,
		_w18888_,
		_w18889_,
		_w18887_,
		_w19161_
	);
	LUT4 #(
		.INIT('h77ef)
	) name13335 (
		_w18888_,
		_w18889_,
		_w18887_,
		_w18890_,
		_w19162_
	);
	LUT3 #(
		.INIT('h31)
	) name13336 (
		_w18886_,
		_w19161_,
		_w19162_,
		_w19163_
	);
	LUT4 #(
		.INIT('hd800)
	) name13337 (
		_w18885_,
		_w19156_,
		_w19160_,
		_w19163_,
		_w19164_
	);
	LUT2 #(
		.INIT('h9)
	) name13338 (
		\u1_L8_reg[18]/NET0131 ,
		_w19164_,
		_w19165_
	);
	LUT4 #(
		.INIT('hc963)
	) name13339 (
		decrypt_pad,
		\u1_R7_reg[4]/NET0131 ,
		\u1_uk_K_r7_reg[47]/NET0131 ,
		\u1_uk_K_r7_reg[54]/NET0131 ,
		_w19166_
	);
	LUT4 #(
		.INIT('hc963)
	) name13340 (
		decrypt_pad,
		\u1_R7_reg[32]/NET0131 ,
		\u1_uk_K_r7_reg[24]/NET0131 ,
		\u1_uk_K_r7_reg[6]/NET0131 ,
		_w19167_
	);
	LUT4 #(
		.INIT('hc963)
	) name13341 (
		decrypt_pad,
		\u1_R7_reg[5]/NET0131 ,
		\u1_uk_K_r7_reg[18]/NET0131 ,
		\u1_uk_K_r7_reg[25]/NET0131 ,
		_w19168_
	);
	LUT4 #(
		.INIT('hc963)
	) name13342 (
		decrypt_pad,
		\u1_R7_reg[1]/NET0131 ,
		\u1_uk_K_r7_reg[20]/NET0131 ,
		\u1_uk_K_r7_reg[27]/NET0131 ,
		_w19169_
	);
	LUT4 #(
		.INIT('hc963)
	) name13343 (
		decrypt_pad,
		\u1_R7_reg[3]/NET0131 ,
		\u1_uk_K_r7_reg[12]/NET0131 ,
		\u1_uk_K_r7_reg[19]/NET0131 ,
		_w19170_
	);
	LUT2 #(
		.INIT('h4)
	) name13344 (
		_w19170_,
		_w19169_,
		_w19171_
	);
	LUT4 #(
		.INIT('hc693)
	) name13345 (
		decrypt_pad,
		\u1_R7_reg[2]/NET0131 ,
		\u1_uk_K_r7_reg[10]/NET0131 ,
		\u1_uk_K_r7_reg[3]/NET0131 ,
		_w19172_
	);
	LUT4 #(
		.INIT('hb705)
	) name13346 (
		_w19172_,
		_w19170_,
		_w19168_,
		_w19169_,
		_w19173_
	);
	LUT3 #(
		.INIT('h08)
	) name13347 (
		_w19170_,
		_w19168_,
		_w19169_,
		_w19174_
	);
	LUT2 #(
		.INIT('h1)
	) name13348 (
		_w19168_,
		_w19169_,
		_w19175_
	);
	LUT4 #(
		.INIT('hccfa)
	) name13349 (
		_w19172_,
		_w19170_,
		_w19168_,
		_w19169_,
		_w19176_
	);
	LUT4 #(
		.INIT('h3120)
	) name13350 (
		_w19167_,
		_w19174_,
		_w19176_,
		_w19173_,
		_w19177_
	);
	LUT2 #(
		.INIT('h2)
	) name13351 (
		_w19166_,
		_w19177_,
		_w19178_
	);
	LUT3 #(
		.INIT('h40)
	) name13352 (
		_w19167_,
		_w19172_,
		_w19170_,
		_w19179_
	);
	LUT4 #(
		.INIT('h4000)
	) name13353 (
		_w19167_,
		_w19172_,
		_w19170_,
		_w19168_,
		_w19180_
	);
	LUT4 #(
		.INIT('hbfee)
	) name13354 (
		_w19167_,
		_w19172_,
		_w19170_,
		_w19168_,
		_w19181_
	);
	LUT2 #(
		.INIT('h4)
	) name13355 (
		_w19181_,
		_w19169_,
		_w19182_
	);
	LUT4 #(
		.INIT('h0020)
	) name13356 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19183_
	);
	LUT4 #(
		.INIT('h0800)
	) name13357 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19184_
	);
	LUT4 #(
		.INIT('hd7df)
	) name13358 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19185_
	);
	LUT3 #(
		.INIT('h0e)
	) name13359 (
		_w19170_,
		_w19183_,
		_w19185_,
		_w19186_
	);
	LUT3 #(
		.INIT('h0e)
	) name13360 (
		_w19182_,
		_w19186_,
		_w19166_,
		_w19187_
	);
	LUT4 #(
		.INIT('h0040)
	) name13361 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19188_
	);
	LUT4 #(
		.INIT('h7cbf)
	) name13362 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19189_
	);
	LUT2 #(
		.INIT('h1)
	) name13363 (
		_w19170_,
		_w19189_,
		_w19190_
	);
	LUT3 #(
		.INIT('h13)
	) name13364 (
		_w19167_,
		_w19170_,
		_w19169_,
		_w19191_
	);
	LUT2 #(
		.INIT('h9)
	) name13365 (
		_w19167_,
		_w19172_,
		_w19192_
	);
	LUT3 #(
		.INIT('h0d)
	) name13366 (
		_w19168_,
		_w19169_,
		_w19166_,
		_w19193_
	);
	LUT3 #(
		.INIT('h80)
	) name13367 (
		_w19192_,
		_w19191_,
		_w19193_,
		_w19194_
	);
	LUT2 #(
		.INIT('h4)
	) name13368 (
		_w19172_,
		_w19170_,
		_w19195_
	);
	LUT4 #(
		.INIT('h0020)
	) name13369 (
		_w19167_,
		_w19172_,
		_w19170_,
		_w19169_,
		_w19196_
	);
	LUT3 #(
		.INIT('h07)
	) name13370 (
		_w19179_,
		_w19175_,
		_w19196_,
		_w19197_
	);
	LUT3 #(
		.INIT('h10)
	) name13371 (
		_w19190_,
		_w19194_,
		_w19197_,
		_w19198_
	);
	LUT4 #(
		.INIT('h5655)
	) name13372 (
		\u1_L7_reg[31]/NET0131 ,
		_w19187_,
		_w19178_,
		_w19198_,
		_w19199_
	);
	LUT4 #(
		.INIT('hc963)
	) name13373 (
		decrypt_pad,
		\u1_R7_reg[24]/NET0131 ,
		\u1_uk_K_r7_reg[16]/NET0131 ,
		\u1_uk_K_r7_reg[23]/P0001 ,
		_w19200_
	);
	LUT4 #(
		.INIT('hc963)
	) name13374 (
		decrypt_pad,
		\u1_R7_reg[22]/NET0131 ,
		\u1_uk_K_r7_reg[1]/NET0131 ,
		\u1_uk_K_r7_reg[8]/NET0131 ,
		_w19201_
	);
	LUT4 #(
		.INIT('hc693)
	) name13375 (
		decrypt_pad,
		\u1_R7_reg[20]/NET0131 ,
		\u1_uk_K_r7_reg[2]/NET0131 ,
		\u1_uk_K_r7_reg[50]/NET0131 ,
		_w19202_
	);
	LUT4 #(
		.INIT('hc963)
	) name13376 (
		decrypt_pad,
		\u1_R7_reg[21]/NET0131 ,
		\u1_uk_K_r7_reg[38]/NET0131 ,
		\u1_uk_K_r7_reg[45]/NET0131 ,
		_w19203_
	);
	LUT4 #(
		.INIT('hc963)
	) name13377 (
		decrypt_pad,
		\u1_R7_reg[25]/NET0131 ,
		\u1_uk_K_r7_reg[35]/NET0131 ,
		\u1_uk_K_r7_reg[42]/NET0131 ,
		_w19204_
	);
	LUT4 #(
		.INIT('ha280)
	) name13378 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19205_
	);
	LUT4 #(
		.INIT('hc963)
	) name13379 (
		decrypt_pad,
		\u1_R7_reg[23]/NET0131 ,
		\u1_uk_K_r7_reg[14]/NET0131 ,
		\u1_uk_K_r7_reg[21]/NET0131 ,
		_w19206_
	);
	LUT4 #(
		.INIT('h4555)
	) name13380 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19207_
	);
	LUT3 #(
		.INIT('h01)
	) name13381 (
		_w19206_,
		_w19207_,
		_w19205_,
		_w19208_
	);
	LUT4 #(
		.INIT('h0004)
	) name13382 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19209_
	);
	LUT4 #(
		.INIT('h1dfb)
	) name13383 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19210_
	);
	LUT2 #(
		.INIT('h1)
	) name13384 (
		_w19201_,
		_w19206_,
		_w19211_
	);
	LUT4 #(
		.INIT('h1000)
	) name13385 (
		_w19201_,
		_w19206_,
		_w19202_,
		_w19204_,
		_w19212_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13386 (
		_w19206_,
		_w19203_,
		_w19210_,
		_w19212_,
		_w19213_
	);
	LUT3 #(
		.INIT('h8a)
	) name13387 (
		_w19200_,
		_w19208_,
		_w19213_,
		_w19214_
	);
	LUT3 #(
		.INIT('h8a)
	) name13388 (
		_w19202_,
		_w19204_,
		_w19203_,
		_w19215_
	);
	LUT3 #(
		.INIT('h54)
	) name13389 (
		_w19201_,
		_w19206_,
		_w19202_,
		_w19216_
	);
	LUT4 #(
		.INIT('h0020)
	) name13390 (
		_w19206_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19217_
	);
	LUT2 #(
		.INIT('h8)
	) name13391 (
		_w19201_,
		_w19206_,
		_w19218_
	);
	LUT4 #(
		.INIT('h0080)
	) name13392 (
		_w19201_,
		_w19206_,
		_w19202_,
		_w19203_,
		_w19219_
	);
	LUT4 #(
		.INIT('h1011)
	) name13393 (
		_w19217_,
		_w19219_,
		_w19215_,
		_w19216_,
		_w19220_
	);
	LUT4 #(
		.INIT('h0080)
	) name13394 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19221_
	);
	LUT4 #(
		.INIT('h0010)
	) name13395 (
		_w19201_,
		_w19206_,
		_w19202_,
		_w19204_,
		_w19222_
	);
	LUT4 #(
		.INIT('h1200)
	) name13396 (
		_w19201_,
		_w19206_,
		_w19202_,
		_w19203_,
		_w19223_
	);
	LUT3 #(
		.INIT('h01)
	) name13397 (
		_w19221_,
		_w19222_,
		_w19223_,
		_w19224_
	);
	LUT3 #(
		.INIT('h15)
	) name13398 (
		_w19200_,
		_w19220_,
		_w19224_,
		_w19225_
	);
	LUT4 #(
		.INIT('hfbdf)
	) name13399 (
		_w19206_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19226_
	);
	LUT2 #(
		.INIT('h1)
	) name13400 (
		_w19201_,
		_w19226_,
		_w19227_
	);
	LUT3 #(
		.INIT('h01)
	) name13401 (
		_w19202_,
		_w19204_,
		_w19203_,
		_w19228_
	);
	LUT4 #(
		.INIT('h7e7f)
	) name13402 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19229_
	);
	LUT4 #(
		.INIT('hef23)
	) name13403 (
		_w19201_,
		_w19206_,
		_w19228_,
		_w19229_,
		_w19230_
	);
	LUT2 #(
		.INIT('h4)
	) name13404 (
		_w19227_,
		_w19230_,
		_w19231_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name13405 (
		\u1_L7_reg[11]/NET0131 ,
		_w19214_,
		_w19225_,
		_w19231_,
		_w19232_
	);
	LUT4 #(
		.INIT('hc963)
	) name13406 (
		decrypt_pad,
		\u1_R7_reg[28]/NET0131 ,
		\u1_uk_K_r7_reg[23]/P0001 ,
		\u1_uk_K_r7_reg[30]/P0001 ,
		_w19233_
	);
	LUT4 #(
		.INIT('hc963)
	) name13407 (
		decrypt_pad,
		\u1_R7_reg[26]/NET0131 ,
		\u1_uk_K_r7_reg[31]/NET0131 ,
		\u1_uk_K_r7_reg[38]/NET0131 ,
		_w19234_
	);
	LUT4 #(
		.INIT('hc963)
	) name13408 (
		decrypt_pad,
		\u1_R7_reg[25]/NET0131 ,
		\u1_uk_K_r7_reg[42]/NET0131 ,
		\u1_uk_K_r7_reg[49]/NET0131 ,
		_w19235_
	);
	LUT4 #(
		.INIT('hc963)
	) name13409 (
		decrypt_pad,
		\u1_R7_reg[29]/NET0131 ,
		\u1_uk_K_r7_reg[15]/NET0131 ,
		\u1_uk_K_r7_reg[22]/NET0131 ,
		_w19236_
	);
	LUT3 #(
		.INIT('hea)
	) name13410 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19237_
	);
	LUT4 #(
		.INIT('hc693)
	) name13411 (
		decrypt_pad,
		\u1_R7_reg[24]/NET0131 ,
		\u1_uk_K_r7_reg[14]/NET0131 ,
		\u1_uk_K_r7_reg[7]/NET0131 ,
		_w19238_
	);
	LUT4 #(
		.INIT('hc963)
	) name13412 (
		decrypt_pad,
		\u1_R7_reg[27]/NET0131 ,
		\u1_uk_K_r7_reg[36]/NET0131 ,
		\u1_uk_K_r7_reg[43]/NET0131 ,
		_w19239_
	);
	LUT3 #(
		.INIT('h70)
	) name13413 (
		_w19234_,
		_w19235_,
		_w19239_,
		_w19240_
	);
	LUT4 #(
		.INIT('h7000)
	) name13414 (
		_w19234_,
		_w19235_,
		_w19238_,
		_w19239_,
		_w19241_
	);
	LUT2 #(
		.INIT('h8)
	) name13415 (
		_w19237_,
		_w19241_,
		_w19242_
	);
	LUT4 #(
		.INIT('h1000)
	) name13416 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19243_
	);
	LUT4 #(
		.INIT('hef3f)
	) name13417 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19244_
	);
	LUT2 #(
		.INIT('h2)
	) name13418 (
		_w19236_,
		_w19238_,
		_w19245_
	);
	LUT4 #(
		.INIT('h0020)
	) name13419 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19246_
	);
	LUT4 #(
		.INIT('hffde)
	) name13420 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19247_
	);
	LUT3 #(
		.INIT('he0)
	) name13421 (
		_w19239_,
		_w19244_,
		_w19247_,
		_w19248_
	);
	LUT3 #(
		.INIT('h8a)
	) name13422 (
		_w19233_,
		_w19242_,
		_w19248_,
		_w19249_
	);
	LUT4 #(
		.INIT('h0072)
	) name13423 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19239_,
		_w19250_
	);
	LUT4 #(
		.INIT('h10f0)
	) name13424 (
		_w19234_,
		_w19235_,
		_w19238_,
		_w19239_,
		_w19251_
	);
	LUT2 #(
		.INIT('h4)
	) name13425 (
		_w19250_,
		_w19251_,
		_w19252_
	);
	LUT4 #(
		.INIT('h0002)
	) name13426 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19253_
	);
	LUT2 #(
		.INIT('h6)
	) name13427 (
		_w19234_,
		_w19238_,
		_w19254_
	);
	LUT3 #(
		.INIT('h8c)
	) name13428 (
		_w19235_,
		_w19236_,
		_w19239_,
		_w19255_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name13429 (
		_w19253_,
		_w19239_,
		_w19254_,
		_w19255_,
		_w19256_
	);
	LUT4 #(
		.INIT('h0008)
	) name13430 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19257_
	);
	LUT4 #(
		.INIT('hfcd7)
	) name13431 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19258_
	);
	LUT4 #(
		.INIT('h0084)
	) name13432 (
		_w19234_,
		_w19235_,
		_w19238_,
		_w19239_,
		_w19259_
	);
	LUT4 #(
		.INIT('h0100)
	) name13433 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19239_,
		_w19260_
	);
	LUT4 #(
		.INIT('h0031)
	) name13434 (
		_w19239_,
		_w19259_,
		_w19258_,
		_w19260_,
		_w19261_
	);
	LUT4 #(
		.INIT('hba00)
	) name13435 (
		_w19233_,
		_w19252_,
		_w19256_,
		_w19261_,
		_w19262_
	);
	LUT3 #(
		.INIT('h65)
	) name13436 (
		\u1_L7_reg[22]/NET0131 ,
		_w19249_,
		_w19262_,
		_w19263_
	);
	LUT4 #(
		.INIT('haa9b)
	) name13437 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19264_
	);
	LUT2 #(
		.INIT('h2)
	) name13438 (
		_w19170_,
		_w19264_,
		_w19265_
	);
	LUT4 #(
		.INIT('h0200)
	) name13439 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19266_
	);
	LUT4 #(
		.INIT('h0809)
	) name13440 (
		_w19167_,
		_w19172_,
		_w19170_,
		_w19169_,
		_w19267_
	);
	LUT3 #(
		.INIT('h80)
	) name13441 (
		_w19172_,
		_w19168_,
		_w19169_,
		_w19268_
	);
	LUT4 #(
		.INIT('h0002)
	) name13442 (
		_w19166_,
		_w19266_,
		_w19267_,
		_w19268_,
		_w19269_
	);
	LUT2 #(
		.INIT('h4)
	) name13443 (
		_w19265_,
		_w19269_,
		_w19270_
	);
	LUT3 #(
		.INIT('h09)
	) name13444 (
		_w19167_,
		_w19168_,
		_w19169_,
		_w19271_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name13445 (
		_w19167_,
		_w19172_,
		_w19170_,
		_w19168_,
		_w19272_
	);
	LUT2 #(
		.INIT('h4)
	) name13446 (
		_w19271_,
		_w19272_,
		_w19273_
	);
	LUT2 #(
		.INIT('h6)
	) name13447 (
		_w19168_,
		_w19169_,
		_w19274_
	);
	LUT3 #(
		.INIT('h82)
	) name13448 (
		_w19167_,
		_w19168_,
		_w19169_,
		_w19275_
	);
	LUT4 #(
		.INIT('h1400)
	) name13449 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19276_
	);
	LUT3 #(
		.INIT('h02)
	) name13450 (
		_w19170_,
		_w19276_,
		_w19275_,
		_w19277_
	);
	LUT3 #(
		.INIT('h01)
	) name13451 (
		_w19184_,
		_w19166_,
		_w19188_,
		_w19278_
	);
	LUT3 #(
		.INIT('he0)
	) name13452 (
		_w19273_,
		_w19277_,
		_w19278_,
		_w19279_
	);
	LUT3 #(
		.INIT('ha9)
	) name13453 (
		\u1_L7_reg[17]/NET0131 ,
		_w19270_,
		_w19279_,
		_w19280_
	);
	LUT4 #(
		.INIT('hc963)
	) name13454 (
		decrypt_pad,
		\u1_R7_reg[12]/NET0131 ,
		\u1_uk_K_r7_reg[13]/NET0131 ,
		\u1_uk_K_r7_reg[20]/NET0131 ,
		_w19281_
	);
	LUT4 #(
		.INIT('hc963)
	) name13455 (
		decrypt_pad,
		\u1_R7_reg[13]/NET0131 ,
		\u1_uk_K_r7_reg[32]/NET0131 ,
		\u1_uk_K_r7_reg[39]/NET0131 ,
		_w19282_
	);
	LUT4 #(
		.INIT('hc963)
	) name13456 (
		decrypt_pad,
		\u1_R7_reg[15]/NET0131 ,
		\u1_uk_K_r7_reg[41]/NET0131 ,
		\u1_uk_K_r7_reg[48]/NET0131 ,
		_w19283_
	);
	LUT4 #(
		.INIT('hc963)
	) name13457 (
		decrypt_pad,
		\u1_R7_reg[14]/NET0131 ,
		\u1_uk_K_r7_reg[33]/NET0131 ,
		\u1_uk_K_r7_reg[40]/NET0131 ,
		_w19284_
	);
	LUT3 #(
		.INIT('h80)
	) name13458 (
		_w19283_,
		_w19284_,
		_w19282_,
		_w19285_
	);
	LUT4 #(
		.INIT('h2000)
	) name13459 (
		_w19283_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19286_
	);
	LUT4 #(
		.INIT('hc693)
	) name13460 (
		decrypt_pad,
		\u1_R7_reg[17]/NET0131 ,
		\u1_uk_K_r7_reg[4]/NET0131 ,
		\u1_uk_K_r7_reg[54]/NET0131 ,
		_w19287_
	);
	LUT4 #(
		.INIT('h0008)
	) name13461 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19288_
	);
	LUT4 #(
		.INIT('hc963)
	) name13462 (
		decrypt_pad,
		\u1_R7_reg[16]/NET0131 ,
		\u1_uk_K_r7_reg[17]/NET0131 ,
		\u1_uk_K_r7_reg[24]/NET0131 ,
		_w19289_
	);
	LUT3 #(
		.INIT('h01)
	) name13463 (
		_w19288_,
		_w19286_,
		_w19289_,
		_w19290_
	);
	LUT2 #(
		.INIT('h2)
	) name13464 (
		_w19287_,
		_w19281_,
		_w19291_
	);
	LUT4 #(
		.INIT('h8002)
	) name13465 (
		_w19283_,
		_w19287_,
		_w19281_,
		_w19282_,
		_w19292_
	);
	LUT3 #(
		.INIT('h01)
	) name13466 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19293_
	);
	LUT4 #(
		.INIT('h0001)
	) name13467 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19294_
	);
	LUT3 #(
		.INIT('h10)
	) name13468 (
		_w19287_,
		_w19281_,
		_w19282_,
		_w19295_
	);
	LUT4 #(
		.INIT('heffe)
	) name13469 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19296_
	);
	LUT4 #(
		.INIT('hbf15)
	) name13470 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19297_
	);
	LUT4 #(
		.INIT('h00c8)
	) name13471 (
		_w19283_,
		_w19296_,
		_w19297_,
		_w19292_,
		_w19298_
	);
	LUT2 #(
		.INIT('h8)
	) name13472 (
		_w19290_,
		_w19298_,
		_w19299_
	);
	LUT3 #(
		.INIT('h01)
	) name13473 (
		_w19287_,
		_w19281_,
		_w19282_,
		_w19300_
	);
	LUT4 #(
		.INIT('h0001)
	) name13474 (
		_w19283_,
		_w19287_,
		_w19281_,
		_w19282_,
		_w19301_
	);
	LUT2 #(
		.INIT('h8)
	) name13475 (
		_w19284_,
		_w19301_,
		_w19302_
	);
	LUT4 #(
		.INIT('h0104)
	) name13476 (
		_w19283_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19303_
	);
	LUT4 #(
		.INIT('h8000)
	) name13477 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19304_
	);
	LUT3 #(
		.INIT('h02)
	) name13478 (
		_w19289_,
		_w19304_,
		_w19303_,
		_w19305_
	);
	LUT4 #(
		.INIT('h0200)
	) name13479 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19306_
	);
	LUT2 #(
		.INIT('h8)
	) name13480 (
		_w19283_,
		_w19281_,
		_w19307_
	);
	LUT4 #(
		.INIT('h2000)
	) name13481 (
		_w19283_,
		_w19287_,
		_w19281_,
		_w19282_,
		_w19308_
	);
	LUT4 #(
		.INIT('h0008)
	) name13482 (
		_w19283_,
		_w19287_,
		_w19281_,
		_w19282_,
		_w19309_
	);
	LUT3 #(
		.INIT('h01)
	) name13483 (
		_w19306_,
		_w19308_,
		_w19309_,
		_w19310_
	);
	LUT3 #(
		.INIT('h40)
	) name13484 (
		_w19302_,
		_w19305_,
		_w19310_,
		_w19311_
	);
	LUT4 #(
		.INIT('h0040)
	) name13485 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19312_
	);
	LUT4 #(
		.INIT('heee4)
	) name13486 (
		_w19283_,
		_w19306_,
		_w19294_,
		_w19312_,
		_w19313_
	);
	LUT2 #(
		.INIT('h4)
	) name13487 (
		_w19284_,
		_w19308_,
		_w19314_
	);
	LUT2 #(
		.INIT('h1)
	) name13488 (
		_w19313_,
		_w19314_,
		_w19315_
	);
	LUT4 #(
		.INIT('ha955)
	) name13489 (
		\u1_L7_reg[20]/NET0131 ,
		_w19299_,
		_w19311_,
		_w19315_,
		_w19316_
	);
	LUT4 #(
		.INIT('h7d7c)
	) name13490 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19317_
	);
	LUT2 #(
		.INIT('h1)
	) name13491 (
		_w19206_,
		_w19317_,
		_w19318_
	);
	LUT4 #(
		.INIT('hc6ff)
	) name13492 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19319_
	);
	LUT2 #(
		.INIT('h2)
	) name13493 (
		_w19206_,
		_w19319_,
		_w19320_
	);
	LUT4 #(
		.INIT('h0012)
	) name13494 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19321_
	);
	LUT3 #(
		.INIT('h01)
	) name13495 (
		_w19221_,
		_w19222_,
		_w19321_,
		_w19322_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name13496 (
		_w19200_,
		_w19320_,
		_w19318_,
		_w19322_,
		_w19323_
	);
	LUT4 #(
		.INIT('h3df2)
	) name13497 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19324_
	);
	LUT4 #(
		.INIT('ha6bf)
	) name13498 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19325_
	);
	LUT4 #(
		.INIT('h0020)
	) name13499 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19326_
	);
	LUT4 #(
		.INIT('h00d8)
	) name13500 (
		_w19206_,
		_w19324_,
		_w19325_,
		_w19326_,
		_w19327_
	);
	LUT4 #(
		.INIT('h4000)
	) name13501 (
		_w19201_,
		_w19206_,
		_w19204_,
		_w19203_,
		_w19328_
	);
	LUT2 #(
		.INIT('h1)
	) name13502 (
		_w19209_,
		_w19328_,
		_w19329_
	);
	LUT3 #(
		.INIT('he0)
	) name13503 (
		_w19200_,
		_w19327_,
		_w19329_,
		_w19330_
	);
	LUT3 #(
		.INIT('h9a)
	) name13504 (
		\u1_L7_reg[29]/NET0131 ,
		_w19323_,
		_w19330_,
		_w19331_
	);
	LUT4 #(
		.INIT('hc963)
	) name13505 (
		decrypt_pad,
		\u1_R7_reg[8]/NET0131 ,
		\u1_uk_K_r7_reg[48]/NET0131 ,
		\u1_uk_K_r7_reg[55]/P0001 ,
		_w19332_
	);
	LUT4 #(
		.INIT('hc963)
	) name13506 (
		decrypt_pad,
		\u1_R7_reg[7]/NET0131 ,
		\u1_uk_K_r7_reg[25]/NET0131 ,
		\u1_uk_K_r7_reg[32]/NET0131 ,
		_w19333_
	);
	LUT4 #(
		.INIT('hc963)
	) name13507 (
		decrypt_pad,
		\u1_R7_reg[5]/NET0131 ,
		\u1_uk_K_r7_reg[40]/NET0131 ,
		\u1_uk_K_r7_reg[47]/NET0131 ,
		_w19334_
	);
	LUT4 #(
		.INIT('hc693)
	) name13508 (
		decrypt_pad,
		\u1_R7_reg[4]/NET0131 ,
		\u1_uk_K_r7_reg[11]/NET0131 ,
		\u1_uk_K_r7_reg[4]/NET0131 ,
		_w19335_
	);
	LUT4 #(
		.INIT('hc693)
	) name13509 (
		decrypt_pad,
		\u1_R7_reg[9]/NET0131 ,
		\u1_uk_K_r7_reg[3]/NET0131 ,
		\u1_uk_K_r7_reg[53]/NET0131 ,
		_w19336_
	);
	LUT4 #(
		.INIT('hc693)
	) name13510 (
		decrypt_pad,
		\u1_R7_reg[6]/NET0131 ,
		\u1_uk_K_r7_reg[13]/NET0131 ,
		\u1_uk_K_r7_reg[6]/NET0131 ,
		_w19337_
	);
	LUT4 #(
		.INIT('h59fb)
	) name13511 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19338_
	);
	LUT2 #(
		.INIT('h1)
	) name13512 (
		_w19333_,
		_w19338_,
		_w19339_
	);
	LUT4 #(
		.INIT('h0034)
	) name13513 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19340_
	);
	LUT4 #(
		.INIT('h0800)
	) name13514 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19341_
	);
	LUT2 #(
		.INIT('h2)
	) name13515 (
		_w19336_,
		_w19337_,
		_w19342_
	);
	LUT4 #(
		.INIT('h0004)
	) name13516 (
		_w19333_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19343_
	);
	LUT4 #(
		.INIT('h4000)
	) name13517 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19344_
	);
	LUT4 #(
		.INIT('h0007)
	) name13518 (
		_w19333_,
		_w19341_,
		_w19343_,
		_w19344_,
		_w19345_
	);
	LUT4 #(
		.INIT('h5455)
	) name13519 (
		_w19332_,
		_w19339_,
		_w19340_,
		_w19345_,
		_w19346_
	);
	LUT4 #(
		.INIT('he6ee)
	) name13520 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19347_
	);
	LUT4 #(
		.INIT('h4044)
	) name13521 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19348_
	);
	LUT3 #(
		.INIT('h51)
	) name13522 (
		_w19333_,
		_w19334_,
		_w19337_,
		_w19349_
	);
	LUT4 #(
		.INIT('hf200)
	) name13523 (
		_w19332_,
		_w19347_,
		_w19348_,
		_w19349_,
		_w19350_
	);
	LUT3 #(
		.INIT('h10)
	) name13524 (
		_w19336_,
		_w19334_,
		_w19337_,
		_w19351_
	);
	LUT4 #(
		.INIT('h0100)
	) name13525 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19352_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name13526 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19353_
	);
	LUT2 #(
		.INIT('h2)
	) name13527 (
		_w19333_,
		_w19353_,
		_w19354_
	);
	LUT4 #(
		.INIT('h0082)
	) name13528 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19355_
	);
	LUT4 #(
		.INIT('h80a0)
	) name13529 (
		_w19333_,
		_w19335_,
		_w19334_,
		_w19337_,
		_w19356_
	);
	LUT3 #(
		.INIT('ha8)
	) name13530 (
		_w19332_,
		_w19355_,
		_w19356_,
		_w19357_
	);
	LUT3 #(
		.INIT('h01)
	) name13531 (
		_w19354_,
		_w19357_,
		_w19350_,
		_w19358_
	);
	LUT3 #(
		.INIT('h65)
	) name13532 (
		\u1_L7_reg[2]/NET0131 ,
		_w19346_,
		_w19358_,
		_w19359_
	);
	LUT4 #(
		.INIT('hfcdf)
	) name13533 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19360_
	);
	LUT2 #(
		.INIT('h1)
	) name13534 (
		_w19206_,
		_w19360_,
		_w19361_
	);
	LUT4 #(
		.INIT('he36f)
	) name13535 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19362_
	);
	LUT4 #(
		.INIT('h0301)
	) name13536 (
		_w19206_,
		_w19209_,
		_w19212_,
		_w19362_,
		_w19363_
	);
	LUT3 #(
		.INIT('h45)
	) name13537 (
		_w19200_,
		_w19361_,
		_w19363_,
		_w19364_
	);
	LUT4 #(
		.INIT('h4000)
	) name13538 (
		_w19201_,
		_w19206_,
		_w19202_,
		_w19204_,
		_w19365_
	);
	LUT4 #(
		.INIT('h5eff)
	) name13539 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19366_
	);
	LUT4 #(
		.INIT('h0d00)
	) name13540 (
		_w19211_,
		_w19215_,
		_w19365_,
		_w19366_,
		_w19367_
	);
	LUT3 #(
		.INIT('h9e)
	) name13541 (
		_w19202_,
		_w19204_,
		_w19203_,
		_w19368_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name13542 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19369_
	);
	LUT4 #(
		.INIT('h2223)
	) name13543 (
		_w19201_,
		_w19206_,
		_w19202_,
		_w19204_,
		_w19370_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name13544 (
		_w19218_,
		_w19368_,
		_w19369_,
		_w19370_,
		_w19371_
	);
	LUT3 #(
		.INIT('hd0)
	) name13545 (
		_w19200_,
		_w19367_,
		_w19371_,
		_w19372_
	);
	LUT3 #(
		.INIT('h65)
	) name13546 (
		\u1_L7_reg[4]/NET0131 ,
		_w19364_,
		_w19372_,
		_w19373_
	);
	LUT4 #(
		.INIT('hc963)
	) name13547 (
		decrypt_pad,
		\u1_R7_reg[32]/NET0131 ,
		\u1_uk_K_r7_reg[43]/NET0131 ,
		\u1_uk_K_r7_reg[50]/NET0131 ,
		_w19374_
	);
	LUT4 #(
		.INIT('hc963)
	) name13548 (
		decrypt_pad,
		\u1_R7_reg[31]/P0001 ,
		\u1_uk_K_r7_reg[37]/NET0131 ,
		\u1_uk_K_r7_reg[44]/NET0131 ,
		_w19375_
	);
	LUT4 #(
		.INIT('hc963)
	) name13549 (
		decrypt_pad,
		\u1_R7_reg[28]/NET0131 ,
		\u1_uk_K_r7_reg[21]/NET0131 ,
		\u1_uk_K_r7_reg[28]/NET0131 ,
		_w19376_
	);
	LUT4 #(
		.INIT('hc693)
	) name13550 (
		decrypt_pad,
		\u1_R7_reg[29]/NET0131 ,
		\u1_uk_K_r7_reg[0]/NET0131 ,
		\u1_uk_K_r7_reg[52]/NET0131 ,
		_w19377_
	);
	LUT4 #(
		.INIT('hc693)
	) name13551 (
		decrypt_pad,
		\u1_R7_reg[1]/NET0131 ,
		\u1_uk_K_r7_reg[16]/NET0131 ,
		\u1_uk_K_r7_reg[9]/NET0131 ,
		_w19378_
	);
	LUT4 #(
		.INIT('hc693)
	) name13552 (
		decrypt_pad,
		\u1_R7_reg[30]/NET0131 ,
		\u1_uk_K_r7_reg[1]/NET0131 ,
		\u1_uk_K_r7_reg[49]/NET0131 ,
		_w19379_
	);
	LUT4 #(
		.INIT('hfcdf)
	) name13553 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19380_
	);
	LUT4 #(
		.INIT('h23a5)
	) name13554 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19381_
	);
	LUT4 #(
		.INIT('h0040)
	) name13555 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19382_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name13556 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19383_
	);
	LUT4 #(
		.INIT('he400)
	) name13557 (
		_w19375_,
		_w19381_,
		_w19380_,
		_w19383_,
		_w19384_
	);
	LUT2 #(
		.INIT('h1)
	) name13558 (
		_w19374_,
		_w19384_,
		_w19385_
	);
	LUT3 #(
		.INIT('h01)
	) name13559 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19386_
	);
	LUT4 #(
		.INIT('h509c)
	) name13560 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19387_
	);
	LUT4 #(
		.INIT('h0800)
	) name13561 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19388_
	);
	LUT4 #(
		.INIT('h001d)
	) name13562 (
		_w19386_,
		_w19375_,
		_w19387_,
		_w19388_,
		_w19389_
	);
	LUT4 #(
		.INIT('h0008)
	) name13563 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19390_
	);
	LUT4 #(
		.INIT('hfff6)
	) name13564 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19391_
	);
	LUT4 #(
		.INIT('h0200)
	) name13565 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19392_
	);
	LUT4 #(
		.INIT('h1000)
	) name13566 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19393_
	);
	LUT4 #(
		.INIT('h0020)
	) name13567 (
		_w19375_,
		_w19392_,
		_w19391_,
		_w19393_,
		_w19394_
	);
	LUT4 #(
		.INIT('h2000)
	) name13568 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19374_,
		_w19395_
	);
	LUT3 #(
		.INIT('h01)
	) name13569 (
		_w19375_,
		_w19382_,
		_w19395_,
		_w19396_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name13570 (
		_w19389_,
		_w19374_,
		_w19394_,
		_w19396_,
		_w19397_
	);
	LUT3 #(
		.INIT('h9a)
	) name13571 (
		\u1_L7_reg[5]/NET0131 ,
		_w19385_,
		_w19397_,
		_w19398_
	);
	LUT4 #(
		.INIT('h0006)
	) name13572 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19399_
	);
	LUT3 #(
		.INIT('h47)
	) name13573 (
		_w19234_,
		_w19235_,
		_w19239_,
		_w19400_
	);
	LUT4 #(
		.INIT('h0051)
	) name13574 (
		_w19233_,
		_w19245_,
		_w19400_,
		_w19399_,
		_w19401_
	);
	LUT3 #(
		.INIT('h10)
	) name13575 (
		_w19234_,
		_w19236_,
		_w19238_,
		_w19402_
	);
	LUT4 #(
		.INIT('h2100)
	) name13576 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19403_
	);
	LUT2 #(
		.INIT('h6)
	) name13577 (
		_w19235_,
		_w19236_,
		_w19404_
	);
	LUT4 #(
		.INIT('h143c)
	) name13578 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19405_
	);
	LUT3 #(
		.INIT('h32)
	) name13579 (
		_w19239_,
		_w19403_,
		_w19405_,
		_w19406_
	);
	LUT2 #(
		.INIT('h8)
	) name13580 (
		_w19401_,
		_w19406_,
		_w19407_
	);
	LUT2 #(
		.INIT('h4)
	) name13581 (
		_w19239_,
		_w19246_,
		_w19408_
	);
	LUT3 #(
		.INIT('h02)
	) name13582 (
		_w19233_,
		_w19243_,
		_w19257_,
		_w19409_
	);
	LUT4 #(
		.INIT('h0240)
	) name13583 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19410_
	);
	LUT4 #(
		.INIT('h33fe)
	) name13584 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19411_
	);
	LUT3 #(
		.INIT('h31)
	) name13585 (
		_w19239_,
		_w19410_,
		_w19411_,
		_w19412_
	);
	LUT3 #(
		.INIT('h40)
	) name13586 (
		_w19408_,
		_w19409_,
		_w19412_,
		_w19413_
	);
	LUT3 #(
		.INIT('ha9)
	) name13587 (
		\u1_L7_reg[12]/NET0131 ,
		_w19407_,
		_w19413_,
		_w19414_
	);
	LUT4 #(
		.INIT('h5515)
	) name13588 (
		_w19333_,
		_w19335_,
		_w19336_,
		_w19334_,
		_w19415_
	);
	LUT3 #(
		.INIT('h40)
	) name13589 (
		_w19335_,
		_w19336_,
		_w19337_,
		_w19416_
	);
	LUT3 #(
		.INIT('h01)
	) name13590 (
		_w19336_,
		_w19334_,
		_w19337_,
		_w19417_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13591 (
		_w19333_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19418_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name13592 (
		_w19351_,
		_w19415_,
		_w19416_,
		_w19418_,
		_w19419_
	);
	LUT4 #(
		.INIT('h0010)
	) name13593 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19420_
	);
	LUT4 #(
		.INIT('h0002)
	) name13594 (
		_w19332_,
		_w19343_,
		_w19344_,
		_w19420_,
		_w19421_
	);
	LUT2 #(
		.INIT('h4)
	) name13595 (
		_w19419_,
		_w19421_,
		_w19422_
	);
	LUT3 #(
		.INIT('h32)
	) name13596 (
		_w19333_,
		_w19335_,
		_w19334_,
		_w19423_
	);
	LUT2 #(
		.INIT('h8)
	) name13597 (
		_w19342_,
		_w19423_,
		_w19424_
	);
	LUT2 #(
		.INIT('h8)
	) name13598 (
		_w19333_,
		_w19335_,
		_w19425_
	);
	LUT3 #(
		.INIT('hb0)
	) name13599 (
		_w19336_,
		_w19334_,
		_w19337_,
		_w19426_
	);
	LUT3 #(
		.INIT('h15)
	) name13600 (
		_w19332_,
		_w19425_,
		_w19426_,
		_w19427_
	);
	LUT4 #(
		.INIT('h5455)
	) name13601 (
		_w19333_,
		_w19335_,
		_w19336_,
		_w19334_,
		_w19428_
	);
	LUT4 #(
		.INIT('h0400)
	) name13602 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19429_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name13603 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19430_
	);
	LUT2 #(
		.INIT('h8)
	) name13604 (
		_w19428_,
		_w19430_,
		_w19431_
	);
	LUT3 #(
		.INIT('h40)
	) name13605 (
		_w19424_,
		_w19427_,
		_w19431_,
		_w19432_
	);
	LUT4 #(
		.INIT('h2000)
	) name13606 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19433_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name13607 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19434_
	);
	LUT3 #(
		.INIT('h09)
	) name13608 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19435_
	);
	LUT3 #(
		.INIT('h02)
	) name13609 (
		_w19335_,
		_w19336_,
		_w19337_,
		_w19436_
	);
	LUT4 #(
		.INIT('h0020)
	) name13610 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19437_
	);
	LUT3 #(
		.INIT('h02)
	) name13611 (
		_w19333_,
		_w19437_,
		_w19435_,
		_w19438_
	);
	LUT3 #(
		.INIT('h40)
	) name13612 (
		_w19424_,
		_w19427_,
		_w19438_,
		_w19439_
	);
	LUT4 #(
		.INIT('h001f)
	) name13613 (
		_w19422_,
		_w19432_,
		_w19434_,
		_w19439_,
		_w19440_
	);
	LUT2 #(
		.INIT('h9)
	) name13614 (
		\u1_L7_reg[13]/NET0131 ,
		_w19440_,
		_w19441_
	);
	LUT4 #(
		.INIT('hc963)
	) name13615 (
		decrypt_pad,
		\u1_R7_reg[19]/NET0131 ,
		\u1_uk_K_r7_reg[44]/NET0131 ,
		\u1_uk_K_r7_reg[51]/NET0131 ,
		_w19442_
	);
	LUT4 #(
		.INIT('hc963)
	) name13616 (
		decrypt_pad,
		\u1_R7_reg[18]/NET0131 ,
		\u1_uk_K_r7_reg[2]/NET0131 ,
		\u1_uk_K_r7_reg[9]/NET0131 ,
		_w19443_
	);
	LUT4 #(
		.INIT('hc693)
	) name13617 (
		decrypt_pad,
		\u1_R7_reg[17]/NET0131 ,
		\u1_uk_K_r7_reg[15]/NET0131 ,
		\u1_uk_K_r7_reg[8]/NET0131 ,
		_w19444_
	);
	LUT4 #(
		.INIT('hc963)
	) name13618 (
		decrypt_pad,
		\u1_R7_reg[21]/NET0131 ,
		\u1_uk_K_r7_reg[29]/NET0131 ,
		\u1_uk_K_r7_reg[36]/NET0131 ,
		_w19445_
	);
	LUT4 #(
		.INIT('hc963)
	) name13619 (
		decrypt_pad,
		\u1_R7_reg[16]/NET0131 ,
		\u1_uk_K_r7_reg[45]/NET0131 ,
		\u1_uk_K_r7_reg[52]/NET0131 ,
		_w19446_
	);
	LUT4 #(
		.INIT('h4000)
	) name13620 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19447_
	);
	LUT2 #(
		.INIT('h4)
	) name13621 (
		_w19445_,
		_w19446_,
		_w19448_
	);
	LUT4 #(
		.INIT('h0100)
	) name13622 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19449_
	);
	LUT4 #(
		.INIT('hb6c7)
	) name13623 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19450_
	);
	LUT3 #(
		.INIT('h04)
	) name13624 (
		_w19443_,
		_w19444_,
		_w19446_,
		_w19451_
	);
	LUT4 #(
		.INIT('h5fb8)
	) name13625 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19452_
	);
	LUT4 #(
		.INIT('h2000)
	) name13626 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19453_
	);
	LUT4 #(
		.INIT('hdffb)
	) name13627 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19454_
	);
	LUT4 #(
		.INIT('he400)
	) name13628 (
		_w19442_,
		_w19450_,
		_w19452_,
		_w19454_,
		_w19455_
	);
	LUT4 #(
		.INIT('hc963)
	) name13629 (
		decrypt_pad,
		\u1_R7_reg[20]/NET0131 ,
		\u1_uk_K_r7_reg[28]/NET0131 ,
		\u1_uk_K_r7_reg[35]/NET0131 ,
		_w19456_
	);
	LUT2 #(
		.INIT('h1)
	) name13630 (
		_w19455_,
		_w19456_,
		_w19457_
	);
	LUT4 #(
		.INIT('ha34f)
	) name13631 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19458_
	);
	LUT2 #(
		.INIT('h2)
	) name13632 (
		_w19442_,
		_w19458_,
		_w19459_
	);
	LUT2 #(
		.INIT('h1)
	) name13633 (
		_w19442_,
		_w19443_,
		_w19460_
	);
	LUT3 #(
		.INIT('hf6)
	) name13634 (
		_w19444_,
		_w19445_,
		_w19446_,
		_w19461_
	);
	LUT2 #(
		.INIT('h2)
	) name13635 (
		_w19460_,
		_w19461_,
		_w19462_
	);
	LUT4 #(
		.INIT('h0600)
	) name13636 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19463_
	);
	LUT3 #(
		.INIT('h8c)
	) name13637 (
		_w19442_,
		_w19443_,
		_w19444_,
		_w19464_
	);
	LUT4 #(
		.INIT('hb000)
	) name13638 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19465_
	);
	LUT3 #(
		.INIT('h45)
	) name13639 (
		_w19463_,
		_w19464_,
		_w19465_,
		_w19466_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name13640 (
		_w19456_,
		_w19459_,
		_w19462_,
		_w19466_,
		_w19467_
	);
	LUT4 #(
		.INIT('h0400)
	) name13641 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19468_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name13642 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19469_
	);
	LUT4 #(
		.INIT('h0020)
	) name13643 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19470_
	);
	LUT4 #(
		.INIT('hffd7)
	) name13644 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19471_
	);
	LUT3 #(
		.INIT('hd8)
	) name13645 (
		_w19442_,
		_w19469_,
		_w19471_,
		_w19472_
	);
	LUT4 #(
		.INIT('h5655)
	) name13646 (
		\u1_L7_reg[14]/NET0131 ,
		_w19457_,
		_w19467_,
		_w19472_,
		_w19473_
	);
	LUT4 #(
		.INIT('h3c3b)
	) name13647 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19474_
	);
	LUT4 #(
		.INIT('h0010)
	) name13648 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19475_
	);
	LUT4 #(
		.INIT('h3302)
	) name13649 (
		_w19375_,
		_w19374_,
		_w19474_,
		_w19475_,
		_w19476_
	);
	LUT4 #(
		.INIT('hdbd6)
	) name13650 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19477_
	);
	LUT2 #(
		.INIT('h1)
	) name13651 (
		_w19375_,
		_w19477_,
		_w19478_
	);
	LUT4 #(
		.INIT('h0200)
	) name13652 (
		_w19379_,
		_w19377_,
		_w19375_,
		_w19378_,
		_w19479_
	);
	LUT4 #(
		.INIT('h2000)
	) name13653 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19480_
	);
	LUT4 #(
		.INIT('h9fbf)
	) name13654 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19481_
	);
	LUT4 #(
		.INIT('h0010)
	) name13655 (
		_w19377_,
		_w19376_,
		_w19375_,
		_w19378_,
		_w19482_
	);
	LUT4 #(
		.INIT('h0100)
	) name13656 (
		_w19390_,
		_w19482_,
		_w19479_,
		_w19481_,
		_w19483_
	);
	LUT4 #(
		.INIT('h0100)
	) name13657 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19484_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name13658 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19485_
	);
	LUT4 #(
		.INIT('h0004)
	) name13659 (
		_w19377_,
		_w19376_,
		_w19375_,
		_w19374_,
		_w19486_
	);
	LUT3 #(
		.INIT('h0d)
	) name13660 (
		_w19375_,
		_w19485_,
		_w19486_,
		_w19487_
	);
	LUT4 #(
		.INIT('h0d00)
	) name13661 (
		_w19374_,
		_w19483_,
		_w19478_,
		_w19487_,
		_w19488_
	);
	LUT3 #(
		.INIT('h65)
	) name13662 (
		\u1_L7_reg[15]/P0001 ,
		_w19476_,
		_w19488_,
		_w19489_
	);
	LUT4 #(
		.INIT('h1001)
	) name13663 (
		_w19206_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19490_
	);
	LUT4 #(
		.INIT('h0200)
	) name13664 (
		_w19206_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19491_
	);
	LUT3 #(
		.INIT('h15)
	) name13665 (
		_w19206_,
		_w19204_,
		_w19203_,
		_w19492_
	);
	LUT3 #(
		.INIT('h8c)
	) name13666 (
		_w19201_,
		_w19202_,
		_w19203_,
		_w19493_
	);
	LUT4 #(
		.INIT('h0045)
	) name13667 (
		_w19200_,
		_w19492_,
		_w19493_,
		_w19491_,
		_w19494_
	);
	LUT4 #(
		.INIT('h2000)
	) name13668 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19495_
	);
	LUT3 #(
		.INIT('h04)
	) name13669 (
		_w19206_,
		_w19202_,
		_w19203_,
		_w19496_
	);
	LUT4 #(
		.INIT('hef00)
	) name13670 (
		_w19201_,
		_w19204_,
		_w19203_,
		_w19200_,
		_w19497_
	);
	LUT3 #(
		.INIT('h10)
	) name13671 (
		_w19496_,
		_w19495_,
		_w19497_,
		_w19498_
	);
	LUT4 #(
		.INIT('hbbcf)
	) name13672 (
		_w19201_,
		_w19202_,
		_w19204_,
		_w19203_,
		_w19499_
	);
	LUT3 #(
		.INIT('h31)
	) name13673 (
		_w19206_,
		_w19321_,
		_w19499_,
		_w19500_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name13674 (
		_w19490_,
		_w19494_,
		_w19498_,
		_w19500_,
		_w19501_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name13675 (
		_w19201_,
		_w19203_,
		_w19212_,
		_w19226_,
		_w19502_
	);
	LUT3 #(
		.INIT('h65)
	) name13676 (
		\u1_L7_reg[19]/P0001 ,
		_w19501_,
		_w19502_,
		_w19503_
	);
	LUT4 #(
		.INIT('h048c)
	) name13677 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19504_
	);
	LUT4 #(
		.INIT('hfda8)
	) name13678 (
		_w19283_,
		_w19293_,
		_w19312_,
		_w19504_,
		_w19505_
	);
	LUT4 #(
		.INIT('h79ff)
	) name13679 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19506_
	);
	LUT3 #(
		.INIT('h45)
	) name13680 (
		_w19289_,
		_w19505_,
		_w19506_,
		_w19507_
	);
	LUT4 #(
		.INIT('hff51)
	) name13681 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19508_
	);
	LUT4 #(
		.INIT('hd4ff)
	) name13682 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19509_
	);
	LUT4 #(
		.INIT('h4000)
	) name13683 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19510_
	);
	LUT4 #(
		.INIT('hbfcf)
	) name13684 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19511_
	);
	LUT4 #(
		.INIT('he400)
	) name13685 (
		_w19283_,
		_w19509_,
		_w19508_,
		_w19511_,
		_w19512_
	);
	LUT4 #(
		.INIT('h8020)
	) name13686 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19513_
	);
	LUT4 #(
		.INIT('h6fdf)
	) name13687 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19514_
	);
	LUT2 #(
		.INIT('h2)
	) name13688 (
		_w19283_,
		_w19514_,
		_w19515_
	);
	LUT4 #(
		.INIT('haabf)
	) name13689 (
		_w19283_,
		_w19284_,
		_w19300_,
		_w19510_,
		_w19516_
	);
	LUT4 #(
		.INIT('h0d00)
	) name13690 (
		_w19289_,
		_w19512_,
		_w19515_,
		_w19516_,
		_w19517_
	);
	LUT3 #(
		.INIT('h65)
	) name13691 (
		\u1_L7_reg[1]/NET0131 ,
		_w19507_,
		_w19517_,
		_w19518_
	);
	LUT4 #(
		.INIT('hfe00)
	) name13692 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19375_,
		_w19519_
	);
	LUT4 #(
		.INIT('h4050)
	) name13693 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19520_
	);
	LUT4 #(
		.INIT('h9d80)
	) name13694 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19521_
	);
	LUT2 #(
		.INIT('h2)
	) name13695 (
		_w19519_,
		_w19521_,
		_w19522_
	);
	LUT3 #(
		.INIT('h01)
	) name13696 (
		_w19375_,
		_w19480_,
		_w19520_,
		_w19523_
	);
	LUT4 #(
		.INIT('h0082)
	) name13697 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19524_
	);
	LUT3 #(
		.INIT('h02)
	) name13698 (
		_w19374_,
		_w19484_,
		_w19524_,
		_w19525_
	);
	LUT3 #(
		.INIT('he0)
	) name13699 (
		_w19522_,
		_w19523_,
		_w19525_,
		_w19526_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name13700 (
		_w19377_,
		_w19376_,
		_w19375_,
		_w19378_,
		_w19527_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name13701 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19528_
	);
	LUT3 #(
		.INIT('h13)
	) name13702 (
		_w19519_,
		_w19527_,
		_w19528_,
		_w19529_
	);
	LUT4 #(
		.INIT('h0200)
	) name13703 (
		_w19379_,
		_w19376_,
		_w19375_,
		_w19378_,
		_w19530_
	);
	LUT4 #(
		.INIT('h00f7)
	) name13704 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19374_,
		_w19531_
	);
	LUT2 #(
		.INIT('h4)
	) name13705 (
		_w19530_,
		_w19531_,
		_w19532_
	);
	LUT2 #(
		.INIT('h4)
	) name13706 (
		_w19377_,
		_w19375_,
		_w19533_
	);
	LUT3 #(
		.INIT('h40)
	) name13707 (
		_w19379_,
		_w19376_,
		_w19378_,
		_w19534_
	);
	LUT4 #(
		.INIT('hffde)
	) name13708 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19535_
	);
	LUT3 #(
		.INIT('hb0)
	) name13709 (
		_w19533_,
		_w19534_,
		_w19535_,
		_w19536_
	);
	LUT3 #(
		.INIT('h40)
	) name13710 (
		_w19529_,
		_w19532_,
		_w19536_,
		_w19537_
	);
	LUT3 #(
		.INIT('ha9)
	) name13711 (
		\u1_L7_reg[21]/NET0131 ,
		_w19526_,
		_w19537_,
		_w19538_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name13712 (
		_w19167_,
		_w19170_,
		_w19168_,
		_w19169_,
		_w19539_
	);
	LUT4 #(
		.INIT('hfdef)
	) name13713 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19540_
	);
	LUT3 #(
		.INIT('h80)
	) name13714 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19541_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name13715 (
		_w19191_,
		_w19541_,
		_w19539_,
		_w19540_,
		_w19542_
	);
	LUT4 #(
		.INIT('h007e)
	) name13716 (
		_w19172_,
		_w19168_,
		_w19169_,
		_w19166_,
		_w19543_
	);
	LUT2 #(
		.INIT('h4)
	) name13717 (
		_w19180_,
		_w19543_,
		_w19544_
	);
	LUT2 #(
		.INIT('h4)
	) name13718 (
		_w19542_,
		_w19544_,
		_w19545_
	);
	LUT3 #(
		.INIT('h14)
	) name13719 (
		_w19167_,
		_w19168_,
		_w19169_,
		_w19546_
	);
	LUT4 #(
		.INIT('h0008)
	) name13720 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19547_
	);
	LUT4 #(
		.INIT('h0004)
	) name13721 (
		_w19170_,
		_w19540_,
		_w19546_,
		_w19547_,
		_w19548_
	);
	LUT3 #(
		.INIT('h40)
	) name13722 (
		_w19167_,
		_w19168_,
		_w19169_,
		_w19549_
	);
	LUT3 #(
		.INIT('h02)
	) name13723 (
		_w19170_,
		_w19184_,
		_w19549_,
		_w19550_
	);
	LUT4 #(
		.INIT('h1030)
	) name13724 (
		_w19179_,
		_w19183_,
		_w19166_,
		_w19175_,
		_w19551_
	);
	LUT3 #(
		.INIT('he0)
	) name13725 (
		_w19548_,
		_w19550_,
		_w19551_,
		_w19552_
	);
	LUT3 #(
		.INIT('he5)
	) name13726 (
		_w19167_,
		_w19168_,
		_w19169_,
		_w19553_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13727 (
		_w19171_,
		_w19195_,
		_w19541_,
		_w19553_,
		_w19554_
	);
	LUT4 #(
		.INIT('h56aa)
	) name13728 (
		\u1_L7_reg[23]/NET0131 ,
		_w19545_,
		_w19552_,
		_w19554_,
		_w19555_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name13729 (
		_w19442_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19556_
	);
	LUT2 #(
		.INIT('h1)
	) name13730 (
		_w19443_,
		_w19556_,
		_w19557_
	);
	LUT2 #(
		.INIT('h2)
	) name13731 (
		_w19442_,
		_w19445_,
		_w19558_
	);
	LUT3 #(
		.INIT('h08)
	) name13732 (
		_w19443_,
		_w19444_,
		_w19446_,
		_w19559_
	);
	LUT4 #(
		.INIT('h0100)
	) name13733 (
		_w19442_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19560_
	);
	LUT4 #(
		.INIT('h1011)
	) name13734 (
		_w19456_,
		_w19560_,
		_w19558_,
		_w19559_,
		_w19561_
	);
	LUT4 #(
		.INIT('h4555)
	) name13735 (
		_w19442_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19562_
	);
	LUT4 #(
		.INIT('h010b)
	) name13736 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19563_
	);
	LUT3 #(
		.INIT('h80)
	) name13737 (
		_w19444_,
		_w19445_,
		_w19446_,
		_w19564_
	);
	LUT4 #(
		.INIT('h2a88)
	) name13738 (
		_w19442_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19565_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name13739 (
		_w19451_,
		_w19562_,
		_w19563_,
		_w19565_,
		_w19566_
	);
	LUT4 #(
		.INIT('h0800)
	) name13740 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19567_
	);
	LUT4 #(
		.INIT('hbf00)
	) name13741 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19456_,
		_w19568_
	);
	LUT2 #(
		.INIT('h4)
	) name13742 (
		_w19567_,
		_w19568_,
		_w19569_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name13743 (
		_w19557_,
		_w19561_,
		_w19566_,
		_w19569_,
		_w19570_
	);
	LUT3 #(
		.INIT('h04)
	) name13744 (
		_w19442_,
		_w19443_,
		_w19444_,
		_w19571_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name13745 (
		_w19442_,
		_w19443_,
		_w19444_,
		_w19445_,
		_w19572_
	);
	LUT4 #(
		.INIT('hf7fd)
	) name13746 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19573_
	);
	LUT4 #(
		.INIT('hf7ed)
	) name13747 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19574_
	);
	LUT4 #(
		.INIT('hf351)
	) name13748 (
		_w19442_,
		_w19446_,
		_w19572_,
		_w19574_,
		_w19575_
	);
	LUT3 #(
		.INIT('h65)
	) name13749 (
		\u1_L7_reg[25]/NET0131 ,
		_w19570_,
		_w19575_,
		_w19576_
	);
	LUT3 #(
		.INIT('h02)
	) name13750 (
		_w19283_,
		_w19306_,
		_w19288_,
		_w19577_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13751 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19578_
	);
	LUT2 #(
		.INIT('h1)
	) name13752 (
		_w19289_,
		_w19578_,
		_w19579_
	);
	LUT4 #(
		.INIT('h0900)
	) name13753 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19580_
	);
	LUT2 #(
		.INIT('h2)
	) name13754 (
		_w19281_,
		_w19284_,
		_w19581_
	);
	LUT4 #(
		.INIT('h0004)
	) name13755 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19582_
	);
	LUT3 #(
		.INIT('h01)
	) name13756 (
		_w19283_,
		_w19580_,
		_w19582_,
		_w19583_
	);
	LUT3 #(
		.INIT('h45)
	) name13757 (
		_w19577_,
		_w19579_,
		_w19583_,
		_w19584_
	);
	LUT3 #(
		.INIT('h54)
	) name13758 (
		_w19281_,
		_w19284_,
		_w19282_,
		_w19585_
	);
	LUT4 #(
		.INIT('h4404)
	) name13759 (
		_w19283_,
		_w19287_,
		_w19281_,
		_w19284_,
		_w19586_
	);
	LUT4 #(
		.INIT('h0002)
	) name13760 (
		_w19283_,
		_w19287_,
		_w19281_,
		_w19282_,
		_w19587_
	);
	LUT4 #(
		.INIT('h0100)
	) name13761 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w19588_
	);
	LUT4 #(
		.INIT('h1011)
	) name13762 (
		_w19587_,
		_w19588_,
		_w19585_,
		_w19586_,
		_w19589_
	);
	LUT4 #(
		.INIT('hf3f7)
	) name13763 (
		_w19283_,
		_w19287_,
		_w19281_,
		_w19282_,
		_w19590_
	);
	LUT4 #(
		.INIT('h0c04)
	) name13764 (
		_w19284_,
		_w19289_,
		_w19510_,
		_w19590_,
		_w19591_
	);
	LUT2 #(
		.INIT('h4)
	) name13765 (
		_w19291_,
		_w19285_,
		_w19592_
	);
	LUT4 #(
		.INIT('h00fd)
	) name13766 (
		_w19281_,
		_w19284_,
		_w19282_,
		_w19289_,
		_w19593_
	);
	LUT3 #(
		.INIT('h10)
	) name13767 (
		_w19306_,
		_w19308_,
		_w19593_,
		_w19594_
	);
	LUT4 #(
		.INIT('h7077)
	) name13768 (
		_w19589_,
		_w19591_,
		_w19592_,
		_w19594_,
		_w19595_
	);
	LUT3 #(
		.INIT('h56)
	) name13769 (
		\u1_L7_reg[26]/NET0131 ,
		_w19584_,
		_w19595_,
		_w19596_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name13770 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19597_
	);
	LUT2 #(
		.INIT('h2)
	) name13771 (
		_w19333_,
		_w19597_,
		_w19598_
	);
	LUT4 #(
		.INIT('hbfae)
	) name13772 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19599_
	);
	LUT2 #(
		.INIT('h1)
	) name13773 (
		_w19333_,
		_w19599_,
		_w19600_
	);
	LUT4 #(
		.INIT('h7737)
	) name13774 (
		_w19333_,
		_w19335_,
		_w19336_,
		_w19334_,
		_w19601_
	);
	LUT3 #(
		.INIT('h32)
	) name13775 (
		_w19337_,
		_w19429_,
		_w19601_,
		_w19602_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name13776 (
		_w19332_,
		_w19600_,
		_w19598_,
		_w19602_,
		_w19603_
	);
	LUT4 #(
		.INIT('hdaff)
	) name13777 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19604_
	);
	LUT2 #(
		.INIT('h1)
	) name13778 (
		_w19333_,
		_w19604_,
		_w19605_
	);
	LUT4 #(
		.INIT('h1145)
	) name13779 (
		_w19333_,
		_w19335_,
		_w19336_,
		_w19334_,
		_w19606_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name13780 (
		_w19333_,
		_w19436_,
		_w19599_,
		_w19606_,
		_w19607_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name13781 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19608_
	);
	LUT4 #(
		.INIT('h2322)
	) name13782 (
		_w19332_,
		_w19605_,
		_w19607_,
		_w19608_,
		_w19609_
	);
	LUT3 #(
		.INIT('h65)
	) name13783 (
		\u1_L7_reg[28]/NET0131 ,
		_w19603_,
		_w19609_,
		_w19610_
	);
	LUT4 #(
		.INIT('h0001)
	) name13784 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19611_
	);
	LUT4 #(
		.INIT('hcffe)
	) name13785 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19612_
	);
	LUT4 #(
		.INIT('hef00)
	) name13786 (
		_w19442_,
		_w19443_,
		_w19446_,
		_w19456_,
		_w19613_
	);
	LUT4 #(
		.INIT('hc400)
	) name13787 (
		_w19442_,
		_w19471_,
		_w19612_,
		_w19613_,
		_w19614_
	);
	LUT4 #(
		.INIT('h00d0)
	) name13788 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19615_
	);
	LUT2 #(
		.INIT('h2)
	) name13789 (
		_w19562_,
		_w19615_,
		_w19616_
	);
	LUT3 #(
		.INIT('h02)
	) name13790 (
		_w19442_,
		_w19449_,
		_w19564_,
		_w19617_
	);
	LUT4 #(
		.INIT('h00fb)
	) name13791 (
		_w19443_,
		_w19444_,
		_w19446_,
		_w19456_,
		_w19618_
	);
	LUT2 #(
		.INIT('h8)
	) name13792 (
		_w19573_,
		_w19618_,
		_w19619_
	);
	LUT4 #(
		.INIT('h0155)
	) name13793 (
		_w19614_,
		_w19616_,
		_w19617_,
		_w19619_,
		_w19620_
	);
	LUT4 #(
		.INIT('hf797)
	) name13794 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19621_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13795 (
		_w19442_,
		_w19448_,
		_w19571_,
		_w19621_,
		_w19622_
	);
	LUT3 #(
		.INIT('h65)
	) name13796 (
		\u1_L7_reg[8]/NET0131 ,
		_w19620_,
		_w19622_,
		_w19623_
	);
	LUT4 #(
		.INIT('hc004)
	) name13797 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19624_
	);
	LUT3 #(
		.INIT('h28)
	) name13798 (
		_w19377_,
		_w19376_,
		_w19378_,
		_w19625_
	);
	LUT4 #(
		.INIT('hf3e2)
	) name13799 (
		_w19386_,
		_w19375_,
		_w19624_,
		_w19625_,
		_w19626_
	);
	LUT4 #(
		.INIT('he6df)
	) name13800 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19627_
	);
	LUT3 #(
		.INIT('h8a)
	) name13801 (
		_w19374_,
		_w19626_,
		_w19627_,
		_w19628_
	);
	LUT4 #(
		.INIT('hf700)
	) name13802 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19375_,
		_w19629_
	);
	LUT3 #(
		.INIT('h4b)
	) name13803 (
		_w19379_,
		_w19377_,
		_w19378_,
		_w19630_
	);
	LUT4 #(
		.INIT('h0800)
	) name13804 (
		_w19379_,
		_w19376_,
		_w19375_,
		_w19378_,
		_w19631_
	);
	LUT4 #(
		.INIT('h0015)
	) name13805 (
		_w19392_,
		_w19629_,
		_w19630_,
		_w19631_,
		_w19632_
	);
	LUT4 #(
		.INIT('h0002)
	) name13806 (
		_w19377_,
		_w19376_,
		_w19378_,
		_w19374_,
		_w19633_
	);
	LUT4 #(
		.INIT('hefb7)
	) name13807 (
		_w19379_,
		_w19377_,
		_w19376_,
		_w19378_,
		_w19634_
	);
	LUT4 #(
		.INIT('h0020)
	) name13808 (
		_w19379_,
		_w19377_,
		_w19375_,
		_w19378_,
		_w19635_
	);
	LUT4 #(
		.INIT('h00ba)
	) name13809 (
		_w19375_,
		_w19633_,
		_w19634_,
		_w19635_,
		_w19636_
	);
	LUT3 #(
		.INIT('he0)
	) name13810 (
		_w19374_,
		_w19632_,
		_w19636_,
		_w19637_
	);
	LUT3 #(
		.INIT('h65)
	) name13811 (
		\u1_L7_reg[27]/NET0131 ,
		_w19628_,
		_w19637_,
		_w19638_
	);
	LUT2 #(
		.INIT('h9)
	) name13812 (
		_w19236_,
		_w19238_,
		_w19639_
	);
	LUT4 #(
		.INIT('hd003)
	) name13813 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19640_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name13814 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19641_
	);
	LUT3 #(
		.INIT('h01)
	) name13815 (
		_w19239_,
		_w19641_,
		_w19640_,
		_w19642_
	);
	LUT4 #(
		.INIT('h0800)
	) name13816 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19643_
	);
	LUT4 #(
		.INIT('hb5bc)
	) name13817 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19644_
	);
	LUT3 #(
		.INIT('h31)
	) name13818 (
		_w19239_,
		_w19643_,
		_w19644_,
		_w19645_
	);
	LUT3 #(
		.INIT('h8a)
	) name13819 (
		_w19233_,
		_w19642_,
		_w19645_,
		_w19646_
	);
	LUT3 #(
		.INIT('h40)
	) name13820 (
		_w19235_,
		_w19236_,
		_w19238_,
		_w19647_
	);
	LUT4 #(
		.INIT('hab89)
	) name13821 (
		_w19239_,
		_w19402_,
		_w19404_,
		_w19647_,
		_w19648_
	);
	LUT4 #(
		.INIT('h7bd7)
	) name13822 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19649_
	);
	LUT4 #(
		.INIT('h00c8)
	) name13823 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19239_,
		_w19650_
	);
	LUT4 #(
		.INIT('h135f)
	) name13824 (
		_w19239_,
		_w19254_,
		_w19246_,
		_w19650_,
		_w19651_
	);
	LUT4 #(
		.INIT('hba00)
	) name13825 (
		_w19233_,
		_w19648_,
		_w19649_,
		_w19651_,
		_w19652_
	);
	LUT3 #(
		.INIT('h65)
	) name13826 (
		\u1_L7_reg[32]/NET0131 ,
		_w19646_,
		_w19652_,
		_w19653_
	);
	LUT4 #(
		.INIT('h0200)
	) name13827 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19654_
	);
	LUT4 #(
		.INIT('h0040)
	) name13828 (
		_w19442_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19655_
	);
	LUT4 #(
		.INIT('h0004)
	) name13829 (
		_w19447_,
		_w19456_,
		_w19655_,
		_w19654_,
		_w19656_
	);
	LUT4 #(
		.INIT('haff3)
	) name13830 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19657_
	);
	LUT4 #(
		.INIT('h2022)
	) name13831 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19658_
	);
	LUT4 #(
		.INIT('hf3af)
	) name13832 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19659_
	);
	LUT3 #(
		.INIT('h10)
	) name13833 (
		_w19456_,
		_w19658_,
		_w19659_,
		_w19660_
	);
	LUT3 #(
		.INIT('h02)
	) name13834 (
		_w19442_,
		_w19449_,
		_w19470_,
		_w19661_
	);
	LUT4 #(
		.INIT('hf800)
	) name13835 (
		_w19656_,
		_w19657_,
		_w19660_,
		_w19661_,
		_w19662_
	);
	LUT4 #(
		.INIT('h4f50)
	) name13836 (
		_w19443_,
		_w19444_,
		_w19445_,
		_w19446_,
		_w19663_
	);
	LUT3 #(
		.INIT('h10)
	) name13837 (
		_w19456_,
		_w19658_,
		_w19663_,
		_w19664_
	);
	LUT4 #(
		.INIT('h0001)
	) name13838 (
		_w19442_,
		_w19453_,
		_w19468_,
		_w19611_,
		_w19665_
	);
	LUT3 #(
		.INIT('he0)
	) name13839 (
		_w19656_,
		_w19664_,
		_w19665_,
		_w19666_
	);
	LUT3 #(
		.INIT('ha9)
	) name13840 (
		\u1_L7_reg[3]/NET0131 ,
		_w19662_,
		_w19666_,
		_w19667_
	);
	LUT4 #(
		.INIT('hc963)
	) name13841 (
		decrypt_pad,
		\u1_R7_reg[11]/NET0131 ,
		\u1_uk_K_r7_reg[11]/NET0131 ,
		\u1_uk_K_r7_reg[18]/NET0131 ,
		_w19668_
	);
	LUT4 #(
		.INIT('hc963)
	) name13842 (
		decrypt_pad,
		\u1_R7_reg[12]/NET0131 ,
		\u1_uk_K_r7_reg[26]/P0001 ,
		\u1_uk_K_r7_reg[33]/NET0131 ,
		_w19669_
	);
	LUT4 #(
		.INIT('hc963)
	) name13843 (
		decrypt_pad,
		\u1_R7_reg[13]/NET0131 ,
		\u1_uk_K_r7_reg[39]/NET0131 ,
		\u1_uk_K_r7_reg[46]/NET0131 ,
		_w19670_
	);
	LUT4 #(
		.INIT('hc963)
	) name13844 (
		decrypt_pad,
		\u1_R7_reg[9]/NET0131 ,
		\u1_uk_K_r7_reg[34]/NET0131 ,
		\u1_uk_K_r7_reg[41]/NET0131 ,
		_w19671_
	);
	LUT4 #(
		.INIT('hc963)
	) name13845 (
		decrypt_pad,
		\u1_R7_reg[10]/NET0131 ,
		\u1_uk_K_r7_reg[10]/NET0131 ,
		\u1_uk_K_r7_reg[17]/NET0131 ,
		_w19672_
	);
	LUT4 #(
		.INIT('hc693)
	) name13846 (
		decrypt_pad,
		\u1_R7_reg[8]/NET0131 ,
		\u1_uk_K_r7_reg[12]/NET0131 ,
		\u1_uk_K_r7_reg[5]/NET0131 ,
		_w19673_
	);
	LUT2 #(
		.INIT('h2)
	) name13847 (
		_w19670_,
		_w19673_,
		_w19674_
	);
	LUT4 #(
		.INIT('h95b5)
	) name13848 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19675_
	);
	LUT4 #(
		.INIT('h0001)
	) name13849 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19676_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name13850 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19677_
	);
	LUT4 #(
		.INIT('h08cc)
	) name13851 (
		_w19669_,
		_w19668_,
		_w19675_,
		_w19677_,
		_w19678_
	);
	LUT2 #(
		.INIT('h1)
	) name13852 (
		_w19671_,
		_w19672_,
		_w19679_
	);
	LUT2 #(
		.INIT('h6)
	) name13853 (
		_w19671_,
		_w19672_,
		_w19680_
	);
	LUT2 #(
		.INIT('h1)
	) name13854 (
		_w19670_,
		_w19673_,
		_w19681_
	);
	LUT2 #(
		.INIT('h8)
	) name13855 (
		_w19670_,
		_w19673_,
		_w19682_
	);
	LUT2 #(
		.INIT('h8)
	) name13856 (
		_w19670_,
		_w19668_,
		_w19683_
	);
	LUT3 #(
		.INIT('h46)
	) name13857 (
		_w19670_,
		_w19673_,
		_w19668_,
		_w19684_
	);
	LUT2 #(
		.INIT('h1)
	) name13858 (
		_w19680_,
		_w19684_,
		_w19685_
	);
	LUT3 #(
		.INIT('h80)
	) name13859 (
		_w19670_,
		_w19671_,
		_w19668_,
		_w19686_
	);
	LUT4 #(
		.INIT('h0660)
	) name13860 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19687_
	);
	LUT3 #(
		.INIT('h45)
	) name13861 (
		_w19669_,
		_w19686_,
		_w19687_,
		_w19688_
	);
	LUT3 #(
		.INIT('h80)
	) name13862 (
		_w19671_,
		_w19672_,
		_w19669_,
		_w19689_
	);
	LUT3 #(
		.INIT('h51)
	) name13863 (
		_w19673_,
		_w19671_,
		_w19672_,
		_w19690_
	);
	LUT4 #(
		.INIT('h0090)
	) name13864 (
		_w19670_,
		_w19671_,
		_w19669_,
		_w19668_,
		_w19691_
	);
	LUT4 #(
		.INIT('h7077)
	) name13865 (
		_w19681_,
		_w19689_,
		_w19690_,
		_w19691_,
		_w19692_
	);
	LUT4 #(
		.INIT('h4500)
	) name13866 (
		_w19678_,
		_w19685_,
		_w19688_,
		_w19692_,
		_w19693_
	);
	LUT2 #(
		.INIT('h9)
	) name13867 (
		\u1_L7_reg[6]/NET0131 ,
		_w19693_,
		_w19694_
	);
	LUT4 #(
		.INIT('hf126)
	) name13868 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19695_
	);
	LUT4 #(
		.INIT('h2880)
	) name13869 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19696_
	);
	LUT4 #(
		.INIT('h5004)
	) name13870 (
		_w19234_,
		_w19235_,
		_w19236_,
		_w19238_,
		_w19697_
	);
	LUT4 #(
		.INIT('h1302)
	) name13871 (
		_w19239_,
		_w19696_,
		_w19697_,
		_w19695_,
		_w19698_
	);
	LUT2 #(
		.INIT('h2)
	) name13872 (
		_w19233_,
		_w19698_,
		_w19699_
	);
	LUT2 #(
		.INIT('h4)
	) name13873 (
		_w19239_,
		_w19696_,
		_w19700_
	);
	LUT2 #(
		.INIT('h2)
	) name13874 (
		_w19233_,
		_w19239_,
		_w19701_
	);
	LUT3 #(
		.INIT('h4c)
	) name13875 (
		_w19235_,
		_w19236_,
		_w19238_,
		_w19702_
	);
	LUT4 #(
		.INIT('h8a00)
	) name13876 (
		_w19234_,
		_w19236_,
		_w19238_,
		_w19239_,
		_w19703_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name13877 (
		_w19240_,
		_w19639_,
		_w19702_,
		_w19703_,
		_w19704_
	);
	LUT3 #(
		.INIT('h45)
	) name13878 (
		_w19253_,
		_w19239_,
		_w19697_,
		_w19705_
	);
	LUT4 #(
		.INIT('h0133)
	) name13879 (
		_w19233_,
		_w19701_,
		_w19704_,
		_w19705_,
		_w19706_
	);
	LUT4 #(
		.INIT('h5556)
	) name13880 (
		\u1_L7_reg[7]/NET0131 ,
		_w19700_,
		_w19706_,
		_w19699_,
		_w19707_
	);
	LUT4 #(
		.INIT('h0df0)
	) name13881 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19708_
	);
	LUT3 #(
		.INIT('h14)
	) name13882 (
		_w19170_,
		_w19168_,
		_w19169_,
		_w19709_
	);
	LUT3 #(
		.INIT('h0e)
	) name13883 (
		_w19191_,
		_w19708_,
		_w19709_,
		_w19710_
	);
	LUT4 #(
		.INIT('h2084)
	) name13884 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19711_
	);
	LUT2 #(
		.INIT('h1)
	) name13885 (
		_w19166_,
		_w19711_,
		_w19712_
	);
	LUT4 #(
		.INIT('h8448)
	) name13886 (
		_w19167_,
		_w19172_,
		_w19168_,
		_w19169_,
		_w19713_
	);
	LUT4 #(
		.INIT('h1030)
	) name13887 (
		_w19167_,
		_w19172_,
		_w19170_,
		_w19169_,
		_w19714_
	);
	LUT4 #(
		.INIT('h2022)
	) name13888 (
		_w19166_,
		_w19266_,
		_w19274_,
		_w19714_,
		_w19715_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name13889 (
		_w19710_,
		_w19712_,
		_w19713_,
		_w19715_,
		_w19716_
	);
	LUT3 #(
		.INIT('h40)
	) name13890 (
		_w19170_,
		_w19168_,
		_w19169_,
		_w19717_
	);
	LUT2 #(
		.INIT('h4)
	) name13891 (
		_w19192_,
		_w19717_,
		_w19718_
	);
	LUT3 #(
		.INIT('h56)
	) name13892 (
		\u1_L7_reg[9]/NET0131 ,
		_w19716_,
		_w19718_,
		_w19719_
	);
	LUT3 #(
		.INIT('h80)
	) name13893 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19720_
	);
	LUT3 #(
		.INIT('h68)
	) name13894 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19721_
	);
	LUT4 #(
		.INIT('h0068)
	) name13895 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19669_,
		_w19722_
	);
	LUT4 #(
		.INIT('h4100)
	) name13896 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19723_
	);
	LUT3 #(
		.INIT('h02)
	) name13897 (
		_w19668_,
		_w19723_,
		_w19722_,
		_w19724_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name13898 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19725_
	);
	LUT3 #(
		.INIT('h20)
	) name13899 (
		_w19673_,
		_w19671_,
		_w19672_,
		_w19726_
	);
	LUT4 #(
		.INIT('h00df)
	) name13900 (
		_w19673_,
		_w19671_,
		_w19672_,
		_w19668_,
		_w19727_
	);
	LUT3 #(
		.INIT('he0)
	) name13901 (
		_w19669_,
		_w19725_,
		_w19727_,
		_w19728_
	);
	LUT2 #(
		.INIT('h1)
	) name13902 (
		_w19724_,
		_w19728_,
		_w19729_
	);
	LUT3 #(
		.INIT('h04)
	) name13903 (
		_w19669_,
		_w19676_,
		_w19725_,
		_w19730_
	);
	LUT4 #(
		.INIT('h0111)
	) name13904 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19668_,
		_w19731_
	);
	LUT3 #(
		.INIT('h01)
	) name13905 (
		_w19672_,
		_w19721_,
		_w19731_,
		_w19732_
	);
	LUT4 #(
		.INIT('h0014)
	) name13906 (
		_w19670_,
		_w19673_,
		_w19672_,
		_w19668_,
		_w19733_
	);
	LUT4 #(
		.INIT('h2000)
	) name13907 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19734_
	);
	LUT2 #(
		.INIT('h1)
	) name13908 (
		_w19733_,
		_w19734_,
		_w19735_
	);
	LUT4 #(
		.INIT('h1311)
	) name13909 (
		_w19669_,
		_w19730_,
		_w19732_,
		_w19735_,
		_w19736_
	);
	LUT3 #(
		.INIT('h65)
	) name13910 (
		\u1_L7_reg[16]/NET0131 ,
		_w19729_,
		_w19736_,
		_w19737_
	);
	LUT4 #(
		.INIT('hfd75)
	) name13911 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19738_
	);
	LUT2 #(
		.INIT('h1)
	) name13912 (
		_w19333_,
		_w19738_,
		_w19739_
	);
	LUT4 #(
		.INIT('h0a20)
	) name13913 (
		_w19333_,
		_w19335_,
		_w19336_,
		_w19334_,
		_w19740_
	);
	LUT3 #(
		.INIT('h02)
	) name13914 (
		_w19332_,
		_w19352_,
		_w19740_,
		_w19741_
	);
	LUT2 #(
		.INIT('h4)
	) name13915 (
		_w19739_,
		_w19741_,
		_w19742_
	);
	LUT4 #(
		.INIT('h1003)
	) name13916 (
		_w19333_,
		_w19335_,
		_w19334_,
		_w19337_,
		_w19743_
	);
	LUT3 #(
		.INIT('h01)
	) name13917 (
		_w19332_,
		_w19433_,
		_w19417_,
		_w19744_
	);
	LUT4 #(
		.INIT('h8000)
	) name13918 (
		_w19333_,
		_w19335_,
		_w19336_,
		_w19334_,
		_w19745_
	);
	LUT2 #(
		.INIT('h1)
	) name13919 (
		_w19341_,
		_w19745_,
		_w19746_
	);
	LUT3 #(
		.INIT('h40)
	) name13920 (
		_w19743_,
		_w19744_,
		_w19746_,
		_w19747_
	);
	LUT4 #(
		.INIT('h1000)
	) name13921 (
		_w19333_,
		_w19335_,
		_w19336_,
		_w19334_,
		_w19748_
	);
	LUT4 #(
		.INIT('h77ef)
	) name13922 (
		_w19335_,
		_w19336_,
		_w19334_,
		_w19337_,
		_w19749_
	);
	LUT3 #(
		.INIT('h31)
	) name13923 (
		_w19333_,
		_w19748_,
		_w19749_,
		_w19750_
	);
	LUT4 #(
		.INIT('ha955)
	) name13924 (
		\u1_L7_reg[18]/NET0131 ,
		_w19742_,
		_w19747_,
		_w19750_,
		_w19751_
	);
	LUT4 #(
		.INIT('h0400)
	) name13925 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19752_
	);
	LUT3 #(
		.INIT('hed)
	) name13926 (
		_w19670_,
		_w19673_,
		_w19672_,
		_w19753_
	);
	LUT3 #(
		.INIT('h10)
	) name13927 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19754_
	);
	LUT4 #(
		.INIT('he2cd)
	) name13928 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19755_
	);
	LUT4 #(
		.INIT('h5054)
	) name13929 (
		_w19669_,
		_w19668_,
		_w19752_,
		_w19755_,
		_w19756_
	);
	LUT2 #(
		.INIT('h8)
	) name13930 (
		_w19679_,
		_w19684_,
		_w19757_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name13931 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19758_
	);
	LUT3 #(
		.INIT('he0)
	) name13932 (
		_w19671_,
		_w19672_,
		_w19668_,
		_w19759_
	);
	LUT4 #(
		.INIT('h0302)
	) name13933 (
		_w19668_,
		_w19674_,
		_w19759_,
		_w19758_,
		_w19760_
	);
	LUT3 #(
		.INIT('ha8)
	) name13934 (
		_w19669_,
		_w19757_,
		_w19760_,
		_w19761_
	);
	LUT4 #(
		.INIT('h1dff)
	) name13935 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19762_
	);
	LUT4 #(
		.INIT('h0024)
	) name13936 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19763_
	);
	LUT4 #(
		.INIT('hcc08)
	) name13937 (
		_w19669_,
		_w19668_,
		_w19762_,
		_w19763_,
		_w19764_
	);
	LUT2 #(
		.INIT('h2)
	) name13938 (
		_w19672_,
		_w19668_,
		_w19765_
	);
	LUT4 #(
		.INIT('h0009)
	) name13939 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19766_
	);
	LUT4 #(
		.INIT('h9db6)
	) name13940 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19767_
	);
	LUT2 #(
		.INIT('h1)
	) name13941 (
		_w19669_,
		_w19668_,
		_w19768_
	);
	LUT4 #(
		.INIT('h7077)
	) name13942 (
		_w19720_,
		_w19765_,
		_w19767_,
		_w19768_,
		_w19769_
	);
	LUT2 #(
		.INIT('h4)
	) name13943 (
		_w19764_,
		_w19769_,
		_w19770_
	);
	LUT4 #(
		.INIT('h5655)
	) name13944 (
		\u1_L7_reg[24]/NET0131 ,
		_w19756_,
		_w19761_,
		_w19770_,
		_w19771_
	);
	LUT4 #(
		.INIT('h0004)
	) name13945 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19772_
	);
	LUT3 #(
		.INIT('h08)
	) name13946 (
		_w19668_,
		_w19753_,
		_w19772_,
		_w19773_
	);
	LUT3 #(
		.INIT('h07)
	) name13947 (
		_w19673_,
		_w19672_,
		_w19668_,
		_w19774_
	);
	LUT2 #(
		.INIT('h4)
	) name13948 (
		_w19754_,
		_w19774_,
		_w19775_
	);
	LUT3 #(
		.INIT('ha8)
	) name13949 (
		_w19669_,
		_w19773_,
		_w19775_,
		_w19776_
	);
	LUT4 #(
		.INIT('h20ac)
	) name13950 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19777_
	);
	LUT4 #(
		.INIT('h8c00)
	) name13951 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19778_
	);
	LUT3 #(
		.INIT('h04)
	) name13952 (
		_w19670_,
		_w19671_,
		_w19672_,
		_w19779_
	);
	LUT4 #(
		.INIT('heee4)
	) name13953 (
		_w19668_,
		_w19777_,
		_w19779_,
		_w19778_,
		_w19780_
	);
	LUT4 #(
		.INIT('h0200)
	) name13954 (
		_w19670_,
		_w19673_,
		_w19671_,
		_w19672_,
		_w19781_
	);
	LUT3 #(
		.INIT('h01)
	) name13955 (
		_w19669_,
		_w19766_,
		_w19781_,
		_w19782_
	);
	LUT2 #(
		.INIT('h4)
	) name13956 (
		_w19780_,
		_w19782_,
		_w19783_
	);
	LUT2 #(
		.INIT('h8)
	) name13957 (
		_w19683_,
		_w19726_,
		_w19784_
	);
	LUT4 #(
		.INIT('h0040)
	) name13958 (
		_w19670_,
		_w19671_,
		_w19672_,
		_w19668_,
		_w19785_
	);
	LUT3 #(
		.INIT('h0d)
	) name13959 (
		_w19689_,
		_w19682_,
		_w19785_,
		_w19786_
	);
	LUT2 #(
		.INIT('h4)
	) name13960 (
		_w19784_,
		_w19786_,
		_w19787_
	);
	LUT4 #(
		.INIT('h56aa)
	) name13961 (
		\u1_L7_reg[30]/NET0131 ,
		_w19776_,
		_w19783_,
		_w19787_,
		_w19788_
	);
	LUT4 #(
		.INIT('hc693)
	) name13962 (
		decrypt_pad,
		\u1_R6_reg[28]/NET0131 ,
		\u1_uk_K_r6_reg[23]/P0001 ,
		\u1_uk_K_r6_reg[30]/P0001 ,
		_w19789_
	);
	LUT4 #(
		.INIT('hc693)
	) name13963 (
		decrypt_pad,
		\u1_R6_reg[26]/NET0131 ,
		\u1_uk_K_r6_reg[31]/NET0131 ,
		\u1_uk_K_r6_reg[38]/NET0131 ,
		_w19790_
	);
	LUT4 #(
		.INIT('hc693)
	) name13964 (
		decrypt_pad,
		\u1_R6_reg[25]/NET0131 ,
		\u1_uk_K_r6_reg[42]/NET0131 ,
		\u1_uk_K_r6_reg[49]/NET0131 ,
		_w19791_
	);
	LUT4 #(
		.INIT('hc693)
	) name13965 (
		decrypt_pad,
		\u1_R6_reg[29]/NET0131 ,
		\u1_uk_K_r6_reg[15]/NET0131 ,
		\u1_uk_K_r6_reg[22]/NET0131 ,
		_w19792_
	);
	LUT3 #(
		.INIT('hea)
	) name13966 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19793_
	);
	LUT4 #(
		.INIT('hc963)
	) name13967 (
		decrypt_pad,
		\u1_R6_reg[24]/NET0131 ,
		\u1_uk_K_r6_reg[14]/NET0131 ,
		\u1_uk_K_r6_reg[7]/NET0131 ,
		_w19794_
	);
	LUT4 #(
		.INIT('hc693)
	) name13968 (
		decrypt_pad,
		\u1_R6_reg[27]/NET0131 ,
		\u1_uk_K_r6_reg[36]/NET0131 ,
		\u1_uk_K_r6_reg[43]/NET0131 ,
		_w19795_
	);
	LUT3 #(
		.INIT('h70)
	) name13969 (
		_w19790_,
		_w19791_,
		_w19795_,
		_w19796_
	);
	LUT4 #(
		.INIT('h7000)
	) name13970 (
		_w19790_,
		_w19791_,
		_w19794_,
		_w19795_,
		_w19797_
	);
	LUT2 #(
		.INIT('h8)
	) name13971 (
		_w19793_,
		_w19797_,
		_w19798_
	);
	LUT4 #(
		.INIT('h1000)
	) name13972 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19799_
	);
	LUT4 #(
		.INIT('hef3f)
	) name13973 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19800_
	);
	LUT2 #(
		.INIT('h2)
	) name13974 (
		_w19792_,
		_w19794_,
		_w19801_
	);
	LUT4 #(
		.INIT('h0020)
	) name13975 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19802_
	);
	LUT4 #(
		.INIT('hffde)
	) name13976 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19803_
	);
	LUT3 #(
		.INIT('he0)
	) name13977 (
		_w19795_,
		_w19800_,
		_w19803_,
		_w19804_
	);
	LUT3 #(
		.INIT('h8a)
	) name13978 (
		_w19789_,
		_w19798_,
		_w19804_,
		_w19805_
	);
	LUT4 #(
		.INIT('h0072)
	) name13979 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19795_,
		_w19806_
	);
	LUT4 #(
		.INIT('h10f0)
	) name13980 (
		_w19790_,
		_w19791_,
		_w19794_,
		_w19795_,
		_w19807_
	);
	LUT2 #(
		.INIT('h4)
	) name13981 (
		_w19806_,
		_w19807_,
		_w19808_
	);
	LUT4 #(
		.INIT('h0002)
	) name13982 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19809_
	);
	LUT2 #(
		.INIT('h6)
	) name13983 (
		_w19790_,
		_w19794_,
		_w19810_
	);
	LUT3 #(
		.INIT('h8c)
	) name13984 (
		_w19791_,
		_w19792_,
		_w19795_,
		_w19811_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name13985 (
		_w19809_,
		_w19795_,
		_w19810_,
		_w19811_,
		_w19812_
	);
	LUT4 #(
		.INIT('h0008)
	) name13986 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19813_
	);
	LUT4 #(
		.INIT('hfcd7)
	) name13987 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19814_
	);
	LUT4 #(
		.INIT('h0084)
	) name13988 (
		_w19790_,
		_w19791_,
		_w19794_,
		_w19795_,
		_w19815_
	);
	LUT4 #(
		.INIT('h0100)
	) name13989 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19795_,
		_w19816_
	);
	LUT4 #(
		.INIT('h0031)
	) name13990 (
		_w19795_,
		_w19815_,
		_w19814_,
		_w19816_,
		_w19817_
	);
	LUT4 #(
		.INIT('hba00)
	) name13991 (
		_w19789_,
		_w19808_,
		_w19812_,
		_w19817_,
		_w19818_
	);
	LUT3 #(
		.INIT('h65)
	) name13992 (
		\u1_L6_reg[22]/NET0131 ,
		_w19805_,
		_w19818_,
		_w19819_
	);
	LUT4 #(
		.INIT('hc693)
	) name13993 (
		decrypt_pad,
		\u1_R6_reg[3]/NET0131 ,
		\u1_uk_K_r6_reg[12]/NET0131 ,
		\u1_uk_K_r6_reg[19]/NET0131 ,
		_w19820_
	);
	LUT4 #(
		.INIT('hc693)
	) name13994 (
		decrypt_pad,
		\u1_R6_reg[4]/NET0131 ,
		\u1_uk_K_r6_reg[47]/NET0131 ,
		\u1_uk_K_r6_reg[54]/NET0131 ,
		_w19821_
	);
	LUT4 #(
		.INIT('hc963)
	) name13995 (
		decrypt_pad,
		\u1_R6_reg[2]/NET0131 ,
		\u1_uk_K_r6_reg[10]/NET0131 ,
		\u1_uk_K_r6_reg[3]/NET0131 ,
		_w19822_
	);
	LUT4 #(
		.INIT('hc693)
	) name13996 (
		decrypt_pad,
		\u1_R6_reg[1]/NET0131 ,
		\u1_uk_K_r6_reg[20]/NET0131 ,
		\u1_uk_K_r6_reg[27]/NET0131 ,
		_w19823_
	);
	LUT4 #(
		.INIT('hc693)
	) name13997 (
		decrypt_pad,
		\u1_R6_reg[5]/NET0131 ,
		\u1_uk_K_r6_reg[18]/NET0131 ,
		\u1_uk_K_r6_reg[25]/NET0131 ,
		_w19824_
	);
	LUT4 #(
		.INIT('hc693)
	) name13998 (
		decrypt_pad,
		\u1_R6_reg[32]/NET0131 ,
		\u1_uk_K_r6_reg[24]/NET0131 ,
		\u1_uk_K_r6_reg[6]/NET0131 ,
		_w19825_
	);
	LUT4 #(
		.INIT('heff4)
	) name13999 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w19826_
	);
	LUT4 #(
		.INIT('h7dbd)
	) name14000 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w19827_
	);
	LUT4 #(
		.INIT('h0133)
	) name14001 (
		_w19821_,
		_w19820_,
		_w19826_,
		_w19827_,
		_w19828_
	);
	LUT3 #(
		.INIT('h04)
	) name14002 (
		_w19824_,
		_w19822_,
		_w19825_,
		_w19829_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name14003 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w19830_
	);
	LUT2 #(
		.INIT('h4)
	) name14004 (
		_w19830_,
		_w19820_,
		_w19831_
	);
	LUT2 #(
		.INIT('h4)
	) name14005 (
		_w19822_,
		_w19820_,
		_w19832_
	);
	LUT3 #(
		.INIT('h8a)
	) name14006 (
		_w19823_,
		_w19822_,
		_w19820_,
		_w19833_
	);
	LUT2 #(
		.INIT('h2)
	) name14007 (
		_w19824_,
		_w19825_,
		_w19834_
	);
	LUT4 #(
		.INIT('h0100)
	) name14008 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w19835_
	);
	LUT4 #(
		.INIT('h04a4)
	) name14009 (
		_w19823_,
		_w19822_,
		_w19825_,
		_w19820_,
		_w19836_
	);
	LUT4 #(
		.INIT('h1011)
	) name14010 (
		_w19835_,
		_w19836_,
		_w19833_,
		_w19834_,
		_w19837_
	);
	LUT3 #(
		.INIT('h8a)
	) name14011 (
		_w19821_,
		_w19831_,
		_w19837_,
		_w19838_
	);
	LUT4 #(
		.INIT('h2800)
	) name14012 (
		_w19823_,
		_w19824_,
		_w19825_,
		_w19820_,
		_w19839_
	);
	LUT2 #(
		.INIT('h2)
	) name14013 (
		_w19822_,
		_w19839_,
		_w19840_
	);
	LUT4 #(
		.INIT('hc040)
	) name14014 (
		_w19823_,
		_w19824_,
		_w19825_,
		_w19820_,
		_w19841_
	);
	LUT3 #(
		.INIT('h02)
	) name14015 (
		_w19823_,
		_w19824_,
		_w19825_,
		_w19842_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name14016 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w19843_
	);
	LUT3 #(
		.INIT('h45)
	) name14017 (
		_w19821_,
		_w19841_,
		_w19843_,
		_w19844_
	);
	LUT2 #(
		.INIT('h4)
	) name14018 (
		_w19823_,
		_w19820_,
		_w19845_
	);
	LUT2 #(
		.INIT('h4)
	) name14019 (
		_w19822_,
		_w19825_,
		_w19846_
	);
	LUT4 #(
		.INIT('h1000)
	) name14020 (
		_w19823_,
		_w19822_,
		_w19825_,
		_w19820_,
		_w19847_
	);
	LUT3 #(
		.INIT('h07)
	) name14021 (
		_w19829_,
		_w19845_,
		_w19847_,
		_w19848_
	);
	LUT3 #(
		.INIT('hb0)
	) name14022 (
		_w19840_,
		_w19844_,
		_w19848_,
		_w19849_
	);
	LUT4 #(
		.INIT('h5655)
	) name14023 (
		\u1_L6_reg[31]/NET0131 ,
		_w19838_,
		_w19828_,
		_w19849_,
		_w19850_
	);
	LUT4 #(
		.INIT('hc693)
	) name14024 (
		decrypt_pad,
		\u1_R6_reg[24]/NET0131 ,
		\u1_uk_K_r6_reg[16]/NET0131 ,
		\u1_uk_K_r6_reg[23]/P0001 ,
		_w19851_
	);
	LUT4 #(
		.INIT('hc693)
	) name14025 (
		decrypt_pad,
		\u1_R6_reg[23]/NET0131 ,
		\u1_uk_K_r6_reg[14]/NET0131 ,
		\u1_uk_K_r6_reg[21]/NET0131 ,
		_w19852_
	);
	LUT4 #(
		.INIT('hc693)
	) name14026 (
		decrypt_pad,
		\u1_R6_reg[21]/NET0131 ,
		\u1_uk_K_r6_reg[38]/NET0131 ,
		\u1_uk_K_r6_reg[45]/NET0131 ,
		_w19853_
	);
	LUT4 #(
		.INIT('hc963)
	) name14027 (
		decrypt_pad,
		\u1_R6_reg[20]/NET0131 ,
		\u1_uk_K_r6_reg[2]/NET0131 ,
		\u1_uk_K_r6_reg[50]/NET0131 ,
		_w19854_
	);
	LUT4 #(
		.INIT('hc693)
	) name14028 (
		decrypt_pad,
		\u1_R6_reg[22]/NET0131 ,
		\u1_uk_K_r6_reg[1]/NET0131 ,
		\u1_uk_K_r6_reg[8]/NET0131 ,
		_w19855_
	);
	LUT4 #(
		.INIT('hc693)
	) name14029 (
		decrypt_pad,
		\u1_R6_reg[25]/NET0131 ,
		\u1_uk_K_r6_reg[35]/NET0131 ,
		\u1_uk_K_r6_reg[42]/NET0131 ,
		_w19856_
	);
	LUT3 #(
		.INIT('hc4)
	) name14030 (
		_w19853_,
		_w19854_,
		_w19856_,
		_w19857_
	);
	LUT4 #(
		.INIT('h57db)
	) name14031 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w19858_
	);
	LUT2 #(
		.INIT('h2)
	) name14032 (
		_w19852_,
		_w19858_,
		_w19859_
	);
	LUT4 #(
		.INIT('he020)
	) name14033 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w19860_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name14034 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w19861_
	);
	LUT3 #(
		.INIT('h01)
	) name14035 (
		_w19852_,
		_w19861_,
		_w19860_,
		_w19862_
	);
	LUT2 #(
		.INIT('h1)
	) name14036 (
		_w19855_,
		_w19852_,
		_w19863_
	);
	LUT4 #(
		.INIT('h0200)
	) name14037 (
		_w19854_,
		_w19855_,
		_w19852_,
		_w19856_,
		_w19864_
	);
	LUT2 #(
		.INIT('h4)
	) name14038 (
		_w19853_,
		_w19864_,
		_w19865_
	);
	LUT4 #(
		.INIT('haaa8)
	) name14039 (
		_w19851_,
		_w19862_,
		_w19859_,
		_w19865_,
		_w19866_
	);
	LUT4 #(
		.INIT('h0028)
	) name14040 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19852_,
		_w19867_
	);
	LUT4 #(
		.INIT('h1000)
	) name14041 (
		_w19853_,
		_w19854_,
		_w19852_,
		_w19856_,
		_w19868_
	);
	LUT4 #(
		.INIT('h0008)
	) name14042 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w19869_
	);
	LUT3 #(
		.INIT('h10)
	) name14043 (
		_w19854_,
		_w19855_,
		_w19852_,
		_w19870_
	);
	LUT3 #(
		.INIT('h01)
	) name14044 (
		_w19869_,
		_w19870_,
		_w19868_,
		_w19871_
	);
	LUT4 #(
		.INIT('haf8c)
	) name14045 (
		_w19853_,
		_w19855_,
		_w19852_,
		_w19856_,
		_w19872_
	);
	LUT3 #(
		.INIT('h8a)
	) name14046 (
		_w19854_,
		_w19855_,
		_w19852_,
		_w19873_
	);
	LUT4 #(
		.INIT('h4000)
	) name14047 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w19874_
	);
	LUT3 #(
		.INIT('h0b)
	) name14048 (
		_w19872_,
		_w19873_,
		_w19874_,
		_w19875_
	);
	LUT4 #(
		.INIT('h00bf)
	) name14049 (
		_w19867_,
		_w19871_,
		_w19875_,
		_w19851_,
		_w19876_
	);
	LUT4 #(
		.INIT('heff7)
	) name14050 (
		_w19853_,
		_w19854_,
		_w19852_,
		_w19856_,
		_w19877_
	);
	LUT2 #(
		.INIT('h1)
	) name14051 (
		_w19855_,
		_w19877_,
		_w19878_
	);
	LUT4 #(
		.INIT('h0002)
	) name14052 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w19879_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name14053 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w19880_
	);
	LUT4 #(
		.INIT('h0001)
	) name14054 (
		_w19854_,
		_w19855_,
		_w19852_,
		_w19856_,
		_w19881_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name14055 (
		_w19853_,
		_w19852_,
		_w19880_,
		_w19881_,
		_w19882_
	);
	LUT2 #(
		.INIT('h4)
	) name14056 (
		_w19878_,
		_w19882_,
		_w19883_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name14057 (
		\u1_L6_reg[11]/NET0131 ,
		_w19876_,
		_w19866_,
		_w19883_,
		_w19884_
	);
	LUT4 #(
		.INIT('hc693)
	) name14058 (
		decrypt_pad,
		\u1_R6_reg[13]/NET0131 ,
		\u1_uk_K_r6_reg[32]/NET0131 ,
		\u1_uk_K_r6_reg[39]/NET0131 ,
		_w19885_
	);
	LUT4 #(
		.INIT('hc693)
	) name14059 (
		decrypt_pad,
		\u1_R6_reg[15]/NET0131 ,
		\u1_uk_K_r6_reg[41]/NET0131 ,
		\u1_uk_K_r6_reg[48]/NET0131 ,
		_w19886_
	);
	LUT4 #(
		.INIT('hc693)
	) name14060 (
		decrypt_pad,
		\u1_R6_reg[12]/NET0131 ,
		\u1_uk_K_r6_reg[13]/NET0131 ,
		\u1_uk_K_r6_reg[20]/NET0131 ,
		_w19887_
	);
	LUT4 #(
		.INIT('hc693)
	) name14061 (
		decrypt_pad,
		\u1_R6_reg[14]/NET0131 ,
		\u1_uk_K_r6_reg[33]/NET0131 ,
		\u1_uk_K_r6_reg[40]/NET0131 ,
		_w19888_
	);
	LUT4 #(
		.INIT('h4000)
	) name14062 (
		_w19887_,
		_w19885_,
		_w19886_,
		_w19888_,
		_w19889_
	);
	LUT4 #(
		.INIT('hc693)
	) name14063 (
		decrypt_pad,
		\u1_R6_reg[16]/NET0131 ,
		\u1_uk_K_r6_reg[17]/NET0131 ,
		\u1_uk_K_r6_reg[24]/NET0131 ,
		_w19890_
	);
	LUT2 #(
		.INIT('h1)
	) name14064 (
		_w19889_,
		_w19890_,
		_w19891_
	);
	LUT4 #(
		.INIT('hc963)
	) name14065 (
		decrypt_pad,
		\u1_R6_reg[17]/NET0131 ,
		\u1_uk_K_r6_reg[4]/NET0131 ,
		\u1_uk_K_r6_reg[54]/NET0131 ,
		_w19892_
	);
	LUT4 #(
		.INIT('h8000)
	) name14066 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19886_,
		_w19893_
	);
	LUT4 #(
		.INIT('h0008)
	) name14067 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w19894_
	);
	LUT2 #(
		.INIT('h4)
	) name14068 (
		_w19885_,
		_w19886_,
		_w19895_
	);
	LUT4 #(
		.INIT('h0100)
	) name14069 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19886_,
		_w19896_
	);
	LUT3 #(
		.INIT('h01)
	) name14070 (
		_w19894_,
		_w19896_,
		_w19893_,
		_w19897_
	);
	LUT2 #(
		.INIT('h2)
	) name14071 (
		_w19887_,
		_w19892_,
		_w19898_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name14072 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w19899_
	);
	LUT2 #(
		.INIT('h4)
	) name14073 (
		_w19887_,
		_w19885_,
		_w19900_
	);
	LUT2 #(
		.INIT('h4)
	) name14074 (
		_w19892_,
		_w19888_,
		_w19901_
	);
	LUT4 #(
		.INIT('h1000)
	) name14075 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w19902_
	);
	LUT4 #(
		.INIT('heffe)
	) name14076 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w19903_
	);
	LUT3 #(
		.INIT('he0)
	) name14077 (
		_w19886_,
		_w19899_,
		_w19903_,
		_w19904_
	);
	LUT3 #(
		.INIT('h80)
	) name14078 (
		_w19891_,
		_w19897_,
		_w19904_,
		_w19905_
	);
	LUT2 #(
		.INIT('h1)
	) name14079 (
		_w19885_,
		_w19886_,
		_w19906_
	);
	LUT4 #(
		.INIT('h0001)
	) name14080 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19886_,
		_w19907_
	);
	LUT4 #(
		.INIT('h7f7e)
	) name14081 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19886_,
		_w19908_
	);
	LUT2 #(
		.INIT('h2)
	) name14082 (
		_w19888_,
		_w19908_,
		_w19909_
	);
	LUT2 #(
		.INIT('h9)
	) name14083 (
		_w19887_,
		_w19885_,
		_w19910_
	);
	LUT4 #(
		.INIT('h0006)
	) name14084 (
		_w19887_,
		_w19885_,
		_w19886_,
		_w19888_,
		_w19911_
	);
	LUT4 #(
		.INIT('h2000)
	) name14085 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19886_,
		_w19912_
	);
	LUT4 #(
		.INIT('h0040)
	) name14086 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w19913_
	);
	LUT2 #(
		.INIT('h4)
	) name14087 (
		_w19887_,
		_w19892_,
		_w19914_
	);
	LUT4 #(
		.INIT('h0400)
	) name14088 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19886_,
		_w19915_
	);
	LUT4 #(
		.INIT('h0004)
	) name14089 (
		_w19912_,
		_w19890_,
		_w19913_,
		_w19915_,
		_w19916_
	);
	LUT3 #(
		.INIT('h10)
	) name14090 (
		_w19911_,
		_w19909_,
		_w19916_,
		_w19917_
	);
	LUT3 #(
		.INIT('hde)
	) name14091 (
		_w19887_,
		_w19892_,
		_w19888_,
		_w19918_
	);
	LUT2 #(
		.INIT('h2)
	) name14092 (
		_w19895_,
		_w19918_,
		_w19919_
	);
	LUT3 #(
		.INIT('h02)
	) name14093 (
		_w19892_,
		_w19886_,
		_w19888_,
		_w19920_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name14094 (
		_w19912_,
		_w19888_,
		_w19900_,
		_w19920_,
		_w19921_
	);
	LUT2 #(
		.INIT('h4)
	) name14095 (
		_w19919_,
		_w19921_,
		_w19922_
	);
	LUT4 #(
		.INIT('ha955)
	) name14096 (
		\u1_L6_reg[20]/NET0131 ,
		_w19905_,
		_w19917_,
		_w19922_,
		_w19923_
	);
	LUT4 #(
		.INIT('hc693)
	) name14097 (
		decrypt_pad,
		\u1_R6_reg[28]/NET0131 ,
		\u1_uk_K_r6_reg[21]/NET0131 ,
		\u1_uk_K_r6_reg[28]/NET0131 ,
		_w19924_
	);
	LUT4 #(
		.INIT('hc963)
	) name14098 (
		decrypt_pad,
		\u1_R6_reg[1]/NET0131 ,
		\u1_uk_K_r6_reg[16]/NET0131 ,
		\u1_uk_K_r6_reg[9]/NET0131 ,
		_w19925_
	);
	LUT4 #(
		.INIT('hc963)
	) name14099 (
		decrypt_pad,
		\u1_R6_reg[29]/NET0131 ,
		\u1_uk_K_r6_reg[0]/NET0131 ,
		\u1_uk_K_r6_reg[52]/NET0131 ,
		_w19926_
	);
	LUT4 #(
		.INIT('hc963)
	) name14100 (
		decrypt_pad,
		\u1_R6_reg[30]/NET0131 ,
		\u1_uk_K_r6_reg[1]/NET0131 ,
		\u1_uk_K_r6_reg[49]/NET0131 ,
		_w19927_
	);
	LUT4 #(
		.INIT('hc693)
	) name14101 (
		decrypt_pad,
		\u1_R6_reg[31]/P0001 ,
		\u1_uk_K_r6_reg[37]/NET0131 ,
		\u1_uk_K_r6_reg[44]/NET0131 ,
		_w19928_
	);
	LUT4 #(
		.INIT('h7b70)
	) name14102 (
		_w19925_,
		_w19926_,
		_w19927_,
		_w19928_,
		_w19929_
	);
	LUT2 #(
		.INIT('h2)
	) name14103 (
		_w19924_,
		_w19929_,
		_w19930_
	);
	LUT4 #(
		.INIT('hf9fb)
	) name14104 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w19931_
	);
	LUT2 #(
		.INIT('h4)
	) name14105 (
		_w19931_,
		_w19928_,
		_w19932_
	);
	LUT3 #(
		.INIT('h0d)
	) name14106 (
		_w19924_,
		_w19925_,
		_w19928_,
		_w19933_
	);
	LUT3 #(
		.INIT('hd8)
	) name14107 (
		_w19925_,
		_w19926_,
		_w19927_,
		_w19934_
	);
	LUT4 #(
		.INIT('hc693)
	) name14108 (
		decrypt_pad,
		\u1_R6_reg[32]/NET0131 ,
		\u1_uk_K_r6_reg[43]/NET0131 ,
		\u1_uk_K_r6_reg[50]/NET0131 ,
		_w19935_
	);
	LUT3 #(
		.INIT('h07)
	) name14109 (
		_w19933_,
		_w19934_,
		_w19935_,
		_w19936_
	);
	LUT3 #(
		.INIT('h10)
	) name14110 (
		_w19932_,
		_w19930_,
		_w19936_,
		_w19937_
	);
	LUT4 #(
		.INIT('h0020)
	) name14111 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w19938_
	);
	LUT4 #(
		.INIT('hcf45)
	) name14112 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w19939_
	);
	LUT3 #(
		.INIT('h02)
	) name14113 (
		_w19928_,
		_w19939_,
		_w19938_,
		_w19940_
	);
	LUT4 #(
		.INIT('h0021)
	) name14114 (
		_w19924_,
		_w19926_,
		_w19927_,
		_w19928_,
		_w19941_
	);
	LUT4 #(
		.INIT('h4000)
	) name14115 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w19942_
	);
	LUT3 #(
		.INIT('h02)
	) name14116 (
		_w19935_,
		_w19942_,
		_w19941_,
		_w19943_
	);
	LUT2 #(
		.INIT('h4)
	) name14117 (
		_w19940_,
		_w19943_,
		_w19944_
	);
	LUT4 #(
		.INIT('h1008)
	) name14118 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w19945_
	);
	LUT4 #(
		.INIT('h0400)
	) name14119 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w19946_
	);
	LUT4 #(
		.INIT('hebf6)
	) name14120 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w19947_
	);
	LUT3 #(
		.INIT('hb1)
	) name14121 (
		_w19928_,
		_w19938_,
		_w19947_,
		_w19948_
	);
	LUT4 #(
		.INIT('h56aa)
	) name14122 (
		\u1_L6_reg[5]/NET0131 ,
		_w19937_,
		_w19944_,
		_w19948_,
		_w19949_
	);
	LUT4 #(
		.INIT('h8400)
	) name14123 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w19950_
	);
	LUT4 #(
		.INIT('hefe7)
	) name14124 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w19951_
	);
	LUT2 #(
		.INIT('h2)
	) name14125 (
		_w19886_,
		_w19951_,
		_w19952_
	);
	LUT3 #(
		.INIT('h31)
	) name14126 (
		_w19885_,
		_w19886_,
		_w19888_,
		_w19953_
	);
	LUT4 #(
		.INIT('h153f)
	) name14127 (
		_w19898_,
		_w19900_,
		_w19920_,
		_w19953_,
		_w19954_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name14128 (
		_w19890_,
		_w19952_,
		_w19950_,
		_w19954_,
		_w19955_
	);
	LUT3 #(
		.INIT('h08)
	) name14129 (
		_w19892_,
		_w19886_,
		_w19888_,
		_w19956_
	);
	LUT4 #(
		.INIT('h0040)
	) name14130 (
		_w19887_,
		_w19892_,
		_w19886_,
		_w19888_,
		_w19957_
	);
	LUT3 #(
		.INIT('ha2)
	) name14131 (
		_w19887_,
		_w19892_,
		_w19888_,
		_w19958_
	);
	LUT4 #(
		.INIT('h0013)
	) name14132 (
		_w19895_,
		_w19907_,
		_w19958_,
		_w19957_,
		_w19959_
	);
	LUT4 #(
		.INIT('hff31)
	) name14133 (
		_w19892_,
		_w19885_,
		_w19886_,
		_w19888_,
		_w19960_
	);
	LUT3 #(
		.INIT('hc4)
	) name14134 (
		_w19887_,
		_w19903_,
		_w19960_,
		_w19961_
	);
	LUT3 #(
		.INIT('h15)
	) name14135 (
		_w19890_,
		_w19959_,
		_w19961_,
		_w19962_
	);
	LUT4 #(
		.INIT('h7bfe)
	) name14136 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w19963_
	);
	LUT2 #(
		.INIT('h1)
	) name14137 (
		_w19886_,
		_w19963_,
		_w19964_
	);
	LUT3 #(
		.INIT('h0d)
	) name14138 (
		_w19912_,
		_w19888_,
		_w19889_,
		_w19965_
	);
	LUT2 #(
		.INIT('h4)
	) name14139 (
		_w19964_,
		_w19965_,
		_w19966_
	);
	LUT4 #(
		.INIT('h5655)
	) name14140 (
		\u1_L6_reg[10]/NET0131 ,
		_w19962_,
		_w19955_,
		_w19966_,
		_w19967_
	);
	LUT4 #(
		.INIT('h0006)
	) name14141 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19968_
	);
	LUT3 #(
		.INIT('h47)
	) name14142 (
		_w19790_,
		_w19791_,
		_w19795_,
		_w19969_
	);
	LUT4 #(
		.INIT('h0051)
	) name14143 (
		_w19789_,
		_w19801_,
		_w19969_,
		_w19968_,
		_w19970_
	);
	LUT3 #(
		.INIT('h10)
	) name14144 (
		_w19790_,
		_w19792_,
		_w19794_,
		_w19971_
	);
	LUT4 #(
		.INIT('h2100)
	) name14145 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19972_
	);
	LUT2 #(
		.INIT('h6)
	) name14146 (
		_w19791_,
		_w19792_,
		_w19973_
	);
	LUT4 #(
		.INIT('h143c)
	) name14147 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19974_
	);
	LUT3 #(
		.INIT('h32)
	) name14148 (
		_w19795_,
		_w19972_,
		_w19974_,
		_w19975_
	);
	LUT2 #(
		.INIT('h8)
	) name14149 (
		_w19970_,
		_w19975_,
		_w19976_
	);
	LUT2 #(
		.INIT('h4)
	) name14150 (
		_w19795_,
		_w19802_,
		_w19977_
	);
	LUT3 #(
		.INIT('h02)
	) name14151 (
		_w19789_,
		_w19799_,
		_w19813_,
		_w19978_
	);
	LUT4 #(
		.INIT('h0240)
	) name14152 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19979_
	);
	LUT4 #(
		.INIT('h33fe)
	) name14153 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w19980_
	);
	LUT3 #(
		.INIT('h31)
	) name14154 (
		_w19795_,
		_w19979_,
		_w19980_,
		_w19981_
	);
	LUT3 #(
		.INIT('h40)
	) name14155 (
		_w19977_,
		_w19978_,
		_w19981_,
		_w19982_
	);
	LUT3 #(
		.INIT('ha9)
	) name14156 (
		\u1_L6_reg[12]/NET0131 ,
		_w19976_,
		_w19982_,
		_w19983_
	);
	LUT4 #(
		.INIT('hc693)
	) name14157 (
		decrypt_pad,
		\u1_R6_reg[20]/NET0131 ,
		\u1_uk_K_r6_reg[28]/NET0131 ,
		\u1_uk_K_r6_reg[35]/NET0131 ,
		_w19984_
	);
	LUT4 #(
		.INIT('hc963)
	) name14158 (
		decrypt_pad,
		\u1_R6_reg[17]/NET0131 ,
		\u1_uk_K_r6_reg[15]/NET0131 ,
		\u1_uk_K_r6_reg[8]/NET0131 ,
		_w19985_
	);
	LUT4 #(
		.INIT('hc693)
	) name14159 (
		decrypt_pad,
		\u1_R6_reg[21]/NET0131 ,
		\u1_uk_K_r6_reg[29]/NET0131 ,
		\u1_uk_K_r6_reg[36]/NET0131 ,
		_w19986_
	);
	LUT2 #(
		.INIT('h6)
	) name14160 (
		_w19985_,
		_w19986_,
		_w19987_
	);
	LUT4 #(
		.INIT('hc693)
	) name14161 (
		decrypt_pad,
		\u1_R6_reg[18]/NET0131 ,
		\u1_uk_K_r6_reg[2]/NET0131 ,
		\u1_uk_K_r6_reg[9]/NET0131 ,
		_w19988_
	);
	LUT4 #(
		.INIT('hc693)
	) name14162 (
		decrypt_pad,
		\u1_R6_reg[16]/NET0131 ,
		\u1_uk_K_r6_reg[45]/NET0131 ,
		\u1_uk_K_r6_reg[52]/NET0131 ,
		_w19989_
	);
	LUT4 #(
		.INIT('h0900)
	) name14163 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w19990_
	);
	LUT4 #(
		.INIT('hc693)
	) name14164 (
		decrypt_pad,
		\u1_R6_reg[19]/NET0131 ,
		\u1_uk_K_r6_reg[44]/NET0131 ,
		\u1_uk_K_r6_reg[51]/NET0131 ,
		_w19991_
	);
	LUT4 #(
		.INIT('h2064)
	) name14165 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w19992_
	);
	LUT3 #(
		.INIT('h01)
	) name14166 (
		_w19991_,
		_w19992_,
		_w19990_,
		_w19993_
	);
	LUT4 #(
		.INIT('hc00a)
	) name14167 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w19994_
	);
	LUT4 #(
		.INIT('hfe00)
	) name14168 (
		_w19985_,
		_w19986_,
		_w19989_,
		_w19991_,
		_w19995_
	);
	LUT2 #(
		.INIT('h4)
	) name14169 (
		_w19994_,
		_w19995_,
		_w19996_
	);
	LUT4 #(
		.INIT('h4002)
	) name14170 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w19997_
	);
	LUT4 #(
		.INIT('h5501)
	) name14171 (
		_w19984_,
		_w19993_,
		_w19996_,
		_w19997_,
		_w19998_
	);
	LUT3 #(
		.INIT('h02)
	) name14172 (
		_w19985_,
		_w19988_,
		_w19989_,
		_w19999_
	);
	LUT4 #(
		.INIT('hd13b)
	) name14173 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20000_
	);
	LUT2 #(
		.INIT('h2)
	) name14174 (
		_w19991_,
		_w20000_,
		_w20001_
	);
	LUT3 #(
		.INIT('h4c)
	) name14175 (
		_w19986_,
		_w19988_,
		_w19989_,
		_w20002_
	);
	LUT3 #(
		.INIT('h0b)
	) name14176 (
		_w19988_,
		_w19989_,
		_w19991_,
		_w20003_
	);
	LUT4 #(
		.INIT('h1000)
	) name14177 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20004_
	);
	LUT4 #(
		.INIT('he9ff)
	) name14178 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20005_
	);
	LUT4 #(
		.INIT('hfb00)
	) name14179 (
		_w19987_,
		_w20003_,
		_w20002_,
		_w20005_,
		_w20006_
	);
	LUT4 #(
		.INIT('h0060)
	) name14180 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20007_
	);
	LUT4 #(
		.INIT('h0200)
	) name14181 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20008_
	);
	LUT4 #(
		.INIT('hfdef)
	) name14182 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20009_
	);
	LUT3 #(
		.INIT('hd1)
	) name14183 (
		_w20007_,
		_w19991_,
		_w20009_,
		_w20010_
	);
	LUT4 #(
		.INIT('h7500)
	) name14184 (
		_w19984_,
		_w20001_,
		_w20006_,
		_w20010_,
		_w20011_
	);
	LUT3 #(
		.INIT('h65)
	) name14185 (
		\u1_L6_reg[14]/NET0131 ,
		_w19998_,
		_w20011_,
		_w20012_
	);
	LUT4 #(
		.INIT('h5f4f)
	) name14186 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20013_
	);
	LUT4 #(
		.INIT('h5b4b)
	) name14187 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20014_
	);
	LUT4 #(
		.INIT('h0002)
	) name14188 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20015_
	);
	LUT4 #(
		.INIT('h3302)
	) name14189 (
		_w19928_,
		_w19935_,
		_w20014_,
		_w20015_,
		_w20016_
	);
	LUT4 #(
		.INIT('h1000)
	) name14190 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20017_
	);
	LUT3 #(
		.INIT('h08)
	) name14191 (
		_w19924_,
		_w19926_,
		_w19927_,
		_w20018_
	);
	LUT4 #(
		.INIT('h0020)
	) name14192 (
		_w19925_,
		_w19926_,
		_w19927_,
		_w19928_,
		_w20019_
	);
	LUT3 #(
		.INIT('h01)
	) name14193 (
		_w20017_,
		_w20018_,
		_w20019_,
		_w20020_
	);
	LUT4 #(
		.INIT('h0800)
	) name14194 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20021_
	);
	LUT4 #(
		.INIT('h0100)
	) name14195 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19928_,
		_w20022_
	);
	LUT2 #(
		.INIT('h1)
	) name14196 (
		_w20021_,
		_w20022_,
		_w20023_
	);
	LUT4 #(
		.INIT('he5be)
	) name14197 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20024_
	);
	LUT4 #(
		.INIT('h0004)
	) name14198 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20025_
	);
	LUT4 #(
		.INIT('hbffb)
	) name14199 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20026_
	);
	LUT4 #(
		.INIT('h0002)
	) name14200 (
		_w19924_,
		_w19926_,
		_w19928_,
		_w19935_,
		_w20027_
	);
	LUT4 #(
		.INIT('h00e4)
	) name14201 (
		_w19928_,
		_w20024_,
		_w20026_,
		_w20027_,
		_w20028_
	);
	LUT4 #(
		.INIT('hd500)
	) name14202 (
		_w19935_,
		_w20020_,
		_w20023_,
		_w20028_,
		_w20029_
	);
	LUT3 #(
		.INIT('h65)
	) name14203 (
		\u1_L6_reg[15]/P0001 ,
		_w20016_,
		_w20029_,
		_w20030_
	);
	LUT4 #(
		.INIT('h0400)
	) name14204 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20031_
	);
	LUT4 #(
		.INIT('hfb05)
	) name14205 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20032_
	);
	LUT4 #(
		.INIT('h00c1)
	) name14206 (
		_w19823_,
		_w19822_,
		_w19825_,
		_w19820_,
		_w20033_
	);
	LUT4 #(
		.INIT('h0200)
	) name14207 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20034_
	);
	LUT4 #(
		.INIT('h7d7f)
	) name14208 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20035_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14209 (
		_w19820_,
		_w20032_,
		_w20033_,
		_w20035_,
		_w20036_
	);
	LUT4 #(
		.INIT('hbbec)
	) name14210 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20037_
	);
	LUT3 #(
		.INIT('h6f)
	) name14211 (
		_w19823_,
		_w19824_,
		_w19825_,
		_w20038_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name14212 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20039_
	);
	LUT4 #(
		.INIT('he400)
	) name14213 (
		_w19820_,
		_w20037_,
		_w20038_,
		_w20039_,
		_w20040_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name14214 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20041_
	);
	LUT4 #(
		.INIT('h0f07)
	) name14215 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20042_
	);
	LUT3 #(
		.INIT('h02)
	) name14216 (
		_w19820_,
		_w20042_,
		_w20041_,
		_w20043_
	);
	LUT4 #(
		.INIT('h0e04)
	) name14217 (
		_w19821_,
		_w20040_,
		_w20043_,
		_w20036_,
		_w20044_
	);
	LUT2 #(
		.INIT('h9)
	) name14218 (
		\u1_L6_reg[17]/NET0131 ,
		_w20044_,
		_w20045_
	);
	LUT4 #(
		.INIT('h2100)
	) name14219 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w20046_
	);
	LUT2 #(
		.INIT('h1)
	) name14220 (
		_w19886_,
		_w20046_,
		_w20047_
	);
	LUT4 #(
		.INIT('hf3f1)
	) name14221 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w20048_
	);
	LUT2 #(
		.INIT('h2)
	) name14222 (
		_w19890_,
		_w20048_,
		_w20049_
	);
	LUT3 #(
		.INIT('h02)
	) name14223 (
		_w19886_,
		_w19902_,
		_w19950_,
		_w20050_
	);
	LUT3 #(
		.INIT('h45)
	) name14224 (
		_w20047_,
		_w20049_,
		_w20050_,
		_w20051_
	);
	LUT4 #(
		.INIT('h2500)
	) name14225 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w20052_
	);
	LUT4 #(
		.INIT('h080c)
	) name14226 (
		_w19892_,
		_w19885_,
		_w19886_,
		_w19888_,
		_w20053_
	);
	LUT4 #(
		.INIT('h080a)
	) name14227 (
		_w19890_,
		_w19958_,
		_w20052_,
		_w20053_,
		_w20054_
	);
	LUT3 #(
		.INIT('h08)
	) name14228 (
		_w19892_,
		_w19885_,
		_w19888_,
		_w20055_
	);
	LUT3 #(
		.INIT('h8a)
	) name14229 (
		_w19887_,
		_w19885_,
		_w19886_,
		_w20056_
	);
	LUT3 #(
		.INIT('h10)
	) name14230 (
		_w19901_,
		_w20055_,
		_w20056_,
		_w20057_
	);
	LUT4 #(
		.INIT('hfdee)
	) name14231 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w20058_
	);
	LUT4 #(
		.INIT('h0301)
	) name14232 (
		_w19886_,
		_w19890_,
		_w19913_,
		_w20058_,
		_w20059_
	);
	LUT3 #(
		.INIT('h45)
	) name14233 (
		_w20054_,
		_w20057_,
		_w20059_,
		_w20060_
	);
	LUT3 #(
		.INIT('h56)
	) name14234 (
		\u1_L6_reg[1]/NET0131 ,
		_w20051_,
		_w20060_,
		_w20061_
	);
	LUT3 #(
		.INIT('h08)
	) name14235 (
		_w19924_,
		_w19925_,
		_w19927_,
		_w20062_
	);
	LUT2 #(
		.INIT('h4)
	) name14236 (
		_w19926_,
		_w19928_,
		_w20063_
	);
	LUT2 #(
		.INIT('h2)
	) name14237 (
		_w20062_,
		_w20063_,
		_w20064_
	);
	LUT4 #(
		.INIT('h00bf)
	) name14238 (
		_w19924_,
		_w19926_,
		_w19927_,
		_w19935_,
		_w20065_
	);
	LUT4 #(
		.INIT('h0040)
	) name14239 (
		_w19924_,
		_w19925_,
		_w19927_,
		_w19928_,
		_w20066_
	);
	LUT2 #(
		.INIT('h2)
	) name14240 (
		_w19926_,
		_w19928_,
		_w20067_
	);
	LUT4 #(
		.INIT('h0010)
	) name14241 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19928_,
		_w20068_
	);
	LUT3 #(
		.INIT('h10)
	) name14242 (
		_w20066_,
		_w20068_,
		_w20065_,
		_w20069_
	);
	LUT4 #(
		.INIT('h0201)
	) name14243 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20070_
	);
	LUT4 #(
		.INIT('hd5df)
	) name14244 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20071_
	);
	LUT3 #(
		.INIT('h31)
	) name14245 (
		_w19928_,
		_w20070_,
		_w20071_,
		_w20072_
	);
	LUT3 #(
		.INIT('h40)
	) name14246 (
		_w20064_,
		_w20069_,
		_w20072_,
		_w20073_
	);
	LUT4 #(
		.INIT('hff02)
	) name14247 (
		_w19924_,
		_w19925_,
		_w19927_,
		_w19928_,
		_w20074_
	);
	LUT4 #(
		.INIT('hfd00)
	) name14248 (
		_w19925_,
		_w19926_,
		_w19927_,
		_w19928_,
		_w20075_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name14249 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20076_
	);
	LUT4 #(
		.INIT('h0eee)
	) name14250 (
		_w20021_,
		_w20074_,
		_w20075_,
		_w20076_,
		_w20077_
	);
	LUT4 #(
		.INIT('h2100)
	) name14251 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20078_
	);
	LUT3 #(
		.INIT('h02)
	) name14252 (
		_w19935_,
		_w20025_,
		_w20078_,
		_w20079_
	);
	LUT2 #(
		.INIT('h4)
	) name14253 (
		_w20077_,
		_w20079_,
		_w20080_
	);
	LUT4 #(
		.INIT('h0100)
	) name14254 (
		_w19924_,
		_w19926_,
		_w19927_,
		_w19928_,
		_w20081_
	);
	LUT3 #(
		.INIT('h07)
	) name14255 (
		_w20067_,
		_w20062_,
		_w20081_,
		_w20082_
	);
	LUT4 #(
		.INIT('ha955)
	) name14256 (
		\u1_L6_reg[21]/NET0131 ,
		_w20073_,
		_w20080_,
		_w20082_,
		_w20083_
	);
	LUT3 #(
		.INIT('hd0)
	) name14257 (
		_w19985_,
		_w19986_,
		_w19991_,
		_w20084_
	);
	LUT4 #(
		.INIT('h3301)
	) name14258 (
		_w19985_,
		_w19988_,
		_w19989_,
		_w19991_,
		_w20085_
	);
	LUT2 #(
		.INIT('h4)
	) name14259 (
		_w20084_,
		_w20085_,
		_w20086_
	);
	LUT2 #(
		.INIT('h4)
	) name14260 (
		_w19986_,
		_w19991_,
		_w20087_
	);
	LUT3 #(
		.INIT('h08)
	) name14261 (
		_w19985_,
		_w19988_,
		_w19989_,
		_w20088_
	);
	LUT4 #(
		.INIT('h0010)
	) name14262 (
		_w19985_,
		_w19986_,
		_w19989_,
		_w19991_,
		_w20089_
	);
	LUT4 #(
		.INIT('h0045)
	) name14263 (
		_w19984_,
		_w20087_,
		_w20088_,
		_w20089_,
		_w20090_
	);
	LUT4 #(
		.INIT('h00bf)
	) name14264 (
		_w19985_,
		_w19986_,
		_w19989_,
		_w19991_,
		_w20091_
	);
	LUT4 #(
		.INIT('h0131)
	) name14265 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20092_
	);
	LUT3 #(
		.INIT('h80)
	) name14266 (
		_w19985_,
		_w19986_,
		_w19989_,
		_w20093_
	);
	LUT4 #(
		.INIT('h7a00)
	) name14267 (
		_w19985_,
		_w19986_,
		_w19989_,
		_w19991_,
		_w20094_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14268 (
		_w19999_,
		_w20091_,
		_w20092_,
		_w20094_,
		_w20095_
	);
	LUT4 #(
		.INIT('h2000)
	) name14269 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20096_
	);
	LUT4 #(
		.INIT('hf700)
	) name14270 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19984_,
		_w20097_
	);
	LUT2 #(
		.INIT('h4)
	) name14271 (
		_w20096_,
		_w20097_,
		_w20098_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14272 (
		_w20086_,
		_w20090_,
		_w20095_,
		_w20098_,
		_w20099_
	);
	LUT4 #(
		.INIT('hdfeb)
	) name14273 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20100_
	);
	LUT4 #(
		.INIT('h0040)
	) name14274 (
		_w19985_,
		_w19988_,
		_w19989_,
		_w19991_,
		_w20101_
	);
	LUT4 #(
		.INIT('h0800)
	) name14275 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20102_
	);
	LUT4 #(
		.INIT('h0031)
	) name14276 (
		_w19991_,
		_w20101_,
		_w20100_,
		_w20102_,
		_w20103_
	);
	LUT3 #(
		.INIT('h65)
	) name14277 (
		\u1_L6_reg[25]/NET0131 ,
		_w20099_,
		_w20103_,
		_w20104_
	);
	LUT4 #(
		.INIT('h0092)
	) name14278 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w20105_
	);
	LUT3 #(
		.INIT('h8c)
	) name14279 (
		_w19887_,
		_w19892_,
		_w19888_,
		_w20106_
	);
	LUT2 #(
		.INIT('h1)
	) name14280 (
		_w19885_,
		_w19890_,
		_w20107_
	);
	LUT4 #(
		.INIT('h5150)
	) name14281 (
		_w19886_,
		_w20106_,
		_w20105_,
		_w20107_,
		_w20108_
	);
	LUT4 #(
		.INIT('h2010)
	) name14282 (
		_w19887_,
		_w19892_,
		_w19885_,
		_w19888_,
		_w20109_
	);
	LUT4 #(
		.INIT('h0f01)
	) name14283 (
		_w19887_,
		_w19885_,
		_w19886_,
		_w19888_,
		_w20110_
	);
	LUT2 #(
		.INIT('h8)
	) name14284 (
		_w20106_,
		_w20110_,
		_w20111_
	);
	LUT3 #(
		.INIT('h40)
	) name14285 (
		_w19887_,
		_w19892_,
		_w19888_,
		_w20112_
	);
	LUT4 #(
		.INIT('h2022)
	) name14286 (
		_w19890_,
		_w19896_,
		_w19906_,
		_w20112_,
		_w20113_
	);
	LUT3 #(
		.INIT('h10)
	) name14287 (
		_w20111_,
		_w20109_,
		_w20113_,
		_w20114_
	);
	LUT3 #(
		.INIT('h80)
	) name14288 (
		_w19885_,
		_w19886_,
		_w19888_,
		_w20115_
	);
	LUT2 #(
		.INIT('h4)
	) name14289 (
		_w19914_,
		_w20115_,
		_w20116_
	);
	LUT4 #(
		.INIT('h00fd)
	) name14290 (
		_w19887_,
		_w19885_,
		_w19888_,
		_w19890_,
		_w20117_
	);
	LUT3 #(
		.INIT('h10)
	) name14291 (
		_w19912_,
		_w19913_,
		_w20117_,
		_w20118_
	);
	LUT2 #(
		.INIT('h4)
	) name14292 (
		_w20116_,
		_w20118_,
		_w20119_
	);
	LUT2 #(
		.INIT('h4)
	) name14293 (
		_w19910_,
		_w19956_,
		_w20120_
	);
	LUT4 #(
		.INIT('h000e)
	) name14294 (
		_w20114_,
		_w20119_,
		_w20120_,
		_w20108_,
		_w20121_
	);
	LUT2 #(
		.INIT('h9)
	) name14295 (
		\u1_L6_reg[26]/NET0131 ,
		_w20121_,
		_w20122_
	);
	LUT4 #(
		.INIT('hc693)
	) name14296 (
		decrypt_pad,
		\u1_R6_reg[8]/NET0131 ,
		\u1_uk_K_r6_reg[48]/NET0131 ,
		\u1_uk_K_r6_reg[55]/P0001 ,
		_w20123_
	);
	LUT4 #(
		.INIT('hc693)
	) name14297 (
		decrypt_pad,
		\u1_R6_reg[7]/NET0131 ,
		\u1_uk_K_r6_reg[25]/NET0131 ,
		\u1_uk_K_r6_reg[32]/NET0131 ,
		_w20124_
	);
	LUT4 #(
		.INIT('hc693)
	) name14298 (
		decrypt_pad,
		\u1_R6_reg[5]/NET0131 ,
		\u1_uk_K_r6_reg[40]/NET0131 ,
		\u1_uk_K_r6_reg[47]/NET0131 ,
		_w20125_
	);
	LUT4 #(
		.INIT('hc963)
	) name14299 (
		decrypt_pad,
		\u1_R6_reg[4]/NET0131 ,
		\u1_uk_K_r6_reg[11]/NET0131 ,
		\u1_uk_K_r6_reg[4]/NET0131 ,
		_w20126_
	);
	LUT4 #(
		.INIT('hc963)
	) name14300 (
		decrypt_pad,
		\u1_R6_reg[9]/NET0131 ,
		\u1_uk_K_r6_reg[3]/NET0131 ,
		\u1_uk_K_r6_reg[53]/NET0131 ,
		_w20127_
	);
	LUT4 #(
		.INIT('hc963)
	) name14301 (
		decrypt_pad,
		\u1_R6_reg[6]/NET0131 ,
		\u1_uk_K_r6_reg[13]/NET0131 ,
		\u1_uk_K_r6_reg[6]/NET0131 ,
		_w20128_
	);
	LUT4 #(
		.INIT('h5fa7)
	) name14302 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20129_
	);
	LUT2 #(
		.INIT('h2)
	) name14303 (
		_w20124_,
		_w20129_,
		_w20130_
	);
	LUT4 #(
		.INIT('hf5fc)
	) name14304 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20131_
	);
	LUT2 #(
		.INIT('h1)
	) name14305 (
		_w20124_,
		_w20131_,
		_w20132_
	);
	LUT2 #(
		.INIT('h4)
	) name14306 (
		_w20128_,
		_w20126_,
		_w20133_
	);
	LUT4 #(
		.INIT('h00bf)
	) name14307 (
		_w20125_,
		_w20126_,
		_w20127_,
		_w20124_,
		_w20134_
	);
	LUT4 #(
		.INIT('h0400)
	) name14308 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20135_
	);
	LUT3 #(
		.INIT('h0d)
	) name14309 (
		_w20133_,
		_w20134_,
		_w20135_,
		_w20136_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name14310 (
		_w20123_,
		_w20132_,
		_w20130_,
		_w20136_,
		_w20137_
	);
	LUT4 #(
		.INIT('hfb7b)
	) name14311 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20138_
	);
	LUT2 #(
		.INIT('h1)
	) name14312 (
		_w20138_,
		_w20124_,
		_w20139_
	);
	LUT4 #(
		.INIT('h5a4f)
	) name14313 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20140_
	);
	LUT4 #(
		.INIT('h4084)
	) name14314 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20141_
	);
	LUT4 #(
		.INIT('h3120)
	) name14315 (
		_w20124_,
		_w20141_,
		_w20131_,
		_w20140_,
		_w20142_
	);
	LUT3 #(
		.INIT('h54)
	) name14316 (
		_w20139_,
		_w20123_,
		_w20142_,
		_w20143_
	);
	LUT3 #(
		.INIT('h65)
	) name14317 (
		\u1_L6_reg[28]/NET0131 ,
		_w20137_,
		_w20143_,
		_w20144_
	);
	LUT4 #(
		.INIT('h779a)
	) name14318 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20145_
	);
	LUT4 #(
		.INIT('h0e02)
	) name14319 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20146_
	);
	LUT4 #(
		.INIT('hf17d)
	) name14320 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20147_
	);
	LUT4 #(
		.INIT('h1000)
	) name14321 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20148_
	);
	LUT4 #(
		.INIT('h00e4)
	) name14322 (
		_w19852_,
		_w20147_,
		_w20145_,
		_w20148_,
		_w20149_
	);
	LUT2 #(
		.INIT('h1)
	) name14323 (
		_w19851_,
		_w20149_,
		_w20150_
	);
	LUT4 #(
		.INIT('hdd7d)
	) name14324 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20151_
	);
	LUT2 #(
		.INIT('h2)
	) name14325 (
		_w19852_,
		_w20151_,
		_w20152_
	);
	LUT3 #(
		.INIT('h48)
	) name14326 (
		_w19854_,
		_w19855_,
		_w19856_,
		_w20153_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name14327 (
		_w19853_,
		_w19855_,
		_w19852_,
		_w19856_,
		_w20154_
	);
	LUT3 #(
		.INIT('h01)
	) name14328 (
		_w20146_,
		_w20154_,
		_w20153_,
		_w20155_
	);
	LUT4 #(
		.INIT('h0004)
	) name14329 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20156_
	);
	LUT4 #(
		.INIT('h2000)
	) name14330 (
		_w19853_,
		_w19855_,
		_w19852_,
		_w19856_,
		_w20157_
	);
	LUT2 #(
		.INIT('h1)
	) name14331 (
		_w20156_,
		_w20157_,
		_w20158_
	);
	LUT4 #(
		.INIT('h5700)
	) name14332 (
		_w19851_,
		_w20152_,
		_w20155_,
		_w20158_,
		_w20159_
	);
	LUT3 #(
		.INIT('h9a)
	) name14333 (
		\u1_L6_reg[29]/NET0131 ,
		_w20150_,
		_w20159_,
		_w20160_
	);
	LUT4 #(
		.INIT('h0122)
	) name14334 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20161_
	);
	LUT2 #(
		.INIT('h1)
	) name14335 (
		_w20124_,
		_w20123_,
		_w20162_
	);
	LUT4 #(
		.INIT('h4000)
	) name14336 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20163_
	);
	LUT4 #(
		.INIT('h0103)
	) name14337 (
		_w20124_,
		_w20123_,
		_w20161_,
		_w20163_,
		_w20164_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name14338 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20165_
	);
	LUT4 #(
		.INIT('h0800)
	) name14339 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20166_
	);
	LUT4 #(
		.INIT('h0010)
	) name14340 (
		_w20125_,
		_w20128_,
		_w20127_,
		_w20124_,
		_w20167_
	);
	LUT4 #(
		.INIT('h000d)
	) name14341 (
		_w20134_,
		_w20165_,
		_w20166_,
		_w20167_,
		_w20168_
	);
	LUT4 #(
		.INIT('h2010)
	) name14342 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20169_
	);
	LUT2 #(
		.INIT('h2)
	) name14343 (
		_w20125_,
		_w20128_,
		_w20170_
	);
	LUT4 #(
		.INIT('ha200)
	) name14344 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20124_,
		_w20171_
	);
	LUT3 #(
		.INIT('h02)
	) name14345 (
		_w20123_,
		_w20171_,
		_w20169_,
		_w20172_
	);
	LUT3 #(
		.INIT('h07)
	) name14346 (
		_w20164_,
		_w20168_,
		_w20172_,
		_w20173_
	);
	LUT4 #(
		.INIT('hbff0)
	) name14347 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20174_
	);
	LUT4 #(
		.INIT('h0b00)
	) name14348 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20175_
	);
	LUT4 #(
		.INIT('h3302)
	) name14349 (
		_w20123_,
		_w20170_,
		_w20174_,
		_w20175_,
		_w20176_
	);
	LUT4 #(
		.INIT('h0004)
	) name14350 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20177_
	);
	LUT4 #(
		.INIT('hdf00)
	) name14351 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20124_,
		_w20178_
	);
	LUT2 #(
		.INIT('h4)
	) name14352 (
		_w20177_,
		_w20178_,
		_w20179_
	);
	LUT3 #(
		.INIT('h0e)
	) name14353 (
		_w20124_,
		_w20176_,
		_w20179_,
		_w20180_
	);
	LUT3 #(
		.INIT('h56)
	) name14354 (
		\u1_L6_reg[2]/NET0131 ,
		_w20173_,
		_w20180_,
		_w20181_
	);
	LUT4 #(
		.INIT('h2000)
	) name14355 (
		_w19854_,
		_w19855_,
		_w19852_,
		_w19856_,
		_w20182_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14356 (
		_w19853_,
		_w19855_,
		_w19856_,
		_w19851_,
		_w20183_
	);
	LUT2 #(
		.INIT('h4)
	) name14357 (
		_w20182_,
		_w20183_,
		_w20184_
	);
	LUT3 #(
		.INIT('h51)
	) name14358 (
		_w19879_,
		_w19863_,
		_w19857_,
		_w20185_
	);
	LUT4 #(
		.INIT('hf070)
	) name14359 (
		_w19853_,
		_w19854_,
		_w19852_,
		_w19856_,
		_w20186_
	);
	LUT4 #(
		.INIT('hbcff)
	) name14360 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20187_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name14361 (
		_w19853_,
		_w19854_,
		_w19852_,
		_w19856_,
		_w20188_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name14362 (
		_w20148_,
		_w20186_,
		_w20187_,
		_w20188_,
		_w20189_
	);
	LUT3 #(
		.INIT('h01)
	) name14363 (
		_w19851_,
		_w19864_,
		_w20156_,
		_w20190_
	);
	LUT4 #(
		.INIT('h7077)
	) name14364 (
		_w20184_,
		_w20185_,
		_w20189_,
		_w20190_,
		_w20191_
	);
	LUT3 #(
		.INIT('h31)
	) name14365 (
		_w19853_,
		_w19854_,
		_w19856_,
		_w20192_
	);
	LUT4 #(
		.INIT('hd060)
	) name14366 (
		_w19853_,
		_w19854_,
		_w19852_,
		_w19856_,
		_w20193_
	);
	LUT4 #(
		.INIT('h070b)
	) name14367 (
		_w19853_,
		_w19854_,
		_w19852_,
		_w19856_,
		_w20194_
	);
	LUT4 #(
		.INIT('h3331)
	) name14368 (
		_w19855_,
		_w19881_,
		_w20194_,
		_w20193_,
		_w20195_
	);
	LUT3 #(
		.INIT('h65)
	) name14369 (
		\u1_L6_reg[4]/NET0131 ,
		_w20191_,
		_w20195_,
		_w20196_
	);
	LUT4 #(
		.INIT('h0201)
	) name14370 (
		_w19853_,
		_w19854_,
		_w19852_,
		_w19856_,
		_w20197_
	);
	LUT4 #(
		.INIT('hf700)
	) name14371 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19852_,
		_w20198_
	);
	LUT4 #(
		.INIT('h8000)
	) name14372 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20199_
	);
	LUT4 #(
		.INIT('h0045)
	) name14373 (
		_w19851_,
		_w20192_,
		_w20198_,
		_w20199_,
		_w20200_
	);
	LUT4 #(
		.INIT('h2010)
	) name14374 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20201_
	);
	LUT3 #(
		.INIT('h04)
	) name14375 (
		_w19868_,
		_w19851_,
		_w20201_,
		_w20202_
	);
	LUT4 #(
		.INIT('h010a)
	) name14376 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19856_,
		_w20203_
	);
	LUT4 #(
		.INIT('h0844)
	) name14377 (
		_w19853_,
		_w19854_,
		_w19855_,
		_w19852_,
		_w20204_
	);
	LUT2 #(
		.INIT('h1)
	) name14378 (
		_w20203_,
		_w20204_,
		_w20205_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name14379 (
		_w20197_,
		_w20200_,
		_w20202_,
		_w20205_,
		_w20206_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name14380 (
		_w19853_,
		_w19855_,
		_w19877_,
		_w19864_,
		_w20207_
	);
	LUT3 #(
		.INIT('h65)
	) name14381 (
		\u1_L6_reg[19]/NET0131 ,
		_w20206_,
		_w20207_,
		_w20208_
	);
	LUT4 #(
		.INIT('hef99)
	) name14382 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20209_
	);
	LUT4 #(
		.INIT('h7dfb)
	) name14383 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20210_
	);
	LUT4 #(
		.INIT('h0233)
	) name14384 (
		_w19821_,
		_w19820_,
		_w20209_,
		_w20210_,
		_w20211_
	);
	LUT4 #(
		.INIT('h1554)
	) name14385 (
		_w19821_,
		_w19823_,
		_w19824_,
		_w19822_,
		_w20212_
	);
	LUT3 #(
		.INIT('h15)
	) name14386 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w20213_
	);
	LUT3 #(
		.INIT('h1d)
	) name14387 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w20214_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name14388 (
		_w19825_,
		_w19820_,
		_w20213_,
		_w20214_,
		_w20215_
	);
	LUT2 #(
		.INIT('h4)
	) name14389 (
		_w19846_,
		_w19839_,
		_w20216_
	);
	LUT4 #(
		.INIT('h002a)
	) name14390 (
		_w19821_,
		_w19829_,
		_w19845_,
		_w20031_,
		_w20217_
	);
	LUT4 #(
		.INIT('h7077)
	) name14391 (
		_w20212_,
		_w20215_,
		_w20216_,
		_w20217_,
		_w20218_
	);
	LUT3 #(
		.INIT('h13)
	) name14392 (
		_w19832_,
		_w19847_,
		_w19842_,
		_w20219_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name14393 (
		\u1_L6_reg[23]/NET0131 ,
		_w20218_,
		_w20211_,
		_w20219_,
		_w20220_
	);
	LUT4 #(
		.INIT('h9f9a)
	) name14394 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20221_
	);
	LUT2 #(
		.INIT('h1)
	) name14395 (
		_w19928_,
		_w20221_,
		_w20222_
	);
	LUT3 #(
		.INIT('hd0)
	) name14396 (
		_w19924_,
		_w19925_,
		_w19928_,
		_w20223_
	);
	LUT4 #(
		.INIT('hbdf3)
	) name14397 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20224_
	);
	LUT3 #(
		.INIT('hb0)
	) name14398 (
		_w20013_,
		_w20223_,
		_w20224_,
		_w20225_
	);
	LUT3 #(
		.INIT('h8a)
	) name14399 (
		_w19935_,
		_w20222_,
		_w20225_,
		_w20226_
	);
	LUT4 #(
		.INIT('hfb00)
	) name14400 (
		_w19925_,
		_w19926_,
		_w19927_,
		_w19928_,
		_w20227_
	);
	LUT4 #(
		.INIT('h23f3)
	) name14401 (
		_w19924_,
		_w19925_,
		_w19926_,
		_w19927_,
		_w20228_
	);
	LUT2 #(
		.INIT('h8)
	) name14402 (
		_w20227_,
		_w20228_,
		_w20229_
	);
	LUT4 #(
		.INIT('h0080)
	) name14403 (
		_w19924_,
		_w19925_,
		_w19927_,
		_w19928_,
		_w20230_
	);
	LUT3 #(
		.INIT('h01)
	) name14404 (
		_w19946_,
		_w20068_,
		_w20230_,
		_w20231_
	);
	LUT4 #(
		.INIT('h1000)
	) name14405 (
		_w19925_,
		_w19926_,
		_w19927_,
		_w19928_,
		_w20232_
	);
	LUT4 #(
		.INIT('h00ab)
	) name14406 (
		_w19928_,
		_w19938_,
		_w19945_,
		_w20232_,
		_w20233_
	);
	LUT4 #(
		.INIT('hba00)
	) name14407 (
		_w19935_,
		_w20229_,
		_w20231_,
		_w20233_,
		_w20234_
	);
	LUT3 #(
		.INIT('h65)
	) name14408 (
		\u1_L6_reg[27]/NET0131 ,
		_w20226_,
		_w20234_,
		_w20235_
	);
	LUT2 #(
		.INIT('h9)
	) name14409 (
		_w19792_,
		_w19794_,
		_w20236_
	);
	LUT4 #(
		.INIT('hd003)
	) name14410 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w20237_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name14411 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w20238_
	);
	LUT3 #(
		.INIT('h01)
	) name14412 (
		_w19795_,
		_w20238_,
		_w20237_,
		_w20239_
	);
	LUT4 #(
		.INIT('h0800)
	) name14413 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w20240_
	);
	LUT4 #(
		.INIT('hb5bc)
	) name14414 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w20241_
	);
	LUT3 #(
		.INIT('h31)
	) name14415 (
		_w19795_,
		_w20240_,
		_w20241_,
		_w20242_
	);
	LUT3 #(
		.INIT('h8a)
	) name14416 (
		_w19789_,
		_w20239_,
		_w20242_,
		_w20243_
	);
	LUT3 #(
		.INIT('h40)
	) name14417 (
		_w19791_,
		_w19792_,
		_w19794_,
		_w20244_
	);
	LUT4 #(
		.INIT('hab89)
	) name14418 (
		_w19795_,
		_w19971_,
		_w19973_,
		_w20244_,
		_w20245_
	);
	LUT4 #(
		.INIT('h7bd7)
	) name14419 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w20246_
	);
	LUT4 #(
		.INIT('h00c8)
	) name14420 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19795_,
		_w20247_
	);
	LUT4 #(
		.INIT('h135f)
	) name14421 (
		_w19795_,
		_w19810_,
		_w19802_,
		_w20247_,
		_w20248_
	);
	LUT4 #(
		.INIT('hba00)
	) name14422 (
		_w19789_,
		_w20245_,
		_w20246_,
		_w20248_,
		_w20249_
	);
	LUT3 #(
		.INIT('h65)
	) name14423 (
		\u1_L6_reg[32]/NET0131 ,
		_w20243_,
		_w20249_,
		_w20250_
	);
	LUT4 #(
		.INIT('hc693)
	) name14424 (
		decrypt_pad,
		\u1_R6_reg[13]/NET0131 ,
		\u1_uk_K_r6_reg[39]/NET0131 ,
		\u1_uk_K_r6_reg[46]/NET0131 ,
		_w20251_
	);
	LUT4 #(
		.INIT('hc693)
	) name14425 (
		decrypt_pad,
		\u1_R6_reg[9]/NET0131 ,
		\u1_uk_K_r6_reg[34]/NET0131 ,
		\u1_uk_K_r6_reg[41]/NET0131 ,
		_w20252_
	);
	LUT4 #(
		.INIT('hc693)
	) name14426 (
		decrypt_pad,
		\u1_R6_reg[11]/NET0131 ,
		\u1_uk_K_r6_reg[11]/NET0131 ,
		\u1_uk_K_r6_reg[18]/NET0131 ,
		_w20253_
	);
	LUT3 #(
		.INIT('h0b)
	) name14427 (
		_w20251_,
		_w20252_,
		_w20253_,
		_w20254_
	);
	LUT4 #(
		.INIT('hc693)
	) name14428 (
		decrypt_pad,
		\u1_R6_reg[10]/NET0131 ,
		\u1_uk_K_r6_reg[10]/NET0131 ,
		\u1_uk_K_r6_reg[17]/NET0131 ,
		_w20255_
	);
	LUT4 #(
		.INIT('hc963)
	) name14429 (
		decrypt_pad,
		\u1_R6_reg[8]/NET0131 ,
		\u1_uk_K_r6_reg[12]/NET0131 ,
		\u1_uk_K_r6_reg[5]/NET0131 ,
		_w20256_
	);
	LUT4 #(
		.INIT('h30bb)
	) name14430 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20257_
	);
	LUT4 #(
		.INIT('h1000)
	) name14431 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20258_
	);
	LUT4 #(
		.INIT('hc693)
	) name14432 (
		decrypt_pad,
		\u1_R6_reg[12]/NET0131 ,
		\u1_uk_K_r6_reg[26]/NET0131 ,
		\u1_uk_K_r6_reg[33]/NET0131 ,
		_w20259_
	);
	LUT4 #(
		.INIT('h5100)
	) name14433 (
		_w20258_,
		_w20254_,
		_w20257_,
		_w20259_,
		_w20260_
	);
	LUT2 #(
		.INIT('h9)
	) name14434 (
		_w20255_,
		_w20252_,
		_w20261_
	);
	LUT3 #(
		.INIT('h46)
	) name14435 (
		_w20251_,
		_w20256_,
		_w20253_,
		_w20262_
	);
	LUT2 #(
		.INIT('h8)
	) name14436 (
		_w20261_,
		_w20262_,
		_w20263_
	);
	LUT4 #(
		.INIT('h0990)
	) name14437 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20264_
	);
	LUT4 #(
		.INIT('h1000)
	) name14438 (
		_w20256_,
		_w20255_,
		_w20252_,
		_w20253_,
		_w20265_
	);
	LUT3 #(
		.INIT('h01)
	) name14439 (
		_w20259_,
		_w20265_,
		_w20264_,
		_w20266_
	);
	LUT2 #(
		.INIT('h2)
	) name14440 (
		_w20251_,
		_w20256_,
		_w20267_
	);
	LUT4 #(
		.INIT('h9b55)
	) name14441 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20268_
	);
	LUT4 #(
		.INIT('h0001)
	) name14442 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20269_
	);
	LUT4 #(
		.INIT('hff5e)
	) name14443 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20270_
	);
	LUT4 #(
		.INIT('h08aa)
	) name14444 (
		_w20253_,
		_w20259_,
		_w20268_,
		_w20270_,
		_w20271_
	);
	LUT4 #(
		.INIT('h00ba)
	) name14445 (
		_w20260_,
		_w20263_,
		_w20266_,
		_w20271_,
		_w20272_
	);
	LUT2 #(
		.INIT('h9)
	) name14446 (
		\u1_L6_reg[6]/NET0131 ,
		_w20272_,
		_w20273_
	);
	LUT4 #(
		.INIT('hf126)
	) name14447 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w20274_
	);
	LUT4 #(
		.INIT('h2880)
	) name14448 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w20275_
	);
	LUT4 #(
		.INIT('h5004)
	) name14449 (
		_w19790_,
		_w19791_,
		_w19792_,
		_w19794_,
		_w20276_
	);
	LUT4 #(
		.INIT('h1302)
	) name14450 (
		_w19795_,
		_w20275_,
		_w20276_,
		_w20274_,
		_w20277_
	);
	LUT2 #(
		.INIT('h2)
	) name14451 (
		_w19789_,
		_w20277_,
		_w20278_
	);
	LUT2 #(
		.INIT('h4)
	) name14452 (
		_w19795_,
		_w20275_,
		_w20279_
	);
	LUT2 #(
		.INIT('h2)
	) name14453 (
		_w19789_,
		_w19795_,
		_w20280_
	);
	LUT3 #(
		.INIT('h4c)
	) name14454 (
		_w19791_,
		_w19792_,
		_w19794_,
		_w20281_
	);
	LUT4 #(
		.INIT('h8a00)
	) name14455 (
		_w19790_,
		_w19792_,
		_w19794_,
		_w19795_,
		_w20282_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name14456 (
		_w19796_,
		_w20236_,
		_w20281_,
		_w20282_,
		_w20283_
	);
	LUT3 #(
		.INIT('h45)
	) name14457 (
		_w19809_,
		_w19795_,
		_w20276_,
		_w20284_
	);
	LUT4 #(
		.INIT('h0133)
	) name14458 (
		_w19789_,
		_w20280_,
		_w20283_,
		_w20284_,
		_w20285_
	);
	LUT4 #(
		.INIT('h5556)
	) name14459 (
		\u1_L6_reg[7]/NET0131 ,
		_w20279_,
		_w20285_,
		_w20278_,
		_w20286_
	);
	LUT4 #(
		.INIT('h008c)
	) name14460 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20287_
	);
	LUT2 #(
		.INIT('h2)
	) name14461 (
		_w20091_,
		_w20287_,
		_w20288_
	);
	LUT4 #(
		.INIT('h0100)
	) name14462 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20289_
	);
	LUT3 #(
		.INIT('h02)
	) name14463 (
		_w19991_,
		_w20093_,
		_w20289_,
		_w20290_
	);
	LUT4 #(
		.INIT('hdfe5)
	) name14464 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20291_
	);
	LUT4 #(
		.INIT('h0155)
	) name14465 (
		_w19984_,
		_w20288_,
		_w20290_,
		_w20291_,
		_w20292_
	);
	LUT4 #(
		.INIT('h0001)
	) name14466 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20293_
	);
	LUT4 #(
		.INIT('hbf00)
	) name14467 (
		_w19985_,
		_w19986_,
		_w19989_,
		_w19991_,
		_w20294_
	);
	LUT4 #(
		.INIT('h4544)
	) name14468 (
		_w20007_,
		_w20003_,
		_w20293_,
		_w20294_,
		_w20295_
	);
	LUT4 #(
		.INIT('hdf97)
	) name14469 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20296_
	);
	LUT4 #(
		.INIT('h5f13)
	) name14470 (
		_w19988_,
		_w19991_,
		_w20089_,
		_w20296_,
		_w20297_
	);
	LUT3 #(
		.INIT('hd0)
	) name14471 (
		_w19984_,
		_w20295_,
		_w20297_,
		_w20298_
	);
	LUT3 #(
		.INIT('h65)
	) name14472 (
		\u1_L6_reg[8]/NET0131 ,
		_w20292_,
		_w20298_,
		_w20299_
	);
	LUT3 #(
		.INIT('h78)
	) name14473 (
		_w20251_,
		_w20256_,
		_w20252_,
		_w20300_
	);
	LUT4 #(
		.INIT('h6979)
	) name14474 (
		_w20251_,
		_w20256_,
		_w20252_,
		_w20253_,
		_w20301_
	);
	LUT4 #(
		.INIT('h2000)
	) name14475 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20302_
	);
	LUT4 #(
		.INIT('h0014)
	) name14476 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20253_,
		_w20303_
	);
	LUT4 #(
		.INIT('h0032)
	) name14477 (
		_w20255_,
		_w20302_,
		_w20301_,
		_w20303_,
		_w20304_
	);
	LUT4 #(
		.INIT('h76dc)
	) name14478 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20305_
	);
	LUT4 #(
		.INIT('h6800)
	) name14479 (
		_w20251_,
		_w20256_,
		_w20252_,
		_w20253_,
		_w20306_
	);
	LUT4 #(
		.INIT('h00f2)
	) name14480 (
		_w20253_,
		_w20269_,
		_w20305_,
		_w20306_,
		_w20307_
	);
	LUT4 #(
		.INIT('h0008)
	) name14481 (
		_w20256_,
		_w20255_,
		_w20252_,
		_w20253_,
		_w20308_
	);
	LUT3 #(
		.INIT('hbe)
	) name14482 (
		_w20251_,
		_w20256_,
		_w20252_,
		_w20309_
	);
	LUT2 #(
		.INIT('h8)
	) name14483 (
		_w20255_,
		_w20253_,
		_w20310_
	);
	LUT3 #(
		.INIT('h45)
	) name14484 (
		_w20308_,
		_w20309_,
		_w20310_,
		_w20311_
	);
	LUT4 #(
		.INIT('hd800)
	) name14485 (
		_w20259_,
		_w20304_,
		_w20307_,
		_w20311_,
		_w20312_
	);
	LUT2 #(
		.INIT('h9)
	) name14486 (
		\u1_L6_reg[16]/NET0131 ,
		_w20312_,
		_w20313_
	);
	LUT2 #(
		.INIT('h1)
	) name14487 (
		_w20255_,
		_w20252_,
		_w20314_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name14488 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20315_
	);
	LUT3 #(
		.INIT('he0)
	) name14489 (
		_w20255_,
		_w20252_,
		_w20253_,
		_w20316_
	);
	LUT4 #(
		.INIT('h0302)
	) name14490 (
		_w20253_,
		_w20267_,
		_w20316_,
		_w20315_,
		_w20317_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name14491 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20318_
	);
	LUT4 #(
		.INIT('h3f15)
	) name14492 (
		_w20253_,
		_w20262_,
		_w20314_,
		_w20318_,
		_w20319_
	);
	LUT3 #(
		.INIT('hed)
	) name14493 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20320_
	);
	LUT4 #(
		.INIT('hec2d)
	) name14494 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20321_
	);
	LUT4 #(
		.INIT('h0040)
	) name14495 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20322_
	);
	LUT4 #(
		.INIT('h0031)
	) name14496 (
		_w20253_,
		_w20259_,
		_w20321_,
		_w20322_,
		_w20323_
	);
	LUT4 #(
		.INIT('h00df)
	) name14497 (
		_w20259_,
		_w20317_,
		_w20319_,
		_w20323_,
		_w20324_
	);
	LUT4 #(
		.INIT('h9bd6)
	) name14498 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20325_
	);
	LUT4 #(
		.INIT('h8000)
	) name14499 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20326_
	);
	LUT4 #(
		.INIT('h5501)
	) name14500 (
		_w20253_,
		_w20259_,
		_w20325_,
		_w20326_,
		_w20327_
	);
	LUT4 #(
		.INIT('h0004)
	) name14501 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20328_
	);
	LUT4 #(
		.INIT('h135f)
	) name14502 (
		_w20251_,
		_w20253_,
		_w20265_,
		_w20328_,
		_w20329_
	);
	LUT2 #(
		.INIT('h4)
	) name14503 (
		_w20327_,
		_w20329_,
		_w20330_
	);
	LUT3 #(
		.INIT('h65)
	) name14504 (
		\u1_L6_reg[24]/NET0131 ,
		_w20324_,
		_w20330_,
		_w20331_
	);
	LUT3 #(
		.INIT('h20)
	) name14505 (
		_w20259_,
		_w20328_,
		_w20320_,
		_w20332_
	);
	LUT3 #(
		.INIT('h10)
	) name14506 (
		_w20251_,
		_w20255_,
		_w20252_,
		_w20333_
	);
	LUT4 #(
		.INIT('h80c0)
	) name14507 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20334_
	);
	LUT4 #(
		.INIT('haaa8)
	) name14508 (
		_w20253_,
		_w20259_,
		_w20334_,
		_w20333_,
		_w20335_
	);
	LUT2 #(
		.INIT('h4)
	) name14509 (
		_w20332_,
		_w20335_,
		_w20336_
	);
	LUT3 #(
		.INIT('h72)
	) name14510 (
		_w20256_,
		_w20255_,
		_w20252_,
		_w20337_
	);
	LUT4 #(
		.INIT('hffd6)
	) name14511 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20338_
	);
	LUT4 #(
		.INIT('h2033)
	) name14512 (
		_w20254_,
		_w20259_,
		_w20337_,
		_w20338_,
		_w20339_
	);
	LUT4 #(
		.INIT('h0072)
	) name14513 (
		_w20251_,
		_w20256_,
		_w20253_,
		_w20259_,
		_w20340_
	);
	LUT4 #(
		.INIT('hf070)
	) name14514 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20253_,
		_w20341_
	);
	LUT3 #(
		.INIT('h20)
	) name14515 (
		_w20300_,
		_w20340_,
		_w20341_,
		_w20342_
	);
	LUT4 #(
		.INIT('h2e3f)
	) name14516 (
		_w20251_,
		_w20256_,
		_w20255_,
		_w20252_,
		_w20343_
	);
	LUT2 #(
		.INIT('h4)
	) name14517 (
		_w20253_,
		_w20259_,
		_w20344_
	);
	LUT2 #(
		.INIT('h4)
	) name14518 (
		_w20343_,
		_w20344_,
		_w20345_
	);
	LUT3 #(
		.INIT('h01)
	) name14519 (
		_w20339_,
		_w20342_,
		_w20345_,
		_w20346_
	);
	LUT3 #(
		.INIT('h9a)
	) name14520 (
		\u1_L6_reg[30]/NET0131 ,
		_w20336_,
		_w20346_,
		_w20347_
	);
	LUT3 #(
		.INIT('h08)
	) name14521 (
		_w19985_,
		_w19986_,
		_w19989_,
		_w20348_
	);
	LUT4 #(
		.INIT('h0002)
	) name14522 (
		_w19984_,
		_w20004_,
		_w20102_,
		_w20348_,
		_w20349_
	);
	LUT4 #(
		.INIT('h4050)
	) name14523 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20350_
	);
	LUT4 #(
		.INIT('h3b0c)
	) name14524 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20351_
	);
	LUT3 #(
		.INIT('h10)
	) name14525 (
		_w19984_,
		_w20350_,
		_w20351_,
		_w20352_
	);
	LUT4 #(
		.INIT('h4000)
	) name14526 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20353_
	);
	LUT4 #(
		.INIT('h0001)
	) name14527 (
		_w19991_,
		_w20008_,
		_w20293_,
		_w20353_,
		_w20354_
	);
	LUT3 #(
		.INIT('he0)
	) name14528 (
		_w20349_,
		_w20352_,
		_w20354_,
		_w20355_
	);
	LUT4 #(
		.INIT('h0c22)
	) name14529 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20356_
	);
	LUT4 #(
		.INIT('h0002)
	) name14530 (
		_w19984_,
		_w20004_,
		_w20102_,
		_w20356_,
		_w20357_
	);
	LUT4 #(
		.INIT('hddf3)
	) name14531 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20358_
	);
	LUT3 #(
		.INIT('h10)
	) name14532 (
		_w19984_,
		_w20350_,
		_w20358_,
		_w20359_
	);
	LUT4 #(
		.INIT('h0040)
	) name14533 (
		_w19985_,
		_w19986_,
		_w19988_,
		_w19989_,
		_w20360_
	);
	LUT3 #(
		.INIT('h02)
	) name14534 (
		_w19991_,
		_w20289_,
		_w20360_,
		_w20361_
	);
	LUT3 #(
		.INIT('he0)
	) name14535 (
		_w20357_,
		_w20359_,
		_w20361_,
		_w20362_
	);
	LUT3 #(
		.INIT('ha9)
	) name14536 (
		\u1_L6_reg[3]/NET0131 ,
		_w20355_,
		_w20362_,
		_w20363_
	);
	LUT4 #(
		.INIT('h9b99)
	) name14537 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20364_
	);
	LUT2 #(
		.INIT('h2)
	) name14538 (
		_w19820_,
		_w20364_,
		_w20365_
	);
	LUT4 #(
		.INIT('h4010)
	) name14539 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20366_
	);
	LUT3 #(
		.INIT('he6)
	) name14540 (
		_w19823_,
		_w19824_,
		_w19825_,
		_w20367_
	);
	LUT4 #(
		.INIT('h0019)
	) name14541 (
		_w19823_,
		_w19824_,
		_w19825_,
		_w19820_,
		_w20368_
	);
	LUT4 #(
		.INIT('h0800)
	) name14542 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20369_
	);
	LUT3 #(
		.INIT('h01)
	) name14543 (
		_w20368_,
		_w20366_,
		_w20369_,
		_w20370_
	);
	LUT3 #(
		.INIT('h45)
	) name14544 (
		_w19821_,
		_w20365_,
		_w20370_,
		_w20371_
	);
	LUT4 #(
		.INIT('hf77f)
	) name14545 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20372_
	);
	LUT2 #(
		.INIT('h1)
	) name14546 (
		_w19820_,
		_w20372_,
		_w20373_
	);
	LUT4 #(
		.INIT('h9060)
	) name14547 (
		_w19823_,
		_w19824_,
		_w19822_,
		_w19825_,
		_w20374_
	);
	LUT4 #(
		.INIT('h0031)
	) name14548 (
		_w19832_,
		_w20034_,
		_w20367_,
		_w20374_,
		_w20375_
	);
	LUT3 #(
		.INIT('h31)
	) name14549 (
		_w19821_,
		_w20373_,
		_w20375_,
		_w20376_
	);
	LUT3 #(
		.INIT('h65)
	) name14550 (
		\u1_L6_reg[9]/NET0131 ,
		_w20371_,
		_w20376_,
		_w20377_
	);
	LUT4 #(
		.INIT('h0109)
	) name14551 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20124_,
		_w20378_
	);
	LUT4 #(
		.INIT('h8000)
	) name14552 (
		_w20125_,
		_w20126_,
		_w20127_,
		_w20124_,
		_w20379_
	);
	LUT3 #(
		.INIT('h01)
	) name14553 (
		_w20125_,
		_w20128_,
		_w20127_,
		_w20380_
	);
	LUT4 #(
		.INIT('hff6e)
	) name14554 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20381_
	);
	LUT4 #(
		.INIT('h0100)
	) name14555 (
		_w20123_,
		_w20163_,
		_w20379_,
		_w20381_,
		_w20382_
	);
	LUT4 #(
		.INIT('h1a00)
	) name14556 (
		_w20125_,
		_w20126_,
		_w20127_,
		_w20124_,
		_w20383_
	);
	LUT4 #(
		.INIT('hcfaf)
	) name14557 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20384_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14558 (
		_w20124_,
		_w20123_,
		_w20177_,
		_w20384_,
		_w20385_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14559 (
		_w20378_,
		_w20382_,
		_w20383_,
		_w20385_,
		_w20386_
	);
	LUT4 #(
		.INIT('h0002)
	) name14560 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20387_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name14561 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w20388_
	);
	LUT4 #(
		.INIT('h0020)
	) name14562 (
		_w20125_,
		_w20126_,
		_w20127_,
		_w20124_,
		_w20389_
	);
	LUT3 #(
		.INIT('h0d)
	) name14563 (
		_w20124_,
		_w20388_,
		_w20389_,
		_w20390_
	);
	LUT3 #(
		.INIT('h65)
	) name14564 (
		\u1_L6_reg[18]/NET0131 ,
		_w20386_,
		_w20390_,
		_w20391_
	);
	LUT4 #(
		.INIT('hc963)
	) name14565 (
		decrypt_pad,
		\u1_R5_reg[4]/NET0131 ,
		\u1_uk_K_r5_reg[11]/NET0131 ,
		\u1_uk_K_r5_reg[33]/NET0131 ,
		_w20392_
	);
	LUT4 #(
		.INIT('hc963)
	) name14566 (
		decrypt_pad,
		\u1_R5_reg[3]/NET0131 ,
		\u1_uk_K_r5_reg[33]/NET0131 ,
		\u1_uk_K_r5_reg[55]/NET0131 ,
		_w20393_
	);
	LUT4 #(
		.INIT('hc963)
	) name14567 (
		decrypt_pad,
		\u1_R5_reg[2]/NET0131 ,
		\u1_uk_K_r5_reg[24]/NET0131 ,
		\u1_uk_K_r5_reg[46]/NET0131 ,
		_w20394_
	);
	LUT4 #(
		.INIT('hc963)
	) name14568 (
		decrypt_pad,
		\u1_R5_reg[1]/NET0131 ,
		\u1_uk_K_r5_reg[41]/NET0131 ,
		\u1_uk_K_r5_reg[6]/NET0131 ,
		_w20395_
	);
	LUT4 #(
		.INIT('hc963)
	) name14569 (
		decrypt_pad,
		\u1_R5_reg[5]/NET0131 ,
		\u1_uk_K_r5_reg[39]/NET0131 ,
		\u1_uk_K_r5_reg[4]/NET0131 ,
		_w20396_
	);
	LUT4 #(
		.INIT('hc693)
	) name14570 (
		decrypt_pad,
		\u1_R5_reg[32]/NET0131 ,
		\u1_uk_K_r5_reg[10]/NET0131 ,
		\u1_uk_K_r5_reg[20]/NET0131 ,
		_w20397_
	);
	LUT4 #(
		.INIT('heff4)
	) name14571 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20398_
	);
	LUT2 #(
		.INIT('h1)
	) name14572 (
		_w20393_,
		_w20398_,
		_w20399_
	);
	LUT2 #(
		.INIT('h1)
	) name14573 (
		_w20396_,
		_w20397_,
		_w20400_
	);
	LUT3 #(
		.INIT('h28)
	) name14574 (
		_w20395_,
		_w20396_,
		_w20397_,
		_w20401_
	);
	LUT4 #(
		.INIT('h4ff3)
	) name14575 (
		_w20393_,
		_w20395_,
		_w20396_,
		_w20397_,
		_w20402_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name14576 (
		_w20393_,
		_w20394_,
		_w20401_,
		_w20402_,
		_w20403_
	);
	LUT3 #(
		.INIT('h45)
	) name14577 (
		_w20392_,
		_w20399_,
		_w20403_,
		_w20404_
	);
	LUT4 #(
		.INIT('hbb8b)
	) name14578 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20405_
	);
	LUT2 #(
		.INIT('h2)
	) name14579 (
		_w20393_,
		_w20405_,
		_w20406_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name14580 (
		_w20393_,
		_w20395_,
		_w20396_,
		_w20394_,
		_w20407_
	);
	LUT2 #(
		.INIT('h2)
	) name14581 (
		_w20393_,
		_w20394_,
		_w20408_
	);
	LUT3 #(
		.INIT('hc4)
	) name14582 (
		_w20393_,
		_w20395_,
		_w20394_,
		_w20409_
	);
	LUT3 #(
		.INIT('h0e)
	) name14583 (
		_w20396_,
		_w20394_,
		_w20397_,
		_w20410_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14584 (
		_w20407_,
		_w20397_,
		_w20409_,
		_w20410_,
		_w20411_
	);
	LUT3 #(
		.INIT('hb0)
	) name14585 (
		_w20406_,
		_w20411_,
		_w20392_,
		_w20412_
	);
	LUT4 #(
		.INIT('h7dbd)
	) name14586 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20413_
	);
	LUT2 #(
		.INIT('h1)
	) name14587 (
		_w20393_,
		_w20413_,
		_w20414_
	);
	LUT3 #(
		.INIT('h20)
	) name14588 (
		_w20393_,
		_w20395_,
		_w20394_,
		_w20415_
	);
	LUT4 #(
		.INIT('h0200)
	) name14589 (
		_w20393_,
		_w20395_,
		_w20394_,
		_w20397_,
		_w20416_
	);
	LUT3 #(
		.INIT('h07)
	) name14590 (
		_w20400_,
		_w20415_,
		_w20416_,
		_w20417_
	);
	LUT2 #(
		.INIT('h4)
	) name14591 (
		_w20414_,
		_w20417_,
		_w20418_
	);
	LUT4 #(
		.INIT('h5655)
	) name14592 (
		\u1_L5_reg[31]/NET0131 ,
		_w20412_,
		_w20404_,
		_w20418_,
		_w20419_
	);
	LUT4 #(
		.INIT('hc693)
	) name14593 (
		decrypt_pad,
		\u1_R5_reg[24]/NET0131 ,
		\u1_uk_K_r5_reg[2]/NET0131 ,
		\u1_uk_K_r5_reg[37]/P0001 ,
		_w20420_
	);
	LUT4 #(
		.INIT('hc693)
	) name14594 (
		decrypt_pad,
		\u1_R5_reg[23]/NET0131 ,
		\u1_uk_K_r5_reg[0]/NET0131 ,
		\u1_uk_K_r5_reg[35]/NET0131 ,
		_w20421_
	);
	LUT4 #(
		.INIT('hc963)
	) name14595 (
		decrypt_pad,
		\u1_R5_reg[22]/NET0131 ,
		\u1_uk_K_r5_reg[22]/NET0131 ,
		\u1_uk_K_r5_reg[42]/NET0131 ,
		_w20422_
	);
	LUT4 #(
		.INIT('hc963)
	) name14596 (
		decrypt_pad,
		\u1_R5_reg[20]/NET0131 ,
		\u1_uk_K_r5_reg[16]/NET0131 ,
		\u1_uk_K_r5_reg[36]/NET0131 ,
		_w20423_
	);
	LUT4 #(
		.INIT('hc963)
	) name14597 (
		decrypt_pad,
		\u1_R5_reg[21]/NET0131 ,
		\u1_uk_K_r5_reg[0]/NET0131 ,
		\u1_uk_K_r5_reg[51]/NET0131 ,
		_w20424_
	);
	LUT4 #(
		.INIT('hc963)
	) name14598 (
		decrypt_pad,
		\u1_R5_reg[25]/NET0131 ,
		\u1_uk_K_r5_reg[1]/NET0131 ,
		\u1_uk_K_r5_reg[21]/NET0131 ,
		_w20425_
	);
	LUT3 #(
		.INIT('h8a)
	) name14599 (
		_w20423_,
		_w20425_,
		_w20424_,
		_w20426_
	);
	LUT4 #(
		.INIT('h1dfb)
	) name14600 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20427_
	);
	LUT2 #(
		.INIT('h2)
	) name14601 (
		_w20421_,
		_w20427_,
		_w20428_
	);
	LUT4 #(
		.INIT('h4555)
	) name14602 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20429_
	);
	LUT4 #(
		.INIT('ha280)
	) name14603 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20430_
	);
	LUT3 #(
		.INIT('h01)
	) name14604 (
		_w20421_,
		_w20430_,
		_w20429_,
		_w20431_
	);
	LUT2 #(
		.INIT('h1)
	) name14605 (
		_w20422_,
		_w20421_,
		_w20432_
	);
	LUT4 #(
		.INIT('h1000)
	) name14606 (
		_w20422_,
		_w20421_,
		_w20423_,
		_w20425_,
		_w20433_
	);
	LUT2 #(
		.INIT('h4)
	) name14607 (
		_w20424_,
		_w20433_,
		_w20434_
	);
	LUT4 #(
		.INIT('haaa8)
	) name14608 (
		_w20420_,
		_w20431_,
		_w20428_,
		_w20434_,
		_w20435_
	);
	LUT4 #(
		.INIT('h0080)
	) name14609 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20436_
	);
	LUT3 #(
		.INIT('h54)
	) name14610 (
		_w20422_,
		_w20421_,
		_w20423_,
		_w20437_
	);
	LUT4 #(
		.INIT('h0010)
	) name14611 (
		_w20422_,
		_w20421_,
		_w20423_,
		_w20425_,
		_w20438_
	);
	LUT4 #(
		.INIT('h000b)
	) name14612 (
		_w20426_,
		_w20437_,
		_w20438_,
		_w20436_,
		_w20439_
	);
	LUT4 #(
		.INIT('h1200)
	) name14613 (
		_w20422_,
		_w20421_,
		_w20423_,
		_w20424_,
		_w20440_
	);
	LUT3 #(
		.INIT('h04)
	) name14614 (
		_w20423_,
		_w20425_,
		_w20424_,
		_w20441_
	);
	LUT4 #(
		.INIT('hff47)
	) name14615 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20442_
	);
	LUT3 #(
		.INIT('h31)
	) name14616 (
		_w20421_,
		_w20440_,
		_w20442_,
		_w20443_
	);
	LUT3 #(
		.INIT('h15)
	) name14617 (
		_w20420_,
		_w20439_,
		_w20443_,
		_w20444_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name14618 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20445_
	);
	LUT4 #(
		.INIT('h888c)
	) name14619 (
		_w20422_,
		_w20421_,
		_w20423_,
		_w20425_,
		_w20446_
	);
	LUT2 #(
		.INIT('h4)
	) name14620 (
		_w20445_,
		_w20446_,
		_w20447_
	);
	LUT3 #(
		.INIT('h20)
	) name14621 (
		_w20423_,
		_w20425_,
		_w20424_,
		_w20448_
	);
	LUT3 #(
		.INIT('hde)
	) name14622 (
		_w20423_,
		_w20425_,
		_w20424_,
		_w20449_
	);
	LUT2 #(
		.INIT('h4)
	) name14623 (
		_w20422_,
		_w20421_,
		_w20450_
	);
	LUT4 #(
		.INIT('hbafe)
	) name14624 (
		_w20422_,
		_w20421_,
		_w20449_,
		_w20441_,
		_w20451_
	);
	LUT2 #(
		.INIT('h4)
	) name14625 (
		_w20447_,
		_w20451_,
		_w20452_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name14626 (
		\u1_L5_reg[11]/NET0131 ,
		_w20444_,
		_w20435_,
		_w20452_,
		_w20453_
	);
	LUT4 #(
		.INIT('hc963)
	) name14627 (
		decrypt_pad,
		\u1_R5_reg[28]/NET0131 ,
		\u1_uk_K_r5_reg[44]/NET0131 ,
		\u1_uk_K_r5_reg[9]/NET0131 ,
		_w20454_
	);
	LUT4 #(
		.INIT('hc693)
	) name14628 (
		decrypt_pad,
		\u1_R5_reg[26]/NET0131 ,
		\u1_uk_K_r5_reg[44]/NET0131 ,
		\u1_uk_K_r5_reg[52]/NET0131 ,
		_w20455_
	);
	LUT4 #(
		.INIT('hc693)
	) name14629 (
		decrypt_pad,
		\u1_R5_reg[25]/NET0131 ,
		\u1_uk_K_r5_reg[28]/NET0131 ,
		\u1_uk_K_r5_reg[8]/NET0131 ,
		_w20456_
	);
	LUT4 #(
		.INIT('hc693)
	) name14630 (
		decrypt_pad,
		\u1_R5_reg[29]/NET0131 ,
		\u1_uk_K_r5_reg[1]/NET0131 ,
		\u1_uk_K_r5_reg[36]/NET0131 ,
		_w20457_
	);
	LUT3 #(
		.INIT('hea)
	) name14631 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20458_
	);
	LUT4 #(
		.INIT('hc963)
	) name14632 (
		decrypt_pad,
		\u1_R5_reg[24]/NET0131 ,
		\u1_uk_K_r5_reg[28]/NET0131 ,
		\u1_uk_K_r5_reg[52]/NET0131 ,
		_w20459_
	);
	LUT4 #(
		.INIT('hc693)
	) name14633 (
		decrypt_pad,
		\u1_R5_reg[27]/NET0131 ,
		\u1_uk_K_r5_reg[22]/NET0131 ,
		\u1_uk_K_r5_reg[2]/NET0131 ,
		_w20460_
	);
	LUT3 #(
		.INIT('h70)
	) name14634 (
		_w20455_,
		_w20456_,
		_w20460_,
		_w20461_
	);
	LUT4 #(
		.INIT('h7000)
	) name14635 (
		_w20455_,
		_w20456_,
		_w20459_,
		_w20460_,
		_w20462_
	);
	LUT2 #(
		.INIT('h8)
	) name14636 (
		_w20458_,
		_w20462_,
		_w20463_
	);
	LUT4 #(
		.INIT('h1000)
	) name14637 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20464_
	);
	LUT4 #(
		.INIT('hef3f)
	) name14638 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20465_
	);
	LUT2 #(
		.INIT('h2)
	) name14639 (
		_w20457_,
		_w20459_,
		_w20466_
	);
	LUT4 #(
		.INIT('h0020)
	) name14640 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20467_
	);
	LUT4 #(
		.INIT('hffde)
	) name14641 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20468_
	);
	LUT3 #(
		.INIT('he0)
	) name14642 (
		_w20460_,
		_w20465_,
		_w20468_,
		_w20469_
	);
	LUT3 #(
		.INIT('h8a)
	) name14643 (
		_w20454_,
		_w20463_,
		_w20469_,
		_w20470_
	);
	LUT4 #(
		.INIT('h0072)
	) name14644 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20460_,
		_w20471_
	);
	LUT4 #(
		.INIT('h10f0)
	) name14645 (
		_w20455_,
		_w20456_,
		_w20459_,
		_w20460_,
		_w20472_
	);
	LUT2 #(
		.INIT('h4)
	) name14646 (
		_w20471_,
		_w20472_,
		_w20473_
	);
	LUT4 #(
		.INIT('h0002)
	) name14647 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20474_
	);
	LUT2 #(
		.INIT('h6)
	) name14648 (
		_w20455_,
		_w20459_,
		_w20475_
	);
	LUT3 #(
		.INIT('h8c)
	) name14649 (
		_w20456_,
		_w20457_,
		_w20460_,
		_w20476_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name14650 (
		_w20474_,
		_w20460_,
		_w20475_,
		_w20476_,
		_w20477_
	);
	LUT4 #(
		.INIT('h0008)
	) name14651 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20478_
	);
	LUT4 #(
		.INIT('hfcd7)
	) name14652 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20479_
	);
	LUT4 #(
		.INIT('h0084)
	) name14653 (
		_w20455_,
		_w20456_,
		_w20459_,
		_w20460_,
		_w20480_
	);
	LUT4 #(
		.INIT('h0100)
	) name14654 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20460_,
		_w20481_
	);
	LUT4 #(
		.INIT('h0031)
	) name14655 (
		_w20460_,
		_w20480_,
		_w20479_,
		_w20481_,
		_w20482_
	);
	LUT4 #(
		.INIT('hba00)
	) name14656 (
		_w20454_,
		_w20473_,
		_w20477_,
		_w20482_,
		_w20483_
	);
	LUT3 #(
		.INIT('h65)
	) name14657 (
		\u1_L5_reg[22]/NET0131 ,
		_w20470_,
		_w20483_,
		_w20484_
	);
	LUT2 #(
		.INIT('h1)
	) name14658 (
		_w20395_,
		_w20394_,
		_w20485_
	);
	LUT4 #(
		.INIT('h0400)
	) name14659 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20486_
	);
	LUT4 #(
		.INIT('hfb05)
	) name14660 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20487_
	);
	LUT4 #(
		.INIT('h5001)
	) name14661 (
		_w20393_,
		_w20395_,
		_w20394_,
		_w20397_,
		_w20488_
	);
	LUT3 #(
		.INIT('h80)
	) name14662 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20489_
	);
	LUT4 #(
		.INIT('h0200)
	) name14663 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20490_
	);
	LUT4 #(
		.INIT('h7d7f)
	) name14664 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20491_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14665 (
		_w20393_,
		_w20487_,
		_w20488_,
		_w20491_,
		_w20492_
	);
	LUT4 #(
		.INIT('hbbec)
	) name14666 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20493_
	);
	LUT3 #(
		.INIT('h6f)
	) name14667 (
		_w20395_,
		_w20396_,
		_w20397_,
		_w20494_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name14668 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20495_
	);
	LUT4 #(
		.INIT('he400)
	) name14669 (
		_w20393_,
		_w20493_,
		_w20494_,
		_w20495_,
		_w20496_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name14670 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20497_
	);
	LUT4 #(
		.INIT('h0f07)
	) name14671 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20498_
	);
	LUT3 #(
		.INIT('h02)
	) name14672 (
		_w20393_,
		_w20498_,
		_w20497_,
		_w20499_
	);
	LUT4 #(
		.INIT('h0e04)
	) name14673 (
		_w20392_,
		_w20496_,
		_w20499_,
		_w20492_,
		_w20500_
	);
	LUT2 #(
		.INIT('h9)
	) name14674 (
		\u1_L5_reg[17]/NET0131 ,
		_w20500_,
		_w20501_
	);
	LUT4 #(
		.INIT('hc963)
	) name14675 (
		decrypt_pad,
		\u1_R5_reg[16]/NET0131 ,
		\u1_uk_K_r5_reg[13]/P0001 ,
		\u1_uk_K_r5_reg[3]/NET0131 ,
		_w20502_
	);
	LUT4 #(
		.INIT('hc693)
	) name14676 (
		decrypt_pad,
		\u1_R5_reg[13]/NET0131 ,
		\u1_uk_K_r5_reg[18]/NET0131 ,
		\u1_uk_K_r5_reg[53]/NET0131 ,
		_w20503_
	);
	LUT4 #(
		.INIT('hc693)
	) name14677 (
		decrypt_pad,
		\u1_R5_reg[15]/NET0131 ,
		\u1_uk_K_r5_reg[27]/NET0131 ,
		\u1_uk_K_r5_reg[5]/NET0131 ,
		_w20504_
	);
	LUT4 #(
		.INIT('hc693)
	) name14678 (
		decrypt_pad,
		\u1_R5_reg[12]/NET0131 ,
		\u1_uk_K_r5_reg[24]/NET0131 ,
		\u1_uk_K_r5_reg[34]/NET0131 ,
		_w20505_
	);
	LUT4 #(
		.INIT('hc963)
	) name14679 (
		decrypt_pad,
		\u1_R5_reg[17]/NET0131 ,
		\u1_uk_K_r5_reg[18]/NET0131 ,
		\u1_uk_K_r5_reg[40]/NET0131 ,
		_w20506_
	);
	LUT4 #(
		.INIT('h0200)
	) name14680 (
		_w20504_,
		_w20503_,
		_w20505_,
		_w20506_,
		_w20507_
	);
	LUT4 #(
		.INIT('hc693)
	) name14681 (
		decrypt_pad,
		\u1_R5_reg[14]/NET0131 ,
		\u1_uk_K_r5_reg[19]/NET0131 ,
		\u1_uk_K_r5_reg[54]/NET0131 ,
		_w20508_
	);
	LUT2 #(
		.INIT('h1)
	) name14682 (
		_w20504_,
		_w20508_,
		_w20509_
	);
	LUT4 #(
		.INIT('h0014)
	) name14683 (
		_w20504_,
		_w20503_,
		_w20505_,
		_w20508_,
		_w20510_
	);
	LUT2 #(
		.INIT('h8)
	) name14684 (
		_w20504_,
		_w20503_,
		_w20511_
	);
	LUT4 #(
		.INIT('h0080)
	) name14685 (
		_w20504_,
		_w20503_,
		_w20505_,
		_w20506_,
		_w20512_
	);
	LUT3 #(
		.INIT('h01)
	) name14686 (
		_w20510_,
		_w20507_,
		_w20512_,
		_w20513_
	);
	LUT4 #(
		.INIT('h0020)
	) name14687 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20514_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name14688 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20515_
	);
	LUT4 #(
		.INIT('h0100)
	) name14689 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20516_
	);
	LUT3 #(
		.INIT('h8c)
	) name14690 (
		_w20504_,
		_w20515_,
		_w20516_,
		_w20517_
	);
	LUT3 #(
		.INIT('h2a)
	) name14691 (
		_w20502_,
		_w20513_,
		_w20517_,
		_w20518_
	);
	LUT4 #(
		.INIT('h0200)
	) name14692 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20519_
	);
	LUT4 #(
		.INIT('h0040)
	) name14693 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20520_
	);
	LUT4 #(
		.INIT('h0002)
	) name14694 (
		_w20504_,
		_w20503_,
		_w20505_,
		_w20506_,
		_w20521_
	);
	LUT3 #(
		.INIT('h01)
	) name14695 (
		_w20520_,
		_w20521_,
		_w20519_,
		_w20522_
	);
	LUT4 #(
		.INIT('ha3af)
	) name14696 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20523_
	);
	LUT2 #(
		.INIT('h1)
	) name14697 (
		_w20504_,
		_w20523_,
		_w20524_
	);
	LUT2 #(
		.INIT('h1)
	) name14698 (
		_w20505_,
		_w20508_,
		_w20525_
	);
	LUT4 #(
		.INIT('h8808)
	) name14699 (
		_w20504_,
		_w20503_,
		_w20505_,
		_w20506_,
		_w20526_
	);
	LUT4 #(
		.INIT('h0001)
	) name14700 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20527_
	);
	LUT3 #(
		.INIT('h0b)
	) name14701 (
		_w20525_,
		_w20526_,
		_w20527_,
		_w20528_
	);
	LUT4 #(
		.INIT('h4555)
	) name14702 (
		_w20502_,
		_w20524_,
		_w20528_,
		_w20522_,
		_w20529_
	);
	LUT4 #(
		.INIT('h0400)
	) name14703 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20530_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name14704 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20531_
	);
	LUT2 #(
		.INIT('h2)
	) name14705 (
		_w20504_,
		_w20531_,
		_w20532_
	);
	LUT3 #(
		.INIT('h02)
	) name14706 (
		_w20505_,
		_w20506_,
		_w20508_,
		_w20533_
	);
	LUT3 #(
		.INIT('h20)
	) name14707 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20534_
	);
	LUT4 #(
		.INIT('h0777)
	) name14708 (
		_w20511_,
		_w20533_,
		_w20509_,
		_w20534_,
		_w20535_
	);
	LUT2 #(
		.INIT('h4)
	) name14709 (
		_w20532_,
		_w20535_,
		_w20536_
	);
	LUT4 #(
		.INIT('h5655)
	) name14710 (
		\u1_L5_reg[20]/NET0131 ,
		_w20529_,
		_w20518_,
		_w20536_,
		_w20537_
	);
	LUT4 #(
		.INIT('hc693)
	) name14711 (
		decrypt_pad,
		\u1_R5_reg[6]/NET0131 ,
		\u1_uk_K_r5_reg[17]/NET0131 ,
		\u1_uk_K_r5_reg[27]/NET0131 ,
		_w20538_
	);
	LUT4 #(
		.INIT('hc963)
	) name14712 (
		decrypt_pad,
		\u1_R5_reg[9]/NET0131 ,
		\u1_uk_K_r5_reg[17]/NET0131 ,
		\u1_uk_K_r5_reg[39]/NET0131 ,
		_w20539_
	);
	LUT4 #(
		.INIT('hc693)
	) name14713 (
		decrypt_pad,
		\u1_R5_reg[5]/NET0131 ,
		\u1_uk_K_r5_reg[26]/NET0131 ,
		\u1_uk_K_r5_reg[4]/NET0131 ,
		_w20540_
	);
	LUT2 #(
		.INIT('h4)
	) name14714 (
		_w20539_,
		_w20540_,
		_w20541_
	);
	LUT4 #(
		.INIT('hc963)
	) name14715 (
		decrypt_pad,
		\u1_R5_reg[4]/NET0131 ,
		\u1_uk_K_r5_reg[25]/NET0131 ,
		\u1_uk_K_r5_reg[47]/NET0131 ,
		_w20542_
	);
	LUT2 #(
		.INIT('h2)
	) name14716 (
		_w20539_,
		_w20540_,
		_w20543_
	);
	LUT4 #(
		.INIT('h0406)
	) name14717 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20544_
	);
	LUT4 #(
		.INIT('hc693)
	) name14718 (
		decrypt_pad,
		\u1_R5_reg[7]/NET0131 ,
		\u1_uk_K_r5_reg[11]/NET0131 ,
		\u1_uk_K_r5_reg[46]/NET0131 ,
		_w20545_
	);
	LUT3 #(
		.INIT('h80)
	) name14719 (
		_w20545_,
		_w20538_,
		_w20542_,
		_w20546_
	);
	LUT4 #(
		.INIT('hc963)
	) name14720 (
		decrypt_pad,
		\u1_R5_reg[8]/NET0131 ,
		\u1_uk_K_r5_reg[12]/P0001 ,
		\u1_uk_K_r5_reg[34]/NET0131 ,
		_w20547_
	);
	LUT4 #(
		.INIT('h0013)
	) name14721 (
		_w20543_,
		_w20544_,
		_w20546_,
		_w20547_,
		_w20548_
	);
	LUT2 #(
		.INIT('h2)
	) name14722 (
		_w20539_,
		_w20542_,
		_w20549_
	);
	LUT4 #(
		.INIT('hf070)
	) name14723 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20550_
	);
	LUT3 #(
		.INIT('h0e)
	) name14724 (
		_w20545_,
		_w20540_,
		_w20538_,
		_w20551_
	);
	LUT4 #(
		.INIT('hff04)
	) name14725 (
		_w20545_,
		_w20539_,
		_w20540_,
		_w20538_,
		_w20552_
	);
	LUT4 #(
		.INIT('h2fdd)
	) name14726 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20553_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name14727 (
		_w20545_,
		_w20550_,
		_w20552_,
		_w20553_,
		_w20554_
	);
	LUT2 #(
		.INIT('h8)
	) name14728 (
		_w20548_,
		_w20554_,
		_w20555_
	);
	LUT4 #(
		.INIT('h51f5)
	) name14729 (
		_w20545_,
		_w20539_,
		_w20538_,
		_w20542_,
		_w20556_
	);
	LUT2 #(
		.INIT('h2)
	) name14730 (
		_w20540_,
		_w20556_,
		_w20557_
	);
	LUT3 #(
		.INIT('h8a)
	) name14731 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20558_
	);
	LUT3 #(
		.INIT('hae)
	) name14732 (
		_w20545_,
		_w20540_,
		_w20538_,
		_w20559_
	);
	LUT2 #(
		.INIT('h9)
	) name14733 (
		_w20539_,
		_w20542_,
		_w20560_
	);
	LUT3 #(
		.INIT('h10)
	) name14734 (
		_w20559_,
		_w20558_,
		_w20560_,
		_w20561_
	);
	LUT3 #(
		.INIT('h01)
	) name14735 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20562_
	);
	LUT4 #(
		.INIT('h0100)
	) name14736 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20563_
	);
	LUT2 #(
		.INIT('h2)
	) name14737 (
		_w20547_,
		_w20563_,
		_w20564_
	);
	LUT3 #(
		.INIT('h10)
	) name14738 (
		_w20561_,
		_w20557_,
		_w20564_,
		_w20565_
	);
	LUT3 #(
		.INIT('h04)
	) name14739 (
		_w20540_,
		_w20538_,
		_w20542_,
		_w20566_
	);
	LUT4 #(
		.INIT('h0010)
	) name14740 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20567_
	);
	LUT4 #(
		.INIT('hf3ef)
	) name14741 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20568_
	);
	LUT3 #(
		.INIT('h0b)
	) name14742 (
		_w20540_,
		_w20538_,
		_w20542_,
		_w20569_
	);
	LUT4 #(
		.INIT('h4404)
	) name14743 (
		_w20545_,
		_w20539_,
		_w20540_,
		_w20538_,
		_w20570_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name14744 (
		_w20545_,
		_w20568_,
		_w20569_,
		_w20570_,
		_w20571_
	);
	LUT4 #(
		.INIT('ha955)
	) name14745 (
		\u1_L5_reg[2]/NET0131 ,
		_w20555_,
		_w20565_,
		_w20571_,
		_w20572_
	);
	LUT4 #(
		.INIT('h3df2)
	) name14746 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20573_
	);
	LUT4 #(
		.INIT('h5140)
	) name14747 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20574_
	);
	LUT4 #(
		.INIT('ha6bf)
	) name14748 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20575_
	);
	LUT4 #(
		.INIT('h0020)
	) name14749 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20576_
	);
	LUT4 #(
		.INIT('h00e4)
	) name14750 (
		_w20421_,
		_w20575_,
		_w20573_,
		_w20576_,
		_w20577_
	);
	LUT2 #(
		.INIT('h1)
	) name14751 (
		_w20420_,
		_w20577_,
		_w20578_
	);
	LUT4 #(
		.INIT('hc6ff)
	) name14752 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20579_
	);
	LUT2 #(
		.INIT('h2)
	) name14753 (
		_w20421_,
		_w20579_,
		_w20580_
	);
	LUT3 #(
		.INIT('h28)
	) name14754 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20581_
	);
	LUT4 #(
		.INIT('hcc04)
	) name14755 (
		_w20422_,
		_w20421_,
		_w20425_,
		_w20424_,
		_w20582_
	);
	LUT3 #(
		.INIT('h01)
	) name14756 (
		_w20574_,
		_w20582_,
		_w20581_,
		_w20583_
	);
	LUT4 #(
		.INIT('h4000)
	) name14757 (
		_w20422_,
		_w20421_,
		_w20425_,
		_w20424_,
		_w20584_
	);
	LUT4 #(
		.INIT('h0004)
	) name14758 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20585_
	);
	LUT2 #(
		.INIT('h1)
	) name14759 (
		_w20584_,
		_w20585_,
		_w20586_
	);
	LUT4 #(
		.INIT('h5700)
	) name14760 (
		_w20420_,
		_w20580_,
		_w20583_,
		_w20586_,
		_w20587_
	);
	LUT3 #(
		.INIT('h9a)
	) name14761 (
		\u1_L5_reg[29]/NET0131 ,
		_w20578_,
		_w20587_,
		_w20588_
	);
	LUT4 #(
		.INIT('hc963)
	) name14762 (
		decrypt_pad,
		\u1_R5_reg[30]/NET0131 ,
		\u1_uk_K_r5_reg[15]/NET0131 ,
		\u1_uk_K_r5_reg[35]/NET0131 ,
		_w20589_
	);
	LUT4 #(
		.INIT('hc963)
	) name14763 (
		decrypt_pad,
		\u1_R5_reg[29]/NET0131 ,
		\u1_uk_K_r5_reg[14]/NET0131 ,
		\u1_uk_K_r5_reg[38]/NET0131 ,
		_w20590_
	);
	LUT4 #(
		.INIT('hc963)
	) name14764 (
		decrypt_pad,
		\u1_R5_reg[1]/NET0131 ,
		\u1_uk_K_r5_reg[30]/NET0131 ,
		\u1_uk_K_r5_reg[50]/NET0131 ,
		_w20591_
	);
	LUT2 #(
		.INIT('h8)
	) name14765 (
		_w20590_,
		_w20591_,
		_w20592_
	);
	LUT4 #(
		.INIT('hc963)
	) name14766 (
		decrypt_pad,
		\u1_R5_reg[28]/NET0131 ,
		\u1_uk_K_r5_reg[42]/NET0131 ,
		\u1_uk_K_r5_reg[7]/NET0131 ,
		_w20593_
	);
	LUT4 #(
		.INIT('h0080)
	) name14767 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20594_
	);
	LUT2 #(
		.INIT('h2)
	) name14768 (
		_w20590_,
		_w20591_,
		_w20595_
	);
	LUT4 #(
		.INIT('h0400)
	) name14769 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20596_
	);
	LUT4 #(
		.INIT('h590c)
	) name14770 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20597_
	);
	LUT4 #(
		.INIT('hc693)
	) name14771 (
		decrypt_pad,
		\u1_R5_reg[31]/P0001 ,
		\u1_uk_K_r5_reg[23]/NET0131 ,
		\u1_uk_K_r5_reg[31]/NET0131 ,
		_w20598_
	);
	LUT4 #(
		.INIT('h00df)
	) name14772 (
		_w20589_,
		_w20590_,
		_w20593_,
		_w20598_,
		_w20599_
	);
	LUT4 #(
		.INIT('h00de)
	) name14773 (
		_w20589_,
		_w20590_,
		_w20593_,
		_w20598_,
		_w20600_
	);
	LUT4 #(
		.INIT('h5510)
	) name14774 (
		_w20594_,
		_w20597_,
		_w20598_,
		_w20600_,
		_w20601_
	);
	LUT4 #(
		.INIT('hc693)
	) name14775 (
		decrypt_pad,
		\u1_R5_reg[32]/NET0131 ,
		\u1_uk_K_r5_reg[29]/NET0131 ,
		\u1_uk_K_r5_reg[9]/NET0131 ,
		_w20602_
	);
	LUT2 #(
		.INIT('h4)
	) name14776 (
		_w20601_,
		_w20602_,
		_w20603_
	);
	LUT4 #(
		.INIT('h0200)
	) name14777 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20604_
	);
	LUT4 #(
		.INIT('hfb00)
	) name14778 (
		_w20590_,
		_w20591_,
		_w20593_,
		_w20598_,
		_w20605_
	);
	LUT3 #(
		.INIT('h02)
	) name14779 (
		_w20589_,
		_w20591_,
		_w20593_,
		_w20606_
	);
	LUT3 #(
		.INIT('h07)
	) name14780 (
		_w20590_,
		_w20591_,
		_w20598_,
		_w20607_
	);
	LUT4 #(
		.INIT('h8acf)
	) name14781 (
		_w20606_,
		_w20604_,
		_w20605_,
		_w20607_,
		_w20608_
	);
	LUT4 #(
		.INIT('h8000)
	) name14782 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20609_
	);
	LUT3 #(
		.INIT('h04)
	) name14783 (
		_w20589_,
		_w20593_,
		_w20598_,
		_w20610_
	);
	LUT3 #(
		.INIT('h01)
	) name14784 (
		_w20596_,
		_w20610_,
		_w20609_,
		_w20611_
	);
	LUT4 #(
		.INIT('h0001)
	) name14785 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20612_
	);
	LUT4 #(
		.INIT('hfff6)
	) name14786 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20613_
	);
	LUT4 #(
		.INIT('h0020)
	) name14787 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20614_
	);
	LUT4 #(
		.INIT('hefd6)
	) name14788 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20615_
	);
	LUT4 #(
		.INIT('h5f13)
	) name14789 (
		_w20595_,
		_w20598_,
		_w20610_,
		_w20615_,
		_w20616_
	);
	LUT4 #(
		.INIT('hba00)
	) name14790 (
		_w20602_,
		_w20608_,
		_w20611_,
		_w20616_,
		_w20617_
	);
	LUT3 #(
		.INIT('h9a)
	) name14791 (
		\u1_L5_reg[5]/NET0131 ,
		_w20603_,
		_w20617_,
		_w20618_
	);
	LUT4 #(
		.INIT('hfcdf)
	) name14792 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20619_
	);
	LUT4 #(
		.INIT('h0302)
	) name14793 (
		_w20421_,
		_w20433_,
		_w20585_,
		_w20619_,
		_w20620_
	);
	LUT2 #(
		.INIT('h1)
	) name14794 (
		_w20420_,
		_w20620_,
		_w20621_
	);
	LUT4 #(
		.INIT('h2802)
	) name14795 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20622_
	);
	LUT4 #(
		.INIT('he36f)
	) name14796 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20623_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name14797 (
		_w20421_,
		_w20420_,
		_w20622_,
		_w20623_,
		_w20624_
	);
	LUT4 #(
		.INIT('ha100)
	) name14798 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20625_
	);
	LUT4 #(
		.INIT('h4000)
	) name14799 (
		_w20422_,
		_w20421_,
		_w20423_,
		_w20425_,
		_w20626_
	);
	LUT4 #(
		.INIT('h000d)
	) name14800 (
		_w20432_,
		_w20426_,
		_w20626_,
		_w20625_,
		_w20627_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name14801 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20628_
	);
	LUT4 #(
		.INIT('h2223)
	) name14802 (
		_w20422_,
		_w20421_,
		_w20423_,
		_w20425_,
		_w20629_
	);
	LUT2 #(
		.INIT('h4)
	) name14803 (
		_w20628_,
		_w20629_,
		_w20630_
	);
	LUT4 #(
		.INIT('h000d)
	) name14804 (
		_w20420_,
		_w20627_,
		_w20624_,
		_w20630_,
		_w20631_
	);
	LUT3 #(
		.INIT('h65)
	) name14805 (
		\u1_L5_reg[4]/NET0131 ,
		_w20621_,
		_w20631_,
		_w20632_
	);
	LUT4 #(
		.INIT('hfdbd)
	) name14806 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20633_
	);
	LUT2 #(
		.INIT('h2)
	) name14807 (
		_w20504_,
		_w20633_,
		_w20634_
	);
	LUT4 #(
		.INIT('h6fff)
	) name14808 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20635_
	);
	LUT4 #(
		.INIT('hf353)
	) name14809 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20636_
	);
	LUT3 #(
		.INIT('h08)
	) name14810 (
		_w20503_,
		_w20505_,
		_w20508_,
		_w20637_
	);
	LUT4 #(
		.INIT('h5515)
	) name14811 (
		_w20504_,
		_w20503_,
		_w20505_,
		_w20508_,
		_w20638_
	);
	LUT3 #(
		.INIT('h8a)
	) name14812 (
		_w20635_,
		_w20636_,
		_w20638_,
		_w20639_
	);
	LUT3 #(
		.INIT('h8a)
	) name14813 (
		_w20502_,
		_w20634_,
		_w20639_,
		_w20640_
	);
	LUT2 #(
		.INIT('h8)
	) name14814 (
		_w20504_,
		_w20508_,
		_w20641_
	);
	LUT4 #(
		.INIT('hf5fc)
	) name14815 (
		_w20504_,
		_w20503_,
		_w20505_,
		_w20506_,
		_w20642_
	);
	LUT2 #(
		.INIT('h1)
	) name14816 (
		_w20641_,
		_w20642_,
		_w20643_
	);
	LUT3 #(
		.INIT('hae)
	) name14817 (
		_w20503_,
		_w20506_,
		_w20508_,
		_w20644_
	);
	LUT2 #(
		.INIT('h8)
	) name14818 (
		_w20504_,
		_w20505_,
		_w20645_
	);
	LUT2 #(
		.INIT('h4)
	) name14819 (
		_w20644_,
		_w20645_,
		_w20646_
	);
	LUT4 #(
		.INIT('h0040)
	) name14820 (
		_w20504_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20647_
	);
	LUT3 #(
		.INIT('h01)
	) name14821 (
		_w20519_,
		_w20637_,
		_w20647_,
		_w20648_
	);
	LUT4 #(
		.INIT('h5455)
	) name14822 (
		_w20502_,
		_w20643_,
		_w20646_,
		_w20648_,
		_w20649_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name14823 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20650_
	);
	LUT2 #(
		.INIT('h1)
	) name14824 (
		_w20504_,
		_w20650_,
		_w20651_
	);
	LUT4 #(
		.INIT('h0800)
	) name14825 (
		_w20504_,
		_w20503_,
		_w20505_,
		_w20508_,
		_w20652_
	);
	LUT3 #(
		.INIT('h07)
	) name14826 (
		_w20511_,
		_w20533_,
		_w20652_,
		_w20653_
	);
	LUT2 #(
		.INIT('h4)
	) name14827 (
		_w20651_,
		_w20653_,
		_w20654_
	);
	LUT4 #(
		.INIT('h5655)
	) name14828 (
		\u1_L5_reg[10]/NET0131 ,
		_w20649_,
		_w20640_,
		_w20654_,
		_w20655_
	);
	LUT4 #(
		.INIT('h0006)
	) name14829 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20656_
	);
	LUT3 #(
		.INIT('h47)
	) name14830 (
		_w20455_,
		_w20456_,
		_w20460_,
		_w20657_
	);
	LUT4 #(
		.INIT('h0051)
	) name14831 (
		_w20454_,
		_w20466_,
		_w20657_,
		_w20656_,
		_w20658_
	);
	LUT3 #(
		.INIT('h10)
	) name14832 (
		_w20455_,
		_w20457_,
		_w20459_,
		_w20659_
	);
	LUT4 #(
		.INIT('h2100)
	) name14833 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20660_
	);
	LUT2 #(
		.INIT('h6)
	) name14834 (
		_w20456_,
		_w20457_,
		_w20661_
	);
	LUT4 #(
		.INIT('h143c)
	) name14835 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20662_
	);
	LUT3 #(
		.INIT('h32)
	) name14836 (
		_w20460_,
		_w20660_,
		_w20662_,
		_w20663_
	);
	LUT2 #(
		.INIT('h8)
	) name14837 (
		_w20658_,
		_w20663_,
		_w20664_
	);
	LUT2 #(
		.INIT('h4)
	) name14838 (
		_w20460_,
		_w20467_,
		_w20665_
	);
	LUT3 #(
		.INIT('h02)
	) name14839 (
		_w20454_,
		_w20464_,
		_w20478_,
		_w20666_
	);
	LUT4 #(
		.INIT('h0240)
	) name14840 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20667_
	);
	LUT4 #(
		.INIT('h33fe)
	) name14841 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20668_
	);
	LUT3 #(
		.INIT('h31)
	) name14842 (
		_w20460_,
		_w20667_,
		_w20668_,
		_w20669_
	);
	LUT3 #(
		.INIT('h40)
	) name14843 (
		_w20665_,
		_w20666_,
		_w20669_,
		_w20670_
	);
	LUT3 #(
		.INIT('ha9)
	) name14844 (
		\u1_L5_reg[12]/NET0131 ,
		_w20664_,
		_w20670_,
		_w20671_
	);
	LUT4 #(
		.INIT('hfe9b)
	) name14845 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20672_
	);
	LUT4 #(
		.INIT('h4000)
	) name14846 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20673_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name14847 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20674_
	);
	LUT4 #(
		.INIT('h0155)
	) name14848 (
		_w20545_,
		_w20547_,
		_w20672_,
		_w20674_,
		_w20675_
	);
	LUT4 #(
		.INIT('hd9ee)
	) name14849 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20676_
	);
	LUT2 #(
		.INIT('h2)
	) name14850 (
		_w20545_,
		_w20676_,
		_w20677_
	);
	LUT2 #(
		.INIT('h8)
	) name14851 (
		_w20551_,
		_w20549_,
		_w20678_
	);
	LUT3 #(
		.INIT('h0b)
	) name14852 (
		_w20541_,
		_w20546_,
		_w20547_,
		_w20679_
	);
	LUT3 #(
		.INIT('h10)
	) name14853 (
		_w20677_,
		_w20678_,
		_w20679_,
		_w20680_
	);
	LUT4 #(
		.INIT('h3210)
	) name14854 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20681_
	);
	LUT3 #(
		.INIT('h08)
	) name14855 (
		_w20539_,
		_w20538_,
		_w20542_,
		_w20682_
	);
	LUT4 #(
		.INIT('hfad8)
	) name14856 (
		_w20545_,
		_w20562_,
		_w20681_,
		_w20682_,
		_w20683_
	);
	LUT4 #(
		.INIT('h0004)
	) name14857 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20684_
	);
	LUT4 #(
		.INIT('h00b0)
	) name14858 (
		_w20550_,
		_w20552_,
		_w20547_,
		_w20684_,
		_w20685_
	);
	LUT3 #(
		.INIT('h20)
	) name14859 (
		_w20674_,
		_w20683_,
		_w20685_,
		_w20686_
	);
	LUT4 #(
		.INIT('h999a)
	) name14860 (
		\u1_L5_reg[13]/NET0131 ,
		_w20675_,
		_w20680_,
		_w20686_,
		_w20687_
	);
	LUT4 #(
		.INIT('hc693)
	) name14861 (
		decrypt_pad,
		\u1_R5_reg[19]/NET0131 ,
		\u1_uk_K_r5_reg[30]/NET0131 ,
		\u1_uk_K_r5_reg[38]/NET0131 ,
		_w20688_
	);
	LUT4 #(
		.INIT('hc963)
	) name14862 (
		decrypt_pad,
		\u1_R5_reg[18]/NET0131 ,
		\u1_uk_K_r5_reg[23]/NET0131 ,
		\u1_uk_K_r5_reg[43]/NET0131 ,
		_w20689_
	);
	LUT4 #(
		.INIT('hc963)
	) name14863 (
		decrypt_pad,
		\u1_R5_reg[17]/NET0131 ,
		\u1_uk_K_r5_reg[29]/NET0131 ,
		\u1_uk_K_r5_reg[49]/NET0131 ,
		_w20690_
	);
	LUT4 #(
		.INIT('hc693)
	) name14864 (
		decrypt_pad,
		\u1_R5_reg[21]/NET0131 ,
		\u1_uk_K_r5_reg[15]/NET0131 ,
		\u1_uk_K_r5_reg[50]/NET0131 ,
		_w20691_
	);
	LUT4 #(
		.INIT('hc693)
	) name14865 (
		decrypt_pad,
		\u1_R5_reg[16]/NET0131 ,
		\u1_uk_K_r5_reg[31]/NET0131 ,
		\u1_uk_K_r5_reg[7]/NET0131 ,
		_w20692_
	);
	LUT4 #(
		.INIT('h4000)
	) name14866 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20693_
	);
	LUT4 #(
		.INIT('h0100)
	) name14867 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20694_
	);
	LUT4 #(
		.INIT('hb6c7)
	) name14868 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20695_
	);
	LUT3 #(
		.INIT('h04)
	) name14869 (
		_w20689_,
		_w20690_,
		_w20692_,
		_w20696_
	);
	LUT4 #(
		.INIT('h5fb8)
	) name14870 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20697_
	);
	LUT4 #(
		.INIT('h2000)
	) name14871 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20698_
	);
	LUT4 #(
		.INIT('hdffb)
	) name14872 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20699_
	);
	LUT4 #(
		.INIT('he400)
	) name14873 (
		_w20688_,
		_w20695_,
		_w20697_,
		_w20699_,
		_w20700_
	);
	LUT4 #(
		.INIT('hc693)
	) name14874 (
		decrypt_pad,
		\u1_R5_reg[20]/NET0131 ,
		\u1_uk_K_r5_reg[14]/NET0131 ,
		\u1_uk_K_r5_reg[49]/NET0131 ,
		_w20701_
	);
	LUT2 #(
		.INIT('h1)
	) name14875 (
		_w20700_,
		_w20701_,
		_w20702_
	);
	LUT4 #(
		.INIT('ha34f)
	) name14876 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20703_
	);
	LUT2 #(
		.INIT('h2)
	) name14877 (
		_w20688_,
		_w20703_,
		_w20704_
	);
	LUT2 #(
		.INIT('h1)
	) name14878 (
		_w20688_,
		_w20689_,
		_w20705_
	);
	LUT3 #(
		.INIT('hf6)
	) name14879 (
		_w20690_,
		_w20691_,
		_w20692_,
		_w20706_
	);
	LUT2 #(
		.INIT('h2)
	) name14880 (
		_w20705_,
		_w20706_,
		_w20707_
	);
	LUT2 #(
		.INIT('h9)
	) name14881 (
		_w20689_,
		_w20690_,
		_w20708_
	);
	LUT4 #(
		.INIT('h0600)
	) name14882 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20709_
	);
	LUT4 #(
		.INIT('h7000)
	) name14883 (
		_w20688_,
		_w20689_,
		_w20691_,
		_w20692_,
		_w20710_
	);
	LUT3 #(
		.INIT('h13)
	) name14884 (
		_w20708_,
		_w20709_,
		_w20710_,
		_w20711_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name14885 (
		_w20701_,
		_w20704_,
		_w20707_,
		_w20711_,
		_w20712_
	);
	LUT4 #(
		.INIT('h0400)
	) name14886 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20713_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name14887 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20714_
	);
	LUT4 #(
		.INIT('h0020)
	) name14888 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20715_
	);
	LUT4 #(
		.INIT('hffd7)
	) name14889 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20716_
	);
	LUT3 #(
		.INIT('hd8)
	) name14890 (
		_w20688_,
		_w20714_,
		_w20716_,
		_w20717_
	);
	LUT4 #(
		.INIT('h5655)
	) name14891 (
		\u1_L5_reg[14]/NET0131 ,
		_w20702_,
		_w20712_,
		_w20717_,
		_w20718_
	);
	LUT4 #(
		.INIT('h33cb)
	) name14892 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20719_
	);
	LUT4 #(
		.INIT('h0100)
	) name14893 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20720_
	);
	LUT4 #(
		.INIT('h0031)
	) name14894 (
		_w20598_,
		_w20602_,
		_w20719_,
		_w20720_,
		_w20721_
	);
	LUT4 #(
		.INIT('hbf00)
	) name14895 (
		_w20589_,
		_w20590_,
		_w20593_,
		_w20602_,
		_w20722_
	);
	LUT2 #(
		.INIT('h4)
	) name14896 (
		_w20590_,
		_w20598_,
		_w20723_
	);
	LUT4 #(
		.INIT('h0100)
	) name14897 (
		_w20590_,
		_w20591_,
		_w20593_,
		_w20598_,
		_w20724_
	);
	LUT4 #(
		.INIT('h0020)
	) name14898 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20598_,
		_w20725_
	);
	LUT4 #(
		.INIT('h2000)
	) name14899 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20726_
	);
	LUT4 #(
		.INIT('hdff7)
	) name14900 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20727_
	);
	LUT4 #(
		.INIT('h1000)
	) name14901 (
		_w20724_,
		_w20725_,
		_w20722_,
		_w20727_,
		_w20728_
	);
	LUT2 #(
		.INIT('h1)
	) name14902 (
		_w20721_,
		_w20728_,
		_w20729_
	);
	LUT4 #(
		.INIT('h0040)
	) name14903 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20730_
	);
	LUT3 #(
		.INIT('h08)
	) name14904 (
		_w20599_,
		_w20613_,
		_w20730_,
		_w20731_
	);
	LUT4 #(
		.INIT('h0010)
	) name14905 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20732_
	);
	LUT3 #(
		.INIT('h04)
	) name14906 (
		_w20594_,
		_w20598_,
		_w20732_,
		_w20733_
	);
	LUT4 #(
		.INIT('h0004)
	) name14907 (
		_w20590_,
		_w20593_,
		_w20598_,
		_w20602_,
		_w20734_
	);
	LUT3 #(
		.INIT('h0e)
	) name14908 (
		_w20731_,
		_w20733_,
		_w20734_,
		_w20735_
	);
	LUT3 #(
		.INIT('h65)
	) name14909 (
		\u1_L5_reg[15]/P0001 ,
		_w20729_,
		_w20735_,
		_w20736_
	);
	LUT3 #(
		.INIT('h51)
	) name14910 (
		_w20421_,
		_w20423_,
		_w20424_,
		_w20737_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name14911 (
		_w20422_,
		_w20421_,
		_w20423_,
		_w20424_,
		_w20738_
	);
	LUT3 #(
		.INIT('h23)
	) name14912 (
		_w20441_,
		_w20737_,
		_w20738_,
		_w20739_
	);
	LUT4 #(
		.INIT('h0510)
	) name14913 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20740_
	);
	LUT4 #(
		.INIT('h2002)
	) name14914 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20741_
	);
	LUT3 #(
		.INIT('h02)
	) name14915 (
		_w20420_,
		_w20741_,
		_w20740_,
		_w20742_
	);
	LUT3 #(
		.INIT('h45)
	) name14916 (
		_w20423_,
		_w20425_,
		_w20424_,
		_w20743_
	);
	LUT2 #(
		.INIT('h2)
	) name14917 (
		_w20738_,
		_w20743_,
		_w20744_
	);
	LUT4 #(
		.INIT('h1001)
	) name14918 (
		_w20421_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20745_
	);
	LUT4 #(
		.INIT('h8000)
	) name14919 (
		_w20422_,
		_w20423_,
		_w20425_,
		_w20424_,
		_w20746_
	);
	LUT3 #(
		.INIT('h01)
	) name14920 (
		_w20420_,
		_w20745_,
		_w20746_,
		_w20747_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14921 (
		_w20739_,
		_w20742_,
		_w20744_,
		_w20747_,
		_w20748_
	);
	LUT2 #(
		.INIT('h8)
	) name14922 (
		_w20432_,
		_w20448_,
		_w20749_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name14923 (
		_w20424_,
		_w20441_,
		_w20450_,
		_w20433_,
		_w20750_
	);
	LUT2 #(
		.INIT('h4)
	) name14924 (
		_w20749_,
		_w20750_,
		_w20751_
	);
	LUT3 #(
		.INIT('h65)
	) name14925 (
		\u1_L5_reg[19]/NET0131 ,
		_w20748_,
		_w20751_,
		_w20752_
	);
	LUT4 #(
		.INIT('hafab)
	) name14926 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20753_
	);
	LUT2 #(
		.INIT('h2)
	) name14927 (
		_w20502_,
		_w20753_,
		_w20754_
	);
	LUT3 #(
		.INIT('h20)
	) name14928 (
		_w20504_,
		_w20519_,
		_w20635_,
		_w20755_
	);
	LUT4 #(
		.INIT('h0800)
	) name14929 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20756_
	);
	LUT3 #(
		.INIT('h01)
	) name14930 (
		_w20504_,
		_w20516_,
		_w20756_,
		_w20757_
	);
	LUT3 #(
		.INIT('h0b)
	) name14931 (
		_w20754_,
		_w20755_,
		_w20757_,
		_w20758_
	);
	LUT3 #(
		.INIT('h40)
	) name14932 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20759_
	);
	LUT4 #(
		.INIT('h5551)
	) name14933 (
		_w20504_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20760_
	);
	LUT2 #(
		.INIT('h4)
	) name14934 (
		_w20759_,
		_w20760_,
		_w20761_
	);
	LUT3 #(
		.INIT('h01)
	) name14935 (
		_w20505_,
		_w20506_,
		_w20508_,
		_w20762_
	);
	LUT3 #(
		.INIT('h02)
	) name14936 (
		_w20504_,
		_w20530_,
		_w20762_,
		_w20763_
	);
	LUT4 #(
		.INIT('h0008)
	) name14937 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20764_
	);
	LUT3 #(
		.INIT('h04)
	) name14938 (
		_w20502_,
		_w20515_,
		_w20764_,
		_w20765_
	);
	LUT4 #(
		.INIT('hdf5d)
	) name14939 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20766_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name14940 (
		_w20502_,
		_w20503_,
		_w20505_,
		_w20508_,
		_w20767_
	);
	LUT4 #(
		.INIT('h3200)
	) name14941 (
		_w20504_,
		_w20756_,
		_w20766_,
		_w20767_,
		_w20768_
	);
	LUT4 #(
		.INIT('h001f)
	) name14942 (
		_w20761_,
		_w20763_,
		_w20765_,
		_w20768_,
		_w20769_
	);
	LUT3 #(
		.INIT('h56)
	) name14943 (
		\u1_L5_reg[1]/NET0131 ,
		_w20758_,
		_w20769_,
		_w20770_
	);
	LUT4 #(
		.INIT('h0002)
	) name14944 (
		_w20590_,
		_w20591_,
		_w20593_,
		_w20598_,
		_w20771_
	);
	LUT3 #(
		.INIT('h01)
	) name14945 (
		_w20602_,
		_w20612_,
		_w20771_,
		_w20772_
	);
	LUT3 #(
		.INIT('h40)
	) name14946 (
		_w20589_,
		_w20591_,
		_w20593_,
		_w20773_
	);
	LUT3 #(
		.INIT('h45)
	) name14947 (
		_w20604_,
		_w20723_,
		_w20773_,
		_w20774_
	);
	LUT4 #(
		.INIT('hf5f1)
	) name14948 (
		_w20590_,
		_w20591_,
		_w20593_,
		_w20598_,
		_w20775_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name14949 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20776_
	);
	LUT4 #(
		.INIT('hf531)
	) name14950 (
		_w20589_,
		_w20598_,
		_w20775_,
		_w20776_,
		_w20777_
	);
	LUT3 #(
		.INIT('h80)
	) name14951 (
		_w20772_,
		_w20774_,
		_w20777_,
		_w20778_
	);
	LUT4 #(
		.INIT('h00ef)
	) name14952 (
		_w20589_,
		_w20591_,
		_w20593_,
		_w20598_,
		_w20779_
	);
	LUT4 #(
		.INIT('hf700)
	) name14953 (
		_w20590_,
		_w20591_,
		_w20593_,
		_w20598_,
		_w20780_
	);
	LUT4 #(
		.INIT('h67ef)
	) name14954 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20781_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name14955 (
		_w20726_,
		_w20779_,
		_w20780_,
		_w20781_,
		_w20782_
	);
	LUT4 #(
		.INIT('h0802)
	) name14956 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20783_
	);
	LUT3 #(
		.INIT('h02)
	) name14957 (
		_w20602_,
		_w20732_,
		_w20783_,
		_w20784_
	);
	LUT2 #(
		.INIT('h4)
	) name14958 (
		_w20782_,
		_w20784_,
		_w20785_
	);
	LUT4 #(
		.INIT('h0100)
	) name14959 (
		_w20589_,
		_w20590_,
		_w20593_,
		_w20598_,
		_w20786_
	);
	LUT3 #(
		.INIT('h07)
	) name14960 (
		_w20592_,
		_w20610_,
		_w20786_,
		_w20787_
	);
	LUT4 #(
		.INIT('ha955)
	) name14961 (
		\u1_L5_reg[21]/NET0131 ,
		_w20778_,
		_w20785_,
		_w20787_,
		_w20788_
	);
	LUT4 #(
		.INIT('hef99)
	) name14962 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20789_
	);
	LUT4 #(
		.INIT('h7dfb)
	) name14963 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20790_
	);
	LUT4 #(
		.INIT('h0455)
	) name14964 (
		_w20393_,
		_w20392_,
		_w20789_,
		_w20790_,
		_w20791_
	);
	LUT3 #(
		.INIT('had)
	) name14965 (
		_w20395_,
		_w20396_,
		_w20397_,
		_w20792_
	);
	LUT2 #(
		.INIT('h2)
	) name14966 (
		_w20408_,
		_w20792_,
		_w20793_
	);
	LUT4 #(
		.INIT('h00fe)
	) name14967 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20392_,
		_w20794_
	);
	LUT4 #(
		.INIT('h0080)
	) name14968 (
		_w20393_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20795_
	);
	LUT3 #(
		.INIT('h10)
	) name14969 (
		_w20489_,
		_w20795_,
		_w20794_,
		_w20796_
	);
	LUT4 #(
		.INIT('h0008)
	) name14970 (
		_w20393_,
		_w20395_,
		_w20396_,
		_w20397_,
		_w20797_
	);
	LUT4 #(
		.INIT('h5400)
	) name14971 (
		_w20393_,
		_w20395_,
		_w20396_,
		_w20397_,
		_w20798_
	);
	LUT3 #(
		.INIT('h23)
	) name14972 (
		_w20485_,
		_w20797_,
		_w20798_,
		_w20799_
	);
	LUT3 #(
		.INIT('ha8)
	) name14973 (
		_w20393_,
		_w20396_,
		_w20394_,
		_w20800_
	);
	LUT2 #(
		.INIT('h8)
	) name14974 (
		_w20401_,
		_w20800_,
		_w20801_
	);
	LUT4 #(
		.INIT('h002a)
	) name14975 (
		_w20392_,
		_w20400_,
		_w20415_,
		_w20486_,
		_w20802_
	);
	LUT4 #(
		.INIT('h7077)
	) name14976 (
		_w20796_,
		_w20799_,
		_w20801_,
		_w20802_,
		_w20803_
	);
	LUT4 #(
		.INIT('haaa9)
	) name14977 (
		\u1_L5_reg[23]/NET0131 ,
		_w20793_,
		_w20803_,
		_w20791_,
		_w20804_
	);
	LUT3 #(
		.INIT('h45)
	) name14978 (
		_w20690_,
		_w20691_,
		_w20692_,
		_w20805_
	);
	LUT3 #(
		.INIT('hc4)
	) name14979 (
		_w20689_,
		_w20690_,
		_w20692_,
		_w20806_
	);
	LUT2 #(
		.INIT('h2)
	) name14980 (
		_w20688_,
		_w20691_,
		_w20807_
	);
	LUT3 #(
		.INIT('h01)
	) name14981 (
		_w20806_,
		_w20805_,
		_w20807_,
		_w20808_
	);
	LUT3 #(
		.INIT('ha2)
	) name14982 (
		_w20688_,
		_w20690_,
		_w20691_,
		_w20809_
	);
	LUT4 #(
		.INIT('h2223)
	) name14983 (
		_w20688_,
		_w20689_,
		_w20690_,
		_w20692_,
		_w20810_
	);
	LUT3 #(
		.INIT('h45)
	) name14984 (
		_w20701_,
		_w20809_,
		_w20810_,
		_w20811_
	);
	LUT4 #(
		.INIT('h4555)
	) name14985 (
		_w20688_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20812_
	);
	LUT4 #(
		.INIT('h010b)
	) name14986 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20813_
	);
	LUT3 #(
		.INIT('h80)
	) name14987 (
		_w20690_,
		_w20691_,
		_w20692_,
		_w20814_
	);
	LUT4 #(
		.INIT('h2a88)
	) name14988 (
		_w20688_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20815_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14989 (
		_w20696_,
		_w20812_,
		_w20813_,
		_w20815_,
		_w20816_
	);
	LUT4 #(
		.INIT('h0800)
	) name14990 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20817_
	);
	LUT4 #(
		.INIT('hbf00)
	) name14991 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20701_,
		_w20818_
	);
	LUT2 #(
		.INIT('h4)
	) name14992 (
		_w20817_,
		_w20818_,
		_w20819_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14993 (
		_w20808_,
		_w20811_,
		_w20816_,
		_w20819_,
		_w20820_
	);
	LUT4 #(
		.INIT('hf7ed)
	) name14994 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20821_
	);
	LUT3 #(
		.INIT('h20)
	) name14995 (
		_w20689_,
		_w20690_,
		_w20692_,
		_w20822_
	);
	LUT4 #(
		.INIT('h2301)
	) name14996 (
		_w20688_,
		_w20693_,
		_w20822_,
		_w20821_,
		_w20823_
	);
	LUT3 #(
		.INIT('h65)
	) name14997 (
		\u1_L5_reg[25]/NET0131 ,
		_w20820_,
		_w20823_,
		_w20824_
	);
	LUT4 #(
		.INIT('h0086)
	) name14998 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20825_
	);
	LUT4 #(
		.INIT('heafa)
	) name14999 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20826_
	);
	LUT4 #(
		.INIT('h0032)
	) name15000 (
		_w20502_,
		_w20504_,
		_w20826_,
		_w20825_,
		_w20827_
	);
	LUT3 #(
		.INIT('h02)
	) name15001 (
		_w20504_,
		_w20520_,
		_w20514_,
		_w20828_
	);
	LUT2 #(
		.INIT('h1)
	) name15002 (
		_w20827_,
		_w20828_,
		_w20829_
	);
	LUT4 #(
		.INIT('hf13f)
	) name15003 (
		_w20504_,
		_w20503_,
		_w20505_,
		_w20506_,
		_w20830_
	);
	LUT2 #(
		.INIT('h2)
	) name15004 (
		_w20508_,
		_w20830_,
		_w20831_
	);
	LUT4 #(
		.INIT('h3fef)
	) name15005 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20832_
	);
	LUT2 #(
		.INIT('h1)
	) name15006 (
		_w20504_,
		_w20832_,
		_w20833_
	);
	LUT4 #(
		.INIT('h0002)
	) name15007 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20508_,
		_w20834_
	);
	LUT3 #(
		.INIT('h02)
	) name15008 (
		_w20502_,
		_w20521_,
		_w20834_,
		_w20835_
	);
	LUT3 #(
		.INIT('h10)
	) name15009 (
		_w20833_,
		_w20831_,
		_w20835_,
		_w20836_
	);
	LUT4 #(
		.INIT('h5545)
	) name15010 (
		_w20502_,
		_w20503_,
		_w20505_,
		_w20508_,
		_w20837_
	);
	LUT2 #(
		.INIT('h4)
	) name15011 (
		_w20512_,
		_w20837_,
		_w20838_
	);
	LUT3 #(
		.INIT('h8a)
	) name15012 (
		_w20503_,
		_w20505_,
		_w20506_,
		_w20839_
	);
	LUT3 #(
		.INIT('h15)
	) name15013 (
		_w20514_,
		_w20641_,
		_w20839_,
		_w20840_
	);
	LUT2 #(
		.INIT('h8)
	) name15014 (
		_w20838_,
		_w20840_,
		_w20841_
	);
	LUT4 #(
		.INIT('h6665)
	) name15015 (
		\u1_L5_reg[26]/NET0131 ,
		_w20829_,
		_w20836_,
		_w20841_,
		_w20842_
	);
	LUT3 #(
		.INIT('h90)
	) name15016 (
		_w20539_,
		_w20540_,
		_w20542_,
		_w20843_
	);
	LUT4 #(
		.INIT('h0040)
	) name15017 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20844_
	);
	LUT3 #(
		.INIT('h8a)
	) name15018 (
		_w20545_,
		_w20538_,
		_w20542_,
		_w20845_
	);
	LUT3 #(
		.INIT('h10)
	) name15019 (
		_w20844_,
		_w20843_,
		_w20845_,
		_w20846_
	);
	LUT4 #(
		.INIT('h5545)
	) name15020 (
		_w20545_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20847_
	);
	LUT4 #(
		.INIT('hff72)
	) name15021 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20848_
	);
	LUT4 #(
		.INIT('hbf72)
	) name15022 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20849_
	);
	LUT2 #(
		.INIT('h8)
	) name15023 (
		_w20847_,
		_w20849_,
		_w20850_
	);
	LUT4 #(
		.INIT('h0220)
	) name15024 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20851_
	);
	LUT2 #(
		.INIT('h2)
	) name15025 (
		_w20547_,
		_w20851_,
		_w20852_
	);
	LUT3 #(
		.INIT('he0)
	) name15026 (
		_w20846_,
		_w20850_,
		_w20852_,
		_w20853_
	);
	LUT4 #(
		.INIT('h32dd)
	) name15027 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20854_
	);
	LUT4 #(
		.INIT('h4e5f)
	) name15028 (
		_w20545_,
		_w20566_,
		_w20848_,
		_w20854_,
		_w20855_
	);
	LUT4 #(
		.INIT('h2010)
	) name15029 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20856_
	);
	LUT3 #(
		.INIT('h01)
	) name15030 (
		_w20547_,
		_w20673_,
		_w20856_,
		_w20857_
	);
	LUT2 #(
		.INIT('h4)
	) name15031 (
		_w20855_,
		_w20857_,
		_w20858_
	);
	LUT3 #(
		.INIT('ha9)
	) name15032 (
		\u1_L5_reg[28]/NET0131 ,
		_w20853_,
		_w20858_,
		_w20859_
	);
	LUT4 #(
		.INIT('h0001)
	) name15033 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20860_
	);
	LUT4 #(
		.INIT('hcffe)
	) name15034 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20861_
	);
	LUT3 #(
		.INIT('h10)
	) name15035 (
		_w20688_,
		_w20689_,
		_w20692_,
		_w20862_
	);
	LUT4 #(
		.INIT('h00c4)
	) name15036 (
		_w20688_,
		_w20716_,
		_w20861_,
		_w20862_,
		_w20863_
	);
	LUT2 #(
		.INIT('h2)
	) name15037 (
		_w20701_,
		_w20863_,
		_w20864_
	);
	LUT4 #(
		.INIT('h00d0)
	) name15038 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20865_
	);
	LUT2 #(
		.INIT('h2)
	) name15039 (
		_w20812_,
		_w20865_,
		_w20866_
	);
	LUT3 #(
		.INIT('h02)
	) name15040 (
		_w20688_,
		_w20694_,
		_w20814_,
		_w20867_
	);
	LUT4 #(
		.INIT('hf7b9)
	) name15041 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20868_
	);
	LUT4 #(
		.INIT('h0155)
	) name15042 (
		_w20701_,
		_w20866_,
		_w20867_,
		_w20868_,
		_w20869_
	);
	LUT4 #(
		.INIT('hf797)
	) name15043 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20870_
	);
	LUT4 #(
		.INIT('hef45)
	) name15044 (
		_w20688_,
		_w20691_,
		_w20822_,
		_w20870_,
		_w20871_
	);
	LUT4 #(
		.INIT('h5655)
	) name15045 (
		\u1_L5_reg[8]/NET0131 ,
		_w20869_,
		_w20864_,
		_w20871_,
		_w20872_
	);
	LUT4 #(
		.INIT('hf32e)
	) name15046 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20873_
	);
	LUT2 #(
		.INIT('h1)
	) name15047 (
		_w20598_,
		_w20873_,
		_w20874_
	);
	LUT4 #(
		.INIT('hef6f)
	) name15048 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20875_
	);
	LUT2 #(
		.INIT('h6)
	) name15049 (
		_w20591_,
		_w20593_,
		_w20876_
	);
	LUT4 #(
		.INIT('hc400)
	) name15050 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20598_,
		_w20877_
	);
	LUT4 #(
		.INIT('h4500)
	) name15051 (
		_w20604_,
		_w20876_,
		_w20877_,
		_w20875_,
		_w20878_
	);
	LUT3 #(
		.INIT('h8a)
	) name15052 (
		_w20602_,
		_w20874_,
		_w20878_,
		_w20879_
	);
	LUT4 #(
		.INIT('hb0b8)
	) name15053 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20880_
	);
	LUT4 #(
		.INIT('hfb00)
	) name15054 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20598_,
		_w20881_
	);
	LUT4 #(
		.INIT('h4544)
	) name15055 (
		_w20602_,
		_w20614_,
		_w20880_,
		_w20881_,
		_w20882_
	);
	LUT4 #(
		.INIT('heff7)
	) name15056 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20593_,
		_w20883_
	);
	LUT2 #(
		.INIT('h1)
	) name15057 (
		_w20598_,
		_w20883_,
		_w20884_
	);
	LUT4 #(
		.INIT('h0080)
	) name15058 (
		_w20589_,
		_w20591_,
		_w20593_,
		_w20598_,
		_w20885_
	);
	LUT3 #(
		.INIT('h54)
	) name15059 (
		_w20602_,
		_w20771_,
		_w20885_,
		_w20886_
	);
	LUT4 #(
		.INIT('h0200)
	) name15060 (
		_w20589_,
		_w20590_,
		_w20591_,
		_w20598_,
		_w20887_
	);
	LUT3 #(
		.INIT('h07)
	) name15061 (
		_w20595_,
		_w20610_,
		_w20887_,
		_w20888_
	);
	LUT4 #(
		.INIT('h0100)
	) name15062 (
		_w20882_,
		_w20884_,
		_w20886_,
		_w20888_,
		_w20889_
	);
	LUT3 #(
		.INIT('h65)
	) name15063 (
		\u1_L5_reg[27]/NET0131 ,
		_w20879_,
		_w20889_,
		_w20890_
	);
	LUT2 #(
		.INIT('h9)
	) name15064 (
		_w20457_,
		_w20459_,
		_w20891_
	);
	LUT4 #(
		.INIT('hd003)
	) name15065 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20892_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name15066 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20893_
	);
	LUT3 #(
		.INIT('h01)
	) name15067 (
		_w20460_,
		_w20893_,
		_w20892_,
		_w20894_
	);
	LUT4 #(
		.INIT('h0800)
	) name15068 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20895_
	);
	LUT4 #(
		.INIT('hb5bc)
	) name15069 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20896_
	);
	LUT3 #(
		.INIT('h31)
	) name15070 (
		_w20460_,
		_w20895_,
		_w20896_,
		_w20897_
	);
	LUT3 #(
		.INIT('h8a)
	) name15071 (
		_w20454_,
		_w20894_,
		_w20897_,
		_w20898_
	);
	LUT3 #(
		.INIT('h40)
	) name15072 (
		_w20456_,
		_w20457_,
		_w20459_,
		_w20899_
	);
	LUT4 #(
		.INIT('hab89)
	) name15073 (
		_w20460_,
		_w20659_,
		_w20661_,
		_w20899_,
		_w20900_
	);
	LUT4 #(
		.INIT('h7bd7)
	) name15074 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20901_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15075 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20460_,
		_w20902_
	);
	LUT4 #(
		.INIT('h135f)
	) name15076 (
		_w20460_,
		_w20475_,
		_w20467_,
		_w20902_,
		_w20903_
	);
	LUT4 #(
		.INIT('hba00)
	) name15077 (
		_w20454_,
		_w20900_,
		_w20901_,
		_w20903_,
		_w20904_
	);
	LUT3 #(
		.INIT('h65)
	) name15078 (
		\u1_L5_reg[32]/NET0131 ,
		_w20898_,
		_w20904_,
		_w20905_
	);
	LUT4 #(
		.INIT('h0200)
	) name15079 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20906_
	);
	LUT4 #(
		.INIT('hbf3f)
	) name15080 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20907_
	);
	LUT3 #(
		.INIT('h20)
	) name15081 (
		_w20701_,
		_w20906_,
		_w20907_,
		_w20908_
	);
	LUT4 #(
		.INIT('h2022)
	) name15082 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20909_
	);
	LUT4 #(
		.INIT('h4f50)
	) name15083 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20910_
	);
	LUT3 #(
		.INIT('h10)
	) name15084 (
		_w20701_,
		_w20909_,
		_w20910_,
		_w20911_
	);
	LUT4 #(
		.INIT('h0001)
	) name15085 (
		_w20688_,
		_w20698_,
		_w20713_,
		_w20860_,
		_w20912_
	);
	LUT3 #(
		.INIT('he0)
	) name15086 (
		_w20908_,
		_w20911_,
		_w20912_,
		_w20913_
	);
	LUT4 #(
		.INIT('hf3af)
	) name15087 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20914_
	);
	LUT3 #(
		.INIT('h10)
	) name15088 (
		_w20701_,
		_w20909_,
		_w20914_,
		_w20915_
	);
	LUT4 #(
		.INIT('haff3)
	) name15089 (
		_w20689_,
		_w20690_,
		_w20691_,
		_w20692_,
		_w20916_
	);
	LUT3 #(
		.INIT('h20)
	) name15090 (
		_w20701_,
		_w20906_,
		_w20916_,
		_w20917_
	);
	LUT3 #(
		.INIT('h02)
	) name15091 (
		_w20688_,
		_w20694_,
		_w20715_,
		_w20918_
	);
	LUT3 #(
		.INIT('he0)
	) name15092 (
		_w20915_,
		_w20917_,
		_w20918_,
		_w20919_
	);
	LUT3 #(
		.INIT('ha9)
	) name15093 (
		\u1_L5_reg[3]/NET0131 ,
		_w20913_,
		_w20919_,
		_w20920_
	);
	LUT4 #(
		.INIT('hc693)
	) name15094 (
		decrypt_pad,
		\u1_R5_reg[13]/NET0131 ,
		\u1_uk_K_r5_reg[25]/NET0131 ,
		\u1_uk_K_r5_reg[3]/NET0131 ,
		_w20921_
	);
	LUT4 #(
		.INIT('hc693)
	) name15095 (
		decrypt_pad,
		\u1_R5_reg[9]/NET0131 ,
		\u1_uk_K_r5_reg[20]/NET0131 ,
		\u1_uk_K_r5_reg[55]/NET0131 ,
		_w20922_
	);
	LUT4 #(
		.INIT('hc963)
	) name15096 (
		decrypt_pad,
		\u1_R5_reg[11]/NET0131 ,
		\u1_uk_K_r5_reg[32]/NET0131 ,
		\u1_uk_K_r5_reg[54]/NET0131 ,
		_w20923_
	);
	LUT3 #(
		.INIT('h0b)
	) name15097 (
		_w20921_,
		_w20922_,
		_w20923_,
		_w20924_
	);
	LUT4 #(
		.INIT('hc693)
	) name15098 (
		decrypt_pad,
		\u1_R5_reg[10]/NET0131 ,
		\u1_uk_K_r5_reg[53]/NET0131 ,
		\u1_uk_K_r5_reg[6]/NET0131 ,
		_w20925_
	);
	LUT4 #(
		.INIT('hc963)
	) name15099 (
		decrypt_pad,
		\u1_R5_reg[8]/NET0131 ,
		\u1_uk_K_r5_reg[26]/NET0131 ,
		\u1_uk_K_r5_reg[48]/NET0131 ,
		_w20926_
	);
	LUT4 #(
		.INIT('h3b0b)
	) name15100 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20927_
	);
	LUT4 #(
		.INIT('h1000)
	) name15101 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20928_
	);
	LUT4 #(
		.INIT('hc693)
	) name15102 (
		decrypt_pad,
		\u1_R5_reg[12]/NET0131 ,
		\u1_uk_K_r5_reg[12]/P0001 ,
		\u1_uk_K_r5_reg[47]/NET0131 ,
		_w20929_
	);
	LUT4 #(
		.INIT('h5100)
	) name15103 (
		_w20928_,
		_w20924_,
		_w20927_,
		_w20929_,
		_w20930_
	);
	LUT2 #(
		.INIT('h8)
	) name15104 (
		_w20921_,
		_w20926_,
		_w20931_
	);
	LUT2 #(
		.INIT('h6)
	) name15105 (
		_w20921_,
		_w20926_,
		_w20932_
	);
	LUT4 #(
		.INIT('h0203)
	) name15106 (
		_w20926_,
		_w20922_,
		_w20925_,
		_w20923_,
		_w20933_
	);
	LUT2 #(
		.INIT('h8)
	) name15107 (
		_w20932_,
		_w20933_,
		_w20934_
	);
	LUT4 #(
		.INIT('h4000)
	) name15108 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20935_
	);
	LUT4 #(
		.INIT('h0400)
	) name15109 (
		_w20926_,
		_w20922_,
		_w20925_,
		_w20923_,
		_w20936_
	);
	LUT3 #(
		.INIT('h01)
	) name15110 (
		_w20929_,
		_w20936_,
		_w20935_,
		_w20937_
	);
	LUT4 #(
		.INIT('h9990)
	) name15111 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20938_
	);
	LUT4 #(
		.INIT('h0990)
	) name15112 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20939_
	);
	LUT4 #(
		.INIT('h2000)
	) name15113 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20940_
	);
	LUT3 #(
		.INIT('h23)
	) name15114 (
		_w20923_,
		_w20939_,
		_w20940_,
		_w20941_
	);
	LUT4 #(
		.INIT('h4555)
	) name15115 (
		_w20930_,
		_w20934_,
		_w20937_,
		_w20941_,
		_w20942_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15116 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20943_
	);
	LUT4 #(
		.INIT('h95b5)
	) name15117 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20944_
	);
	LUT4 #(
		.INIT('h0001)
	) name15118 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20945_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name15119 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20946_
	);
	LUT4 #(
		.INIT('h08aa)
	) name15120 (
		_w20923_,
		_w20929_,
		_w20944_,
		_w20946_,
		_w20947_
	);
	LUT3 #(
		.INIT('h56)
	) name15121 (
		\u1_L5_reg[6]/NET0131 ,
		_w20942_,
		_w20947_,
		_w20948_
	);
	LUT4 #(
		.INIT('hf126)
	) name15122 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20949_
	);
	LUT4 #(
		.INIT('h2880)
	) name15123 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20950_
	);
	LUT4 #(
		.INIT('h5004)
	) name15124 (
		_w20455_,
		_w20456_,
		_w20457_,
		_w20459_,
		_w20951_
	);
	LUT4 #(
		.INIT('h1302)
	) name15125 (
		_w20460_,
		_w20950_,
		_w20951_,
		_w20949_,
		_w20952_
	);
	LUT2 #(
		.INIT('h2)
	) name15126 (
		_w20454_,
		_w20952_,
		_w20953_
	);
	LUT2 #(
		.INIT('h4)
	) name15127 (
		_w20460_,
		_w20950_,
		_w20954_
	);
	LUT2 #(
		.INIT('h2)
	) name15128 (
		_w20454_,
		_w20460_,
		_w20955_
	);
	LUT3 #(
		.INIT('h4c)
	) name15129 (
		_w20456_,
		_w20457_,
		_w20459_,
		_w20956_
	);
	LUT4 #(
		.INIT('h8a00)
	) name15130 (
		_w20455_,
		_w20457_,
		_w20459_,
		_w20460_,
		_w20957_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name15131 (
		_w20461_,
		_w20891_,
		_w20956_,
		_w20957_,
		_w20958_
	);
	LUT3 #(
		.INIT('h45)
	) name15132 (
		_w20474_,
		_w20460_,
		_w20951_,
		_w20959_
	);
	LUT4 #(
		.INIT('h0133)
	) name15133 (
		_w20454_,
		_w20955_,
		_w20958_,
		_w20959_,
		_w20960_
	);
	LUT4 #(
		.INIT('h5556)
	) name15134 (
		\u1_L5_reg[7]/NET0131 ,
		_w20954_,
		_w20960_,
		_w20953_,
		_w20961_
	);
	LUT4 #(
		.INIT('h9b99)
	) name15135 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20962_
	);
	LUT2 #(
		.INIT('h2)
	) name15136 (
		_w20393_,
		_w20962_,
		_w20963_
	);
	LUT4 #(
		.INIT('h4010)
	) name15137 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20964_
	);
	LUT3 #(
		.INIT('he6)
	) name15138 (
		_w20395_,
		_w20396_,
		_w20397_,
		_w20965_
	);
	LUT4 #(
		.INIT('h0141)
	) name15139 (
		_w20393_,
		_w20395_,
		_w20396_,
		_w20397_,
		_w20966_
	);
	LUT4 #(
		.INIT('h0800)
	) name15140 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20967_
	);
	LUT3 #(
		.INIT('h01)
	) name15141 (
		_w20966_,
		_w20964_,
		_w20967_,
		_w20968_
	);
	LUT3 #(
		.INIT('h45)
	) name15142 (
		_w20392_,
		_w20963_,
		_w20968_,
		_w20969_
	);
	LUT4 #(
		.INIT('hf77f)
	) name15143 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20970_
	);
	LUT2 #(
		.INIT('h1)
	) name15144 (
		_w20393_,
		_w20970_,
		_w20971_
	);
	LUT4 #(
		.INIT('h9060)
	) name15145 (
		_w20395_,
		_w20396_,
		_w20394_,
		_w20397_,
		_w20972_
	);
	LUT4 #(
		.INIT('h0031)
	) name15146 (
		_w20408_,
		_w20490_,
		_w20965_,
		_w20972_,
		_w20973_
	);
	LUT3 #(
		.INIT('h31)
	) name15147 (
		_w20392_,
		_w20971_,
		_w20973_,
		_w20974_
	);
	LUT3 #(
		.INIT('h65)
	) name15148 (
		\u1_L5_reg[9]/NET0131 ,
		_w20969_,
		_w20974_,
		_w20975_
	);
	LUT3 #(
		.INIT('h80)
	) name15149 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20976_
	);
	LUT4 #(
		.INIT('h6979)
	) name15150 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20923_,
		_w20977_
	);
	LUT2 #(
		.INIT('h1)
	) name15151 (
		_w20925_,
		_w20977_,
		_w20978_
	);
	LUT4 #(
		.INIT('h0014)
	) name15152 (
		_w20921_,
		_w20926_,
		_w20925_,
		_w20923_,
		_w20979_
	);
	LUT3 #(
		.INIT('h02)
	) name15153 (
		_w20929_,
		_w20940_,
		_w20979_,
		_w20980_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name15154 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20981_
	);
	LUT2 #(
		.INIT('h1)
	) name15155 (
		_w20923_,
		_w20981_,
		_w20982_
	);
	LUT4 #(
		.INIT('h6800)
	) name15156 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20923_,
		_w20983_
	);
	LUT3 #(
		.INIT('h01)
	) name15157 (
		_w20929_,
		_w20945_,
		_w20983_,
		_w20984_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15158 (
		_w20978_,
		_w20980_,
		_w20982_,
		_w20984_,
		_w20985_
	);
	LUT4 #(
		.INIT('hbeff)
	) name15159 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w20986_
	);
	LUT4 #(
		.INIT('h0020)
	) name15160 (
		_w20926_,
		_w20922_,
		_w20925_,
		_w20923_,
		_w20987_
	);
	LUT3 #(
		.INIT('h0d)
	) name15161 (
		_w20923_,
		_w20986_,
		_w20987_,
		_w20988_
	);
	LUT3 #(
		.INIT('h65)
	) name15162 (
		\u1_L5_reg[16]/NET0131 ,
		_w20985_,
		_w20988_,
		_w20989_
	);
	LUT4 #(
		.INIT('h2028)
	) name15163 (
		_w20545_,
		_w20539_,
		_w20540_,
		_w20542_,
		_w20990_
	);
	LUT4 #(
		.INIT('he4ff)
	) name15164 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20991_
	);
	LUT4 #(
		.INIT('h0032)
	) name15165 (
		_w20545_,
		_w20567_,
		_w20991_,
		_w20990_,
		_w20992_
	);
	LUT4 #(
		.INIT('h0043)
	) name15166 (
		_w20545_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20993_
	);
	LUT4 #(
		.INIT('h6000)
	) name15167 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20994_
	);
	LUT4 #(
		.INIT('h8000)
	) name15168 (
		_w20545_,
		_w20539_,
		_w20540_,
		_w20542_,
		_w20995_
	);
	LUT4 #(
		.INIT('h0001)
	) name15169 (
		_w20562_,
		_w20995_,
		_w20994_,
		_w20993_,
		_w20996_
	);
	LUT4 #(
		.INIT('h0040)
	) name15170 (
		_w20545_,
		_w20539_,
		_w20540_,
		_w20542_,
		_w20997_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name15171 (
		_w20539_,
		_w20540_,
		_w20538_,
		_w20542_,
		_w20998_
	);
	LUT3 #(
		.INIT('h31)
	) name15172 (
		_w20545_,
		_w20997_,
		_w20998_,
		_w20999_
	);
	LUT4 #(
		.INIT('hd800)
	) name15173 (
		_w20547_,
		_w20992_,
		_w20996_,
		_w20999_,
		_w21000_
	);
	LUT2 #(
		.INIT('h9)
	) name15174 (
		\u1_L5_reg[18]/NET0131 ,
		_w21000_,
		_w21001_
	);
	LUT4 #(
		.INIT('h1df2)
	) name15175 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w21002_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15176 (
		_w20923_,
		_w20932_,
		_w20933_,
		_w21002_,
		_w21003_
	);
	LUT2 #(
		.INIT('h2)
	) name15177 (
		_w20929_,
		_w21003_,
		_w21004_
	);
	LUT3 #(
		.INIT('hed)
	) name15178 (
		_w20921_,
		_w20926_,
		_w20925_,
		_w21005_
	);
	LUT4 #(
		.INIT('he2cd)
	) name15179 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w21006_
	);
	LUT4 #(
		.INIT('h0400)
	) name15180 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w21007_
	);
	LUT4 #(
		.INIT('h3302)
	) name15181 (
		_w20923_,
		_w20929_,
		_w21006_,
		_w21007_,
		_w21008_
	);
	LUT4 #(
		.INIT('h0009)
	) name15182 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w21009_
	);
	LUT3 #(
		.INIT('h04)
	) name15183 (
		_w20929_,
		_w20943_,
		_w21009_,
		_w21010_
	);
	LUT3 #(
		.INIT('h51)
	) name15184 (
		_w20923_,
		_w20929_,
		_w20938_,
		_w21011_
	);
	LUT2 #(
		.INIT('h2)
	) name15185 (
		_w20925_,
		_w20923_,
		_w21012_
	);
	LUT3 #(
		.INIT('hd0)
	) name15186 (
		_w20921_,
		_w20922_,
		_w20923_,
		_w21013_
	);
	LUT4 #(
		.INIT('h0026)
	) name15187 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w21014_
	);
	LUT4 #(
		.INIT('h0777)
	) name15188 (
		_w20976_,
		_w21012_,
		_w21013_,
		_w21014_,
		_w21015_
	);
	LUT4 #(
		.INIT('h4500)
	) name15189 (
		_w21008_,
		_w21010_,
		_w21011_,
		_w21015_,
		_w21016_
	);
	LUT3 #(
		.INIT('h65)
	) name15190 (
		\u1_L5_reg[24]/NET0131 ,
		_w21004_,
		_w21016_,
		_w21017_
	);
	LUT3 #(
		.INIT('h04)
	) name15191 (
		_w20921_,
		_w20922_,
		_w20925_,
		_w21018_
	);
	LUT4 #(
		.INIT('h8c00)
	) name15192 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w21019_
	);
	LUT3 #(
		.INIT('h01)
	) name15193 (
		_w20929_,
		_w21019_,
		_w21018_,
		_w21020_
	);
	LUT4 #(
		.INIT('h0004)
	) name15194 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w21021_
	);
	LUT4 #(
		.INIT('haa2a)
	) name15195 (
		_w20923_,
		_w20929_,
		_w21005_,
		_w21021_,
		_w21022_
	);
	LUT2 #(
		.INIT('h4)
	) name15196 (
		_w21020_,
		_w21022_,
		_w21023_
	);
	LUT4 #(
		.INIT('hdd02)
	) name15197 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20925_,
		_w21024_
	);
	LUT4 #(
		.INIT('hf450)
	) name15198 (
		_w20921_,
		_w20926_,
		_w20922_,
		_w20923_,
		_w21025_
	);
	LUT3 #(
		.INIT('h01)
	) name15199 (
		_w20929_,
		_w21024_,
		_w21025_,
		_w21026_
	);
	LUT3 #(
		.INIT('h23)
	) name15200 (
		_w20926_,
		_w20925_,
		_w20929_,
		_w21027_
	);
	LUT3 #(
		.INIT('h04)
	) name15201 (
		_w20921_,
		_w20922_,
		_w20923_,
		_w21028_
	);
	LUT2 #(
		.INIT('h4)
	) name15202 (
		_w21027_,
		_w21028_,
		_w21029_
	);
	LUT4 #(
		.INIT('h8880)
	) name15203 (
		_w20926_,
		_w20925_,
		_w20923_,
		_w20929_,
		_w21030_
	);
	LUT3 #(
		.INIT('h80)
	) name15204 (
		_w20922_,
		_w20925_,
		_w20929_,
		_w21031_
	);
	LUT4 #(
		.INIT('h8acf)
	) name15205 (
		_w20931_,
		_w21013_,
		_w21030_,
		_w21031_,
		_w21032_
	);
	LUT3 #(
		.INIT('h10)
	) name15206 (
		_w21026_,
		_w21029_,
		_w21032_,
		_w21033_
	);
	LUT3 #(
		.INIT('h9a)
	) name15207 (
		\u1_L5_reg[30]/NET0131 ,
		_w21023_,
		_w21033_,
		_w21034_
	);
	LUT4 #(
		.INIT('hc963)
	) name15208 (
		decrypt_pad,
		\u1_R4_reg[28]/NET0131 ,
		\u1_uk_K_r4_reg[31]/P0001 ,
		\u1_uk_K_r4_reg[50]/NET0131 ,
		_w21035_
	);
	LUT4 #(
		.INIT('hc693)
	) name15209 (
		decrypt_pad,
		\u1_R4_reg[24]/NET0131 ,
		\u1_uk_K_r4_reg[38]/NET0131 ,
		\u1_uk_K_r4_reg[42]/NET0131 ,
		_w21036_
	);
	LUT4 #(
		.INIT('hc693)
	) name15210 (
		decrypt_pad,
		\u1_R4_reg[26]/NET0131 ,
		\u1_uk_K_r4_reg[30]/NET0131 ,
		\u1_uk_K_r4_reg[7]/NET0131 ,
		_w21037_
	);
	LUT4 #(
		.INIT('hc693)
	) name15211 (
		decrypt_pad,
		\u1_R4_reg[25]/NET0131 ,
		\u1_uk_K_r4_reg[14]/NET0131 ,
		\u1_uk_K_r4_reg[22]/NET0131 ,
		_w21038_
	);
	LUT4 #(
		.INIT('hc963)
	) name15212 (
		decrypt_pad,
		\u1_R4_reg[27]/NET0131 ,
		\u1_uk_K_r4_reg[16]/NET0131 ,
		\u1_uk_K_r4_reg[8]/NET0131 ,
		_w21039_
	);
	LUT4 #(
		.INIT('hc693)
	) name15213 (
		decrypt_pad,
		\u1_R4_reg[29]/NET0131 ,
		\u1_uk_K_r4_reg[42]/NET0131 ,
		\u1_uk_K_r4_reg[50]/NET0131 ,
		_w21040_
	);
	LUT4 #(
		.INIT('hfc3a)
	) name15214 (
		_w21040_,
		_w21038_,
		_w21037_,
		_w21039_,
		_w21041_
	);
	LUT2 #(
		.INIT('h2)
	) name15215 (
		_w21036_,
		_w21041_,
		_w21042_
	);
	LUT4 #(
		.INIT('h0100)
	) name15216 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21043_
	);
	LUT2 #(
		.INIT('h6)
	) name15217 (
		_w21036_,
		_w21037_,
		_w21044_
	);
	LUT3 #(
		.INIT('h8a)
	) name15218 (
		_w21040_,
		_w21038_,
		_w21039_,
		_w21045_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name15219 (
		_w21043_,
		_w21039_,
		_w21044_,
		_w21045_,
		_w21046_
	);
	LUT4 #(
		.INIT('h0100)
	) name15220 (
		_w21040_,
		_w21038_,
		_w21037_,
		_w21039_,
		_w21047_
	);
	LUT4 #(
		.INIT('h0082)
	) name15221 (
		_w21038_,
		_w21036_,
		_w21037_,
		_w21039_,
		_w21048_
	);
	LUT2 #(
		.INIT('h1)
	) name15222 (
		_w21047_,
		_w21048_,
		_w21049_
	);
	LUT4 #(
		.INIT('hba00)
	) name15223 (
		_w21035_,
		_w21042_,
		_w21046_,
		_w21049_,
		_w21050_
	);
	LUT4 #(
		.INIT('hf47c)
	) name15224 (
		_w21035_,
		_w21040_,
		_w21038_,
		_w21037_,
		_w21051_
	);
	LUT4 #(
		.INIT('h0600)
	) name15225 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21052_
	);
	LUT4 #(
		.INIT('hcc08)
	) name15226 (
		_w21036_,
		_w21039_,
		_w21051_,
		_w21052_,
		_w21053_
	);
	LUT2 #(
		.INIT('h2)
	) name15227 (
		_w21040_,
		_w21036_,
		_w21054_
	);
	LUT4 #(
		.INIT('hf700)
	) name15228 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21055_
	);
	LUT3 #(
		.INIT('h20)
	) name15229 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21056_
	);
	LUT4 #(
		.INIT('h0028)
	) name15230 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21039_,
		_w21057_
	);
	LUT4 #(
		.INIT('h0200)
	) name15231 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21058_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name15232 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21059_
	);
	LUT4 #(
		.INIT('h20aa)
	) name15233 (
		_w21035_,
		_w21055_,
		_w21057_,
		_w21059_,
		_w21060_
	);
	LUT2 #(
		.INIT('h1)
	) name15234 (
		_w21053_,
		_w21060_,
		_w21061_
	);
	LUT3 #(
		.INIT('h95)
	) name15235 (
		\u1_L4_reg[22]/NET0131 ,
		_w21050_,
		_w21061_,
		_w21062_
	);
	LUT4 #(
		.INIT('hc693)
	) name15236 (
		decrypt_pad,
		\u1_R4_reg[4]/NET0131 ,
		\u1_uk_K_r4_reg[19]/NET0131 ,
		\u1_uk_K_r4_reg[25]/NET0131 ,
		_w21063_
	);
	LUT4 #(
		.INIT('hc693)
	) name15237 (
		decrypt_pad,
		\u1_R4_reg[3]/NET0131 ,
		\u1_uk_K_r4_reg[41]/NET0131 ,
		\u1_uk_K_r4_reg[47]/NET0131 ,
		_w21064_
	);
	LUT4 #(
		.INIT('hc693)
	) name15238 (
		decrypt_pad,
		\u1_R4_reg[5]/NET0131 ,
		\u1_uk_K_r4_reg[47]/NET0131 ,
		\u1_uk_K_r4_reg[53]/NET0131 ,
		_w21065_
	);
	LUT4 #(
		.INIT('hc693)
	) name15239 (
		decrypt_pad,
		\u1_R4_reg[1]/NET0131 ,
		\u1_uk_K_r4_reg[17]/NET0131 ,
		\u1_uk_K_r4_reg[55]/NET0131 ,
		_w21066_
	);
	LUT4 #(
		.INIT('hc963)
	) name15240 (
		decrypt_pad,
		\u1_R4_reg[2]/NET0131 ,
		\u1_uk_K_r4_reg[13]/NET0131 ,
		\u1_uk_K_r4_reg[32]/NET0131 ,
		_w21067_
	);
	LUT4 #(
		.INIT('hc963)
	) name15241 (
		decrypt_pad,
		\u1_R4_reg[32]/NET0131 ,
		\u1_uk_K_r4_reg[34]/NET0131 ,
		\u1_uk_K_r4_reg[53]/NET0131 ,
		_w21068_
	);
	LUT4 #(
		.INIT('hfd0d)
	) name15242 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21069_
	);
	LUT2 #(
		.INIT('h2)
	) name15243 (
		_w21064_,
		_w21069_,
		_w21070_
	);
	LUT2 #(
		.INIT('h4)
	) name15244 (
		_w21068_,
		_w21065_,
		_w21071_
	);
	LUT2 #(
		.INIT('h2)
	) name15245 (
		_w21064_,
		_w21067_,
		_w21072_
	);
	LUT3 #(
		.INIT('hd0)
	) name15246 (
		_w21064_,
		_w21067_,
		_w21066_,
		_w21073_
	);
	LUT2 #(
		.INIT('h2)
	) name15247 (
		_w21071_,
		_w21073_,
		_w21074_
	);
	LUT3 #(
		.INIT('h02)
	) name15248 (
		_w21067_,
		_w21068_,
		_w21066_,
		_w21075_
	);
	LUT4 #(
		.INIT('h0004)
	) name15249 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21076_
	);
	LUT3 #(
		.INIT('h40)
	) name15250 (
		_w21064_,
		_w21068_,
		_w21066_,
		_w21077_
	);
	LUT3 #(
		.INIT('h01)
	) name15251 (
		_w21076_,
		_w21077_,
		_w21075_,
		_w21078_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15252 (
		_w21063_,
		_w21070_,
		_w21074_,
		_w21078_,
		_w21079_
	);
	LUT4 #(
		.INIT('heef6)
	) name15253 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21080_
	);
	LUT2 #(
		.INIT('h1)
	) name15254 (
		_w21064_,
		_w21080_,
		_w21081_
	);
	LUT3 #(
		.INIT('h60)
	) name15255 (
		_w21068_,
		_w21065_,
		_w21066_,
		_w21082_
	);
	LUT4 #(
		.INIT('h7c3f)
	) name15256 (
		_w21064_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21083_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name15257 (
		_w21064_,
		_w21067_,
		_w21082_,
		_w21083_,
		_w21084_
	);
	LUT3 #(
		.INIT('h45)
	) name15258 (
		_w21063_,
		_w21081_,
		_w21084_,
		_w21085_
	);
	LUT3 #(
		.INIT('h80)
	) name15259 (
		_w21068_,
		_w21065_,
		_w21066_,
		_w21086_
	);
	LUT4 #(
		.INIT('h0020)
	) name15260 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21087_
	);
	LUT4 #(
		.INIT('h7adf)
	) name15261 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21088_
	);
	LUT2 #(
		.INIT('h1)
	) name15262 (
		_w21064_,
		_w21088_,
		_w21089_
	);
	LUT4 #(
		.INIT('h0020)
	) name15263 (
		_w21064_,
		_w21067_,
		_w21068_,
		_w21066_,
		_w21090_
	);
	LUT2 #(
		.INIT('h2)
	) name15264 (
		_w21064_,
		_w21065_,
		_w21091_
	);
	LUT3 #(
		.INIT('h13)
	) name15265 (
		_w21075_,
		_w21090_,
		_w21091_,
		_w21092_
	);
	LUT2 #(
		.INIT('h4)
	) name15266 (
		_w21089_,
		_w21092_,
		_w21093_
	);
	LUT4 #(
		.INIT('h5655)
	) name15267 (
		\u1_L4_reg[31]/NET0131 ,
		_w21085_,
		_w21079_,
		_w21093_,
		_w21094_
	);
	LUT4 #(
		.INIT('hc693)
	) name15268 (
		decrypt_pad,
		\u1_R4_reg[24]/NET0131 ,
		\u1_uk_K_r4_reg[43]/NET0131 ,
		\u1_uk_K_r4_reg[51]/NET0131 ,
		_w21095_
	);
	LUT4 #(
		.INIT('hc693)
	) name15269 (
		decrypt_pad,
		\u1_R4_reg[22]/NET0131 ,
		\u1_uk_K_r4_reg[28]/NET0131 ,
		\u1_uk_K_r4_reg[36]/NET0131 ,
		_w21096_
	);
	LUT4 #(
		.INIT('hc693)
	) name15270 (
		decrypt_pad,
		\u1_R4_reg[20]/NET0131 ,
		\u1_uk_K_r4_reg[22]/NET0131 ,
		\u1_uk_K_r4_reg[30]/NET0131 ,
		_w21097_
	);
	LUT4 #(
		.INIT('hc963)
	) name15271 (
		decrypt_pad,
		\u1_R4_reg[21]/NET0131 ,
		\u1_uk_K_r4_reg[14]/NET0131 ,
		\u1_uk_K_r4_reg[37]/NET0131 ,
		_w21098_
	);
	LUT4 #(
		.INIT('hc963)
	) name15272 (
		decrypt_pad,
		\u1_R4_reg[25]/NET0131 ,
		\u1_uk_K_r4_reg[15]/NET0131 ,
		\u1_uk_K_r4_reg[7]/NET0131 ,
		_w21099_
	);
	LUT4 #(
		.INIT('hd080)
	) name15273 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21100_
	);
	LUT4 #(
		.INIT('hc693)
	) name15274 (
		decrypt_pad,
		\u1_R4_reg[23]/NET0131 ,
		\u1_uk_K_r4_reg[45]/NET0131 ,
		\u1_uk_K_r4_reg[49]/NET0131 ,
		_w21101_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name15275 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21102_
	);
	LUT3 #(
		.INIT('h01)
	) name15276 (
		_w21101_,
		_w21102_,
		_w21100_,
		_w21103_
	);
	LUT4 #(
		.INIT('h0002)
	) name15277 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21104_
	);
	LUT4 #(
		.INIT('h27fd)
	) name15278 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21105_
	);
	LUT4 #(
		.INIT('h0008)
	) name15279 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21101_,
		_w21106_
	);
	LUT2 #(
		.INIT('h4)
	) name15280 (
		_w21098_,
		_w21106_,
		_w21107_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name15281 (
		_w21098_,
		_w21101_,
		_w21105_,
		_w21106_,
		_w21108_
	);
	LUT3 #(
		.INIT('h8a)
	) name15282 (
		_w21095_,
		_w21103_,
		_w21108_,
		_w21109_
	);
	LUT4 #(
		.INIT('h0060)
	) name15283 (
		_w21097_,
		_w21096_,
		_w21098_,
		_w21101_,
		_w21110_
	);
	LUT4 #(
		.INIT('hf010)
	) name15284 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21111_
	);
	LUT3 #(
		.INIT('hd0)
	) name15285 (
		_w21097_,
		_w21096_,
		_w21101_,
		_w21112_
	);
	LUT2 #(
		.INIT('h4)
	) name15286 (
		_w21111_,
		_w21112_,
		_w21113_
	);
	LUT4 #(
		.INIT('h0200)
	) name15287 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21114_
	);
	LUT4 #(
		.INIT('h0002)
	) name15288 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21101_,
		_w21115_
	);
	LUT4 #(
		.INIT('h0080)
	) name15289 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21116_
	);
	LUT3 #(
		.INIT('h01)
	) name15290 (
		_w21114_,
		_w21115_,
		_w21116_,
		_w21117_
	);
	LUT4 #(
		.INIT('h5455)
	) name15291 (
		_w21095_,
		_w21113_,
		_w21110_,
		_w21117_,
		_w21118_
	);
	LUT3 #(
		.INIT('h04)
	) name15292 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21119_
	);
	LUT4 #(
		.INIT('h0004)
	) name15293 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21120_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name15294 (
		_w21098_,
		_w21101_,
		_w21115_,
		_w21119_,
		_w21121_
	);
	LUT4 #(
		.INIT('h0001)
	) name15295 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21101_,
		_w21122_
	);
	LUT3 #(
		.INIT('hb0)
	) name15296 (
		_w21097_,
		_w21099_,
		_w21101_,
		_w21123_
	);
	LUT4 #(
		.INIT('hc5c4)
	) name15297 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21124_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name15298 (
		_w21098_,
		_w21122_,
		_w21123_,
		_w21124_,
		_w21125_
	);
	LUT2 #(
		.INIT('h8)
	) name15299 (
		_w21121_,
		_w21125_,
		_w21126_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name15300 (
		\u1_L4_reg[11]/P0001 ,
		_w21118_,
		_w21109_,
		_w21126_,
		_w21127_
	);
	LUT4 #(
		.INIT('hc963)
	) name15301 (
		decrypt_pad,
		\u1_R4_reg[13]/NET0131 ,
		\u1_uk_K_r4_reg[10]/NET0131 ,
		\u1_uk_K_r4_reg[4]/NET0131 ,
		_w21128_
	);
	LUT4 #(
		.INIT('hc693)
	) name15302 (
		decrypt_pad,
		\u1_R4_reg[17]/NET0131 ,
		\u1_uk_K_r4_reg[26]/NET0131 ,
		\u1_uk_K_r4_reg[32]/NET0131 ,
		_w21129_
	);
	LUT4 #(
		.INIT('hc693)
	) name15303 (
		decrypt_pad,
		\u1_R4_reg[12]/NET0131 ,
		\u1_uk_K_r4_reg[10]/NET0131 ,
		\u1_uk_K_r4_reg[48]/NET0131 ,
		_w21130_
	);
	LUT4 #(
		.INIT('hc693)
	) name15304 (
		decrypt_pad,
		\u1_R4_reg[15]/NET0131 ,
		\u1_uk_K_r4_reg[13]/NET0131 ,
		\u1_uk_K_r4_reg[19]/NET0131 ,
		_w21131_
	);
	LUT4 #(
		.INIT('h7e00)
	) name15305 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21131_,
		_w21132_
	);
	LUT4 #(
		.INIT('hc963)
	) name15306 (
		decrypt_pad,
		\u1_R4_reg[14]/NET0131 ,
		\u1_uk_K_r4_reg[11]/NET0131 ,
		\u1_uk_K_r4_reg[5]/NET0131 ,
		_w21133_
	);
	LUT3 #(
		.INIT('h40)
	) name15307 (
		_w21129_,
		_w21130_,
		_w21133_,
		_w21134_
	);
	LUT3 #(
		.INIT('h0d)
	) name15308 (
		_w21129_,
		_w21128_,
		_w21131_,
		_w21135_
	);
	LUT3 #(
		.INIT('h45)
	) name15309 (
		_w21132_,
		_w21134_,
		_w21135_,
		_w21136_
	);
	LUT2 #(
		.INIT('h1)
	) name15310 (
		_w21129_,
		_w21130_,
		_w21137_
	);
	LUT3 #(
		.INIT('h10)
	) name15311 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21138_
	);
	LUT3 #(
		.INIT('h01)
	) name15312 (
		_w21129_,
		_w21130_,
		_w21133_,
		_w21139_
	);
	LUT4 #(
		.INIT('h0001)
	) name15313 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21140_
	);
	LUT4 #(
		.INIT('heffe)
	) name15314 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21141_
	);
	LUT4 #(
		.INIT('h0008)
	) name15315 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21142_
	);
	LUT4 #(
		.INIT('hc963)
	) name15316 (
		decrypt_pad,
		\u1_R4_reg[16]/NET0131 ,
		\u1_uk_K_r4_reg[27]/P0001 ,
		\u1_uk_K_r4_reg[46]/NET0131 ,
		_w21143_
	);
	LUT3 #(
		.INIT('h80)
	) name15317 (
		_w21128_,
		_w21133_,
		_w21131_,
		_w21144_
	);
	LUT4 #(
		.INIT('h4000)
	) name15318 (
		_w21130_,
		_w21128_,
		_w21133_,
		_w21131_,
		_w21145_
	);
	LUT4 #(
		.INIT('h0002)
	) name15319 (
		_w21141_,
		_w21143_,
		_w21145_,
		_w21142_,
		_w21146_
	);
	LUT2 #(
		.INIT('h4)
	) name15320 (
		_w21136_,
		_w21146_,
		_w21147_
	);
	LUT4 #(
		.INIT('h0001)
	) name15321 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21131_,
		_w21148_
	);
	LUT2 #(
		.INIT('h8)
	) name15322 (
		_w21133_,
		_w21148_,
		_w21149_
	);
	LUT2 #(
		.INIT('h2)
	) name15323 (
		_w21129_,
		_w21130_,
		_w21150_
	);
	LUT4 #(
		.INIT('h0200)
	) name15324 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21131_,
		_w21151_
	);
	LUT4 #(
		.INIT('h4000)
	) name15325 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21131_,
		_w21152_
	);
	LUT3 #(
		.INIT('h02)
	) name15326 (
		_w21143_,
		_w21152_,
		_w21151_,
		_w21153_
	);
	LUT4 #(
		.INIT('h0020)
	) name15327 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21154_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name15328 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21155_
	);
	LUT4 #(
		.INIT('h0006)
	) name15329 (
		_w21130_,
		_w21128_,
		_w21133_,
		_w21131_,
		_w21156_
	);
	LUT2 #(
		.INIT('h2)
	) name15330 (
		_w21155_,
		_w21156_,
		_w21157_
	);
	LUT3 #(
		.INIT('h40)
	) name15331 (
		_w21149_,
		_w21153_,
		_w21157_,
		_w21158_
	);
	LUT4 #(
		.INIT('h0400)
	) name15332 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21159_
	);
	LUT4 #(
		.INIT('hfcb8)
	) name15333 (
		_w21140_,
		_w21131_,
		_w21154_,
		_w21159_,
		_w21160_
	);
	LUT2 #(
		.INIT('h4)
	) name15334 (
		_w21133_,
		_w21152_,
		_w21161_
	);
	LUT2 #(
		.INIT('h1)
	) name15335 (
		_w21160_,
		_w21161_,
		_w21162_
	);
	LUT4 #(
		.INIT('ha955)
	) name15336 (
		\u1_L4_reg[20]/NET0131 ,
		_w21147_,
		_w21158_,
		_w21162_,
		_w21163_
	);
	LUT4 #(
		.INIT('hc963)
	) name15337 (
		decrypt_pad,
		\u1_R4_reg[28]/NET0131 ,
		\u1_uk_K_r4_reg[1]/NET0131 ,
		\u1_uk_K_r4_reg[52]/NET0131 ,
		_w21164_
	);
	LUT4 #(
		.INIT('hc693)
	) name15338 (
		decrypt_pad,
		\u1_R4_reg[30]/NET0131 ,
		\u1_uk_K_r4_reg[21]/NET0131 ,
		\u1_uk_K_r4_reg[29]/NET0131 ,
		_w21165_
	);
	LUT4 #(
		.INIT('hc963)
	) name15339 (
		decrypt_pad,
		\u1_R4_reg[29]/NET0131 ,
		\u1_uk_K_r4_reg[28]/NET0131 ,
		\u1_uk_K_r4_reg[51]/NET0131 ,
		_w21166_
	);
	LUT4 #(
		.INIT('hc693)
	) name15340 (
		decrypt_pad,
		\u1_R4_reg[1]/NET0131 ,
		\u1_uk_K_r4_reg[36]/NET0131 ,
		\u1_uk_K_r4_reg[44]/NET0131 ,
		_w21167_
	);
	LUT4 #(
		.INIT('hc963)
	) name15341 (
		decrypt_pad,
		\u1_R4_reg[31]/P0001 ,
		\u1_uk_K_r4_reg[45]/NET0131 ,
		\u1_uk_K_r4_reg[9]/NET0131 ,
		_w21168_
	);
	LUT2 #(
		.INIT('h1)
	) name15342 (
		_w21165_,
		_w21168_,
		_w21169_
	);
	LUT4 #(
		.INIT('h7d4c)
	) name15343 (
		_w21166_,
		_w21165_,
		_w21167_,
		_w21168_,
		_w21170_
	);
	LUT2 #(
		.INIT('h2)
	) name15344 (
		_w21164_,
		_w21170_,
		_w21171_
	);
	LUT4 #(
		.INIT('h0020)
	) name15345 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21172_
	);
	LUT4 #(
		.INIT('heedf)
	) name15346 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21173_
	);
	LUT3 #(
		.INIT('h0b)
	) name15347 (
		_w21164_,
		_w21165_,
		_w21167_,
		_w21174_
	);
	LUT3 #(
		.INIT('h0b)
	) name15348 (
		_w21166_,
		_w21167_,
		_w21168_,
		_w21175_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15349 (
		_w21173_,
		_w21168_,
		_w21174_,
		_w21175_,
		_w21176_
	);
	LUT4 #(
		.INIT('hc693)
	) name15350 (
		decrypt_pad,
		\u1_R4_reg[32]/NET0131 ,
		\u1_uk_K_r4_reg[15]/NET0131 ,
		\u1_uk_K_r4_reg[23]/P0001 ,
		_w21177_
	);
	LUT3 #(
		.INIT('h0b)
	) name15351 (
		_w21171_,
		_w21176_,
		_w21177_,
		_w21178_
	);
	LUT4 #(
		.INIT('h0008)
	) name15352 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21179_
	);
	LUT4 #(
		.INIT('hf531)
	) name15353 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21180_
	);
	LUT3 #(
		.INIT('h02)
	) name15354 (
		_w21168_,
		_w21180_,
		_w21179_,
		_w21181_
	);
	LUT4 #(
		.INIT('h4000)
	) name15355 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21182_
	);
	LUT4 #(
		.INIT('h0001)
	) name15356 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21168_,
		_w21183_
	);
	LUT2 #(
		.INIT('h1)
	) name15357 (
		_w21182_,
		_w21183_,
		_w21184_
	);
	LUT3 #(
		.INIT('h8a)
	) name15358 (
		_w21177_,
		_w21181_,
		_w21184_,
		_w21185_
	);
	LUT4 #(
		.INIT('h0240)
	) name15359 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21186_
	);
	LUT4 #(
		.INIT('h0001)
	) name15360 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21187_
	);
	LUT4 #(
		.INIT('h1000)
	) name15361 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21188_
	);
	LUT4 #(
		.INIT('hedbe)
	) name15362 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21189_
	);
	LUT2 #(
		.INIT('h2)
	) name15363 (
		_w21168_,
		_w21189_,
		_w21190_
	);
	LUT3 #(
		.INIT('h08)
	) name15364 (
		_w21164_,
		_w21166_,
		_w21167_,
		_w21191_
	);
	LUT3 #(
		.INIT('h20)
	) name15365 (
		_w21164_,
		_w21166_,
		_w21177_,
		_w21192_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15366 (
		_w21165_,
		_w21168_,
		_w21191_,
		_w21192_,
		_w21193_
	);
	LUT2 #(
		.INIT('h4)
	) name15367 (
		_w21190_,
		_w21193_,
		_w21194_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name15368 (
		\u1_L4_reg[5]/NET0131 ,
		_w21178_,
		_w21185_,
		_w21194_,
		_w21195_
	);
	LUT4 #(
		.INIT('h4404)
	) name15369 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21196_
	);
	LUT3 #(
		.INIT('h01)
	) name15370 (
		_w21131_,
		_w21154_,
		_w21196_,
		_w21197_
	);
	LUT3 #(
		.INIT('h04)
	) name15371 (
		_w21138_,
		_w21131_,
		_w21142_,
		_w21198_
	);
	LUT4 #(
		.INIT('h8200)
	) name15372 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21199_
	);
	LUT4 #(
		.INIT('haa02)
	) name15373 (
		_w21143_,
		_w21197_,
		_w21198_,
		_w21199_,
		_w21200_
	);
	LUT4 #(
		.INIT('h0008)
	) name15374 (
		_w21129_,
		_w21130_,
		_w21133_,
		_w21131_,
		_w21201_
	);
	LUT3 #(
		.INIT('h08)
	) name15375 (
		_w21130_,
		_w21128_,
		_w21133_,
		_w21202_
	);
	LUT3 #(
		.INIT('h01)
	) name15376 (
		_w21148_,
		_w21201_,
		_w21202_,
		_w21203_
	);
	LUT4 #(
		.INIT('h0200)
	) name15377 (
		_w21129_,
		_w21130_,
		_w21133_,
		_w21131_,
		_w21204_
	);
	LUT2 #(
		.INIT('h2)
	) name15378 (
		_w21129_,
		_w21133_,
		_w21205_
	);
	LUT3 #(
		.INIT('h20)
	) name15379 (
		_w21130_,
		_w21128_,
		_w21131_,
		_w21206_
	);
	LUT3 #(
		.INIT('h45)
	) name15380 (
		_w21204_,
		_w21205_,
		_w21206_,
		_w21207_
	);
	LUT4 #(
		.INIT('h1333)
	) name15381 (
		_w21141_,
		_w21143_,
		_w21203_,
		_w21207_,
		_w21208_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name15382 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21209_
	);
	LUT2 #(
		.INIT('h1)
	) name15383 (
		_w21131_,
		_w21209_,
		_w21210_
	);
	LUT3 #(
		.INIT('h23)
	) name15384 (
		_w21133_,
		_w21145_,
		_w21152_,
		_w21211_
	);
	LUT2 #(
		.INIT('h4)
	) name15385 (
		_w21210_,
		_w21211_,
		_w21212_
	);
	LUT4 #(
		.INIT('h5655)
	) name15386 (
		\u1_L4_reg[10]/NET0131 ,
		_w21200_,
		_w21208_,
		_w21212_,
		_w21213_
	);
	LUT3 #(
		.INIT('h09)
	) name15387 (
		_w21040_,
		_w21038_,
		_w21039_,
		_w21214_
	);
	LUT4 #(
		.INIT('h0004)
	) name15388 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21215_
	);
	LUT3 #(
		.INIT('h27)
	) name15389 (
		_w21038_,
		_w21037_,
		_w21039_,
		_w21216_
	);
	LUT4 #(
		.INIT('h0031)
	) name15390 (
		_w21054_,
		_w21215_,
		_w21216_,
		_w21214_,
		_w21217_
	);
	LUT3 #(
		.INIT('h04)
	) name15391 (
		_w21040_,
		_w21036_,
		_w21037_,
		_w21218_
	);
	LUT4 #(
		.INIT('h2010)
	) name15392 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21219_
	);
	LUT3 #(
		.INIT('h08)
	) name15393 (
		_w21036_,
		_w21037_,
		_w21039_,
		_w21220_
	);
	LUT4 #(
		.INIT('h0001)
	) name15394 (
		_w21035_,
		_w21043_,
		_w21219_,
		_w21220_,
		_w21221_
	);
	LUT2 #(
		.INIT('h9)
	) name15395 (
		_w21040_,
		_w21036_,
		_w21222_
	);
	LUT4 #(
		.INIT('h4050)
	) name15396 (
		_w21038_,
		_w21036_,
		_w21037_,
		_w21039_,
		_w21223_
	);
	LUT4 #(
		.INIT('h0400)
	) name15397 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21224_
	);
	LUT4 #(
		.INIT('h2022)
	) name15398 (
		_w21035_,
		_w21224_,
		_w21222_,
		_w21223_,
		_w21225_
	);
	LUT4 #(
		.INIT('h0028)
	) name15399 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21226_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name15400 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21227_
	);
	LUT3 #(
		.INIT('h31)
	) name15401 (
		_w21039_,
		_w21226_,
		_w21227_,
		_w21228_
	);
	LUT4 #(
		.INIT('h0777)
	) name15402 (
		_w21217_,
		_w21221_,
		_w21225_,
		_w21228_,
		_w21229_
	);
	LUT2 #(
		.INIT('h6)
	) name15403 (
		\u1_L4_reg[12]/NET0131 ,
		_w21229_,
		_w21230_
	);
	LUT4 #(
		.INIT('hc693)
	) name15404 (
		decrypt_pad,
		\u1_R4_reg[20]/NET0131 ,
		\u1_uk_K_r4_reg[0]/P0001 ,
		\u1_uk_K_r4_reg[8]/NET0131 ,
		_w21231_
	);
	LUT4 #(
		.INIT('hc693)
	) name15405 (
		decrypt_pad,
		\u1_R4_reg[19]/NET0131 ,
		\u1_uk_K_r4_reg[16]/NET0131 ,
		\u1_uk_K_r4_reg[52]/NET0131 ,
		_w21232_
	);
	LUT4 #(
		.INIT('hc693)
	) name15406 (
		decrypt_pad,
		\u1_R4_reg[18]/NET0131 ,
		\u1_uk_K_r4_reg[29]/NET0131 ,
		\u1_uk_K_r4_reg[37]/NET0131 ,
		_w21233_
	);
	LUT4 #(
		.INIT('hc963)
	) name15407 (
		decrypt_pad,
		\u1_R4_reg[16]/NET0131 ,
		\u1_uk_K_r4_reg[21]/NET0131 ,
		\u1_uk_K_r4_reg[44]/NET0131 ,
		_w21234_
	);
	LUT4 #(
		.INIT('hc693)
	) name15408 (
		decrypt_pad,
		\u1_R4_reg[21]/NET0131 ,
		\u1_uk_K_r4_reg[1]/NET0131 ,
		\u1_uk_K_r4_reg[9]/NET0131 ,
		_w21235_
	);
	LUT4 #(
		.INIT('hc693)
	) name15409 (
		decrypt_pad,
		\u1_R4_reg[17]/NET0131 ,
		\u1_uk_K_r4_reg[35]/NET0131 ,
		\u1_uk_K_r4_reg[43]/NET0131 ,
		_w21236_
	);
	LUT3 #(
		.INIT('h02)
	) name15410 (
		_w21234_,
		_w21235_,
		_w21236_,
		_w21237_
	);
	LUT4 #(
		.INIT('h0002)
	) name15411 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21238_
	);
	LUT4 #(
		.INIT('h0800)
	) name15412 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21239_
	);
	LUT3 #(
		.INIT('h04)
	) name15413 (
		_w21234_,
		_w21235_,
		_w21236_,
		_w21240_
	);
	LUT4 #(
		.INIT('hc7b9)
	) name15414 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21241_
	);
	LUT3 #(
		.INIT('h10)
	) name15415 (
		_w21234_,
		_w21233_,
		_w21236_,
		_w21242_
	);
	LUT4 #(
		.INIT('h7a6e)
	) name15416 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21243_
	);
	LUT4 #(
		.INIT('h0180)
	) name15417 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21244_
	);
	LUT4 #(
		.INIT('h00d8)
	) name15418 (
		_w21232_,
		_w21243_,
		_w21241_,
		_w21244_,
		_w21245_
	);
	LUT2 #(
		.INIT('h1)
	) name15419 (
		_w21231_,
		_w21245_,
		_w21246_
	);
	LUT4 #(
		.INIT('h95b3)
	) name15420 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21247_
	);
	LUT2 #(
		.INIT('h4)
	) name15421 (
		_w21247_,
		_w21232_,
		_w21248_
	);
	LUT2 #(
		.INIT('h9)
	) name15422 (
		_w21233_,
		_w21236_,
		_w21249_
	);
	LUT4 #(
		.INIT('h0220)
	) name15423 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21250_
	);
	LUT4 #(
		.INIT('h0888)
	) name15424 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21232_,
		_w21251_
	);
	LUT3 #(
		.INIT('h13)
	) name15425 (
		_w21249_,
		_w21250_,
		_w21251_,
		_w21252_
	);
	LUT3 #(
		.INIT('h8a)
	) name15426 (
		_w21231_,
		_w21248_,
		_w21252_,
		_w21253_
	);
	LUT4 #(
		.INIT('h0010)
	) name15427 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21254_
	);
	LUT4 #(
		.INIT('h0200)
	) name15428 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21255_
	);
	LUT3 #(
		.INIT('h02)
	) name15429 (
		_w21232_,
		_w21255_,
		_w21254_,
		_w21256_
	);
	LUT3 #(
		.INIT('h40)
	) name15430 (
		_w21234_,
		_w21235_,
		_w21236_,
		_w21257_
	);
	LUT3 #(
		.INIT('hbe)
	) name15431 (
		_w21234_,
		_w21235_,
		_w21236_,
		_w21258_
	);
	LUT2 #(
		.INIT('h2)
	) name15432 (
		_w21231_,
		_w21233_,
		_w21259_
	);
	LUT4 #(
		.INIT('h1040)
	) name15433 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21260_
	);
	LUT4 #(
		.INIT('h1011)
	) name15434 (
		_w21232_,
		_w21260_,
		_w21258_,
		_w21259_,
		_w21261_
	);
	LUT2 #(
		.INIT('h1)
	) name15435 (
		_w21256_,
		_w21261_,
		_w21262_
	);
	LUT4 #(
		.INIT('h5556)
	) name15436 (
		\u1_L4_reg[14]/NET0131 ,
		_w21253_,
		_w21262_,
		_w21246_,
		_w21263_
	);
	LUT4 #(
		.INIT('h7773)
	) name15437 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21264_
	);
	LUT4 #(
		.INIT('h6673)
	) name15438 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21265_
	);
	LUT4 #(
		.INIT('h0002)
	) name15439 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21266_
	);
	LUT4 #(
		.INIT('h3302)
	) name15440 (
		_w21168_,
		_w21177_,
		_w21265_,
		_w21266_,
		_w21267_
	);
	LUT4 #(
		.INIT('h0040)
	) name15441 (
		_w21166_,
		_w21165_,
		_w21167_,
		_w21168_,
		_w21268_
	);
	LUT4 #(
		.INIT('hf7b7)
	) name15442 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21269_
	);
	LUT4 #(
		.INIT('h0100)
	) name15443 (
		_w21164_,
		_w21166_,
		_w21167_,
		_w21168_,
		_w21270_
	);
	LUT4 #(
		.INIT('h2000)
	) name15444 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21271_
	);
	LUT4 #(
		.INIT('h0100)
	) name15445 (
		_w21270_,
		_w21268_,
		_w21271_,
		_w21269_,
		_w21272_
	);
	LUT3 #(
		.INIT('h02)
	) name15446 (
		_w21164_,
		_w21166_,
		_w21177_,
		_w21273_
	);
	LUT4 #(
		.INIT('hfbbf)
	) name15447 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21274_
	);
	LUT4 #(
		.INIT('h00df)
	) name15448 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21168_,
		_w21275_
	);
	LUT4 #(
		.INIT('h1000)
	) name15449 (
		_w21187_,
		_w21273_,
		_w21275_,
		_w21274_,
		_w21276_
	);
	LUT4 #(
		.INIT('h0100)
	) name15450 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21277_
	);
	LUT3 #(
		.INIT('h02)
	) name15451 (
		_w21168_,
		_w21182_,
		_w21277_,
		_w21278_
	);
	LUT4 #(
		.INIT('hddd0)
	) name15452 (
		_w21177_,
		_w21272_,
		_w21276_,
		_w21278_,
		_w21279_
	);
	LUT3 #(
		.INIT('h65)
	) name15453 (
		\u1_L4_reg[15]/P0001 ,
		_w21267_,
		_w21279_,
		_w21280_
	);
	LUT4 #(
		.INIT('h084c)
	) name15454 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21281_
	);
	LUT4 #(
		.INIT('hfbc8)
	) name15455 (
		_w21139_,
		_w21131_,
		_w21159_,
		_w21281_,
		_w21282_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name15456 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21283_
	);
	LUT3 #(
		.INIT('h45)
	) name15457 (
		_w21143_,
		_w21282_,
		_w21283_,
		_w21284_
	);
	LUT4 #(
		.INIT('hdf4f)
	) name15458 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21285_
	);
	LUT4 #(
		.INIT('h4000)
	) name15459 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21286_
	);
	LUT4 #(
		.INIT('hbcff)
	) name15460 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21287_
	);
	LUT4 #(
		.INIT('h02aa)
	) name15461 (
		_w21143_,
		_w21131_,
		_w21285_,
		_w21287_,
		_w21288_
	);
	LUT4 #(
		.INIT('h6dff)
	) name15462 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21289_
	);
	LUT2 #(
		.INIT('h2)
	) name15463 (
		_w21131_,
		_w21289_,
		_w21290_
	);
	LUT2 #(
		.INIT('h4)
	) name15464 (
		_w21131_,
		_w21286_,
		_w21291_
	);
	LUT4 #(
		.INIT('hf5f1)
	) name15465 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21292_
	);
	LUT2 #(
		.INIT('h8)
	) name15466 (
		_w21143_,
		_w21131_,
		_w21293_
	);
	LUT4 #(
		.INIT('h7077)
	) name15467 (
		_w21133_,
		_w21148_,
		_w21292_,
		_w21293_,
		_w21294_
	);
	LUT4 #(
		.INIT('h0100)
	) name15468 (
		_w21290_,
		_w21291_,
		_w21288_,
		_w21294_,
		_w21295_
	);
	LUT3 #(
		.INIT('h65)
	) name15469 (
		\u1_L4_reg[1]/NET0131 ,
		_w21284_,
		_w21295_,
		_w21296_
	);
	LUT4 #(
		.INIT('h0040)
	) name15470 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21297_
	);
	LUT4 #(
		.INIT('hcc9d)
	) name15471 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21298_
	);
	LUT2 #(
		.INIT('h2)
	) name15472 (
		_w21064_,
		_w21298_,
		_w21299_
	);
	LUT4 #(
		.INIT('h0400)
	) name15473 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21300_
	);
	LUT4 #(
		.INIT('h4041)
	) name15474 (
		_w21064_,
		_w21067_,
		_w21068_,
		_w21066_,
		_w21301_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15475 (
		_w21063_,
		_w21067_,
		_w21065_,
		_w21066_,
		_w21302_
	);
	LUT3 #(
		.INIT('h10)
	) name15476 (
		_w21301_,
		_w21300_,
		_w21302_,
		_w21303_
	);
	LUT4 #(
		.INIT('h01c3)
	) name15477 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21304_
	);
	LUT4 #(
		.INIT('h0200)
	) name15478 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21305_
	);
	LUT4 #(
		.INIT('h2ff3)
	) name15479 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21306_
	);
	LUT4 #(
		.INIT('he4ee)
	) name15480 (
		_w21064_,
		_w21304_,
		_w21305_,
		_w21306_,
		_w21307_
	);
	LUT4 #(
		.INIT('h0800)
	) name15481 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21308_
	);
	LUT3 #(
		.INIT('h01)
	) name15482 (
		_w21063_,
		_w21087_,
		_w21308_,
		_w21309_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15483 (
		_w21299_,
		_w21303_,
		_w21307_,
		_w21309_,
		_w21310_
	);
	LUT2 #(
		.INIT('h6)
	) name15484 (
		\u1_L4_reg[17]/NET0131 ,
		_w21310_,
		_w21311_
	);
	LUT4 #(
		.INIT('h080a)
	) name15485 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21312_
	);
	LUT3 #(
		.INIT('h01)
	) name15486 (
		_w21168_,
		_w21271_,
		_w21312_,
		_w21313_
	);
	LUT4 #(
		.INIT('h8381)
	) name15487 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21314_
	);
	LUT4 #(
		.INIT('hbf00)
	) name15488 (
		_w21164_,
		_w21166_,
		_w21167_,
		_w21168_,
		_w21315_
	);
	LUT2 #(
		.INIT('h4)
	) name15489 (
		_w21314_,
		_w21315_,
		_w21316_
	);
	LUT4 #(
		.INIT('h0090)
	) name15490 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21317_
	);
	LUT3 #(
		.INIT('h02)
	) name15491 (
		_w21177_,
		_w21277_,
		_w21317_,
		_w21318_
	);
	LUT3 #(
		.INIT('he0)
	) name15492 (
		_w21313_,
		_w21316_,
		_w21318_,
		_w21319_
	);
	LUT4 #(
		.INIT('hde56)
	) name15493 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21320_
	);
	LUT2 #(
		.INIT('h2)
	) name15494 (
		_w21168_,
		_w21320_,
		_w21321_
	);
	LUT4 #(
		.INIT('h00bf)
	) name15495 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21177_,
		_w21322_
	);
	LUT2 #(
		.INIT('h4)
	) name15496 (
		_w21172_,
		_w21322_,
		_w21323_
	);
	LUT2 #(
		.INIT('h8)
	) name15497 (
		_w21164_,
		_w21167_,
		_w21324_
	);
	LUT3 #(
		.INIT('hdc)
	) name15498 (
		_w21166_,
		_w21165_,
		_w21168_,
		_w21325_
	);
	LUT2 #(
		.INIT('h2)
	) name15499 (
		_w21324_,
		_w21325_,
		_w21326_
	);
	LUT2 #(
		.INIT('h1)
	) name15500 (
		_w21164_,
		_w21168_,
		_w21327_
	);
	LUT3 #(
		.INIT('h35)
	) name15501 (
		_w21166_,
		_w21165_,
		_w21167_,
		_w21328_
	);
	LUT3 #(
		.INIT('h51)
	) name15502 (
		_w21187_,
		_w21327_,
		_w21328_,
		_w21329_
	);
	LUT4 #(
		.INIT('h1000)
	) name15503 (
		_w21321_,
		_w21326_,
		_w21323_,
		_w21329_,
		_w21330_
	);
	LUT3 #(
		.INIT('ha9)
	) name15504 (
		\u1_L4_reg[21]/NET0131 ,
		_w21319_,
		_w21330_,
		_w21331_
	);
	LUT4 #(
		.INIT('h67a8)
	) name15505 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21332_
	);
	LUT4 #(
		.INIT('hfa77)
	) name15506 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21333_
	);
	LUT4 #(
		.INIT('hd3ff)
	) name15507 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21334_
	);
	LUT4 #(
		.INIT('hd800)
	) name15508 (
		_w21232_,
		_w21332_,
		_w21333_,
		_w21334_,
		_w21335_
	);
	LUT2 #(
		.INIT('h2)
	) name15509 (
		_w21231_,
		_w21335_,
		_w21336_
	);
	LUT3 #(
		.INIT('hb0)
	) name15510 (
		_w21235_,
		_w21236_,
		_w21232_,
		_w21337_
	);
	LUT4 #(
		.INIT('h3301)
	) name15511 (
		_w21234_,
		_w21233_,
		_w21236_,
		_w21232_,
		_w21338_
	);
	LUT2 #(
		.INIT('h4)
	) name15512 (
		_w21337_,
		_w21338_,
		_w21339_
	);
	LUT4 #(
		.INIT('h4000)
	) name15513 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21340_
	);
	LUT4 #(
		.INIT('hafdd)
	) name15514 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21341_
	);
	LUT3 #(
		.INIT('h32)
	) name15515 (
		_w21232_,
		_w21340_,
		_w21341_,
		_w21342_
	);
	LUT4 #(
		.INIT('hdfef)
	) name15516 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21343_
	);
	LUT4 #(
		.INIT('hdfeb)
	) name15517 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21344_
	);
	LUT4 #(
		.INIT('h0008)
	) name15518 (
		_w21234_,
		_w21233_,
		_w21236_,
		_w21232_,
		_w21345_
	);
	LUT4 #(
		.INIT('h0301)
	) name15519 (
		_w21232_,
		_w21239_,
		_w21345_,
		_w21344_,
		_w21346_
	);
	LUT4 #(
		.INIT('hba00)
	) name15520 (
		_w21231_,
		_w21339_,
		_w21342_,
		_w21346_,
		_w21347_
	);
	LUT3 #(
		.INIT('h65)
	) name15521 (
		\u1_L4_reg[25]/NET0131 ,
		_w21336_,
		_w21347_,
		_w21348_
	);
	LUT4 #(
		.INIT('hc693)
	) name15522 (
		decrypt_pad,
		\u1_R4_reg[8]/NET0131 ,
		\u1_uk_K_r4_reg[20]/NET0131 ,
		\u1_uk_K_r4_reg[26]/NET0131 ,
		_w21349_
	);
	LUT4 #(
		.INIT('hc963)
	) name15523 (
		decrypt_pad,
		\u1_R4_reg[7]/NET0131 ,
		\u1_uk_K_r4_reg[3]/NET0131 ,
		\u1_uk_K_r4_reg[54]/NET0131 ,
		_w21350_
	);
	LUT4 #(
		.INIT('hc693)
	) name15524 (
		decrypt_pad,
		\u1_R4_reg[5]/NET0131 ,
		\u1_uk_K_r4_reg[12]/NET0131 ,
		\u1_uk_K_r4_reg[18]/NET0131 ,
		_w21351_
	);
	LUT4 #(
		.INIT('hc693)
	) name15525 (
		decrypt_pad,
		\u1_R4_reg[4]/NET0131 ,
		\u1_uk_K_r4_reg[33]/NET0131 ,
		\u1_uk_K_r4_reg[39]/NET0131 ,
		_w21352_
	);
	LUT4 #(
		.INIT('hc693)
	) name15526 (
		decrypt_pad,
		\u1_R4_reg[9]/NET0131 ,
		\u1_uk_K_r4_reg[25]/NET0131 ,
		\u1_uk_K_r4_reg[6]/NET0131 ,
		_w21353_
	);
	LUT4 #(
		.INIT('hc693)
	) name15527 (
		decrypt_pad,
		\u1_R4_reg[6]/NET0131 ,
		\u1_uk_K_r4_reg[3]/NET0131 ,
		\u1_uk_K_r4_reg[41]/NET0131 ,
		_w21354_
	);
	LUT4 #(
		.INIT('h59fb)
	) name15528 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21355_
	);
	LUT2 #(
		.INIT('h1)
	) name15529 (
		_w21350_,
		_w21355_,
		_w21356_
	);
	LUT4 #(
		.INIT('h0034)
	) name15530 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21357_
	);
	LUT4 #(
		.INIT('h0800)
	) name15531 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21358_
	);
	LUT4 #(
		.INIT('h0004)
	) name15532 (
		_w21350_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21359_
	);
	LUT4 #(
		.INIT('h4000)
	) name15533 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21360_
	);
	LUT4 #(
		.INIT('h0007)
	) name15534 (
		_w21350_,
		_w21358_,
		_w21359_,
		_w21360_,
		_w21361_
	);
	LUT4 #(
		.INIT('h5455)
	) name15535 (
		_w21349_,
		_w21356_,
		_w21357_,
		_w21361_,
		_w21362_
	);
	LUT4 #(
		.INIT('he6ee)
	) name15536 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21363_
	);
	LUT4 #(
		.INIT('h4044)
	) name15537 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21364_
	);
	LUT3 #(
		.INIT('h51)
	) name15538 (
		_w21350_,
		_w21351_,
		_w21354_,
		_w21365_
	);
	LUT4 #(
		.INIT('hf200)
	) name15539 (
		_w21349_,
		_w21363_,
		_w21364_,
		_w21365_,
		_w21366_
	);
	LUT4 #(
		.INIT('h0002)
	) name15540 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21367_
	);
	LUT4 #(
		.INIT('h80a0)
	) name15541 (
		_w21350_,
		_w21352_,
		_w21351_,
		_w21354_,
		_w21368_
	);
	LUT4 #(
		.INIT('h0080)
	) name15542 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21369_
	);
	LUT4 #(
		.INIT('haaa8)
	) name15543 (
		_w21349_,
		_w21367_,
		_w21368_,
		_w21369_,
		_w21370_
	);
	LUT3 #(
		.INIT('ha2)
	) name15544 (
		_w21352_,
		_w21351_,
		_w21354_,
		_w21371_
	);
	LUT3 #(
		.INIT('h45)
	) name15545 (
		_w21352_,
		_w21351_,
		_w21354_,
		_w21372_
	);
	LUT3 #(
		.INIT('h8a)
	) name15546 (
		_w21350_,
		_w21352_,
		_w21353_,
		_w21373_
	);
	LUT3 #(
		.INIT('h10)
	) name15547 (
		_w21372_,
		_w21371_,
		_w21373_,
		_w21374_
	);
	LUT3 #(
		.INIT('h01)
	) name15548 (
		_w21370_,
		_w21374_,
		_w21366_,
		_w21375_
	);
	LUT3 #(
		.INIT('h65)
	) name15549 (
		\u1_L4_reg[2]/NET0131 ,
		_w21362_,
		_w21375_,
		_w21376_
	);
	LUT3 #(
		.INIT('h02)
	) name15550 (
		_w21131_,
		_w21142_,
		_w21154_,
		_w21377_
	);
	LUT4 #(
		.INIT('h0094)
	) name15551 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21378_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name15552 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21379_
	);
	LUT4 #(
		.INIT('h0302)
	) name15553 (
		_w21143_,
		_w21131_,
		_w21378_,
		_w21379_,
		_w21380_
	);
	LUT2 #(
		.INIT('h1)
	) name15554 (
		_w21377_,
		_w21380_,
		_w21381_
	);
	LUT3 #(
		.INIT('h8d)
	) name15555 (
		_w21128_,
		_w21133_,
		_w21131_,
		_w21382_
	);
	LUT4 #(
		.INIT('h0c04)
	) name15556 (
		_w21137_,
		_w21143_,
		_w21286_,
		_w21382_,
		_w21383_
	);
	LUT4 #(
		.INIT('h7775)
	) name15557 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21133_,
		_w21384_
	);
	LUT3 #(
		.INIT('h0d)
	) name15558 (
		_w21130_,
		_w21133_,
		_w21131_,
		_w21385_
	);
	LUT4 #(
		.INIT('hdddf)
	) name15559 (
		_w21129_,
		_w21130_,
		_w21128_,
		_w21131_,
		_w21386_
	);
	LUT4 #(
		.INIT('hcf45)
	) name15560 (
		_w21133_,
		_w21384_,
		_w21385_,
		_w21386_,
		_w21387_
	);
	LUT2 #(
		.INIT('h2)
	) name15561 (
		_w21144_,
		_w21150_,
		_w21388_
	);
	LUT4 #(
		.INIT('h00fd)
	) name15562 (
		_w21130_,
		_w21128_,
		_w21133_,
		_w21143_,
		_w21389_
	);
	LUT3 #(
		.INIT('h10)
	) name15563 (
		_w21154_,
		_w21152_,
		_w21389_,
		_w21390_
	);
	LUT4 #(
		.INIT('h7077)
	) name15564 (
		_w21383_,
		_w21387_,
		_w21388_,
		_w21390_,
		_w21391_
	);
	LUT3 #(
		.INIT('h56)
	) name15565 (
		\u1_L4_reg[26]/NET0131 ,
		_w21381_,
		_w21391_,
		_w21392_
	);
	LUT2 #(
		.INIT('h1)
	) name15566 (
		_w21352_,
		_w21354_,
		_w21393_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name15567 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21394_
	);
	LUT2 #(
		.INIT('h2)
	) name15568 (
		_w21350_,
		_w21394_,
		_w21395_
	);
	LUT4 #(
		.INIT('hbfae)
	) name15569 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21396_
	);
	LUT2 #(
		.INIT('h1)
	) name15570 (
		_w21350_,
		_w21396_,
		_w21397_
	);
	LUT2 #(
		.INIT('h8)
	) name15571 (
		_w21350_,
		_w21352_,
		_w21398_
	);
	LUT4 #(
		.INIT('h7737)
	) name15572 (
		_w21350_,
		_w21352_,
		_w21353_,
		_w21351_,
		_w21399_
	);
	LUT4 #(
		.INIT('h0400)
	) name15573 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21400_
	);
	LUT3 #(
		.INIT('h0e)
	) name15574 (
		_w21354_,
		_w21399_,
		_w21400_,
		_w21401_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15575 (
		_w21349_,
		_w21397_,
		_w21395_,
		_w21401_,
		_w21402_
	);
	LUT4 #(
		.INIT('hdaff)
	) name15576 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21403_
	);
	LUT2 #(
		.INIT('h1)
	) name15577 (
		_w21350_,
		_w21403_,
		_w21404_
	);
	LUT3 #(
		.INIT('h02)
	) name15578 (
		_w21352_,
		_w21353_,
		_w21354_,
		_w21405_
	);
	LUT4 #(
		.INIT('h1145)
	) name15579 (
		_w21350_,
		_w21352_,
		_w21353_,
		_w21351_,
		_w21406_
	);
	LUT4 #(
		.INIT('h7077)
	) name15580 (
		_w21350_,
		_w21396_,
		_w21405_,
		_w21406_,
		_w21407_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name15581 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21408_
	);
	LUT4 #(
		.INIT('h2322)
	) name15582 (
		_w21349_,
		_w21404_,
		_w21407_,
		_w21408_,
		_w21409_
	);
	LUT3 #(
		.INIT('h65)
	) name15583 (
		\u1_L4_reg[28]/NET0131 ,
		_w21402_,
		_w21409_,
		_w21410_
	);
	LUT4 #(
		.INIT('h67dc)
	) name15584 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21411_
	);
	LUT4 #(
		.INIT('hd2f7)
	) name15585 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21412_
	);
	LUT4 #(
		.INIT('h0040)
	) name15586 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21413_
	);
	LUT4 #(
		.INIT('h00e4)
	) name15587 (
		_w21101_,
		_w21412_,
		_w21411_,
		_w21413_,
		_w21414_
	);
	LUT2 #(
		.INIT('h1)
	) name15588 (
		_w21095_,
		_w21414_,
		_w21415_
	);
	LUT4 #(
		.INIT('h9aff)
	) name15589 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21416_
	);
	LUT2 #(
		.INIT('h2)
	) name15590 (
		_w21101_,
		_w21416_,
		_w21417_
	);
	LUT4 #(
		.INIT('h6f6e)
	) name15591 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21418_
	);
	LUT2 #(
		.INIT('h1)
	) name15592 (
		_w21101_,
		_w21418_,
		_w21419_
	);
	LUT4 #(
		.INIT('h0010)
	) name15593 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21420_
	);
	LUT4 #(
		.INIT('h0001)
	) name15594 (
		_w21115_,
		_w21116_,
		_w21120_,
		_w21420_,
		_w21421_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15595 (
		_w21095_,
		_w21419_,
		_w21417_,
		_w21421_,
		_w21422_
	);
	LUT4 #(
		.INIT('h2000)
	) name15596 (
		_w21099_,
		_w21096_,
		_w21098_,
		_w21101_,
		_w21423_
	);
	LUT2 #(
		.INIT('h1)
	) name15597 (
		_w21104_,
		_w21423_,
		_w21424_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name15598 (
		\u1_L4_reg[29]/NET0131 ,
		_w21422_,
		_w21415_,
		_w21424_,
		_w21425_
	);
	LUT4 #(
		.INIT('hefcc)
	) name15599 (
		_w21099_,
		_w21096_,
		_w21098_,
		_w21101_,
		_w21426_
	);
	LUT2 #(
		.INIT('h1)
	) name15600 (
		_w21097_,
		_w21426_,
		_w21427_
	);
	LUT4 #(
		.INIT('h0010)
	) name15601 (
		_w21099_,
		_w21096_,
		_w21098_,
		_w21101_,
		_w21428_
	);
	LUT3 #(
		.INIT('h80)
	) name15602 (
		_w21099_,
		_w21096_,
		_w21098_,
		_w21429_
	);
	LUT4 #(
		.INIT('h0800)
	) name15603 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21101_,
		_w21430_
	);
	LUT4 #(
		.INIT('h0002)
	) name15604 (
		_w21095_,
		_w21428_,
		_w21430_,
		_w21429_,
		_w21431_
	);
	LUT2 #(
		.INIT('h4)
	) name15605 (
		_w21427_,
		_w21431_,
		_w21432_
	);
	LUT4 #(
		.INIT('hdf00)
	) name15606 (
		_w21097_,
		_w21099_,
		_w21098_,
		_w21101_,
		_w21433_
	);
	LUT4 #(
		.INIT('hfb7b)
	) name15607 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21434_
	);
	LUT2 #(
		.INIT('h8)
	) name15608 (
		_w21433_,
		_w21434_,
		_w21435_
	);
	LUT3 #(
		.INIT('h10)
	) name15609 (
		_w21097_,
		_w21099_,
		_w21098_,
		_w21436_
	);
	LUT3 #(
		.INIT('h01)
	) name15610 (
		_w21101_,
		_w21413_,
		_w21436_,
		_w21437_
	);
	LUT3 #(
		.INIT('h01)
	) name15611 (
		_w21095_,
		_w21104_,
		_w21106_,
		_w21438_
	);
	LUT3 #(
		.INIT('he0)
	) name15612 (
		_w21435_,
		_w21437_,
		_w21438_,
		_w21439_
	);
	LUT4 #(
		.INIT('h9e00)
	) name15613 (
		_w21097_,
		_w21099_,
		_w21098_,
		_w21101_,
		_w21440_
	);
	LUT4 #(
		.INIT('h007d)
	) name15614 (
		_w21097_,
		_w21099_,
		_w21098_,
		_w21101_,
		_w21441_
	);
	LUT4 #(
		.INIT('h3331)
	) name15615 (
		_w21096_,
		_w21122_,
		_w21441_,
		_w21440_,
		_w21442_
	);
	LUT4 #(
		.INIT('ha955)
	) name15616 (
		\u1_L4_reg[4]/NET0131 ,
		_w21432_,
		_w21439_,
		_w21442_,
		_w21443_
	);
	LUT3 #(
		.INIT('h10)
	) name15617 (
		_w21353_,
		_w21351_,
		_w21354_,
		_w21444_
	);
	LUT4 #(
		.INIT('h5515)
	) name15618 (
		_w21350_,
		_w21352_,
		_w21353_,
		_w21351_,
		_w21445_
	);
	LUT3 #(
		.INIT('h40)
	) name15619 (
		_w21352_,
		_w21353_,
		_w21354_,
		_w21446_
	);
	LUT4 #(
		.INIT('haaa8)
	) name15620 (
		_w21350_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21447_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15621 (
		_w21444_,
		_w21445_,
		_w21446_,
		_w21447_,
		_w21448_
	);
	LUT4 #(
		.INIT('h0010)
	) name15622 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21449_
	);
	LUT4 #(
		.INIT('h0002)
	) name15623 (
		_w21349_,
		_w21359_,
		_w21360_,
		_w21449_,
		_w21450_
	);
	LUT2 #(
		.INIT('h4)
	) name15624 (
		_w21448_,
		_w21450_,
		_w21451_
	);
	LUT3 #(
		.INIT('hc8)
	) name15625 (
		_w21350_,
		_w21353_,
		_w21351_,
		_w21452_
	);
	LUT2 #(
		.INIT('h8)
	) name15626 (
		_w21393_,
		_w21452_,
		_w21453_
	);
	LUT3 #(
		.INIT('hb0)
	) name15627 (
		_w21353_,
		_w21351_,
		_w21354_,
		_w21454_
	);
	LUT3 #(
		.INIT('h15)
	) name15628 (
		_w21349_,
		_w21398_,
		_w21454_,
		_w21455_
	);
	LUT3 #(
		.INIT('h10)
	) name15629 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21456_
	);
	LUT4 #(
		.INIT('h0001)
	) name15630 (
		_w21350_,
		_w21367_,
		_w21400_,
		_w21456_,
		_w21457_
	);
	LUT3 #(
		.INIT('h40)
	) name15631 (
		_w21453_,
		_w21455_,
		_w21457_,
		_w21458_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name15632 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21459_
	);
	LUT4 #(
		.INIT('h0929)
	) name15633 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21460_
	);
	LUT2 #(
		.INIT('h2)
	) name15634 (
		_w21350_,
		_w21460_,
		_w21461_
	);
	LUT3 #(
		.INIT('h40)
	) name15635 (
		_w21453_,
		_w21455_,
		_w21461_,
		_w21462_
	);
	LUT4 #(
		.INIT('h001f)
	) name15636 (
		_w21451_,
		_w21458_,
		_w21459_,
		_w21462_,
		_w21463_
	);
	LUT2 #(
		.INIT('h9)
	) name15637 (
		\u1_L4_reg[13]/NET0131 ,
		_w21463_,
		_w21464_
	);
	LUT4 #(
		.INIT('h4010)
	) name15638 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21465_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15639 (
		_w21095_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21466_
	);
	LUT4 #(
		.INIT('h2000)
	) name15640 (
		_w21097_,
		_w21096_,
		_w21098_,
		_w21101_,
		_w21467_
	);
	LUT4 #(
		.INIT('h040a)
	) name15641 (
		_w21097_,
		_w21099_,
		_w21098_,
		_w21101_,
		_w21468_
	);
	LUT4 #(
		.INIT('h0100)
	) name15642 (
		_w21120_,
		_w21467_,
		_w21468_,
		_w21466_,
		_w21469_
	);
	LUT4 #(
		.INIT('h4e55)
	) name15643 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21470_
	);
	LUT2 #(
		.INIT('h2)
	) name15644 (
		_w21101_,
		_w21470_,
		_w21471_
	);
	LUT4 #(
		.INIT('h0041)
	) name15645 (
		_w21097_,
		_w21099_,
		_w21098_,
		_w21101_,
		_w21472_
	);
	LUT4 #(
		.INIT('h8000)
	) name15646 (
		_w21097_,
		_w21099_,
		_w21096_,
		_w21098_,
		_w21473_
	);
	LUT3 #(
		.INIT('h01)
	) name15647 (
		_w21095_,
		_w21473_,
		_w21472_,
		_w21474_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15648 (
		_w21465_,
		_w21469_,
		_w21471_,
		_w21474_,
		_w21475_
	);
	LUT2 #(
		.INIT('h2)
	) name15649 (
		_w21121_,
		_w21107_,
		_w21476_
	);
	LUT3 #(
		.INIT('h65)
	) name15650 (
		\u1_L4_reg[19]/P0001 ,
		_w21475_,
		_w21476_,
		_w21477_
	);
	LUT3 #(
		.INIT('he3)
	) name15651 (
		_w21068_,
		_w21065_,
		_w21066_,
		_w21478_
	);
	LUT4 #(
		.INIT('hfcc7)
	) name15652 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21479_
	);
	LUT3 #(
		.INIT('ha8)
	) name15653 (
		_w21063_,
		_w21064_,
		_w21479_,
		_w21480_
	);
	LUT3 #(
		.INIT('h7e)
	) name15654 (
		_w21067_,
		_w21065_,
		_w21066_,
		_w21481_
	);
	LUT2 #(
		.INIT('h4)
	) name15655 (
		_w21064_,
		_w21067_,
		_w21482_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name15656 (
		_w21064_,
		_w21067_,
		_w21068_,
		_w21065_,
		_w21483_
	);
	LUT4 #(
		.INIT('h0200)
	) name15657 (
		_w21064_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21484_
	);
	LUT4 #(
		.INIT('h4555)
	) name15658 (
		_w21063_,
		_w21064_,
		_w21068_,
		_w21066_,
		_w21485_
	);
	LUT4 #(
		.INIT('h4000)
	) name15659 (
		_w21484_,
		_w21485_,
		_w21481_,
		_w21483_,
		_w21486_
	);
	LUT2 #(
		.INIT('h1)
	) name15660 (
		_w21480_,
		_w21486_,
		_w21487_
	);
	LUT3 #(
		.INIT('ha8)
	) name15661 (
		_w21064_,
		_w21067_,
		_w21065_,
		_w21488_
	);
	LUT2 #(
		.INIT('h8)
	) name15662 (
		_w21082_,
		_w21488_,
		_w21489_
	);
	LUT3 #(
		.INIT('h07)
	) name15663 (
		_w21075_,
		_w21091_,
		_w21297_,
		_w21490_
	);
	LUT3 #(
		.INIT('h8a)
	) name15664 (
		_w21063_,
		_w21489_,
		_w21490_,
		_w21491_
	);
	LUT4 #(
		.INIT('hfbef)
	) name15665 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21492_
	);
	LUT2 #(
		.INIT('h1)
	) name15666 (
		_w21064_,
		_w21492_,
		_w21493_
	);
	LUT2 #(
		.INIT('h4)
	) name15667 (
		_w21067_,
		_w21484_,
		_w21494_
	);
	LUT3 #(
		.INIT('h15)
	) name15668 (
		_w21090_,
		_w21086_,
		_w21482_,
		_w21495_
	);
	LUT3 #(
		.INIT('h10)
	) name15669 (
		_w21493_,
		_w21494_,
		_w21495_,
		_w21496_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name15670 (
		\u1_L4_reg[23]/NET0131 ,
		_w21487_,
		_w21491_,
		_w21496_,
		_w21497_
	);
	LUT4 #(
		.INIT('hba76)
	) name15671 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21498_
	);
	LUT2 #(
		.INIT('h1)
	) name15672 (
		_w21168_,
		_w21498_,
		_w21499_
	);
	LUT3 #(
		.INIT('hd0)
	) name15673 (
		_w21164_,
		_w21167_,
		_w21168_,
		_w21500_
	);
	LUT4 #(
		.INIT('hbcdf)
	) name15674 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21501_
	);
	LUT3 #(
		.INIT('hb0)
	) name15675 (
		_w21264_,
		_w21500_,
		_w21501_,
		_w21502_
	);
	LUT3 #(
		.INIT('h8a)
	) name15676 (
		_w21177_,
		_w21499_,
		_w21502_,
		_w21503_
	);
	LUT4 #(
		.INIT('hfd00)
	) name15677 (
		_w21166_,
		_w21165_,
		_w21167_,
		_w21168_,
		_w21504_
	);
	LUT4 #(
		.INIT('h0cbf)
	) name15678 (
		_w21164_,
		_w21166_,
		_w21165_,
		_w21167_,
		_w21505_
	);
	LUT2 #(
		.INIT('h8)
	) name15679 (
		_w21504_,
		_w21505_,
		_w21506_
	);
	LUT4 #(
		.INIT('h0080)
	) name15680 (
		_w21164_,
		_w21165_,
		_w21167_,
		_w21168_,
		_w21507_
	);
	LUT4 #(
		.INIT('h0004)
	) name15681 (
		_w21164_,
		_w21166_,
		_w21167_,
		_w21168_,
		_w21508_
	);
	LUT3 #(
		.INIT('h01)
	) name15682 (
		_w21188_,
		_w21508_,
		_w21507_,
		_w21509_
	);
	LUT3 #(
		.INIT('h45)
	) name15683 (
		_w21177_,
		_w21506_,
		_w21509_,
		_w21510_
	);
	LUT2 #(
		.INIT('h4)
	) name15684 (
		_w21168_,
		_w21186_,
		_w21511_
	);
	LUT4 #(
		.INIT('h0400)
	) name15685 (
		_w21166_,
		_w21165_,
		_w21167_,
		_w21168_,
		_w21512_
	);
	LUT3 #(
		.INIT('h07)
	) name15686 (
		_w21169_,
		_w21191_,
		_w21512_,
		_w21513_
	);
	LUT2 #(
		.INIT('h4)
	) name15687 (
		_w21511_,
		_w21513_,
		_w21514_
	);
	LUT4 #(
		.INIT('h5655)
	) name15688 (
		\u1_L4_reg[27]/NET0131 ,
		_w21503_,
		_w21510_,
		_w21514_,
		_w21515_
	);
	LUT4 #(
		.INIT('h4000)
	) name15689 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21516_
	);
	LUT3 #(
		.INIT('h09)
	) name15690 (
		_w21040_,
		_w21036_,
		_w21037_,
		_w21517_
	);
	LUT4 #(
		.INIT('h2012)
	) name15691 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21518_
	);
	LUT4 #(
		.INIT('h00fb)
	) name15692 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21039_,
		_w21519_
	);
	LUT4 #(
		.INIT('h0189)
	) name15693 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21520_
	);
	LUT4 #(
		.INIT('hbf00)
	) name15694 (
		_w21040_,
		_w21036_,
		_w21037_,
		_w21039_,
		_w21521_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15695 (
		_w21518_,
		_w21519_,
		_w21520_,
		_w21521_,
		_w21522_
	);
	LUT3 #(
		.INIT('ha8)
	) name15696 (
		_w21035_,
		_w21516_,
		_w21522_,
		_w21523_
	);
	LUT4 #(
		.INIT('h79bf)
	) name15697 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21524_
	);
	LUT4 #(
		.INIT('h5057)
	) name15698 (
		_w21039_,
		_w21056_,
		_w21218_,
		_w21214_,
		_w21525_
	);
	LUT4 #(
		.INIT('h008c)
	) name15699 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21039_,
		_w21526_
	);
	LUT4 #(
		.INIT('h135f)
	) name15700 (
		_w21039_,
		_w21044_,
		_w21058_,
		_w21526_,
		_w21527_
	);
	LUT4 #(
		.INIT('hea00)
	) name15701 (
		_w21035_,
		_w21524_,
		_w21525_,
		_w21527_,
		_w21528_
	);
	LUT3 #(
		.INIT('h65)
	) name15702 (
		\u1_L4_reg[32]/NET0131 ,
		_w21523_,
		_w21528_,
		_w21529_
	);
	LUT4 #(
		.INIT('hc693)
	) name15703 (
		decrypt_pad,
		\u1_R4_reg[11]/P0001 ,
		\u1_uk_K_r4_reg[40]/NET0131 ,
		\u1_uk_K_r4_reg[46]/NET0131 ,
		_w21530_
	);
	LUT4 #(
		.INIT('hc963)
	) name15704 (
		decrypt_pad,
		\u1_R4_reg[12]/NET0131 ,
		\u1_uk_K_r4_reg[4]/NET0131 ,
		\u1_uk_K_r4_reg[55]/NET0131 ,
		_w21531_
	);
	LUT4 #(
		.INIT('hc693)
	) name15705 (
		decrypt_pad,
		\u1_R4_reg[13]/NET0131 ,
		\u1_uk_K_r4_reg[11]/NET0131 ,
		\u1_uk_K_r4_reg[17]/NET0131 ,
		_w21532_
	);
	LUT4 #(
		.INIT('hc963)
	) name15706 (
		decrypt_pad,
		\u1_R4_reg[9]/NET0131 ,
		\u1_uk_K_r4_reg[12]/NET0131 ,
		\u1_uk_K_r4_reg[6]/NET0131 ,
		_w21533_
	);
	LUT4 #(
		.INIT('hc693)
	) name15707 (
		decrypt_pad,
		\u1_R4_reg[8]/NET0131 ,
		\u1_uk_K_r4_reg[34]/NET0131 ,
		\u1_uk_K_r4_reg[40]/NET0131 ,
		_w21534_
	);
	LUT4 #(
		.INIT('hc963)
	) name15708 (
		decrypt_pad,
		\u1_R4_reg[10]/NET0131 ,
		\u1_uk_K_r4_reg[20]/NET0131 ,
		\u1_uk_K_r4_reg[39]/NET0131 ,
		_w21535_
	);
	LUT4 #(
		.INIT('h95b5)
	) name15709 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21536_
	);
	LUT2 #(
		.INIT('h1)
	) name15710 (
		_w21532_,
		_w21534_,
		_w21537_
	);
	LUT4 #(
		.INIT('h0001)
	) name15711 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21538_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name15712 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21539_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15713 (
		_w21531_,
		_w21530_,
		_w21536_,
		_w21539_,
		_w21540_
	);
	LUT2 #(
		.INIT('h8)
	) name15714 (
		_w21532_,
		_w21534_,
		_w21541_
	);
	LUT2 #(
		.INIT('h6)
	) name15715 (
		_w21532_,
		_w21534_,
		_w21542_
	);
	LUT4 #(
		.INIT('h000d)
	) name15716 (
		_w21530_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21543_
	);
	LUT4 #(
		.INIT('h0020)
	) name15717 (
		_w21530_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21544_
	);
	LUT4 #(
		.INIT('h4000)
	) name15718 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21545_
	);
	LUT4 #(
		.INIT('h0103)
	) name15719 (
		_w21542_,
		_w21544_,
		_w21545_,
		_w21543_,
		_w21546_
	);
	LUT3 #(
		.INIT('h20)
	) name15720 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21547_
	);
	LUT4 #(
		.INIT('h2000)
	) name15721 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21548_
	);
	LUT4 #(
		.INIT('h9990)
	) name15722 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21549_
	);
	LUT4 #(
		.INIT('h0990)
	) name15723 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21550_
	);
	LUT3 #(
		.INIT('h0b)
	) name15724 (
		_w21530_,
		_w21548_,
		_w21550_,
		_w21551_
	);
	LUT3 #(
		.INIT('h80)
	) name15725 (
		_w21531_,
		_w21533_,
		_w21535_,
		_w21552_
	);
	LUT3 #(
		.INIT('h80)
	) name15726 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21553_
	);
	LUT4 #(
		.INIT('h7b5b)
	) name15727 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21554_
	);
	LUT2 #(
		.INIT('h2)
	) name15728 (
		_w21531_,
		_w21530_,
		_w21555_
	);
	LUT4 #(
		.INIT('h7077)
	) name15729 (
		_w21537_,
		_w21552_,
		_w21554_,
		_w21555_,
		_w21556_
	);
	LUT4 #(
		.INIT('hea00)
	) name15730 (
		_w21531_,
		_w21546_,
		_w21551_,
		_w21556_,
		_w21557_
	);
	LUT3 #(
		.INIT('h65)
	) name15731 (
		\u1_L4_reg[6]/NET0131 ,
		_w21540_,
		_w21557_,
		_w21558_
	);
	LUT4 #(
		.INIT('h00a4)
	) name15732 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21559_
	);
	LUT2 #(
		.INIT('h2)
	) name15733 (
		_w21039_,
		_w21559_,
		_w21560_
	);
	LUT3 #(
		.INIT('h21)
	) name15734 (
		_w21038_,
		_w21036_,
		_w21037_,
		_w21561_
	);
	LUT3 #(
		.INIT('h48)
	) name15735 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21562_
	);
	LUT4 #(
		.INIT('h00bf)
	) name15736 (
		_w21040_,
		_w21036_,
		_w21037_,
		_w21039_,
		_w21563_
	);
	LUT3 #(
		.INIT('h10)
	) name15737 (
		_w21562_,
		_w21561_,
		_w21563_,
		_w21564_
	);
	LUT4 #(
		.INIT('h6800)
	) name15738 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21565_
	);
	LUT2 #(
		.INIT('h2)
	) name15739 (
		_w21035_,
		_w21565_,
		_w21566_
	);
	LUT4 #(
		.INIT('h4800)
	) name15740 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21037_,
		_w21567_
	);
	LUT4 #(
		.INIT('hdf00)
	) name15741 (
		_w21040_,
		_w21038_,
		_w21036_,
		_w21039_,
		_w21568_
	);
	LUT4 #(
		.INIT('h5455)
	) name15742 (
		_w21035_,
		_w21517_,
		_w21567_,
		_w21568_,
		_w21569_
	);
	LUT4 #(
		.INIT('h001f)
	) name15743 (
		_w21560_,
		_w21564_,
		_w21566_,
		_w21569_,
		_w21570_
	);
	LUT2 #(
		.INIT('h4)
	) name15744 (
		_w21039_,
		_w21565_,
		_w21571_
	);
	LUT2 #(
		.INIT('h2)
	) name15745 (
		_w21035_,
		_w21039_,
		_w21572_
	);
	LUT4 #(
		.INIT('h00ba)
	) name15746 (
		_w21043_,
		_w21039_,
		_w21559_,
		_w21572_,
		_w21573_
	);
	LUT2 #(
		.INIT('h1)
	) name15747 (
		_w21571_,
		_w21573_,
		_w21574_
	);
	LUT3 #(
		.INIT('h65)
	) name15748 (
		\u1_L4_reg[7]/NET0131 ,
		_w21570_,
		_w21574_,
		_w21575_
	);
	LUT4 #(
		.INIT('hff76)
	) name15749 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21576_
	);
	LUT3 #(
		.INIT('h02)
	) name15750 (
		_w21234_,
		_w21233_,
		_w21232_,
		_w21577_
	);
	LUT4 #(
		.INIT('h0031)
	) name15751 (
		_w21232_,
		_w21260_,
		_w21576_,
		_w21577_,
		_w21578_
	);
	LUT2 #(
		.INIT('h2)
	) name15752 (
		_w21231_,
		_w21578_,
		_w21579_
	);
	LUT4 #(
		.INIT('h8000)
	) name15753 (
		_w21234_,
		_w21235_,
		_w21236_,
		_w21232_,
		_w21580_
	);
	LUT3 #(
		.INIT('h04)
	) name15754 (
		_w21242_,
		_w21343_,
		_w21580_,
		_w21581_
	);
	LUT4 #(
		.INIT('hbb73)
	) name15755 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21582_
	);
	LUT3 #(
		.INIT('h72)
	) name15756 (
		_w21232_,
		_w21238_,
		_w21582_,
		_w21583_
	);
	LUT4 #(
		.INIT('hcbbf)
	) name15757 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21584_
	);
	LUT4 #(
		.INIT('haf23)
	) name15758 (
		_w21235_,
		_w21232_,
		_w21345_,
		_w21584_,
		_w21585_
	);
	LUT4 #(
		.INIT('hea00)
	) name15759 (
		_w21231_,
		_w21581_,
		_w21583_,
		_w21585_,
		_w21586_
	);
	LUT3 #(
		.INIT('h65)
	) name15760 (
		\u1_L4_reg[8]/NET0131 ,
		_w21579_,
		_w21586_,
		_w21587_
	);
	LUT4 #(
		.INIT('h3dc3)
	) name15761 (
		_w21530_,
		_w21532_,
		_w21534_,
		_w21533_,
		_w21588_
	);
	LUT4 #(
		.INIT('h0110)
	) name15762 (
		_w21530_,
		_w21532_,
		_w21534_,
		_w21535_,
		_w21589_
	);
	LUT4 #(
		.INIT('h0074)
	) name15763 (
		_w21547_,
		_w21535_,
		_w21588_,
		_w21589_,
		_w21590_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name15764 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21591_
	);
	LUT4 #(
		.INIT('h2880)
	) name15765 (
		_w21530_,
		_w21532_,
		_w21534_,
		_w21533_,
		_w21592_
	);
	LUT4 #(
		.INIT('h0032)
	) name15766 (
		_w21530_,
		_w21538_,
		_w21591_,
		_w21592_,
		_w21593_
	);
	LUT4 #(
		.INIT('hbeff)
	) name15767 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21594_
	);
	LUT4 #(
		.INIT('h0400)
	) name15768 (
		_w21530_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21595_
	);
	LUT3 #(
		.INIT('h0d)
	) name15769 (
		_w21530_,
		_w21594_,
		_w21595_,
		_w21596_
	);
	LUT4 #(
		.INIT('he400)
	) name15770 (
		_w21531_,
		_w21593_,
		_w21590_,
		_w21596_,
		_w21597_
	);
	LUT2 #(
		.INIT('h9)
	) name15771 (
		\u1_L4_reg[16]/NET0131 ,
		_w21597_,
		_w21598_
	);
	LUT2 #(
		.INIT('h4)
	) name15772 (
		_w21530_,
		_w21549_,
		_w21599_
	);
	LUT4 #(
		.INIT('h1dff)
	) name15773 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21600_
	);
	LUT2 #(
		.INIT('h2)
	) name15774 (
		_w21530_,
		_w21600_,
		_w21601_
	);
	LUT2 #(
		.INIT('h2)
	) name15775 (
		_w21530_,
		_w21535_,
		_w21602_
	);
	LUT3 #(
		.INIT('h0d)
	) name15776 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21603_
	);
	LUT4 #(
		.INIT('h0777)
	) name15777 (
		_w21542_,
		_w21543_,
		_w21602_,
		_w21603_,
		_w21604_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15778 (
		_w21531_,
		_w21601_,
		_w21599_,
		_w21604_,
		_w21605_
	);
	LUT4 #(
		.INIT('he2cd)
	) name15779 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21606_
	);
	LUT4 #(
		.INIT('h0400)
	) name15780 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21607_
	);
	LUT4 #(
		.INIT('h5504)
	) name15781 (
		_w21531_,
		_w21530_,
		_w21606_,
		_w21607_,
		_w21608_
	);
	LUT4 #(
		.INIT('h0009)
	) name15782 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21609_
	);
	LUT4 #(
		.INIT('h9db6)
	) name15783 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21610_
	);
	LUT2 #(
		.INIT('h1)
	) name15784 (
		_w21531_,
		_w21530_,
		_w21611_
	);
	LUT2 #(
		.INIT('h4)
	) name15785 (
		_w21610_,
		_w21611_,
		_w21612_
	);
	LUT3 #(
		.INIT('hdb)
	) name15786 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21613_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name15787 (
		_w21530_,
		_w21535_,
		_w21553_,
		_w21613_,
		_w21614_
	);
	LUT3 #(
		.INIT('h10)
	) name15788 (
		_w21608_,
		_w21612_,
		_w21614_,
		_w21615_
	);
	LUT3 #(
		.INIT('h65)
	) name15789 (
		\u1_L4_reg[24]/NET0131 ,
		_w21605_,
		_w21615_,
		_w21616_
	);
	LUT4 #(
		.INIT('h0200)
	) name15790 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21617_
	);
	LUT3 #(
		.INIT('h01)
	) name15791 (
		_w21531_,
		_w21609_,
		_w21617_,
		_w21618_
	);
	LUT2 #(
		.INIT('h8)
	) name15792 (
		_w21534_,
		_w21535_,
		_w21619_
	);
	LUT4 #(
		.INIT('h73af)
	) name15793 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21620_
	);
	LUT4 #(
		.INIT('hdf53)
	) name15794 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21621_
	);
	LUT3 #(
		.INIT('hd8)
	) name15795 (
		_w21530_,
		_w21620_,
		_w21621_,
		_w21622_
	);
	LUT4 #(
		.INIT('heed9)
	) name15796 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21623_
	);
	LUT4 #(
		.INIT('h23ef)
	) name15797 (
		_w21532_,
		_w21534_,
		_w21533_,
		_w21535_,
		_w21624_
	);
	LUT4 #(
		.INIT('ha820)
	) name15798 (
		_w21531_,
		_w21530_,
		_w21624_,
		_w21623_,
		_w21625_
	);
	LUT3 #(
		.INIT('h07)
	) name15799 (
		_w21618_,
		_w21622_,
		_w21625_,
		_w21626_
	);
	LUT3 #(
		.INIT('h08)
	) name15800 (
		_w21530_,
		_w21532_,
		_w21533_,
		_w21627_
	);
	LUT2 #(
		.INIT('h8)
	) name15801 (
		_w21619_,
		_w21627_,
		_w21628_
	);
	LUT4 #(
		.INIT('h1000)
	) name15802 (
		_w21530_,
		_w21532_,
		_w21533_,
		_w21535_,
		_w21629_
	);
	LUT3 #(
		.INIT('h0b)
	) name15803 (
		_w21541_,
		_w21552_,
		_w21629_,
		_w21630_
	);
	LUT2 #(
		.INIT('h4)
	) name15804 (
		_w21628_,
		_w21630_,
		_w21631_
	);
	LUT3 #(
		.INIT('h9a)
	) name15805 (
		\u1_L4_reg[30]/NET0131 ,
		_w21626_,
		_w21631_,
		_w21632_
	);
	LUT4 #(
		.INIT('he6f7)
	) name15806 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21633_
	);
	LUT4 #(
		.INIT('hf7df)
	) name15807 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21634_
	);
	LUT4 #(
		.INIT('hb100)
	) name15808 (
		_w21232_,
		_w21257_,
		_w21633_,
		_w21634_,
		_w21635_
	);
	LUT2 #(
		.INIT('h2)
	) name15809 (
		_w21231_,
		_w21635_,
		_w21636_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name15810 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21637_
	);
	LUT4 #(
		.INIT('h00d0)
	) name15811 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21638_
	);
	LUT4 #(
		.INIT('h2e26)
	) name15812 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21639_
	);
	LUT4 #(
		.INIT('h3210)
	) name15813 (
		_w21232_,
		_w21638_,
		_w21639_,
		_w21637_,
		_w21640_
	);
	LUT4 #(
		.INIT('hfd7e)
	) name15814 (
		_w21234_,
		_w21235_,
		_w21233_,
		_w21236_,
		_w21641_
	);
	LUT2 #(
		.INIT('h1)
	) name15815 (
		_w21232_,
		_w21641_,
		_w21642_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15816 (
		_w21233_,
		_w21232_,
		_w21240_,
		_w21237_,
		_w21643_
	);
	LUT4 #(
		.INIT('h0e00)
	) name15817 (
		_w21231_,
		_w21640_,
		_w21642_,
		_w21643_,
		_w21644_
	);
	LUT3 #(
		.INIT('h65)
	) name15818 (
		\u1_L4_reg[3]/NET0131 ,
		_w21636_,
		_w21644_,
		_w21645_
	);
	LUT4 #(
		.INIT('h8228)
	) name15819 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21646_
	);
	LUT3 #(
		.INIT('hbc)
	) name15820 (
		_w21068_,
		_w21065_,
		_w21066_,
		_w21647_
	);
	LUT4 #(
		.INIT('h0031)
	) name15821 (
		_w21072_,
		_w21300_,
		_w21647_,
		_w21646_,
		_w21648_
	);
	LUT4 #(
		.INIT('h9fff)
	) name15822 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21649_
	);
	LUT2 #(
		.INIT('h1)
	) name15823 (
		_w21064_,
		_w21649_,
		_w21650_
	);
	LUT4 #(
		.INIT('h4550)
	) name15824 (
		_w21064_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21651_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name15825 (
		_w21064_,
		_w21067_,
		_w21065_,
		_w21066_,
		_w21652_
	);
	LUT4 #(
		.INIT('hbf7d)
	) name15826 (
		_w21067_,
		_w21068_,
		_w21065_,
		_w21066_,
		_w21653_
	);
	LUT4 #(
		.INIT('hec00)
	) name15827 (
		_w21478_,
		_w21651_,
		_w21652_,
		_w21653_,
		_w21654_
	);
	LUT4 #(
		.INIT('h3210)
	) name15828 (
		_w21063_,
		_w21650_,
		_w21654_,
		_w21648_,
		_w21655_
	);
	LUT2 #(
		.INIT('h9)
	) name15829 (
		\u1_L4_reg[9]/NET0131 ,
		_w21655_,
		_w21656_
	);
	LUT4 #(
		.INIT('h0a20)
	) name15830 (
		_w21350_,
		_w21352_,
		_w21353_,
		_w21351_,
		_w21657_
	);
	LUT3 #(
		.INIT('he4)
	) name15831 (
		_w21353_,
		_w21351_,
		_w21354_,
		_w21658_
	);
	LUT3 #(
		.INIT('h74)
	) name15832 (
		_w21350_,
		_w21352_,
		_w21354_,
		_w21659_
	);
	LUT4 #(
		.INIT('h8a88)
	) name15833 (
		_w21349_,
		_w21657_,
		_w21658_,
		_w21659_,
		_w21660_
	);
	LUT4 #(
		.INIT('h8000)
	) name15834 (
		_w21350_,
		_w21352_,
		_w21353_,
		_w21351_,
		_w21661_
	);
	LUT4 #(
		.INIT('hdffc)
	) name15835 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21662_
	);
	LUT4 #(
		.INIT('h1003)
	) name15836 (
		_w21350_,
		_w21352_,
		_w21351_,
		_w21354_,
		_w21663_
	);
	LUT4 #(
		.INIT('h0100)
	) name15837 (
		_w21358_,
		_w21661_,
		_w21663_,
		_w21662_,
		_w21664_
	);
	LUT4 #(
		.INIT('h1000)
	) name15838 (
		_w21350_,
		_w21352_,
		_w21353_,
		_w21351_,
		_w21665_
	);
	LUT4 #(
		.INIT('h77ef)
	) name15839 (
		_w21352_,
		_w21353_,
		_w21351_,
		_w21354_,
		_w21666_
	);
	LUT3 #(
		.INIT('h31)
	) name15840 (
		_w21350_,
		_w21665_,
		_w21666_,
		_w21667_
	);
	LUT4 #(
		.INIT('h0e00)
	) name15841 (
		_w21349_,
		_w21664_,
		_w21660_,
		_w21667_,
		_w21668_
	);
	LUT2 #(
		.INIT('h9)
	) name15842 (
		\u1_L4_reg[18]/NET0131 ,
		_w21668_,
		_w21669_
	);
	LUT4 #(
		.INIT('hffda)
	) name15843 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w21670_
	);
	LUT2 #(
		.INIT('h1)
	) name15844 (
		_w5834_,
		_w21670_,
		_w21671_
	);
	LUT3 #(
		.INIT('h60)
	) name15845 (
		_w5832_,
		_w5829_,
		_w5834_,
		_w21672_
	);
	LUT2 #(
		.INIT('h2)
	) name15846 (
		_w5832_,
		_w5834_,
		_w21673_
	);
	LUT4 #(
		.INIT('h4404)
	) name15847 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5834_,
		_w21674_
	);
	LUT2 #(
		.INIT('h4)
	) name15848 (
		_w21672_,
		_w21674_,
		_w21675_
	);
	LUT2 #(
		.INIT('h4)
	) name15849 (
		_w5832_,
		_w5834_,
		_w21676_
	);
	LUT3 #(
		.INIT('hce)
	) name15850 (
		_w5827_,
		_w5832_,
		_w5834_,
		_w21677_
	);
	LUT2 #(
		.INIT('h8)
	) name15851 (
		_w5834_,
		_w5839_,
		_w21678_
	);
	LUT4 #(
		.INIT('h7707)
	) name15852 (
		_w5834_,
		_w5839_,
		_w5846_,
		_w21677_,
		_w21679_
	);
	LUT4 #(
		.INIT('h5455)
	) name15853 (
		_w5840_,
		_w21671_,
		_w21675_,
		_w21679_,
		_w21680_
	);
	LUT4 #(
		.INIT('hadfd)
	) name15854 (
		_w5828_,
		_w5827_,
		_w5829_,
		_w5834_,
		_w21681_
	);
	LUT2 #(
		.INIT('h1)
	) name15855 (
		_w5832_,
		_w21681_,
		_w21682_
	);
	LUT4 #(
		.INIT('hccaf)
	) name15856 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w21683_
	);
	LUT4 #(
		.INIT('h1110)
	) name15857 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w21684_
	);
	LUT3 #(
		.INIT('h08)
	) name15858 (
		_w5828_,
		_w5827_,
		_w5834_,
		_w21685_
	);
	LUT4 #(
		.INIT('h000d)
	) name15859 (
		_w5834_,
		_w21683_,
		_w21684_,
		_w21685_,
		_w21686_
	);
	LUT3 #(
		.INIT('h8a)
	) name15860 (
		_w5840_,
		_w21682_,
		_w21686_,
		_w21687_
	);
	LUT4 #(
		.INIT('h6ff3)
	) name15861 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w21688_
	);
	LUT2 #(
		.INIT('h1)
	) name15862 (
		_w5834_,
		_w21688_,
		_w21689_
	);
	LUT3 #(
		.INIT('h20)
	) name15863 (
		_w5832_,
		_w5829_,
		_w5834_,
		_w21690_
	);
	LUT4 #(
		.INIT('h0200)
	) name15864 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5834_,
		_w21691_
	);
	LUT3 #(
		.INIT('h07)
	) name15865 (
		_w5841_,
		_w21690_,
		_w21691_,
		_w21692_
	);
	LUT2 #(
		.INIT('h4)
	) name15866 (
		_w21689_,
		_w21692_,
		_w21693_
	);
	LUT4 #(
		.INIT('h5655)
	) name15867 (
		\u1_L3_reg[31]/NET0131 ,
		_w21687_,
		_w21680_,
		_w21693_,
		_w21694_
	);
	LUT4 #(
		.INIT('hc693)
	) name15868 (
		decrypt_pad,
		\u1_R3_reg[24]/NET0131 ,
		\u1_uk_K_r3_reg[29]/NET0131 ,
		\u1_uk_K_r3_reg[38]/NET0131 ,
		_w21695_
	);
	LUT4 #(
		.INIT('hc693)
	) name15869 (
		decrypt_pad,
		\u1_R3_reg[22]/NET0131 ,
		\u1_uk_K_r3_reg[14]/NET0131 ,
		\u1_uk_K_r3_reg[50]/NET0131 ,
		_w21696_
	);
	LUT4 #(
		.INIT('hc693)
	) name15870 (
		decrypt_pad,
		\u1_R3_reg[21]/NET0131 ,
		\u1_uk_K_r3_reg[23]/NET0131 ,
		\u1_uk_K_r3_reg[28]/NET0131 ,
		_w21697_
	);
	LUT4 #(
		.INIT('hc963)
	) name15871 (
		decrypt_pad,
		\u1_R3_reg[20]/NET0131 ,
		\u1_uk_K_r3_reg[44]/NET0131 ,
		\u1_uk_K_r3_reg[8]/NET0131 ,
		_w21698_
	);
	LUT4 #(
		.INIT('hc963)
	) name15872 (
		decrypt_pad,
		\u1_R3_reg[25]/NET0131 ,
		\u1_uk_K_r3_reg[29]/NET0131 ,
		\u1_uk_K_r3_reg[52]/NET0131 ,
		_w21699_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name15873 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21700_
	);
	LUT3 #(
		.INIT('h80)
	) name15874 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21701_
	);
	LUT4 #(
		.INIT('hc693)
	) name15875 (
		decrypt_pad,
		\u1_R3_reg[23]/NET0131 ,
		\u1_uk_K_r3_reg[31]/NET0131 ,
		\u1_uk_K_r3_reg[8]/NET0131 ,
		_w21702_
	);
	LUT4 #(
		.INIT('h00bf)
	) name15876 (
		_w21698_,
		_w21696_,
		_w21697_,
		_w21702_,
		_w21703_
	);
	LUT3 #(
		.INIT('h10)
	) name15877 (
		_w21701_,
		_w21700_,
		_w21703_,
		_w21704_
	);
	LUT4 #(
		.INIT('h0002)
	) name15878 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21705_
	);
	LUT4 #(
		.INIT('h27fd)
	) name15879 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21706_
	);
	LUT2 #(
		.INIT('h1)
	) name15880 (
		_w21696_,
		_w21702_,
		_w21707_
	);
	LUT4 #(
		.INIT('h0008)
	) name15881 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21702_,
		_w21708_
	);
	LUT2 #(
		.INIT('h4)
	) name15882 (
		_w21697_,
		_w21708_,
		_w21709_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name15883 (
		_w21697_,
		_w21702_,
		_w21706_,
		_w21708_,
		_w21710_
	);
	LUT3 #(
		.INIT('h8a)
	) name15884 (
		_w21695_,
		_w21704_,
		_w21710_,
		_w21711_
	);
	LUT3 #(
		.INIT('h04)
	) name15885 (
		_w21698_,
		_w21699_,
		_w21697_,
		_w21712_
	);
	LUT4 #(
		.INIT('hfa1a)
	) name15886 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21713_
	);
	LUT2 #(
		.INIT('h4)
	) name15887 (
		_w21713_,
		_w21702_,
		_w21714_
	);
	LUT4 #(
		.INIT('h0060)
	) name15888 (
		_w21698_,
		_w21696_,
		_w21697_,
		_w21702_,
		_w21715_
	);
	LUT4 #(
		.INIT('h0200)
	) name15889 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21716_
	);
	LUT4 #(
		.INIT('h0002)
	) name15890 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21702_,
		_w21717_
	);
	LUT4 #(
		.INIT('h0080)
	) name15891 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21718_
	);
	LUT4 #(
		.INIT('h0001)
	) name15892 (
		_w21716_,
		_w21717_,
		_w21718_,
		_w21715_,
		_w21719_
	);
	LUT3 #(
		.INIT('h45)
	) name15893 (
		_w21695_,
		_w21714_,
		_w21719_,
		_w21720_
	);
	LUT4 #(
		.INIT('h0100)
	) name15894 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21721_
	);
	LUT4 #(
		.INIT('h7e7f)
	) name15895 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21722_
	);
	LUT2 #(
		.INIT('h2)
	) name15896 (
		_w21702_,
		_w21722_,
		_w21723_
	);
	LUT3 #(
		.INIT('h01)
	) name15897 (
		_w21698_,
		_w21699_,
		_w21697_,
		_w21724_
	);
	LUT2 #(
		.INIT('h8)
	) name15898 (
		_w21707_,
		_w21724_,
		_w21725_
	);
	LUT3 #(
		.INIT('h20)
	) name15899 (
		_w21698_,
		_w21699_,
		_w21697_,
		_w21726_
	);
	LUT4 #(
		.INIT('hbabf)
	) name15900 (
		_w21696_,
		_w21712_,
		_w21702_,
		_w21726_,
		_w21727_
	);
	LUT3 #(
		.INIT('h10)
	) name15901 (
		_w21723_,
		_w21725_,
		_w21727_,
		_w21728_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name15902 (
		\u1_L3_reg[11]/NET0131 ,
		_w21720_,
		_w21711_,
		_w21728_,
		_w21729_
	);
	LUT4 #(
		.INIT('hc693)
	) name15903 (
		decrypt_pad,
		\u1_R3_reg[28]/NET0131 ,
		\u1_uk_K_r3_reg[36]/NET0131 ,
		\u1_uk_K_r3_reg[45]/NET0131 ,
		_w21730_
	);
	LUT4 #(
		.INIT('hc693)
	) name15904 (
		decrypt_pad,
		\u1_R3_reg[26]/NET0131 ,
		\u1_uk_K_r3_reg[16]/NET0131 ,
		\u1_uk_K_r3_reg[21]/NET0131 ,
		_w21731_
	);
	LUT4 #(
		.INIT('hc693)
	) name15905 (
		decrypt_pad,
		\u1_R3_reg[25]/NET0131 ,
		\u1_uk_K_r3_reg[0]/NET0131 ,
		\u1_uk_K_r3_reg[36]/NET0131 ,
		_w21732_
	);
	LUT4 #(
		.INIT('hc693)
	) name15906 (
		decrypt_pad,
		\u1_R3_reg[29]/NET0131 ,
		\u1_uk_K_r3_reg[28]/NET0131 ,
		\u1_uk_K_r3_reg[9]/NET0131 ,
		_w21733_
	);
	LUT3 #(
		.INIT('hea)
	) name15907 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21734_
	);
	LUT4 #(
		.INIT('hc963)
	) name15908 (
		decrypt_pad,
		\u1_R3_reg[24]/NET0131 ,
		\u1_uk_K_r3_reg[1]/NET0131 ,
		\u1_uk_K_r3_reg[51]/NET0131 ,
		_w21735_
	);
	LUT4 #(
		.INIT('hc963)
	) name15909 (
		decrypt_pad,
		\u1_R3_reg[27]/NET0131 ,
		\u1_uk_K_r3_reg[30]/NET0131 ,
		\u1_uk_K_r3_reg[49]/NET0131 ,
		_w21736_
	);
	LUT3 #(
		.INIT('h70)
	) name15910 (
		_w21731_,
		_w21732_,
		_w21736_,
		_w21737_
	);
	LUT4 #(
		.INIT('h7000)
	) name15911 (
		_w21731_,
		_w21732_,
		_w21735_,
		_w21736_,
		_w21738_
	);
	LUT2 #(
		.INIT('h8)
	) name15912 (
		_w21734_,
		_w21738_,
		_w21739_
	);
	LUT4 #(
		.INIT('h1000)
	) name15913 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21740_
	);
	LUT4 #(
		.INIT('hef3f)
	) name15914 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21741_
	);
	LUT2 #(
		.INIT('h2)
	) name15915 (
		_w21733_,
		_w21735_,
		_w21742_
	);
	LUT4 #(
		.INIT('h0020)
	) name15916 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21743_
	);
	LUT4 #(
		.INIT('hffde)
	) name15917 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21744_
	);
	LUT3 #(
		.INIT('he0)
	) name15918 (
		_w21736_,
		_w21741_,
		_w21744_,
		_w21745_
	);
	LUT3 #(
		.INIT('h8a)
	) name15919 (
		_w21730_,
		_w21739_,
		_w21745_,
		_w21746_
	);
	LUT4 #(
		.INIT('h0072)
	) name15920 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21736_,
		_w21747_
	);
	LUT4 #(
		.INIT('h10f0)
	) name15921 (
		_w21731_,
		_w21732_,
		_w21735_,
		_w21736_,
		_w21748_
	);
	LUT2 #(
		.INIT('h4)
	) name15922 (
		_w21747_,
		_w21748_,
		_w21749_
	);
	LUT4 #(
		.INIT('h0002)
	) name15923 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21750_
	);
	LUT2 #(
		.INIT('h6)
	) name15924 (
		_w21731_,
		_w21735_,
		_w21751_
	);
	LUT3 #(
		.INIT('h8c)
	) name15925 (
		_w21732_,
		_w21733_,
		_w21736_,
		_w21752_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name15926 (
		_w21750_,
		_w21736_,
		_w21751_,
		_w21752_,
		_w21753_
	);
	LUT4 #(
		.INIT('h0008)
	) name15927 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21754_
	);
	LUT4 #(
		.INIT('hfcd7)
	) name15928 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21755_
	);
	LUT4 #(
		.INIT('h0084)
	) name15929 (
		_w21731_,
		_w21732_,
		_w21735_,
		_w21736_,
		_w21756_
	);
	LUT4 #(
		.INIT('h0100)
	) name15930 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21736_,
		_w21757_
	);
	LUT4 #(
		.INIT('h0031)
	) name15931 (
		_w21736_,
		_w21756_,
		_w21755_,
		_w21757_,
		_w21758_
	);
	LUT4 #(
		.INIT('hba00)
	) name15932 (
		_w21730_,
		_w21749_,
		_w21753_,
		_w21758_,
		_w21759_
	);
	LUT3 #(
		.INIT('h65)
	) name15933 (
		\u1_L3_reg[22]/NET0131 ,
		_w21746_,
		_w21759_,
		_w21760_
	);
	LUT4 #(
		.INIT('hc693)
	) name15934 (
		decrypt_pad,
		\u1_R3_reg[16]/NET0131 ,
		\u1_uk_K_r3_reg[32]/NET0131 ,
		\u1_uk_K_r3_reg[41]/NET0131 ,
		_w21761_
	);
	LUT4 #(
		.INIT('hc693)
	) name15935 (
		decrypt_pad,
		\u1_R3_reg[12]/NET0131 ,
		\u1_uk_K_r3_reg[53]/NET0131 ,
		\u1_uk_K_r3_reg[5]/NET0131 ,
		_w21762_
	);
	LUT4 #(
		.INIT('hc693)
	) name15936 (
		decrypt_pad,
		\u1_R3_reg[17]/NET0131 ,
		\u1_uk_K_r3_reg[12]/NET0131 ,
		\u1_uk_K_r3_reg[46]/NET0131 ,
		_w21763_
	);
	LUT4 #(
		.INIT('hc963)
	) name15937 (
		decrypt_pad,
		\u1_R3_reg[13]/NET0131 ,
		\u1_uk_K_r3_reg[24]/NET0131 ,
		\u1_uk_K_r3_reg[47]/NET0131 ,
		_w21764_
	);
	LUT4 #(
		.INIT('hc693)
	) name15938 (
		decrypt_pad,
		\u1_R3_reg[15]/NET0131 ,
		\u1_uk_K_r3_reg[24]/NET0131 ,
		\u1_uk_K_r3_reg[33]/NET0131 ,
		_w21765_
	);
	LUT4 #(
		.INIT('h0080)
	) name15939 (
		_w21762_,
		_w21764_,
		_w21765_,
		_w21763_,
		_w21766_
	);
	LUT4 #(
		.INIT('hc963)
	) name15940 (
		decrypt_pad,
		\u1_R3_reg[14]/NET0131 ,
		\u1_uk_K_r3_reg[25]/NET0131 ,
		\u1_uk_K_r3_reg[48]/NET0131 ,
		_w21767_
	);
	LUT2 #(
		.INIT('h4)
	) name15941 (
		_w21762_,
		_w21763_,
		_w21768_
	);
	LUT4 #(
		.INIT('h0400)
	) name15942 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21769_
	);
	LUT2 #(
		.INIT('h1)
	) name15943 (
		_w21766_,
		_w21769_,
		_w21770_
	);
	LUT4 #(
		.INIT('h1000)
	) name15944 (
		_w21762_,
		_w21764_,
		_w21765_,
		_w21763_,
		_w21771_
	);
	LUT2 #(
		.INIT('h8)
	) name15945 (
		_w21762_,
		_w21763_,
		_w21772_
	);
	LUT4 #(
		.INIT('h8000)
	) name15946 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21773_
	);
	LUT2 #(
		.INIT('h1)
	) name15947 (
		_w21771_,
		_w21773_,
		_w21774_
	);
	LUT3 #(
		.INIT('h01)
	) name15948 (
		_w21762_,
		_w21764_,
		_w21763_,
		_w21775_
	);
	LUT2 #(
		.INIT('h4)
	) name15949 (
		_w21765_,
		_w21767_,
		_w21776_
	);
	LUT2 #(
		.INIT('h4)
	) name15950 (
		_w21762_,
		_w21764_,
		_w21777_
	);
	LUT4 #(
		.INIT('h0006)
	) name15951 (
		_w21762_,
		_w21764_,
		_w21765_,
		_w21767_,
		_w21778_
	);
	LUT3 #(
		.INIT('h07)
	) name15952 (
		_w21775_,
		_w21776_,
		_w21778_,
		_w21779_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15953 (
		_w21761_,
		_w21770_,
		_w21774_,
		_w21779_,
		_w21780_
	);
	LUT4 #(
		.INIT('hcc5f)
	) name15954 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21781_
	);
	LUT2 #(
		.INIT('h1)
	) name15955 (
		_w21765_,
		_w21781_,
		_w21782_
	);
	LUT4 #(
		.INIT('h0040)
	) name15956 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21783_
	);
	LUT2 #(
		.INIT('h8)
	) name15957 (
		_w21765_,
		_w21767_,
		_w21784_
	);
	LUT4 #(
		.INIT('h4000)
	) name15958 (
		_w21762_,
		_w21764_,
		_w21765_,
		_w21767_,
		_w21785_
	);
	LUT2 #(
		.INIT('h1)
	) name15959 (
		_w21783_,
		_w21785_,
		_w21786_
	);
	LUT3 #(
		.INIT('h72)
	) name15960 (
		_w21764_,
		_w21765_,
		_w21767_,
		_w21787_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name15961 (
		_w21772_,
		_w21787_,
		_w21775_,
		_w21776_,
		_w21788_
	);
	LUT4 #(
		.INIT('h00bf)
	) name15962 (
		_w21782_,
		_w21786_,
		_w21788_,
		_w21761_,
		_w21789_
	);
	LUT3 #(
		.INIT('h01)
	) name15963 (
		_w21762_,
		_w21767_,
		_w21763_,
		_w21790_
	);
	LUT4 #(
		.INIT('h0020)
	) name15964 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21791_
	);
	LUT4 #(
		.INIT('hffde)
	) name15965 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21792_
	);
	LUT2 #(
		.INIT('h2)
	) name15966 (
		_w21765_,
		_w21792_,
		_w21793_
	);
	LUT3 #(
		.INIT('h10)
	) name15967 (
		_w21765_,
		_w21767_,
		_w21763_,
		_w21794_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name15968 (
		_w21777_,
		_w21767_,
		_w21794_,
		_w21766_,
		_w21795_
	);
	LUT2 #(
		.INIT('h4)
	) name15969 (
		_w21793_,
		_w21795_,
		_w21796_
	);
	LUT4 #(
		.INIT('h5655)
	) name15970 (
		\u1_L3_reg[20]/NET0131 ,
		_w21789_,
		_w21780_,
		_w21796_,
		_w21797_
	);
	LUT4 #(
		.INIT('hdaff)
	) name15971 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21798_
	);
	LUT4 #(
		.INIT('h9aff)
	) name15972 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21799_
	);
	LUT2 #(
		.INIT('h2)
	) name15973 (
		_w21702_,
		_w21799_,
		_w21800_
	);
	LUT4 #(
		.INIT('h6f6e)
	) name15974 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21801_
	);
	LUT2 #(
		.INIT('h1)
	) name15975 (
		_w21702_,
		_w21801_,
		_w21802_
	);
	LUT4 #(
		.INIT('hffeb)
	) name15976 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21803_
	);
	LUT3 #(
		.INIT('h10)
	) name15977 (
		_w21717_,
		_w21718_,
		_w21803_,
		_w21804_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15978 (
		_w21695_,
		_w21800_,
		_w21802_,
		_w21804_,
		_w21805_
	);
	LUT4 #(
		.INIT('h67dc)
	) name15979 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21806_
	);
	LUT2 #(
		.INIT('h2)
	) name15980 (
		_w21702_,
		_w21806_,
		_w21807_
	);
	LUT4 #(
		.INIT('h0040)
	) name15981 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21808_
	);
	LUT4 #(
		.INIT('h0032)
	) name15982 (
		_w21702_,
		_w21708_,
		_w21798_,
		_w21808_,
		_w21809_
	);
	LUT4 #(
		.INIT('h2000)
	) name15983 (
		_w21699_,
		_w21696_,
		_w21697_,
		_w21702_,
		_w21810_
	);
	LUT2 #(
		.INIT('h1)
	) name15984 (
		_w21705_,
		_w21810_,
		_w21811_
	);
	LUT4 #(
		.INIT('hba00)
	) name15985 (
		_w21695_,
		_w21807_,
		_w21809_,
		_w21811_,
		_w21812_
	);
	LUT3 #(
		.INIT('h9a)
	) name15986 (
		\u1_L3_reg[29]/NET0131 ,
		_w21805_,
		_w21812_,
		_w21813_
	);
	LUT4 #(
		.INIT('hc963)
	) name15987 (
		decrypt_pad,
		\u1_R3_reg[8]/NET0131 ,
		\u1_uk_K_r3_reg[40]/NET0131 ,
		\u1_uk_K_r3_reg[6]/NET0131 ,
		_w21814_
	);
	LUT4 #(
		.INIT('hc963)
	) name15988 (
		decrypt_pad,
		\u1_R3_reg[7]/NET0131 ,
		\u1_uk_K_r3_reg[17]/NET0131 ,
		\u1_uk_K_r3_reg[40]/NET0131 ,
		_w21815_
	);
	LUT4 #(
		.INIT('hc963)
	) name15989 (
		decrypt_pad,
		\u1_R3_reg[5]/NET0131 ,
		\u1_uk_K_r3_reg[32]/NET0131 ,
		\u1_uk_K_r3_reg[55]/NET0131 ,
		_w21816_
	);
	LUT4 #(
		.INIT('hc693)
	) name15990 (
		decrypt_pad,
		\u1_R3_reg[4]/NET0131 ,
		\u1_uk_K_r3_reg[19]/NET0131 ,
		\u1_uk_K_r3_reg[53]/NET0131 ,
		_w21817_
	);
	LUT4 #(
		.INIT('hc693)
	) name15991 (
		decrypt_pad,
		\u1_R3_reg[9]/NET0131 ,
		\u1_uk_K_r3_reg[11]/NET0131 ,
		\u1_uk_K_r3_reg[20]/NET0131 ,
		_w21818_
	);
	LUT4 #(
		.INIT('hc693)
	) name15992 (
		decrypt_pad,
		\u1_R3_reg[6]/NET0131 ,
		\u1_uk_K_r3_reg[46]/NET0131 ,
		\u1_uk_K_r3_reg[55]/NET0131 ,
		_w21819_
	);
	LUT4 #(
		.INIT('h59fb)
	) name15993 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21820_
	);
	LUT2 #(
		.INIT('h1)
	) name15994 (
		_w21815_,
		_w21820_,
		_w21821_
	);
	LUT4 #(
		.INIT('h0034)
	) name15995 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21822_
	);
	LUT4 #(
		.INIT('h0800)
	) name15996 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21823_
	);
	LUT2 #(
		.INIT('h2)
	) name15997 (
		_w21818_,
		_w21819_,
		_w21824_
	);
	LUT4 #(
		.INIT('h0004)
	) name15998 (
		_w21815_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21825_
	);
	LUT4 #(
		.INIT('h4000)
	) name15999 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21826_
	);
	LUT4 #(
		.INIT('h0007)
	) name16000 (
		_w21815_,
		_w21823_,
		_w21825_,
		_w21826_,
		_w21827_
	);
	LUT4 #(
		.INIT('h5455)
	) name16001 (
		_w21814_,
		_w21821_,
		_w21822_,
		_w21827_,
		_w21828_
	);
	LUT4 #(
		.INIT('he6ee)
	) name16002 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21829_
	);
	LUT4 #(
		.INIT('h4044)
	) name16003 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21830_
	);
	LUT3 #(
		.INIT('h51)
	) name16004 (
		_w21815_,
		_w21816_,
		_w21819_,
		_w21831_
	);
	LUT4 #(
		.INIT('hf200)
	) name16005 (
		_w21814_,
		_w21829_,
		_w21830_,
		_w21831_,
		_w21832_
	);
	LUT3 #(
		.INIT('h10)
	) name16006 (
		_w21818_,
		_w21816_,
		_w21819_,
		_w21833_
	);
	LUT4 #(
		.INIT('h0100)
	) name16007 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21834_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name16008 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21835_
	);
	LUT2 #(
		.INIT('h2)
	) name16009 (
		_w21815_,
		_w21835_,
		_w21836_
	);
	LUT4 #(
		.INIT('h0082)
	) name16010 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21837_
	);
	LUT4 #(
		.INIT('h80a0)
	) name16011 (
		_w21815_,
		_w21817_,
		_w21816_,
		_w21819_,
		_w21838_
	);
	LUT3 #(
		.INIT('ha8)
	) name16012 (
		_w21814_,
		_w21837_,
		_w21838_,
		_w21839_
	);
	LUT3 #(
		.INIT('h01)
	) name16013 (
		_w21836_,
		_w21839_,
		_w21832_,
		_w21840_
	);
	LUT3 #(
		.INIT('h65)
	) name16014 (
		\u1_L3_reg[2]/NET0131 ,
		_w21828_,
		_w21840_,
		_w21841_
	);
	LUT4 #(
		.INIT('h0800)
	) name16015 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21702_,
		_w21842_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name16016 (
		_w21695_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21843_
	);
	LUT3 #(
		.INIT('h10)
	) name16017 (
		_w21721_,
		_w21842_,
		_w21843_,
		_w21844_
	);
	LUT4 #(
		.INIT('hd97b)
	) name16018 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21845_
	);
	LUT2 #(
		.INIT('h2)
	) name16019 (
		_w21702_,
		_w21845_,
		_w21846_
	);
	LUT3 #(
		.INIT('h01)
	) name16020 (
		_w21695_,
		_w21705_,
		_w21708_,
		_w21847_
	);
	LUT3 #(
		.INIT('h45)
	) name16021 (
		_w21844_,
		_w21846_,
		_w21847_,
		_w21848_
	);
	LUT4 #(
		.INIT('heebf)
	) name16022 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21849_
	);
	LUT3 #(
		.INIT('h01)
	) name16023 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21850_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name16024 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w21851_
	);
	LUT4 #(
		.INIT('h3210)
	) name16025 (
		_w21695_,
		_w21850_,
		_w21849_,
		_w21851_,
		_w21852_
	);
	LUT4 #(
		.INIT('h007d)
	) name16026 (
		_w21698_,
		_w21699_,
		_w21697_,
		_w21702_,
		_w21853_
	);
	LUT3 #(
		.INIT('hbe)
	) name16027 (
		_w21698_,
		_w21699_,
		_w21697_,
		_w21854_
	);
	LUT4 #(
		.INIT('h9e00)
	) name16028 (
		_w21698_,
		_w21699_,
		_w21697_,
		_w21702_,
		_w21855_
	);
	LUT3 #(
		.INIT('h02)
	) name16029 (
		_w21696_,
		_w21855_,
		_w21853_,
		_w21856_
	);
	LUT3 #(
		.INIT('h0e)
	) name16030 (
		_w21702_,
		_w21852_,
		_w21856_,
		_w21857_
	);
	LUT3 #(
		.INIT('h65)
	) name16031 (
		\u1_L3_reg[4]/NET0131 ,
		_w21848_,
		_w21857_,
		_w21858_
	);
	LUT4 #(
		.INIT('hc693)
	) name16032 (
		decrypt_pad,
		\u1_R3_reg[29]/NET0131 ,
		\u1_uk_K_r3_reg[37]/NET0131 ,
		\u1_uk_K_r3_reg[42]/NET0131 ,
		_w21859_
	);
	LUT4 #(
		.INIT('hc693)
	) name16033 (
		decrypt_pad,
		\u1_R3_reg[1]/NET0131 ,
		\u1_uk_K_r3_reg[22]/NET0131 ,
		\u1_uk_K_r3_reg[31]/NET0131 ,
		_w21860_
	);
	LUT4 #(
		.INIT('hc963)
	) name16034 (
		decrypt_pad,
		\u1_R3_reg[30]/NET0131 ,
		\u1_uk_K_r3_reg[43]/NET0131 ,
		\u1_uk_K_r3_reg[7]/NET0131 ,
		_w21861_
	);
	LUT4 #(
		.INIT('hc963)
	) name16035 (
		decrypt_pad,
		\u1_R3_reg[28]/NET0131 ,
		\u1_uk_K_r3_reg[15]/NET0131 ,
		\u1_uk_K_r3_reg[38]/NET0131 ,
		_w21862_
	);
	LUT2 #(
		.INIT('h4)
	) name16036 (
		_w21861_,
		_w21862_,
		_w21863_
	);
	LUT4 #(
		.INIT('h0400)
	) name16037 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21864_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16038 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21865_
	);
	LUT4 #(
		.INIT('hc963)
	) name16039 (
		decrypt_pad,
		\u1_R3_reg[31]/P0001 ,
		\u1_uk_K_r3_reg[0]/NET0131 ,
		\u1_uk_K_r3_reg[50]/NET0131 ,
		_w21866_
	);
	LUT3 #(
		.INIT('h10)
	) name16040 (
		_w21865_,
		_w21864_,
		_w21866_,
		_w21867_
	);
	LUT4 #(
		.INIT('h0001)
	) name16041 (
		_w21861_,
		_w21862_,
		_w21859_,
		_w21866_,
		_w21868_
	);
	LUT4 #(
		.INIT('h2000)
	) name16042 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21869_
	);
	LUT4 #(
		.INIT('hc693)
	) name16043 (
		decrypt_pad,
		\u1_R3_reg[32]/NET0131 ,
		\u1_uk_K_r3_reg[1]/NET0131 ,
		\u1_uk_K_r3_reg[37]/NET0131 ,
		_w21870_
	);
	LUT3 #(
		.INIT('h04)
	) name16044 (
		_w21869_,
		_w21870_,
		_w21868_,
		_w21871_
	);
	LUT4 #(
		.INIT('h0008)
	) name16045 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21872_
	);
	LUT4 #(
		.INIT('hfb00)
	) name16046 (
		_w21862_,
		_w21860_,
		_w21859_,
		_w21866_,
		_w21873_
	);
	LUT3 #(
		.INIT('h02)
	) name16047 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21874_
	);
	LUT3 #(
		.INIT('h07)
	) name16048 (
		_w21860_,
		_w21859_,
		_w21866_,
		_w21875_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16049 (
		_w21872_,
		_w21873_,
		_w21874_,
		_w21875_,
		_w21876_
	);
	LUT3 #(
		.INIT('hb0)
	) name16050 (
		_w21860_,
		_w21859_,
		_w21866_,
		_w21877_
	);
	LUT4 #(
		.INIT('h8000)
	) name16051 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21878_
	);
	LUT4 #(
		.INIT('h0301)
	) name16052 (
		_w21863_,
		_w21870_,
		_w21878_,
		_w21877_,
		_w21879_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16053 (
		_w21867_,
		_w21871_,
		_w21876_,
		_w21879_,
		_w21880_
	);
	LUT4 #(
		.INIT('h00f7)
	) name16054 (
		_w21861_,
		_w21862_,
		_w21859_,
		_w21866_,
		_w21881_
	);
	LUT2 #(
		.INIT('h1)
	) name16055 (
		_w21866_,
		_w21870_,
		_w21882_
	);
	LUT3 #(
		.INIT('h54)
	) name16056 (
		_w21864_,
		_w21881_,
		_w21882_,
		_w21883_
	);
	LUT4 #(
		.INIT('h0001)
	) name16057 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21884_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name16058 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21885_
	);
	LUT4 #(
		.INIT('h0020)
	) name16059 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21886_
	);
	LUT4 #(
		.INIT('h0040)
	) name16060 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21887_
	);
	LUT4 #(
		.INIT('h0008)
	) name16061 (
		_w21866_,
		_w21885_,
		_w21886_,
		_w21887_,
		_w21888_
	);
	LUT2 #(
		.INIT('h1)
	) name16062 (
		_w21883_,
		_w21888_,
		_w21889_
	);
	LUT3 #(
		.INIT('ha9)
	) name16063 (
		\u1_L3_reg[5]/NET0131 ,
		_w21880_,
		_w21889_,
		_w21890_
	);
	LUT4 #(
		.INIT('hfb5d)
	) name16064 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21891_
	);
	LUT4 #(
		.INIT('h6fff)
	) name16065 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21892_
	);
	LUT3 #(
		.INIT('h02)
	) name16066 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21893_
	);
	LUT4 #(
		.INIT('hfdbb)
	) name16067 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21894_
	);
	LUT4 #(
		.INIT('hc480)
	) name16068 (
		_w21765_,
		_w21892_,
		_w21894_,
		_w21891_,
		_w21895_
	);
	LUT2 #(
		.INIT('h2)
	) name16069 (
		_w21761_,
		_w21895_,
		_w21896_
	);
	LUT4 #(
		.INIT('hb4b1)
	) name16070 (
		_w21764_,
		_w21765_,
		_w21767_,
		_w21763_,
		_w21897_
	);
	LUT2 #(
		.INIT('h2)
	) name16071 (
		_w21762_,
		_w21897_,
		_w21898_
	);
	LUT4 #(
		.INIT('hafee)
	) name16072 (
		_w21762_,
		_w21764_,
		_w21765_,
		_w21763_,
		_w21899_
	);
	LUT3 #(
		.INIT('h54)
	) name16073 (
		_w21783_,
		_w21784_,
		_w21899_,
		_w21900_
	);
	LUT3 #(
		.INIT('h45)
	) name16074 (
		_w21761_,
		_w21898_,
		_w21900_,
		_w21901_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name16075 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w21902_
	);
	LUT2 #(
		.INIT('h1)
	) name16076 (
		_w21765_,
		_w21902_,
		_w21903_
	);
	LUT3 #(
		.INIT('h23)
	) name16077 (
		_w21767_,
		_w21785_,
		_w21766_,
		_w21904_
	);
	LUT2 #(
		.INIT('h4)
	) name16078 (
		_w21903_,
		_w21904_,
		_w21905_
	);
	LUT4 #(
		.INIT('h5655)
	) name16079 (
		\u1_L3_reg[10]/NET0131 ,
		_w21901_,
		_w21896_,
		_w21905_,
		_w21906_
	);
	LUT4 #(
		.INIT('h0006)
	) name16080 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21907_
	);
	LUT3 #(
		.INIT('h47)
	) name16081 (
		_w21731_,
		_w21732_,
		_w21736_,
		_w21908_
	);
	LUT4 #(
		.INIT('h0051)
	) name16082 (
		_w21730_,
		_w21742_,
		_w21908_,
		_w21907_,
		_w21909_
	);
	LUT3 #(
		.INIT('h10)
	) name16083 (
		_w21731_,
		_w21733_,
		_w21735_,
		_w21910_
	);
	LUT4 #(
		.INIT('h2100)
	) name16084 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21911_
	);
	LUT2 #(
		.INIT('h6)
	) name16085 (
		_w21732_,
		_w21733_,
		_w21912_
	);
	LUT4 #(
		.INIT('h143c)
	) name16086 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21913_
	);
	LUT3 #(
		.INIT('h32)
	) name16087 (
		_w21736_,
		_w21911_,
		_w21913_,
		_w21914_
	);
	LUT2 #(
		.INIT('h8)
	) name16088 (
		_w21909_,
		_w21914_,
		_w21915_
	);
	LUT2 #(
		.INIT('h4)
	) name16089 (
		_w21736_,
		_w21743_,
		_w21916_
	);
	LUT3 #(
		.INIT('h02)
	) name16090 (
		_w21730_,
		_w21740_,
		_w21754_,
		_w21917_
	);
	LUT4 #(
		.INIT('h0240)
	) name16091 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21918_
	);
	LUT4 #(
		.INIT('h33fe)
	) name16092 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w21919_
	);
	LUT3 #(
		.INIT('h31)
	) name16093 (
		_w21736_,
		_w21918_,
		_w21919_,
		_w21920_
	);
	LUT3 #(
		.INIT('h40)
	) name16094 (
		_w21916_,
		_w21917_,
		_w21920_,
		_w21921_
	);
	LUT3 #(
		.INIT('ha9)
	) name16095 (
		\u1_L3_reg[12]/NET0131 ,
		_w21915_,
		_w21921_,
		_w21922_
	);
	LUT4 #(
		.INIT('hc693)
	) name16096 (
		decrypt_pad,
		\u1_R3_reg[19]/NET0131 ,
		\u1_uk_K_r3_reg[2]/NET0131 ,
		\u1_uk_K_r3_reg[7]/NET0131 ,
		_w21923_
	);
	LUT4 #(
		.INIT('hc693)
	) name16097 (
		decrypt_pad,
		\u1_R3_reg[18]/NET0131 ,
		\u1_uk_K_r3_reg[15]/NET0131 ,
		\u1_uk_K_r3_reg[51]/NET0131 ,
		_w21924_
	);
	LUT4 #(
		.INIT('hc963)
	) name16098 (
		decrypt_pad,
		\u1_R3_reg[21]/NET0131 ,
		\u1_uk_K_r3_reg[23]/NET0131 ,
		\u1_uk_K_r3_reg[42]/NET0131 ,
		_w21925_
	);
	LUT4 #(
		.INIT('hc693)
	) name16099 (
		decrypt_pad,
		\u1_R3_reg[16]/NET0131 ,
		\u1_uk_K_r3_reg[30]/NET0131 ,
		\u1_uk_K_r3_reg[35]/NET0131 ,
		_w21926_
	);
	LUT4 #(
		.INIT('hc693)
	) name16100 (
		decrypt_pad,
		\u1_R3_reg[17]/NET0131 ,
		\u1_uk_K_r3_reg[21]/NET0131 ,
		\u1_uk_K_r3_reg[2]/NET0131 ,
		_w21927_
	);
	LUT4 #(
		.INIT('h0040)
	) name16101 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21928_
	);
	LUT4 #(
		.INIT('hefbf)
	) name16102 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21929_
	);
	LUT3 #(
		.INIT('h04)
	) name16103 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21930_
	);
	LUT4 #(
		.INIT('h0001)
	) name16104 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21931_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name16105 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21932_
	);
	LUT3 #(
		.INIT('h40)
	) name16106 (
		_w21923_,
		_w21929_,
		_w21932_,
		_w21933_
	);
	LUT4 #(
		.INIT('h0200)
	) name16107 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21934_
	);
	LUT4 #(
		.INIT('hfdef)
	) name16108 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21935_
	);
	LUT4 #(
		.INIT('hdf00)
	) name16109 (
		_w21926_,
		_w21925_,
		_w21927_,
		_w21923_,
		_w21936_
	);
	LUT2 #(
		.INIT('h8)
	) name16110 (
		_w21926_,
		_w21925_,
		_w21937_
	);
	LUT4 #(
		.INIT('hb7b3)
	) name16111 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21938_
	);
	LUT3 #(
		.INIT('h80)
	) name16112 (
		_w21936_,
		_w21935_,
		_w21938_,
		_w21939_
	);
	LUT3 #(
		.INIT('he6)
	) name16113 (
		_w21924_,
		_w21927_,
		_w21923_,
		_w21940_
	);
	LUT2 #(
		.INIT('h2)
	) name16114 (
		_w21937_,
		_w21940_,
		_w21941_
	);
	LUT4 #(
		.INIT('h0020)
	) name16115 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21942_
	);
	LUT4 #(
		.INIT('hc963)
	) name16116 (
		decrypt_pad,
		\u1_R3_reg[20]/NET0131 ,
		\u1_uk_K_r3_reg[22]/NET0131 ,
		\u1_uk_K_r3_reg[45]/NET0131 ,
		_w21943_
	);
	LUT3 #(
		.INIT('h10)
	) name16117 (
		_w21934_,
		_w21942_,
		_w21943_,
		_w21944_
	);
	LUT4 #(
		.INIT('h0e00)
	) name16118 (
		_w21933_,
		_w21939_,
		_w21941_,
		_w21944_,
		_w21945_
	);
	LUT4 #(
		.INIT('h0800)
	) name16119 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21946_
	);
	LUT4 #(
		.INIT('h0002)
	) name16120 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21947_
	);
	LUT4 #(
		.INIT('hc7b9)
	) name16121 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21948_
	);
	LUT3 #(
		.INIT('h40)
	) name16122 (
		_w21923_,
		_w21929_,
		_w21948_,
		_w21949_
	);
	LUT4 #(
		.INIT('h8091)
	) name16123 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21950_
	);
	LUT3 #(
		.INIT('h10)
	) name16124 (
		_w21926_,
		_w21924_,
		_w21927_,
		_w21951_
	);
	LUT4 #(
		.INIT('hef00)
	) name16125 (
		_w21926_,
		_w21924_,
		_w21927_,
		_w21923_,
		_w21952_
	);
	LUT3 #(
		.INIT('h20)
	) name16126 (
		_w21935_,
		_w21950_,
		_w21952_,
		_w21953_
	);
	LUT4 #(
		.INIT('h0100)
	) name16127 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21954_
	);
	LUT4 #(
		.INIT('h0080)
	) name16128 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w21955_
	);
	LUT3 #(
		.INIT('h01)
	) name16129 (
		_w21943_,
		_w21955_,
		_w21954_,
		_w21956_
	);
	LUT3 #(
		.INIT('he0)
	) name16130 (
		_w21949_,
		_w21953_,
		_w21956_,
		_w21957_
	);
	LUT3 #(
		.INIT('ha9)
	) name16131 (
		\u1_L3_reg[14]/NET0131 ,
		_w21945_,
		_w21957_,
		_w21958_
	);
	LUT4 #(
		.INIT('h32cf)
	) name16132 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21959_
	);
	LUT4 #(
		.INIT('h0004)
	) name16133 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21960_
	);
	LUT4 #(
		.INIT('h0031)
	) name16134 (
		_w21866_,
		_w21870_,
		_w21959_,
		_w21960_,
		_w21961_
	);
	LUT4 #(
		.INIT('hbf00)
	) name16135 (
		_w21861_,
		_w21862_,
		_w21859_,
		_w21870_,
		_w21962_
	);
	LUT4 #(
		.INIT('h0100)
	) name16136 (
		_w21862_,
		_w21860_,
		_w21859_,
		_w21866_,
		_w21963_
	);
	LUT4 #(
		.INIT('h0008)
	) name16137 (
		_w21861_,
		_w21860_,
		_w21859_,
		_w21866_,
		_w21964_
	);
	LUT4 #(
		.INIT('h0080)
	) name16138 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21965_
	);
	LUT4 #(
		.INIT('hfd7f)
	) name16139 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21966_
	);
	LUT4 #(
		.INIT('h1000)
	) name16140 (
		_w21963_,
		_w21964_,
		_w21962_,
		_w21966_,
		_w21967_
	);
	LUT2 #(
		.INIT('h1)
	) name16141 (
		_w21961_,
		_w21967_,
		_w21968_
	);
	LUT4 #(
		.INIT('h1000)
	) name16142 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21969_
	);
	LUT3 #(
		.INIT('h08)
	) name16143 (
		_w21881_,
		_w21885_,
		_w21969_,
		_w21970_
	);
	LUT4 #(
		.INIT('h0010)
	) name16144 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w21971_
	);
	LUT3 #(
		.INIT('h04)
	) name16145 (
		_w21869_,
		_w21866_,
		_w21971_,
		_w21972_
	);
	LUT4 #(
		.INIT('h0002)
	) name16146 (
		_w21862_,
		_w21859_,
		_w21866_,
		_w21870_,
		_w21973_
	);
	LUT3 #(
		.INIT('h0e)
	) name16147 (
		_w21970_,
		_w21972_,
		_w21973_,
		_w21974_
	);
	LUT3 #(
		.INIT('h65)
	) name16148 (
		\u1_L3_reg[15]/P0001 ,
		_w21968_,
		_w21974_,
		_w21975_
	);
	LUT4 #(
		.INIT('h5515)
	) name16149 (
		_w21815_,
		_w21817_,
		_w21818_,
		_w21816_,
		_w21976_
	);
	LUT3 #(
		.INIT('h40)
	) name16150 (
		_w21817_,
		_w21818_,
		_w21819_,
		_w21977_
	);
	LUT3 #(
		.INIT('h01)
	) name16151 (
		_w21818_,
		_w21816_,
		_w21819_,
		_w21978_
	);
	LUT4 #(
		.INIT('haaa8)
	) name16152 (
		_w21815_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21979_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16153 (
		_w21833_,
		_w21976_,
		_w21977_,
		_w21979_,
		_w21980_
	);
	LUT4 #(
		.INIT('h0010)
	) name16154 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21981_
	);
	LUT4 #(
		.INIT('h0002)
	) name16155 (
		_w21814_,
		_w21825_,
		_w21826_,
		_w21981_,
		_w21982_
	);
	LUT2 #(
		.INIT('h4)
	) name16156 (
		_w21980_,
		_w21982_,
		_w21983_
	);
	LUT3 #(
		.INIT('h32)
	) name16157 (
		_w21815_,
		_w21817_,
		_w21816_,
		_w21984_
	);
	LUT2 #(
		.INIT('h8)
	) name16158 (
		_w21824_,
		_w21984_,
		_w21985_
	);
	LUT2 #(
		.INIT('h8)
	) name16159 (
		_w21815_,
		_w21817_,
		_w21986_
	);
	LUT3 #(
		.INIT('hb0)
	) name16160 (
		_w21818_,
		_w21816_,
		_w21819_,
		_w21987_
	);
	LUT3 #(
		.INIT('h15)
	) name16161 (
		_w21814_,
		_w21986_,
		_w21987_,
		_w21988_
	);
	LUT4 #(
		.INIT('h5455)
	) name16162 (
		_w21815_,
		_w21817_,
		_w21818_,
		_w21816_,
		_w21989_
	);
	LUT4 #(
		.INIT('h0400)
	) name16163 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21990_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name16164 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21991_
	);
	LUT2 #(
		.INIT('h8)
	) name16165 (
		_w21989_,
		_w21991_,
		_w21992_
	);
	LUT3 #(
		.INIT('h40)
	) name16166 (
		_w21985_,
		_w21988_,
		_w21992_,
		_w21993_
	);
	LUT4 #(
		.INIT('h2000)
	) name16167 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21994_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name16168 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21995_
	);
	LUT3 #(
		.INIT('h09)
	) name16169 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21996_
	);
	LUT3 #(
		.INIT('h02)
	) name16170 (
		_w21817_,
		_w21818_,
		_w21819_,
		_w21997_
	);
	LUT4 #(
		.INIT('h0020)
	) name16171 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w21998_
	);
	LUT3 #(
		.INIT('h02)
	) name16172 (
		_w21815_,
		_w21998_,
		_w21996_,
		_w21999_
	);
	LUT3 #(
		.INIT('h40)
	) name16173 (
		_w21985_,
		_w21988_,
		_w21999_,
		_w22000_
	);
	LUT4 #(
		.INIT('h001f)
	) name16174 (
		_w21983_,
		_w21993_,
		_w21995_,
		_w22000_,
		_w22001_
	);
	LUT2 #(
		.INIT('h9)
	) name16175 (
		\u1_L3_reg[13]/NET0131 ,
		_w22001_,
		_w22002_
	);
	LUT4 #(
		.INIT('h4e55)
	) name16176 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w22003_
	);
	LUT4 #(
		.INIT('h8000)
	) name16177 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w22004_
	);
	LUT4 #(
		.INIT('h0e04)
	) name16178 (
		_w21702_,
		_w21854_,
		_w22004_,
		_w22003_,
		_w22005_
	);
	LUT2 #(
		.INIT('h1)
	) name16179 (
		_w21695_,
		_w22005_,
		_w22006_
	);
	LUT4 #(
		.INIT('h4010)
	) name16180 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w22007_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name16181 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w22008_
	);
	LUT3 #(
		.INIT('h02)
	) name16182 (
		_w21698_,
		_w21697_,
		_w21702_,
		_w22009_
	);
	LUT4 #(
		.INIT('hfcfb)
	) name16183 (
		_w21698_,
		_w21699_,
		_w21696_,
		_w21697_,
		_w22010_
	);
	LUT4 #(
		.INIT('h0d00)
	) name16184 (
		_w21702_,
		_w22008_,
		_w22009_,
		_w22010_,
		_w22011_
	);
	LUT3 #(
		.INIT('h8a)
	) name16185 (
		_w21695_,
		_w22007_,
		_w22011_,
		_w22012_
	);
	LUT2 #(
		.INIT('h2)
	) name16186 (
		_w21727_,
		_w21709_,
		_w22013_
	);
	LUT4 #(
		.INIT('h5655)
	) name16187 (
		\u1_L3_reg[19]/NET0131 ,
		_w22012_,
		_w22006_,
		_w22013_,
		_w22014_
	);
	LUT4 #(
		.INIT('h220a)
	) name16188 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w22015_
	);
	LUT4 #(
		.INIT('hfda8)
	) name16189 (
		_w21765_,
		_w21790_,
		_w21791_,
		_w22015_,
		_w22016_
	);
	LUT4 #(
		.INIT('h7bf7)
	) name16190 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w22017_
	);
	LUT3 #(
		.INIT('h45)
	) name16191 (
		_w21761_,
		_w22016_,
		_w22017_,
		_w22018_
	);
	LUT4 #(
		.INIT('hb3fb)
	) name16192 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w22019_
	);
	LUT4 #(
		.INIT('h0080)
	) name16193 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w22020_
	);
	LUT4 #(
		.INIT('hef6f)
	) name16194 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w22021_
	);
	LUT4 #(
		.INIT('h04cc)
	) name16195 (
		_w21765_,
		_w21761_,
		_w22019_,
		_w22021_,
		_w22022_
	);
	LUT4 #(
		.INIT('h6fbf)
	) name16196 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w22023_
	);
	LUT2 #(
		.INIT('h2)
	) name16197 (
		_w21765_,
		_w22023_,
		_w22024_
	);
	LUT4 #(
		.INIT('hccfd)
	) name16198 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w22025_
	);
	LUT2 #(
		.INIT('h8)
	) name16199 (
		_w21765_,
		_w21761_,
		_w22026_
	);
	LUT2 #(
		.INIT('h4)
	) name16200 (
		_w22025_,
		_w22026_,
		_w22027_
	);
	LUT4 #(
		.INIT('haabf)
	) name16201 (
		_w21765_,
		_w21767_,
		_w21775_,
		_w22020_,
		_w22028_
	);
	LUT4 #(
		.INIT('h0100)
	) name16202 (
		_w22024_,
		_w22027_,
		_w22022_,
		_w22028_,
		_w22029_
	);
	LUT3 #(
		.INIT('h65)
	) name16203 (
		\u1_L3_reg[1]/NET0131 ,
		_w22018_,
		_w22029_,
		_w22030_
	);
	LUT4 #(
		.INIT('h4000)
	) name16204 (
		_w5828_,
		_w5827_,
		_w5829_,
		_w5834_,
		_w22031_
	);
	LUT4 #(
		.INIT('h0013)
	) name16205 (
		_w5841_,
		_w5847_,
		_w21690_,
		_w22031_,
		_w22032_
	);
	LUT3 #(
		.INIT('h8a)
	) name16206 (
		_w5840_,
		_w21678_,
		_w22032_,
		_w22033_
	);
	LUT4 #(
		.INIT('h4080)
	) name16207 (
		_w5828_,
		_w5832_,
		_w5829_,
		_w5834_,
		_w22034_
	);
	LUT3 #(
		.INIT('h04)
	) name16208 (
		_w5828_,
		_w5827_,
		_w5829_,
		_w22035_
	);
	LUT4 #(
		.INIT('h0400)
	) name16209 (
		_w5828_,
		_w5827_,
		_w5829_,
		_w5834_,
		_w22036_
	);
	LUT3 #(
		.INIT('h01)
	) name16210 (
		_w5827_,
		_w5832_,
		_w5829_,
		_w22037_
	);
	LUT4 #(
		.INIT('h0001)
	) name16211 (
		_w5851_,
		_w21685_,
		_w22037_,
		_w22036_,
		_w22038_
	);
	LUT3 #(
		.INIT('h45)
	) name16212 (
		_w5840_,
		_w22034_,
		_w22038_,
		_w22039_
	);
	LUT4 #(
		.INIT('hee9b)
	) name16213 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w22040_
	);
	LUT2 #(
		.INIT('h4)
	) name16214 (
		_w5834_,
		_w5840_,
		_w22041_
	);
	LUT2 #(
		.INIT('h4)
	) name16215 (
		_w22040_,
		_w22041_,
		_w22042_
	);
	LUT4 #(
		.INIT('hfef7)
	) name16216 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w22043_
	);
	LUT2 #(
		.INIT('h1)
	) name16217 (
		_w5834_,
		_w22043_,
		_w22044_
	);
	LUT2 #(
		.INIT('h8)
	) name16218 (
		_w5830_,
		_w21673_,
		_w22045_
	);
	LUT3 #(
		.INIT('h13)
	) name16219 (
		_w21676_,
		_w21691_,
		_w22035_,
		_w22046_
	);
	LUT4 #(
		.INIT('h0100)
	) name16220 (
		_w22044_,
		_w22045_,
		_w22042_,
		_w22046_,
		_w22047_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name16221 (
		\u1_L3_reg[23]/NET0131 ,
		_w22039_,
		_w22033_,
		_w22047_,
		_w22048_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name16222 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w22049_
	);
	LUT2 #(
		.INIT('h2)
	) name16223 (
		_w21815_,
		_w22049_,
		_w22050_
	);
	LUT4 #(
		.INIT('hbfae)
	) name16224 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w22051_
	);
	LUT2 #(
		.INIT('h1)
	) name16225 (
		_w21815_,
		_w22051_,
		_w22052_
	);
	LUT4 #(
		.INIT('h7737)
	) name16226 (
		_w21815_,
		_w21817_,
		_w21818_,
		_w21816_,
		_w22053_
	);
	LUT3 #(
		.INIT('h32)
	) name16227 (
		_w21819_,
		_w21990_,
		_w22053_,
		_w22054_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name16228 (
		_w21814_,
		_w22052_,
		_w22050_,
		_w22054_,
		_w22055_
	);
	LUT4 #(
		.INIT('hdaff)
	) name16229 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w22056_
	);
	LUT2 #(
		.INIT('h1)
	) name16230 (
		_w21815_,
		_w22056_,
		_w22057_
	);
	LUT4 #(
		.INIT('h1145)
	) name16231 (
		_w21815_,
		_w21817_,
		_w21818_,
		_w21816_,
		_w22058_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name16232 (
		_w21815_,
		_w21997_,
		_w22051_,
		_w22058_,
		_w22059_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name16233 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w22060_
	);
	LUT4 #(
		.INIT('h2322)
	) name16234 (
		_w21814_,
		_w22057_,
		_w22059_,
		_w22060_,
		_w22061_
	);
	LUT3 #(
		.INIT('h65)
	) name16235 (
		\u1_L3_reg[28]/NET0131 ,
		_w22055_,
		_w22061_,
		_w22062_
	);
	LUT4 #(
		.INIT('h00f7)
	) name16236 (
		_w21926_,
		_w21925_,
		_w21927_,
		_w21923_,
		_w22063_
	);
	LUT4 #(
		.INIT('h7f00)
	) name16237 (
		_w21926_,
		_w21925_,
		_w21927_,
		_w21923_,
		_w22064_
	);
	LUT4 #(
		.INIT('hefa8)
	) name16238 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22065_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name16239 (
		_w21951_,
		_w22063_,
		_w22064_,
		_w22065_,
		_w22066_
	);
	LUT4 #(
		.INIT('hd3ff)
	) name16240 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22067_
	);
	LUT3 #(
		.INIT('h8a)
	) name16241 (
		_w21943_,
		_w22066_,
		_w22067_,
		_w22068_
	);
	LUT3 #(
		.INIT('hb0)
	) name16242 (
		_w21926_,
		_w21925_,
		_w21923_,
		_w22069_
	);
	LUT4 #(
		.INIT('h5022)
	) name16243 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22070_
	);
	LUT3 #(
		.INIT('hb0)
	) name16244 (
		_w21925_,
		_w21927_,
		_w21923_,
		_w22071_
	);
	LUT4 #(
		.INIT('h3301)
	) name16245 (
		_w21926_,
		_w21924_,
		_w21927_,
		_w21923_,
		_w22072_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16246 (
		_w22069_,
		_w22070_,
		_w22071_,
		_w22072_,
		_w22073_
	);
	LUT4 #(
		.INIT('hdfeb)
	) name16247 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22074_
	);
	LUT4 #(
		.INIT('h0008)
	) name16248 (
		_w21926_,
		_w21924_,
		_w21927_,
		_w21923_,
		_w22075_
	);
	LUT4 #(
		.INIT('h0031)
	) name16249 (
		_w21923_,
		_w21946_,
		_w22074_,
		_w22075_,
		_w22076_
	);
	LUT3 #(
		.INIT('he0)
	) name16250 (
		_w21943_,
		_w22073_,
		_w22076_,
		_w22077_
	);
	LUT3 #(
		.INIT('h65)
	) name16251 (
		\u1_L3_reg[25]/NET0131 ,
		_w22068_,
		_w22077_,
		_w22078_
	);
	LUT4 #(
		.INIT('hff76)
	) name16252 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22079_
	);
	LUT3 #(
		.INIT('h02)
	) name16253 (
		_w21926_,
		_w21924_,
		_w21923_,
		_w22080_
	);
	LUT4 #(
		.INIT('h00c4)
	) name16254 (
		_w21923_,
		_w21929_,
		_w22079_,
		_w22080_,
		_w22081_
	);
	LUT2 #(
		.INIT('h2)
	) name16255 (
		_w21943_,
		_w22081_,
		_w22082_
	);
	LUT4 #(
		.INIT('h4404)
	) name16256 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22083_
	);
	LUT4 #(
		.INIT('haf23)
	) name16257 (
		_w21947_,
		_w22063_,
		_w22064_,
		_w22083_,
		_w22084_
	);
	LUT4 #(
		.INIT('hdaef)
	) name16258 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22085_
	);
	LUT4 #(
		.INIT('hcbbf)
	) name16259 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22086_
	);
	LUT3 #(
		.INIT('hb1)
	) name16260 (
		_w21923_,
		_w21942_,
		_w22086_,
		_w22087_
	);
	LUT4 #(
		.INIT('hba00)
	) name16261 (
		_w21943_,
		_w22084_,
		_w22085_,
		_w22087_,
		_w22088_
	);
	LUT3 #(
		.INIT('h65)
	) name16262 (
		\u1_L3_reg[8]/NET0131 ,
		_w22082_,
		_w22088_,
		_w22089_
	);
	LUT4 #(
		.INIT('hc3ee)
	) name16263 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w22090_
	);
	LUT2 #(
		.INIT('h1)
	) name16264 (
		_w21866_,
		_w22090_,
		_w22091_
	);
	LUT4 #(
		.INIT('h3233)
	) name16265 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w22092_
	);
	LUT3 #(
		.INIT('h2a)
	) name16266 (
		_w21862_,
		_w21860_,
		_w21859_,
		_w22093_
	);
	LUT4 #(
		.INIT('hd500)
	) name16267 (
		_w21862_,
		_w21860_,
		_w21859_,
		_w21866_,
		_w22094_
	);
	LUT4 #(
		.INIT('hdfa7)
	) name16268 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w22095_
	);
	LUT3 #(
		.INIT('hb0)
	) name16269 (
		_w22092_,
		_w22094_,
		_w22095_,
		_w22096_
	);
	LUT3 #(
		.INIT('h8a)
	) name16270 (
		_w21870_,
		_w22091_,
		_w22096_,
		_w22097_
	);
	LUT4 #(
		.INIT('hf9bf)
	) name16271 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w22098_
	);
	LUT2 #(
		.INIT('h1)
	) name16272 (
		_w21866_,
		_w22098_,
		_w22099_
	);
	LUT4 #(
		.INIT('ha2f0)
	) name16273 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w22100_
	);
	LUT4 #(
		.INIT('hef00)
	) name16274 (
		_w21861_,
		_w21860_,
		_w21859_,
		_w21866_,
		_w22101_
	);
	LUT4 #(
		.INIT('h4544)
	) name16275 (
		_w21870_,
		_w21886_,
		_w22100_,
		_w22101_,
		_w22102_
	);
	LUT4 #(
		.INIT('h0200)
	) name16276 (
		_w21861_,
		_w21860_,
		_w21859_,
		_w21866_,
		_w22103_
	);
	LUT4 #(
		.INIT('h0010)
	) name16277 (
		_w21862_,
		_w21860_,
		_w21859_,
		_w21866_,
		_w22104_
	);
	LUT2 #(
		.INIT('h8)
	) name16278 (
		_w21862_,
		_w21860_,
		_w22105_
	);
	LUT4 #(
		.INIT('h0080)
	) name16279 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21866_,
		_w22106_
	);
	LUT4 #(
		.INIT('h2223)
	) name16280 (
		_w21870_,
		_w22103_,
		_w22104_,
		_w22106_,
		_w22107_
	);
	LUT3 #(
		.INIT('h10)
	) name16281 (
		_w22102_,
		_w22099_,
		_w22107_,
		_w22108_
	);
	LUT3 #(
		.INIT('h65)
	) name16282 (
		\u1_L3_reg[27]/NET0131 ,
		_w22097_,
		_w22108_,
		_w22109_
	);
	LUT2 #(
		.INIT('h9)
	) name16283 (
		_w21733_,
		_w21735_,
		_w22110_
	);
	LUT4 #(
		.INIT('hd003)
	) name16284 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w22111_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name16285 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w22112_
	);
	LUT3 #(
		.INIT('h01)
	) name16286 (
		_w21736_,
		_w22112_,
		_w22111_,
		_w22113_
	);
	LUT4 #(
		.INIT('h0800)
	) name16287 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w22114_
	);
	LUT4 #(
		.INIT('hb5bc)
	) name16288 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w22115_
	);
	LUT3 #(
		.INIT('h31)
	) name16289 (
		_w21736_,
		_w22114_,
		_w22115_,
		_w22116_
	);
	LUT3 #(
		.INIT('h8a)
	) name16290 (
		_w21730_,
		_w22113_,
		_w22116_,
		_w22117_
	);
	LUT3 #(
		.INIT('h40)
	) name16291 (
		_w21732_,
		_w21733_,
		_w21735_,
		_w22118_
	);
	LUT4 #(
		.INIT('hab89)
	) name16292 (
		_w21736_,
		_w21910_,
		_w21912_,
		_w22118_,
		_w22119_
	);
	LUT4 #(
		.INIT('h7bd7)
	) name16293 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w22120_
	);
	LUT4 #(
		.INIT('h00c8)
	) name16294 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21736_,
		_w22121_
	);
	LUT4 #(
		.INIT('h135f)
	) name16295 (
		_w21736_,
		_w21751_,
		_w21743_,
		_w22121_,
		_w22122_
	);
	LUT4 #(
		.INIT('hba00)
	) name16296 (
		_w21730_,
		_w22119_,
		_w22120_,
		_w22122_,
		_w22123_
	);
	LUT3 #(
		.INIT('h65)
	) name16297 (
		\u1_L3_reg[32]/NET0131 ,
		_w22117_,
		_w22123_,
		_w22124_
	);
	LUT3 #(
		.INIT('h2e)
	) name16298 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w22125_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name16299 (
		_w21930_,
		_w21936_,
		_w22063_,
		_w22125_,
		_w22126_
	);
	LUT4 #(
		.INIT('h00d0)
	) name16300 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22127_
	);
	LUT2 #(
		.INIT('h1)
	) name16301 (
		_w21943_,
		_w22127_,
		_w22128_
	);
	LUT4 #(
		.INIT('he6f7)
	) name16302 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21927_,
		_w22129_
	);
	LUT2 #(
		.INIT('h2)
	) name16303 (
		_w21923_,
		_w22129_,
		_w22130_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name16304 (
		_w21926_,
		_w21925_,
		_w21924_,
		_w21923_,
		_w22131_
	);
	LUT4 #(
		.INIT('h3010)
	) name16305 (
		_w21927_,
		_w21942_,
		_w21943_,
		_w22131_,
		_w22132_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16306 (
		_w22126_,
		_w22128_,
		_w22130_,
		_w22132_,
		_w22133_
	);
	LUT4 #(
		.INIT('h0001)
	) name16307 (
		_w21923_,
		_w21931_,
		_w21934_,
		_w21955_,
		_w22134_
	);
	LUT3 #(
		.INIT('h02)
	) name16308 (
		_w21923_,
		_w21928_,
		_w21947_,
		_w22135_
	);
	LUT2 #(
		.INIT('h1)
	) name16309 (
		_w22134_,
		_w22135_,
		_w22136_
	);
	LUT3 #(
		.INIT('h56)
	) name16310 (
		\u1_L3_reg[3]/NET0131 ,
		_w22133_,
		_w22136_,
		_w22137_
	);
	LUT4 #(
		.INIT('hf126)
	) name16311 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w22138_
	);
	LUT4 #(
		.INIT('h2880)
	) name16312 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w22139_
	);
	LUT4 #(
		.INIT('h5004)
	) name16313 (
		_w21731_,
		_w21732_,
		_w21733_,
		_w21735_,
		_w22140_
	);
	LUT4 #(
		.INIT('h1302)
	) name16314 (
		_w21736_,
		_w22139_,
		_w22140_,
		_w22138_,
		_w22141_
	);
	LUT2 #(
		.INIT('h2)
	) name16315 (
		_w21730_,
		_w22141_,
		_w22142_
	);
	LUT2 #(
		.INIT('h4)
	) name16316 (
		_w21736_,
		_w22139_,
		_w22143_
	);
	LUT2 #(
		.INIT('h2)
	) name16317 (
		_w21730_,
		_w21736_,
		_w22144_
	);
	LUT3 #(
		.INIT('h4c)
	) name16318 (
		_w21732_,
		_w21733_,
		_w21735_,
		_w22145_
	);
	LUT4 #(
		.INIT('h8a00)
	) name16319 (
		_w21731_,
		_w21733_,
		_w21735_,
		_w21736_,
		_w22146_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name16320 (
		_w21737_,
		_w22110_,
		_w22145_,
		_w22146_,
		_w22147_
	);
	LUT3 #(
		.INIT('h45)
	) name16321 (
		_w21750_,
		_w21736_,
		_w22140_,
		_w22148_
	);
	LUT4 #(
		.INIT('h0133)
	) name16322 (
		_w21730_,
		_w22144_,
		_w22147_,
		_w22148_,
		_w22149_
	);
	LUT4 #(
		.INIT('h5556)
	) name16323 (
		\u1_L3_reg[7]/NET0131 ,
		_w22143_,
		_w22149_,
		_w22142_,
		_w22150_
	);
	LUT4 #(
		.INIT('hc693)
	) name16324 (
		decrypt_pad,
		\u1_R3_reg[11]/NET0131 ,
		\u1_uk_K_r3_reg[26]/NET0131 ,
		\u1_uk_K_r3_reg[3]/NET0131 ,
		_w22151_
	);
	LUT4 #(
		.INIT('hc963)
	) name16325 (
		decrypt_pad,
		\u1_R3_reg[12]/NET0131 ,
		\u1_uk_K_r3_reg[18]/NET0131 ,
		\u1_uk_K_r3_reg[41]/NET0131 ,
		_w22152_
	);
	LUT4 #(
		.INIT('hc693)
	) name16326 (
		decrypt_pad,
		\u1_R3_reg[13]/NET0131 ,
		\u1_uk_K_r3_reg[54]/NET0131 ,
		\u1_uk_K_r3_reg[6]/NET0131 ,
		_w22153_
	);
	LUT4 #(
		.INIT('hc693)
	) name16327 (
		decrypt_pad,
		\u1_R3_reg[9]/NET0131 ,
		\u1_uk_K_r3_reg[17]/NET0131 ,
		\u1_uk_K_r3_reg[26]/NET0131 ,
		_w22154_
	);
	LUT4 #(
		.INIT('hc693)
	) name16328 (
		decrypt_pad,
		\u1_R3_reg[10]/NET0131 ,
		\u1_uk_K_r3_reg[25]/NET0131 ,
		\u1_uk_K_r3_reg[34]/NET0131 ,
		_w22155_
	);
	LUT4 #(
		.INIT('hc693)
	) name16329 (
		decrypt_pad,
		\u1_R3_reg[8]/NET0131 ,
		\u1_uk_K_r3_reg[20]/NET0131 ,
		\u1_uk_K_r3_reg[54]/NET0131 ,
		_w22156_
	);
	LUT2 #(
		.INIT('h2)
	) name16330 (
		_w22153_,
		_w22156_,
		_w22157_
	);
	LUT4 #(
		.INIT('h995d)
	) name16331 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22158_
	);
	LUT4 #(
		.INIT('h0001)
	) name16332 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22159_
	);
	LUT4 #(
		.INIT('hdfde)
	) name16333 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22160_
	);
	LUT4 #(
		.INIT('h08cc)
	) name16334 (
		_w22152_,
		_w22151_,
		_w22158_,
		_w22160_,
		_w22161_
	);
	LUT3 #(
		.INIT('h0b)
	) name16335 (
		_w22153_,
		_w22154_,
		_w22151_,
		_w22162_
	);
	LUT4 #(
		.INIT('h22f3)
	) name16336 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22163_
	);
	LUT4 #(
		.INIT('h0040)
	) name16337 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22164_
	);
	LUT4 #(
		.INIT('haa08)
	) name16338 (
		_w22152_,
		_w22162_,
		_w22163_,
		_w22164_,
		_w22165_
	);
	LUT2 #(
		.INIT('h1)
	) name16339 (
		_w22154_,
		_w22155_,
		_w22166_
	);
	LUT2 #(
		.INIT('h6)
	) name16340 (
		_w22154_,
		_w22155_,
		_w22167_
	);
	LUT2 #(
		.INIT('h8)
	) name16341 (
		_w22153_,
		_w22156_,
		_w22168_
	);
	LUT3 #(
		.INIT('h52)
	) name16342 (
		_w22153_,
		_w22151_,
		_w22156_,
		_w22169_
	);
	LUT2 #(
		.INIT('h1)
	) name16343 (
		_w22167_,
		_w22169_,
		_w22170_
	);
	LUT3 #(
		.INIT('h02)
	) name16344 (
		_w22151_,
		_w22155_,
		_w22156_,
		_w22171_
	);
	LUT4 #(
		.INIT('h1428)
	) name16345 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22172_
	);
	LUT3 #(
		.INIT('h45)
	) name16346 (
		_w22152_,
		_w22171_,
		_w22172_,
		_w22173_
	);
	LUT4 #(
		.INIT('h0045)
	) name16347 (
		_w22165_,
		_w22170_,
		_w22173_,
		_w22161_,
		_w22174_
	);
	LUT2 #(
		.INIT('h9)
	) name16348 (
		\u1_L3_reg[6]/NET0131 ,
		_w22174_,
		_w22175_
	);
	LUT4 #(
		.INIT('h9060)
	) name16349 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w22176_
	);
	LUT3 #(
		.INIT('h43)
	) name16350 (
		_w5828_,
		_w5827_,
		_w5829_,
		_w22177_
	);
	LUT4 #(
		.INIT('h0015)
	) name16351 (
		_w5850_,
		_w21676_,
		_w22177_,
		_w22176_,
		_w22178_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name16352 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w22179_
	);
	LUT2 #(
		.INIT('h1)
	) name16353 (
		_w5834_,
		_w22179_,
		_w22180_
	);
	LUT4 #(
		.INIT('hcc3b)
	) name16354 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w22181_
	);
	LUT4 #(
		.INIT('hd7ef)
	) name16355 (
		_w5828_,
		_w5827_,
		_w5832_,
		_w5829_,
		_w22182_
	);
	LUT4 #(
		.INIT('h8d00)
	) name16356 (
		_w5834_,
		_w22181_,
		_w22177_,
		_w22182_,
		_w22183_
	);
	LUT4 #(
		.INIT('h3210)
	) name16357 (
		_w5840_,
		_w22180_,
		_w22183_,
		_w22178_,
		_w22184_
	);
	LUT2 #(
		.INIT('h9)
	) name16358 (
		\u1_L3_reg[9]/NET0131 ,
		_w22184_,
		_w22185_
	);
	LUT3 #(
		.INIT('h80)
	) name16359 (
		_w22153_,
		_w22154_,
		_w22156_,
		_w22186_
	);
	LUT2 #(
		.INIT('h4)
	) name16360 (
		_w22153_,
		_w22156_,
		_w22187_
	);
	LUT4 #(
		.INIT('h669d)
	) name16361 (
		_w22153_,
		_w22154_,
		_w22151_,
		_w22156_,
		_w22188_
	);
	LUT2 #(
		.INIT('h1)
	) name16362 (
		_w22155_,
		_w22188_,
		_w22189_
	);
	LUT4 #(
		.INIT('h0110)
	) name16363 (
		_w22153_,
		_w22151_,
		_w22155_,
		_w22156_,
		_w22190_
	);
	LUT4 #(
		.INIT('h0080)
	) name16364 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22191_
	);
	LUT3 #(
		.INIT('h02)
	) name16365 (
		_w22152_,
		_w22191_,
		_w22190_,
		_w22192_
	);
	LUT4 #(
		.INIT('h77d8)
	) name16366 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22193_
	);
	LUT2 #(
		.INIT('h1)
	) name16367 (
		_w22151_,
		_w22193_,
		_w22194_
	);
	LUT4 #(
		.INIT('h6080)
	) name16368 (
		_w22153_,
		_w22154_,
		_w22151_,
		_w22156_,
		_w22195_
	);
	LUT3 #(
		.INIT('h01)
	) name16369 (
		_w22152_,
		_w22159_,
		_w22195_,
		_w22196_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16370 (
		_w22189_,
		_w22192_,
		_w22194_,
		_w22196_,
		_w22197_
	);
	LUT4 #(
		.INIT('hb0e0)
	) name16371 (
		_w22153_,
		_w22154_,
		_w22151_,
		_w22156_,
		_w22198_
	);
	LUT2 #(
		.INIT('h8)
	) name16372 (
		_w22155_,
		_w22156_,
		_w22199_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name16373 (
		_w22154_,
		_w22151_,
		_w22155_,
		_w22156_,
		_w22200_
	);
	LUT2 #(
		.INIT('h4)
	) name16374 (
		_w22198_,
		_w22200_,
		_w22201_
	);
	LUT3 #(
		.INIT('h56)
	) name16375 (
		\u1_L3_reg[16]/NET0131 ,
		_w22197_,
		_w22201_,
		_w22202_
	);
	LUT4 #(
		.INIT('hfd75)
	) name16376 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w22203_
	);
	LUT2 #(
		.INIT('h1)
	) name16377 (
		_w21815_,
		_w22203_,
		_w22204_
	);
	LUT4 #(
		.INIT('h0a20)
	) name16378 (
		_w21815_,
		_w21817_,
		_w21818_,
		_w21816_,
		_w22205_
	);
	LUT3 #(
		.INIT('h02)
	) name16379 (
		_w21814_,
		_w21834_,
		_w22205_,
		_w22206_
	);
	LUT2 #(
		.INIT('h4)
	) name16380 (
		_w22204_,
		_w22206_,
		_w22207_
	);
	LUT4 #(
		.INIT('h1003)
	) name16381 (
		_w21815_,
		_w21817_,
		_w21816_,
		_w21819_,
		_w22208_
	);
	LUT3 #(
		.INIT('h01)
	) name16382 (
		_w21814_,
		_w21994_,
		_w21978_,
		_w22209_
	);
	LUT4 #(
		.INIT('h8000)
	) name16383 (
		_w21815_,
		_w21817_,
		_w21818_,
		_w21816_,
		_w22210_
	);
	LUT2 #(
		.INIT('h1)
	) name16384 (
		_w21823_,
		_w22210_,
		_w22211_
	);
	LUT3 #(
		.INIT('h40)
	) name16385 (
		_w22208_,
		_w22209_,
		_w22211_,
		_w22212_
	);
	LUT4 #(
		.INIT('h1000)
	) name16386 (
		_w21815_,
		_w21817_,
		_w21818_,
		_w21816_,
		_w22213_
	);
	LUT4 #(
		.INIT('h77ef)
	) name16387 (
		_w21817_,
		_w21818_,
		_w21816_,
		_w21819_,
		_w22214_
	);
	LUT3 #(
		.INIT('h31)
	) name16388 (
		_w21815_,
		_w22213_,
		_w22214_,
		_w22215_
	);
	LUT4 #(
		.INIT('ha955)
	) name16389 (
		\u1_L3_reg[18]/NET0131 ,
		_w22207_,
		_w22212_,
		_w22215_,
		_w22216_
	);
	LUT3 #(
		.INIT('hf9)
	) name16390 (
		_w22153_,
		_w22155_,
		_w22156_,
		_w22217_
	);
	LUT3 #(
		.INIT('h04)
	) name16391 (
		_w22153_,
		_w22154_,
		_w22156_,
		_w22218_
	);
	LUT4 #(
		.INIT('hcfa1)
	) name16392 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22219_
	);
	LUT4 #(
		.INIT('h1000)
	) name16393 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22220_
	);
	LUT4 #(
		.INIT('h5504)
	) name16394 (
		_w22152_,
		_w22151_,
		_w22219_,
		_w22220_,
		_w22221_
	);
	LUT3 #(
		.INIT('h32)
	) name16395 (
		_w22154_,
		_w22151_,
		_w22155_,
		_w22222_
	);
	LUT3 #(
		.INIT('h04)
	) name16396 (
		_w22154_,
		_w22151_,
		_w22155_,
		_w22223_
	);
	LUT4 #(
		.INIT('h5510)
	) name16397 (
		_w22157_,
		_w22187_,
		_w22222_,
		_w22223_,
		_w22224_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name16398 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22225_
	);
	LUT4 #(
		.INIT('h3f15)
	) name16399 (
		_w22151_,
		_w22166_,
		_w22169_,
		_w22225_,
		_w22226_
	);
	LUT3 #(
		.INIT('h8a)
	) name16400 (
		_w22152_,
		_w22224_,
		_w22226_,
		_w22227_
	);
	LUT4 #(
		.INIT('hb95e)
	) name16401 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22228_
	);
	LUT2 #(
		.INIT('h1)
	) name16402 (
		_w22152_,
		_w22151_,
		_w22229_
	);
	LUT2 #(
		.INIT('h4)
	) name16403 (
		_w22228_,
		_w22229_,
		_w22230_
	);
	LUT3 #(
		.INIT('he7)
	) name16404 (
		_w22153_,
		_w22154_,
		_w22156_,
		_w22231_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name16405 (
		_w22151_,
		_w22155_,
		_w22186_,
		_w22231_,
		_w22232_
	);
	LUT2 #(
		.INIT('h4)
	) name16406 (
		_w22230_,
		_w22232_,
		_w22233_
	);
	LUT4 #(
		.INIT('h5655)
	) name16407 (
		\u1_L3_reg[24]/NET0131 ,
		_w22227_,
		_w22221_,
		_w22233_,
		_w22234_
	);
	LUT3 #(
		.INIT('h15)
	) name16408 (
		_w22151_,
		_w22155_,
		_w22156_,
		_w22235_
	);
	LUT2 #(
		.INIT('h4)
	) name16409 (
		_w22218_,
		_w22235_,
		_w22236_
	);
	LUT4 #(
		.INIT('h0100)
	) name16410 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22237_
	);
	LUT3 #(
		.INIT('h08)
	) name16411 (
		_w22151_,
		_w22217_,
		_w22237_,
		_w22238_
	);
	LUT3 #(
		.INIT('ha8)
	) name16412 (
		_w22152_,
		_w22236_,
		_w22238_,
		_w22239_
	);
	LUT4 #(
		.INIT('hf052)
	) name16413 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22240_
	);
	LUT4 #(
		.INIT('hd4c4)
	) name16414 (
		_w22153_,
		_w22154_,
		_w22151_,
		_w22156_,
		_w22241_
	);
	LUT2 #(
		.INIT('h1)
	) name16415 (
		_w22240_,
		_w22241_,
		_w22242_
	);
	LUT4 #(
		.INIT('h4bfb)
	) name16416 (
		_w22153_,
		_w22154_,
		_w22155_,
		_w22156_,
		_w22243_
	);
	LUT3 #(
		.INIT('h51)
	) name16417 (
		_w22152_,
		_w22151_,
		_w22243_,
		_w22244_
	);
	LUT2 #(
		.INIT('h4)
	) name16418 (
		_w22242_,
		_w22244_,
		_w22245_
	);
	LUT3 #(
		.INIT('h20)
	) name16419 (
		_w22153_,
		_w22154_,
		_w22151_,
		_w22246_
	);
	LUT2 #(
		.INIT('h8)
	) name16420 (
		_w22199_,
		_w22246_,
		_w22247_
	);
	LUT4 #(
		.INIT('h0400)
	) name16421 (
		_w22153_,
		_w22154_,
		_w22151_,
		_w22155_,
		_w22248_
	);
	LUT3 #(
		.INIT('h80)
	) name16422 (
		_w22152_,
		_w22154_,
		_w22155_,
		_w22249_
	);
	LUT3 #(
		.INIT('h23)
	) name16423 (
		_w22168_,
		_w22248_,
		_w22249_,
		_w22250_
	);
	LUT2 #(
		.INIT('h4)
	) name16424 (
		_w22247_,
		_w22250_,
		_w22251_
	);
	LUT4 #(
		.INIT('h56aa)
	) name16425 (
		\u1_L3_reg[30]/NET0131 ,
		_w22239_,
		_w22245_,
		_w22251_,
		_w22252_
	);
	LUT4 #(
		.INIT('hc963)
	) name16426 (
		decrypt_pad,
		\u1_R2_reg[28]/NET0131 ,
		\u1_uk_K_r2_reg[0]/NET0131 ,
		\u1_uk_K_r2_reg[22]/NET0131 ,
		_w22253_
	);
	LUT4 #(
		.INIT('hc693)
	) name16427 (
		decrypt_pad,
		\u1_R2_reg[26]/NET0131 ,
		\u1_uk_K_r2_reg[2]/NET0131 ,
		\u1_uk_K_r2_reg[35]/NET0131 ,
		_w22254_
	);
	LUT4 #(
		.INIT('hc693)
	) name16428 (
		decrypt_pad,
		\u1_R2_reg[25]/NET0131 ,
		\u1_uk_K_r2_reg[45]/NET0131 ,
		\u1_uk_K_r2_reg[50]/NET0131 ,
		_w22255_
	);
	LUT4 #(
		.INIT('hc693)
	) name16429 (
		decrypt_pad,
		\u1_R2_reg[29]/NET0131 ,
		\u1_uk_K_r2_reg[14]/NET0131 ,
		\u1_uk_K_r2_reg[23]/NET0131 ,
		_w22256_
	);
	LUT3 #(
		.INIT('hea)
	) name16430 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22257_
	);
	LUT4 #(
		.INIT('hc963)
	) name16431 (
		decrypt_pad,
		\u1_R2_reg[24]/NET0131 ,
		\u1_uk_K_r2_reg[15]/NET0131 ,
		\u1_uk_K_r2_reg[37]/NET0131 ,
		_w22258_
	);
	LUT4 #(
		.INIT('hc693)
	) name16432 (
		decrypt_pad,
		\u1_R2_reg[27]/NET0131 ,
		\u1_uk_K_r2_reg[35]/NET0131 ,
		\u1_uk_K_r2_reg[44]/NET0131 ,
		_w22259_
	);
	LUT3 #(
		.INIT('h70)
	) name16433 (
		_w22254_,
		_w22255_,
		_w22259_,
		_w22260_
	);
	LUT4 #(
		.INIT('h7000)
	) name16434 (
		_w22254_,
		_w22255_,
		_w22258_,
		_w22259_,
		_w22261_
	);
	LUT2 #(
		.INIT('h8)
	) name16435 (
		_w22257_,
		_w22261_,
		_w22262_
	);
	LUT4 #(
		.INIT('h1000)
	) name16436 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22263_
	);
	LUT4 #(
		.INIT('hef3f)
	) name16437 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22264_
	);
	LUT2 #(
		.INIT('h2)
	) name16438 (
		_w22256_,
		_w22258_,
		_w22265_
	);
	LUT4 #(
		.INIT('h0020)
	) name16439 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22266_
	);
	LUT4 #(
		.INIT('hffde)
	) name16440 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22267_
	);
	LUT3 #(
		.INIT('he0)
	) name16441 (
		_w22259_,
		_w22264_,
		_w22267_,
		_w22268_
	);
	LUT3 #(
		.INIT('h8a)
	) name16442 (
		_w22253_,
		_w22262_,
		_w22268_,
		_w22269_
	);
	LUT4 #(
		.INIT('h0072)
	) name16443 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22259_,
		_w22270_
	);
	LUT4 #(
		.INIT('h10f0)
	) name16444 (
		_w22254_,
		_w22255_,
		_w22258_,
		_w22259_,
		_w22271_
	);
	LUT2 #(
		.INIT('h4)
	) name16445 (
		_w22270_,
		_w22271_,
		_w22272_
	);
	LUT4 #(
		.INIT('h0002)
	) name16446 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22273_
	);
	LUT2 #(
		.INIT('h6)
	) name16447 (
		_w22254_,
		_w22258_,
		_w22274_
	);
	LUT3 #(
		.INIT('h8c)
	) name16448 (
		_w22255_,
		_w22256_,
		_w22259_,
		_w22275_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name16449 (
		_w22273_,
		_w22259_,
		_w22274_,
		_w22275_,
		_w22276_
	);
	LUT4 #(
		.INIT('h0008)
	) name16450 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22277_
	);
	LUT4 #(
		.INIT('hfcd7)
	) name16451 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22278_
	);
	LUT4 #(
		.INIT('h0084)
	) name16452 (
		_w22254_,
		_w22255_,
		_w22258_,
		_w22259_,
		_w22279_
	);
	LUT4 #(
		.INIT('h0100)
	) name16453 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22259_,
		_w22280_
	);
	LUT4 #(
		.INIT('h0031)
	) name16454 (
		_w22259_,
		_w22279_,
		_w22278_,
		_w22280_,
		_w22281_
	);
	LUT4 #(
		.INIT('hba00)
	) name16455 (
		_w22253_,
		_w22272_,
		_w22276_,
		_w22281_,
		_w22282_
	);
	LUT3 #(
		.INIT('h65)
	) name16456 (
		\u1_L2_reg[22]/NET0131 ,
		_w22269_,
		_w22282_,
		_w22283_
	);
	LUT4 #(
		.INIT('hc693)
	) name16457 (
		decrypt_pad,
		\u1_R2_reg[4]/NET0131 ,
		\u1_uk_K_r2_reg[48]/NET0131 ,
		\u1_uk_K_r2_reg[53]/P0001 ,
		_w22284_
	);
	LUT4 #(
		.INIT('hc693)
	) name16458 (
		decrypt_pad,
		\u1_R2_reg[32]/NET0131 ,
		\u1_uk_K_r2_reg[25]/NET0131 ,
		\u1_uk_K_r2_reg[5]/NET0131 ,
		_w22285_
	);
	LUT4 #(
		.INIT('hc963)
	) name16459 (
		decrypt_pad,
		\u1_R2_reg[1]/NET0131 ,
		\u1_uk_K_r2_reg[26]/NET0131 ,
		\u1_uk_K_r2_reg[46]/NET0131 ,
		_w22286_
	);
	LUT4 #(
		.INIT('hc963)
	) name16460 (
		decrypt_pad,
		\u1_R2_reg[2]/NET0131 ,
		\u1_uk_K_r2_reg[41]/NET0131 ,
		\u1_uk_K_r2_reg[4]/NET0131 ,
		_w22287_
	);
	LUT4 #(
		.INIT('hc693)
	) name16461 (
		decrypt_pad,
		\u1_R2_reg[5]/NET0131 ,
		\u1_uk_K_r2_reg[19]/NET0131 ,
		\u1_uk_K_r2_reg[24]/NET0131 ,
		_w22288_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name16462 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22289_
	);
	LUT2 #(
		.INIT('h1)
	) name16463 (
		_w22288_,
		_w22285_,
		_w22290_
	);
	LUT4 #(
		.INIT('hc693)
	) name16464 (
		decrypt_pad,
		\u1_R2_reg[3]/NET0131 ,
		\u1_uk_K_r2_reg[13]/NET0131 ,
		\u1_uk_K_r2_reg[18]/NET0131 ,
		_w22291_
	);
	LUT2 #(
		.INIT('h4)
	) name16465 (
		_w22287_,
		_w22291_,
		_w22292_
	);
	LUT3 #(
		.INIT('hb0)
	) name16466 (
		_w22287_,
		_w22291_,
		_w22286_,
		_w22293_
	);
	LUT3 #(
		.INIT('h01)
	) name16467 (
		_w22290_,
		_w22293_,
		_w22289_,
		_w22294_
	);
	LUT3 #(
		.INIT('h02)
	) name16468 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22295_
	);
	LUT4 #(
		.INIT('hfd31)
	) name16469 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22296_
	);
	LUT4 #(
		.INIT('h300a)
	) name16470 (
		_w22287_,
		_w22291_,
		_w22285_,
		_w22286_,
		_w22297_
	);
	LUT3 #(
		.INIT('h0d)
	) name16471 (
		_w22291_,
		_w22296_,
		_w22297_,
		_w22298_
	);
	LUT3 #(
		.INIT('h8a)
	) name16472 (
		_w22284_,
		_w22294_,
		_w22298_,
		_w22299_
	);
	LUT3 #(
		.INIT('he6)
	) name16473 (
		_w22287_,
		_w22285_,
		_w22286_,
		_w22300_
	);
	LUT3 #(
		.INIT('h51)
	) name16474 (
		_w22291_,
		_w22288_,
		_w22286_,
		_w22301_
	);
	LUT2 #(
		.INIT('h4)
	) name16475 (
		_w22300_,
		_w22301_,
		_w22302_
	);
	LUT2 #(
		.INIT('h8)
	) name16476 (
		_w22287_,
		_w22291_,
		_w22303_
	);
	LUT3 #(
		.INIT('h60)
	) name16477 (
		_w22288_,
		_w22285_,
		_w22286_,
		_w22304_
	);
	LUT4 #(
		.INIT('h7c3f)
	) name16478 (
		_w22291_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22305_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name16479 (
		_w22287_,
		_w22291_,
		_w22304_,
		_w22305_,
		_w22306_
	);
	LUT2 #(
		.INIT('h2)
	) name16480 (
		_w22291_,
		_w22286_,
		_w22307_
	);
	LUT3 #(
		.INIT('had)
	) name16481 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22308_
	);
	LUT4 #(
		.INIT('h8000)
	) name16482 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22309_
	);
	LUT4 #(
		.INIT('h0008)
	) name16483 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22310_
	);
	LUT4 #(
		.INIT('h6ef7)
	) name16484 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22311_
	);
	LUT4 #(
		.INIT('hfda8)
	) name16485 (
		_w22291_,
		_w22286_,
		_w22308_,
		_w22311_,
		_w22312_
	);
	LUT4 #(
		.INIT('hba00)
	) name16486 (
		_w22284_,
		_w22302_,
		_w22306_,
		_w22312_,
		_w22313_
	);
	LUT3 #(
		.INIT('h65)
	) name16487 (
		\u1_L2_reg[31]/NET0131 ,
		_w22299_,
		_w22313_,
		_w22314_
	);
	LUT4 #(
		.INIT('hc693)
	) name16488 (
		decrypt_pad,
		\u1_R2_reg[24]/NET0131 ,
		\u1_uk_K_r2_reg[15]/NET0131 ,
		\u1_uk_K_r2_reg[52]/NET0131 ,
		_w22315_
	);
	LUT4 #(
		.INIT('hc963)
	) name16489 (
		decrypt_pad,
		\u1_R2_reg[23]/NET0131 ,
		\u1_uk_K_r2_reg[22]/NET0131 ,
		\u1_uk_K_r2_reg[44]/NET0131 ,
		_w22316_
	);
	LUT4 #(
		.INIT('hc963)
	) name16490 (
		decrypt_pad,
		\u1_R2_reg[21]/NET0131 ,
		\u1_uk_K_r2_reg[42]/NET0131 ,
		\u1_uk_K_r2_reg[9]/NET0131 ,
		_w22317_
	);
	LUT4 #(
		.INIT('hc963)
	) name16491 (
		decrypt_pad,
		\u1_R2_reg[20]/NET0131 ,
		\u1_uk_K_r2_reg[31]/NET0131 ,
		\u1_uk_K_r2_reg[49]/NET0131 ,
		_w22318_
	);
	LUT4 #(
		.INIT('hc693)
	) name16492 (
		decrypt_pad,
		\u1_R2_reg[22]/NET0131 ,
		\u1_uk_K_r2_reg[0]/NET0131 ,
		\u1_uk_K_r2_reg[9]/NET0131 ,
		_w22319_
	);
	LUT4 #(
		.INIT('hc693)
	) name16493 (
		decrypt_pad,
		\u1_R2_reg[25]/NET0131 ,
		\u1_uk_K_r2_reg[38]/NET0131 ,
		\u1_uk_K_r2_reg[43]/NET0131 ,
		_w22320_
	);
	LUT3 #(
		.INIT('hc4)
	) name16494 (
		_w22317_,
		_w22318_,
		_w22320_,
		_w22321_
	);
	LUT4 #(
		.INIT('h57db)
	) name16495 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22322_
	);
	LUT2 #(
		.INIT('h2)
	) name16496 (
		_w22316_,
		_w22322_,
		_w22323_
	);
	LUT4 #(
		.INIT('he020)
	) name16497 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22324_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name16498 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22325_
	);
	LUT3 #(
		.INIT('h01)
	) name16499 (
		_w22316_,
		_w22325_,
		_w22324_,
		_w22326_
	);
	LUT2 #(
		.INIT('h1)
	) name16500 (
		_w22319_,
		_w22316_,
		_w22327_
	);
	LUT4 #(
		.INIT('h0200)
	) name16501 (
		_w22318_,
		_w22319_,
		_w22316_,
		_w22320_,
		_w22328_
	);
	LUT2 #(
		.INIT('h4)
	) name16502 (
		_w22317_,
		_w22328_,
		_w22329_
	);
	LUT4 #(
		.INIT('haaa8)
	) name16503 (
		_w22315_,
		_w22326_,
		_w22323_,
		_w22329_,
		_w22330_
	);
	LUT4 #(
		.INIT('h0028)
	) name16504 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22316_,
		_w22331_
	);
	LUT4 #(
		.INIT('h1000)
	) name16505 (
		_w22317_,
		_w22318_,
		_w22316_,
		_w22320_,
		_w22332_
	);
	LUT4 #(
		.INIT('h0008)
	) name16506 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22333_
	);
	LUT3 #(
		.INIT('h10)
	) name16507 (
		_w22318_,
		_w22319_,
		_w22316_,
		_w22334_
	);
	LUT3 #(
		.INIT('h01)
	) name16508 (
		_w22333_,
		_w22334_,
		_w22332_,
		_w22335_
	);
	LUT4 #(
		.INIT('haf8c)
	) name16509 (
		_w22317_,
		_w22319_,
		_w22316_,
		_w22320_,
		_w22336_
	);
	LUT3 #(
		.INIT('h8a)
	) name16510 (
		_w22318_,
		_w22319_,
		_w22316_,
		_w22337_
	);
	LUT4 #(
		.INIT('h4000)
	) name16511 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22338_
	);
	LUT3 #(
		.INIT('h0b)
	) name16512 (
		_w22336_,
		_w22337_,
		_w22338_,
		_w22339_
	);
	LUT4 #(
		.INIT('h00bf)
	) name16513 (
		_w22331_,
		_w22335_,
		_w22339_,
		_w22315_,
		_w22340_
	);
	LUT4 #(
		.INIT('heff7)
	) name16514 (
		_w22317_,
		_w22318_,
		_w22316_,
		_w22320_,
		_w22341_
	);
	LUT2 #(
		.INIT('h1)
	) name16515 (
		_w22319_,
		_w22341_,
		_w22342_
	);
	LUT4 #(
		.INIT('h0002)
	) name16516 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22343_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name16517 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22344_
	);
	LUT4 #(
		.INIT('h0001)
	) name16518 (
		_w22318_,
		_w22319_,
		_w22316_,
		_w22320_,
		_w22345_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name16519 (
		_w22317_,
		_w22316_,
		_w22344_,
		_w22345_,
		_w22346_
	);
	LUT2 #(
		.INIT('h4)
	) name16520 (
		_w22342_,
		_w22346_,
		_w22347_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name16521 (
		\u1_L2_reg[11]/NET0131 ,
		_w22340_,
		_w22330_,
		_w22347_,
		_w22348_
	);
	LUT4 #(
		.INIT('hc963)
	) name16522 (
		decrypt_pad,
		\u1_R2_reg[13]/NET0131 ,
		\u1_uk_K_r2_reg[13]/NET0131 ,
		\u1_uk_K_r2_reg[33]/NET0131 ,
		_w22349_
	);
	LUT4 #(
		.INIT('hc963)
	) name16523 (
		decrypt_pad,
		\u1_R2_reg[12]/NET0131 ,
		\u1_uk_K_r2_reg[19]/NET0131 ,
		\u1_uk_K_r2_reg[39]/NET0131 ,
		_w22350_
	);
	LUT4 #(
		.INIT('hc963)
	) name16524 (
		decrypt_pad,
		\u1_R2_reg[17]/NET0131 ,
		\u1_uk_K_r2_reg[3]/NET0131 ,
		\u1_uk_K_r2_reg[55]/NET0131 ,
		_w22351_
	);
	LUT4 #(
		.INIT('hc693)
	) name16525 (
		decrypt_pad,
		\u1_R2_reg[15]/NET0131 ,
		\u1_uk_K_r2_reg[10]/NET0131 ,
		\u1_uk_K_r2_reg[47]/NET0131 ,
		_w22352_
	);
	LUT4 #(
		.INIT('h2aa8)
	) name16526 (
		_w22352_,
		_w22350_,
		_w22349_,
		_w22351_,
		_w22353_
	);
	LUT4 #(
		.INIT('hc693)
	) name16527 (
		decrypt_pad,
		\u1_R2_reg[14]/NET0131 ,
		\u1_uk_K_r2_reg[34]/NET0131 ,
		\u1_uk_K_r2_reg[39]/NET0131 ,
		_w22354_
	);
	LUT3 #(
		.INIT('h08)
	) name16528 (
		_w22350_,
		_w22354_,
		_w22351_,
		_w22355_
	);
	LUT3 #(
		.INIT('h45)
	) name16529 (
		_w22352_,
		_w22349_,
		_w22351_,
		_w22356_
	);
	LUT3 #(
		.INIT('h45)
	) name16530 (
		_w22353_,
		_w22355_,
		_w22356_,
		_w22357_
	);
	LUT3 #(
		.INIT('h01)
	) name16531 (
		_w22350_,
		_w22354_,
		_w22351_,
		_w22358_
	);
	LUT4 #(
		.INIT('h0001)
	) name16532 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22359_
	);
	LUT3 #(
		.INIT('h04)
	) name16533 (
		_w22350_,
		_w22349_,
		_w22351_,
		_w22360_
	);
	LUT4 #(
		.INIT('hffbe)
	) name16534 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22361_
	);
	LUT4 #(
		.INIT('h0200)
	) name16535 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22362_
	);
	LUT4 #(
		.INIT('hc693)
	) name16536 (
		decrypt_pad,
		\u1_R2_reg[16]/NET0131 ,
		\u1_uk_K_r2_reg[18]/NET0131 ,
		\u1_uk_K_r2_reg[55]/NET0131 ,
		_w22363_
	);
	LUT3 #(
		.INIT('h80)
	) name16537 (
		_w22352_,
		_w22349_,
		_w22354_,
		_w22364_
	);
	LUT4 #(
		.INIT('h2000)
	) name16538 (
		_w22352_,
		_w22350_,
		_w22349_,
		_w22354_,
		_w22365_
	);
	LUT4 #(
		.INIT('h0002)
	) name16539 (
		_w22361_,
		_w22363_,
		_w22365_,
		_w22362_,
		_w22366_
	);
	LUT2 #(
		.INIT('h4)
	) name16540 (
		_w22357_,
		_w22366_,
		_w22367_
	);
	LUT4 #(
		.INIT('h0001)
	) name16541 (
		_w22352_,
		_w22350_,
		_w22349_,
		_w22351_,
		_w22368_
	);
	LUT4 #(
		.INIT('h3ffe)
	) name16542 (
		_w22352_,
		_w22350_,
		_w22349_,
		_w22351_,
		_w22369_
	);
	LUT2 #(
		.INIT('h2)
	) name16543 (
		_w22354_,
		_w22369_,
		_w22370_
	);
	LUT2 #(
		.INIT('h2)
	) name16544 (
		_w22350_,
		_w22349_,
		_w22371_
	);
	LUT4 #(
		.INIT('h0014)
	) name16545 (
		_w22352_,
		_w22350_,
		_w22349_,
		_w22354_,
		_w22372_
	);
	LUT2 #(
		.INIT('h2)
	) name16546 (
		_w22363_,
		_w22372_,
		_w22373_
	);
	LUT4 #(
		.INIT('h0400)
	) name16547 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22374_
	);
	LUT4 #(
		.INIT('h0080)
	) name16548 (
		_w22352_,
		_w22350_,
		_w22349_,
		_w22351_,
		_w22375_
	);
	LUT2 #(
		.INIT('h4)
	) name16549 (
		_w22350_,
		_w22351_,
		_w22376_
	);
	LUT4 #(
		.INIT('h0200)
	) name16550 (
		_w22352_,
		_w22350_,
		_w22349_,
		_w22351_,
		_w22377_
	);
	LUT3 #(
		.INIT('h01)
	) name16551 (
		_w22374_,
		_w22375_,
		_w22377_,
		_w22378_
	);
	LUT3 #(
		.INIT('h40)
	) name16552 (
		_w22370_,
		_w22373_,
		_w22378_,
		_w22379_
	);
	LUT4 #(
		.INIT('h0020)
	) name16553 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22380_
	);
	LUT4 #(
		.INIT('heee4)
	) name16554 (
		_w22352_,
		_w22374_,
		_w22359_,
		_w22380_,
		_w22381_
	);
	LUT2 #(
		.INIT('h4)
	) name16555 (
		_w22354_,
		_w22375_,
		_w22382_
	);
	LUT2 #(
		.INIT('h1)
	) name16556 (
		_w22381_,
		_w22382_,
		_w22383_
	);
	LUT4 #(
		.INIT('ha955)
	) name16557 (
		\u1_L2_reg[20]/NET0131 ,
		_w22367_,
		_w22379_,
		_w22383_,
		_w22384_
	);
	LUT4 #(
		.INIT('hc693)
	) name16558 (
		decrypt_pad,
		\u1_R2_reg[32]/NET0131 ,
		\u1_uk_K_r2_reg[42]/NET0131 ,
		\u1_uk_K_r2_reg[51]/NET0131 ,
		_w22385_
	);
	LUT4 #(
		.INIT('hc963)
	) name16559 (
		decrypt_pad,
		\u1_R2_reg[30]/NET0131 ,
		\u1_uk_K_r2_reg[2]/NET0131 ,
		\u1_uk_K_r2_reg[52]/NET0131 ,
		_w22386_
	);
	LUT4 #(
		.INIT('hc963)
	) name16560 (
		decrypt_pad,
		\u1_R2_reg[28]/NET0131 ,
		\u1_uk_K_r2_reg[29]/NET0131 ,
		\u1_uk_K_r2_reg[51]/NET0131 ,
		_w22387_
	);
	LUT4 #(
		.INIT('hc963)
	) name16561 (
		decrypt_pad,
		\u1_R2_reg[1]/NET0131 ,
		\u1_uk_K_r2_reg[45]/NET0131 ,
		\u1_uk_K_r2_reg[8]/NET0131 ,
		_w22388_
	);
	LUT4 #(
		.INIT('hc963)
	) name16562 (
		decrypt_pad,
		\u1_R2_reg[29]/NET0131 ,
		\u1_uk_K_r2_reg[1]/NET0131 ,
		\u1_uk_K_r2_reg[23]/NET0131 ,
		_w22389_
	);
	LUT4 #(
		.INIT('h0800)
	) name16563 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22390_
	);
	LUT4 #(
		.INIT('hc963)
	) name16564 (
		decrypt_pad,
		\u1_R2_reg[31]/P0001 ,
		\u1_uk_K_r2_reg[14]/NET0131 ,
		\u1_uk_K_r2_reg[36]/NET0131 ,
		_w22391_
	);
	LUT4 #(
		.INIT('h4555)
	) name16565 (
		_w22391_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22392_
	);
	LUT4 #(
		.INIT('h4554)
	) name16566 (
		_w22391_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22393_
	);
	LUT2 #(
		.INIT('h2)
	) name16567 (
		_w22387_,
		_w22386_,
		_w22394_
	);
	LUT2 #(
		.INIT('h4)
	) name16568 (
		_w22388_,
		_w22389_,
		_w22395_
	);
	LUT4 #(
		.INIT('h070d)
	) name16569 (
		_w22391_,
		_w22394_,
		_w22393_,
		_w22395_,
		_w22396_
	);
	LUT3 #(
		.INIT('ha8)
	) name16570 (
		_w22385_,
		_w22390_,
		_w22396_,
		_w22397_
	);
	LUT4 #(
		.INIT('h1000)
	) name16571 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22398_
	);
	LUT4 #(
		.INIT('haaa2)
	) name16572 (
		_w22391_,
		_w22388_,
		_w22389_,
		_w22387_,
		_w22399_
	);
	LUT3 #(
		.INIT('h10)
	) name16573 (
		_w22388_,
		_w22387_,
		_w22386_,
		_w22400_
	);
	LUT3 #(
		.INIT('h15)
	) name16574 (
		_w22391_,
		_w22388_,
		_w22389_,
		_w22401_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16575 (
		_w22398_,
		_w22399_,
		_w22400_,
		_w22401_,
		_w22402_
	);
	LUT3 #(
		.INIT('h04)
	) name16576 (
		_w22391_,
		_w22387_,
		_w22386_,
		_w22403_
	);
	LUT3 #(
		.INIT('h2a)
	) name16577 (
		_w22388_,
		_w22387_,
		_w22386_,
		_w22404_
	);
	LUT4 #(
		.INIT('h8040)
	) name16578 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22405_
	);
	LUT2 #(
		.INIT('h1)
	) name16579 (
		_w22403_,
		_w22405_,
		_w22406_
	);
	LUT3 #(
		.INIT('h51)
	) name16580 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22407_
	);
	LUT4 #(
		.INIT('hae22)
	) name16581 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22408_
	);
	LUT4 #(
		.INIT('h0420)
	) name16582 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22409_
	);
	LUT4 #(
		.INIT('h0200)
	) name16583 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22410_
	);
	LUT4 #(
		.INIT('h0001)
	) name16584 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22411_
	);
	LUT4 #(
		.INIT('hf9de)
	) name16585 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22412_
	);
	LUT4 #(
		.INIT('h31f5)
	) name16586 (
		_w22391_,
		_w22403_,
		_w22412_,
		_w22395_,
		_w22413_
	);
	LUT4 #(
		.INIT('hba00)
	) name16587 (
		_w22385_,
		_w22402_,
		_w22406_,
		_w22413_,
		_w22414_
	);
	LUT3 #(
		.INIT('h9a)
	) name16588 (
		\u1_L2_reg[5]/NET0131 ,
		_w22397_,
		_w22414_,
		_w22415_
	);
	LUT3 #(
		.INIT('h02)
	) name16589 (
		_w22352_,
		_w22360_,
		_w22362_,
		_w22416_
	);
	LUT4 #(
		.INIT('h00a2)
	) name16590 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22417_
	);
	LUT3 #(
		.INIT('h01)
	) name16591 (
		_w22352_,
		_w22374_,
		_w22417_,
		_w22418_
	);
	LUT4 #(
		.INIT('h6fff)
	) name16592 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22419_
	);
	LUT4 #(
		.INIT('h02aa)
	) name16593 (
		_w22363_,
		_w22416_,
		_w22418_,
		_w22419_,
		_w22420_
	);
	LUT3 #(
		.INIT('h08)
	) name16594 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22421_
	);
	LUT4 #(
		.INIT('h0400)
	) name16595 (
		_w22352_,
		_w22350_,
		_w22354_,
		_w22351_,
		_w22422_
	);
	LUT3 #(
		.INIT('h01)
	) name16596 (
		_w22368_,
		_w22421_,
		_w22422_,
		_w22423_
	);
	LUT3 #(
		.INIT('h8a)
	) name16597 (
		_w22352_,
		_w22354_,
		_w22351_,
		_w22424_
	);
	LUT4 #(
		.INIT('h0200)
	) name16598 (
		_w22352_,
		_w22350_,
		_w22354_,
		_w22351_,
		_w22425_
	);
	LUT3 #(
		.INIT('h07)
	) name16599 (
		_w22371_,
		_w22424_,
		_w22425_,
		_w22426_
	);
	LUT4 #(
		.INIT('h1333)
	) name16600 (
		_w22361_,
		_w22363_,
		_w22423_,
		_w22426_,
		_w22427_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name16601 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22428_
	);
	LUT2 #(
		.INIT('h1)
	) name16602 (
		_w22352_,
		_w22428_,
		_w22429_
	);
	LUT3 #(
		.INIT('h0b)
	) name16603 (
		_w22354_,
		_w22375_,
		_w22365_,
		_w22430_
	);
	LUT2 #(
		.INIT('h4)
	) name16604 (
		_w22429_,
		_w22430_,
		_w22431_
	);
	LUT4 #(
		.INIT('h5655)
	) name16605 (
		\u1_L2_reg[10]/NET0131 ,
		_w22427_,
		_w22420_,
		_w22431_,
		_w22432_
	);
	LUT4 #(
		.INIT('h0006)
	) name16606 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22433_
	);
	LUT3 #(
		.INIT('h47)
	) name16607 (
		_w22254_,
		_w22255_,
		_w22259_,
		_w22434_
	);
	LUT4 #(
		.INIT('h0051)
	) name16608 (
		_w22253_,
		_w22265_,
		_w22434_,
		_w22433_,
		_w22435_
	);
	LUT3 #(
		.INIT('h10)
	) name16609 (
		_w22254_,
		_w22256_,
		_w22258_,
		_w22436_
	);
	LUT4 #(
		.INIT('h2100)
	) name16610 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22437_
	);
	LUT2 #(
		.INIT('h6)
	) name16611 (
		_w22255_,
		_w22256_,
		_w22438_
	);
	LUT4 #(
		.INIT('h143c)
	) name16612 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22439_
	);
	LUT3 #(
		.INIT('h32)
	) name16613 (
		_w22259_,
		_w22437_,
		_w22439_,
		_w22440_
	);
	LUT2 #(
		.INIT('h8)
	) name16614 (
		_w22435_,
		_w22440_,
		_w22441_
	);
	LUT2 #(
		.INIT('h4)
	) name16615 (
		_w22259_,
		_w22266_,
		_w22442_
	);
	LUT3 #(
		.INIT('h02)
	) name16616 (
		_w22253_,
		_w22263_,
		_w22277_,
		_w22443_
	);
	LUT4 #(
		.INIT('h0240)
	) name16617 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22444_
	);
	LUT4 #(
		.INIT('h33fe)
	) name16618 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22445_
	);
	LUT3 #(
		.INIT('h31)
	) name16619 (
		_w22259_,
		_w22444_,
		_w22445_,
		_w22446_
	);
	LUT3 #(
		.INIT('h40)
	) name16620 (
		_w22442_,
		_w22443_,
		_w22446_,
		_w22447_
	);
	LUT3 #(
		.INIT('ha9)
	) name16621 (
		\u1_L2_reg[12]/NET0131 ,
		_w22441_,
		_w22447_,
		_w22448_
	);
	LUT4 #(
		.INIT('hc693)
	) name16622 (
		decrypt_pad,
		\u1_R2_reg[20]/NET0131 ,
		\u1_uk_K_r2_reg[31]/NET0131 ,
		\u1_uk_K_r2_reg[36]/NET0131 ,
		_w22449_
	);
	LUT4 #(
		.INIT('hc963)
	) name16623 (
		decrypt_pad,
		\u1_R2_reg[19]/NET0131 ,
		\u1_uk_K_r2_reg[21]/NET0131 ,
		\u1_uk_K_r2_reg[43]/NET0131 ,
		_w22450_
	);
	LUT4 #(
		.INIT('hc693)
	) name16624 (
		decrypt_pad,
		\u1_R2_reg[18]/NET0131 ,
		\u1_uk_K_r2_reg[1]/NET0131 ,
		\u1_uk_K_r2_reg[38]/NET0131 ,
		_w22451_
	);
	LUT4 #(
		.INIT('hc693)
	) name16625 (
		decrypt_pad,
		\u1_R2_reg[16]/NET0131 ,
		\u1_uk_K_r2_reg[16]/NET0131 ,
		\u1_uk_K_r2_reg[49]/NET0131 ,
		_w22452_
	);
	LUT4 #(
		.INIT('hc693)
	) name16626 (
		decrypt_pad,
		\u1_R2_reg[21]/NET0131 ,
		\u1_uk_K_r2_reg[28]/NET0131 ,
		\u1_uk_K_r2_reg[37]/NET0131 ,
		_w22453_
	);
	LUT4 #(
		.INIT('hc963)
	) name16627 (
		decrypt_pad,
		\u1_R2_reg[17]/NET0131 ,
		\u1_uk_K_r2_reg[16]/NET0131 ,
		\u1_uk_K_r2_reg[7]/NET0131 ,
		_w22454_
	);
	LUT3 #(
		.INIT('h02)
	) name16628 (
		_w22452_,
		_w22453_,
		_w22454_,
		_w22455_
	);
	LUT4 #(
		.INIT('h0002)
	) name16629 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22456_
	);
	LUT4 #(
		.INIT('h0800)
	) name16630 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22457_
	);
	LUT3 #(
		.INIT('h04)
	) name16631 (
		_w22452_,
		_w22453_,
		_w22454_,
		_w22458_
	);
	LUT4 #(
		.INIT('hc7b9)
	) name16632 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22459_
	);
	LUT3 #(
		.INIT('h10)
	) name16633 (
		_w22452_,
		_w22451_,
		_w22454_,
		_w22460_
	);
	LUT4 #(
		.INIT('h7a6e)
	) name16634 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22461_
	);
	LUT4 #(
		.INIT('h0180)
	) name16635 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22462_
	);
	LUT4 #(
		.INIT('h00d8)
	) name16636 (
		_w22450_,
		_w22461_,
		_w22459_,
		_w22462_,
		_w22463_
	);
	LUT2 #(
		.INIT('h1)
	) name16637 (
		_w22449_,
		_w22463_,
		_w22464_
	);
	LUT4 #(
		.INIT('h95b3)
	) name16638 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22465_
	);
	LUT2 #(
		.INIT('h4)
	) name16639 (
		_w22465_,
		_w22450_,
		_w22466_
	);
	LUT2 #(
		.INIT('h9)
	) name16640 (
		_w22451_,
		_w22454_,
		_w22467_
	);
	LUT4 #(
		.INIT('h0220)
	) name16641 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22468_
	);
	LUT4 #(
		.INIT('h0888)
	) name16642 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22450_,
		_w22469_
	);
	LUT3 #(
		.INIT('h13)
	) name16643 (
		_w22467_,
		_w22468_,
		_w22469_,
		_w22470_
	);
	LUT3 #(
		.INIT('h8a)
	) name16644 (
		_w22449_,
		_w22466_,
		_w22470_,
		_w22471_
	);
	LUT4 #(
		.INIT('h0010)
	) name16645 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22472_
	);
	LUT4 #(
		.INIT('h0200)
	) name16646 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22473_
	);
	LUT3 #(
		.INIT('h02)
	) name16647 (
		_w22450_,
		_w22473_,
		_w22472_,
		_w22474_
	);
	LUT3 #(
		.INIT('h40)
	) name16648 (
		_w22452_,
		_w22453_,
		_w22454_,
		_w22475_
	);
	LUT3 #(
		.INIT('hbe)
	) name16649 (
		_w22452_,
		_w22453_,
		_w22454_,
		_w22476_
	);
	LUT2 #(
		.INIT('h2)
	) name16650 (
		_w22449_,
		_w22451_,
		_w22477_
	);
	LUT4 #(
		.INIT('h1040)
	) name16651 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22478_
	);
	LUT4 #(
		.INIT('h1011)
	) name16652 (
		_w22450_,
		_w22478_,
		_w22476_,
		_w22477_,
		_w22479_
	);
	LUT2 #(
		.INIT('h1)
	) name16653 (
		_w22474_,
		_w22479_,
		_w22480_
	);
	LUT4 #(
		.INIT('h5556)
	) name16654 (
		\u1_L2_reg[14]/NET0131 ,
		_w22471_,
		_w22480_,
		_w22464_,
		_w22481_
	);
	LUT4 #(
		.INIT('hfe3c)
	) name16655 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22482_
	);
	LUT2 #(
		.INIT('h1)
	) name16656 (
		_w22291_,
		_w22482_,
		_w22483_
	);
	LUT4 #(
		.INIT('h35f3)
	) name16657 (
		_w22287_,
		_w22291_,
		_w22288_,
		_w22286_,
		_w22484_
	);
	LUT4 #(
		.INIT('h0501)
	) name16658 (
		_w22284_,
		_w22285_,
		_w22310_,
		_w22484_,
		_w22485_
	);
	LUT4 #(
		.INIT('h0040)
	) name16659 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22486_
	);
	LUT4 #(
		.INIT('hf0b5)
	) name16660 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22487_
	);
	LUT2 #(
		.INIT('h2)
	) name16661 (
		_w22291_,
		_w22487_,
		_w22488_
	);
	LUT4 #(
		.INIT('h1000)
	) name16662 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22489_
	);
	LUT4 #(
		.INIT('h2021)
	) name16663 (
		_w22287_,
		_w22291_,
		_w22285_,
		_w22286_,
		_w22490_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name16664 (
		_w22284_,
		_w22287_,
		_w22288_,
		_w22286_,
		_w22491_
	);
	LUT3 #(
		.INIT('h10)
	) name16665 (
		_w22490_,
		_w22489_,
		_w22491_,
		_w22492_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16666 (
		_w22483_,
		_w22485_,
		_w22488_,
		_w22492_,
		_w22493_
	);
	LUT3 #(
		.INIT('he0)
	) name16667 (
		_w22287_,
		_w22288_,
		_w22286_,
		_w22494_
	);
	LUT4 #(
		.INIT('h004c)
	) name16668 (
		_w22287_,
		_w22291_,
		_w22288_,
		_w22285_,
		_w22495_
	);
	LUT2 #(
		.INIT('h8)
	) name16669 (
		_w22494_,
		_w22495_,
		_w22496_
	);
	LUT3 #(
		.INIT('h56)
	) name16670 (
		\u1_L2_reg[17]/NET0131 ,
		_w22493_,
		_w22496_,
		_w22497_
	);
	LUT4 #(
		.INIT('hccfd)
	) name16671 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22498_
	);
	LUT4 #(
		.INIT('h6fbf)
	) name16672 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22499_
	);
	LUT4 #(
		.INIT('h08aa)
	) name16673 (
		_w22352_,
		_w22363_,
		_w22498_,
		_w22499_,
		_w22500_
	);
	LUT4 #(
		.INIT('h220a)
	) name16674 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22501_
	);
	LUT4 #(
		.INIT('hfda8)
	) name16675 (
		_w22352_,
		_w22358_,
		_w22380_,
		_w22501_,
		_w22502_
	);
	LUT4 #(
		.INIT('h7bf7)
	) name16676 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22503_
	);
	LUT3 #(
		.INIT('h45)
	) name16677 (
		_w22363_,
		_w22502_,
		_w22503_,
		_w22504_
	);
	LUT4 #(
		.INIT('hb3fb)
	) name16678 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22505_
	);
	LUT4 #(
		.INIT('h0080)
	) name16679 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22506_
	);
	LUT4 #(
		.INIT('hef6f)
	) name16680 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22507_
	);
	LUT4 #(
		.INIT('h04cc)
	) name16681 (
		_w22352_,
		_w22363_,
		_w22505_,
		_w22507_,
		_w22508_
	);
	LUT2 #(
		.INIT('h1)
	) name16682 (
		_w22352_,
		_w22351_,
		_w22509_
	);
	LUT2 #(
		.INIT('h4)
	) name16683 (
		_w22507_,
		_w22509_,
		_w22510_
	);
	LUT2 #(
		.INIT('h1)
	) name16684 (
		_w22508_,
		_w22510_,
		_w22511_
	);
	LUT4 #(
		.INIT('h5655)
	) name16685 (
		\u1_L2_reg[1]/NET0131 ,
		_w22504_,
		_w22500_,
		_w22511_,
		_w22512_
	);
	LUT2 #(
		.INIT('h4)
	) name16686 (
		_w22391_,
		_w22388_,
		_w22513_
	);
	LUT4 #(
		.INIT('h0400)
	) name16687 (
		_w22391_,
		_w22388_,
		_w22389_,
		_w22386_,
		_w22514_
	);
	LUT3 #(
		.INIT('h08)
	) name16688 (
		_w22389_,
		_w22387_,
		_w22386_,
		_w22515_
	);
	LUT4 #(
		.INIT('h0002)
	) name16689 (
		_w22391_,
		_w22388_,
		_w22389_,
		_w22387_,
		_w22516_
	);
	LUT4 #(
		.INIT('h0002)
	) name16690 (
		_w22385_,
		_w22514_,
		_w22515_,
		_w22516_,
		_w22517_
	);
	LUT4 #(
		.INIT('h0400)
	) name16691 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22518_
	);
	LUT4 #(
		.INIT('h2000)
	) name16692 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22519_
	);
	LUT4 #(
		.INIT('hdbff)
	) name16693 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22520_
	);
	LUT4 #(
		.INIT('h3d39)
	) name16694 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22521_
	);
	LUT4 #(
		.INIT('h0010)
	) name16695 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22522_
	);
	LUT4 #(
		.INIT('h0051)
	) name16696 (
		_w22385_,
		_w22391_,
		_w22521_,
		_w22522_,
		_w22523_
	);
	LUT3 #(
		.INIT('h07)
	) name16697 (
		_w22517_,
		_w22520_,
		_w22523_,
		_w22524_
	);
	LUT4 #(
		.INIT('hfff6)
	) name16698 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22525_
	);
	LUT3 #(
		.INIT('h20)
	) name16699 (
		_w22392_,
		_w22518_,
		_w22525_,
		_w22526_
	);
	LUT4 #(
		.INIT('h0002)
	) name16700 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22527_
	);
	LUT3 #(
		.INIT('h02)
	) name16701 (
		_w22391_,
		_w22390_,
		_w22527_,
		_w22528_
	);
	LUT2 #(
		.INIT('h1)
	) name16702 (
		_w22385_,
		_w22391_,
		_w22529_
	);
	LUT4 #(
		.INIT('h0100)
	) name16703 (
		_w22385_,
		_w22391_,
		_w22389_,
		_w22387_,
		_w22530_
	);
	LUT3 #(
		.INIT('h0e)
	) name16704 (
		_w22526_,
		_w22528_,
		_w22530_,
		_w22531_
	);
	LUT3 #(
		.INIT('h65)
	) name16705 (
		\u1_L2_reg[15]/P0001 ,
		_w22524_,
		_w22531_,
		_w22532_
	);
	LUT4 #(
		.INIT('haa2a)
	) name16706 (
		_w22391_,
		_w22388_,
		_w22389_,
		_w22387_,
		_w22533_
	);
	LUT4 #(
		.INIT('h3fdd)
	) name16707 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22534_
	);
	LUT4 #(
		.INIT('h5545)
	) name16708 (
		_w22391_,
		_w22388_,
		_w22387_,
		_w22386_,
		_w22535_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name16709 (
		_w22519_,
		_w22533_,
		_w22534_,
		_w22535_,
		_w22536_
	);
	LUT4 #(
		.INIT('h4100)
	) name16710 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22537_
	);
	LUT3 #(
		.INIT('h02)
	) name16711 (
		_w22385_,
		_w22527_,
		_w22537_,
		_w22538_
	);
	LUT2 #(
		.INIT('h4)
	) name16712 (
		_w22536_,
		_w22538_,
		_w22539_
	);
	LUT4 #(
		.INIT('h002e)
	) name16713 (
		_w22391_,
		_w22388_,
		_w22387_,
		_w22386_,
		_w22540_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name16714 (
		_w22391_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22541_
	);
	LUT3 #(
		.INIT('h10)
	) name16715 (
		_w22407_,
		_w22540_,
		_w22541_,
		_w22542_
	);
	LUT2 #(
		.INIT('h1)
	) name16716 (
		_w22385_,
		_w22398_,
		_w22543_
	);
	LUT3 #(
		.INIT('h70)
	) name16717 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22544_
	);
	LUT3 #(
		.INIT('ha8)
	) name16718 (
		_w22391_,
		_w22389_,
		_w22386_,
		_w22545_
	);
	LUT3 #(
		.INIT('h15)
	) name16719 (
		_w22411_,
		_w22544_,
		_w22545_,
		_w22546_
	);
	LUT3 #(
		.INIT('h40)
	) name16720 (
		_w22542_,
		_w22543_,
		_w22546_,
		_w22547_
	);
	LUT4 #(
		.INIT('h0002)
	) name16721 (
		_w22391_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22548_
	);
	LUT3 #(
		.INIT('h07)
	) name16722 (
		_w22513_,
		_w22515_,
		_w22548_,
		_w22549_
	);
	LUT4 #(
		.INIT('ha955)
	) name16723 (
		\u1_L2_reg[21]/NET0131 ,
		_w22539_,
		_w22547_,
		_w22549_,
		_w22550_
	);
	LUT4 #(
		.INIT('h67a8)
	) name16724 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22551_
	);
	LUT4 #(
		.INIT('hfa77)
	) name16725 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22552_
	);
	LUT4 #(
		.INIT('hd3ff)
	) name16726 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22553_
	);
	LUT4 #(
		.INIT('hd800)
	) name16727 (
		_w22450_,
		_w22551_,
		_w22552_,
		_w22553_,
		_w22554_
	);
	LUT2 #(
		.INIT('h2)
	) name16728 (
		_w22449_,
		_w22554_,
		_w22555_
	);
	LUT3 #(
		.INIT('hb0)
	) name16729 (
		_w22453_,
		_w22454_,
		_w22450_,
		_w22556_
	);
	LUT4 #(
		.INIT('h3301)
	) name16730 (
		_w22452_,
		_w22451_,
		_w22454_,
		_w22450_,
		_w22557_
	);
	LUT2 #(
		.INIT('h4)
	) name16731 (
		_w22556_,
		_w22557_,
		_w22558_
	);
	LUT4 #(
		.INIT('h4000)
	) name16732 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22559_
	);
	LUT4 #(
		.INIT('hafdd)
	) name16733 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22560_
	);
	LUT3 #(
		.INIT('h32)
	) name16734 (
		_w22450_,
		_w22559_,
		_w22560_,
		_w22561_
	);
	LUT4 #(
		.INIT('hdfef)
	) name16735 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22562_
	);
	LUT4 #(
		.INIT('hdfeb)
	) name16736 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22563_
	);
	LUT4 #(
		.INIT('h0008)
	) name16737 (
		_w22452_,
		_w22451_,
		_w22454_,
		_w22450_,
		_w22564_
	);
	LUT4 #(
		.INIT('h0301)
	) name16738 (
		_w22450_,
		_w22457_,
		_w22564_,
		_w22563_,
		_w22565_
	);
	LUT4 #(
		.INIT('hba00)
	) name16739 (
		_w22449_,
		_w22558_,
		_w22561_,
		_w22565_,
		_w22566_
	);
	LUT3 #(
		.INIT('h65)
	) name16740 (
		\u1_L2_reg[25]/NET0131 ,
		_w22555_,
		_w22566_,
		_w22567_
	);
	LUT3 #(
		.INIT('h02)
	) name16741 (
		_w22352_,
		_w22374_,
		_w22362_,
		_w22568_
	);
	LUT4 #(
		.INIT('h0806)
	) name16742 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22569_
	);
	LUT4 #(
		.INIT('hefcc)
	) name16743 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22570_
	);
	LUT4 #(
		.INIT('h0504)
	) name16744 (
		_w22352_,
		_w22363_,
		_w22569_,
		_w22570_,
		_w22571_
	);
	LUT2 #(
		.INIT('h1)
	) name16745 (
		_w22568_,
		_w22571_,
		_w22572_
	);
	LUT4 #(
		.INIT('h0002)
	) name16746 (
		_w22352_,
		_w22350_,
		_w22349_,
		_w22351_,
		_w22573_
	);
	LUT4 #(
		.INIT('h0004)
	) name16747 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22574_
	);
	LUT4 #(
		.INIT('h0002)
	) name16748 (
		_w22363_,
		_w22506_,
		_w22573_,
		_w22574_,
		_w22575_
	);
	LUT4 #(
		.INIT('h54ff)
	) name16749 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22351_,
		_w22576_
	);
	LUT3 #(
		.INIT('h51)
	) name16750 (
		_w22352_,
		_w22350_,
		_w22354_,
		_w22577_
	);
	LUT4 #(
		.INIT('hcdff)
	) name16751 (
		_w22352_,
		_w22350_,
		_w22349_,
		_w22351_,
		_w22578_
	);
	LUT4 #(
		.INIT('hcf45)
	) name16752 (
		_w22354_,
		_w22576_,
		_w22577_,
		_w22578_,
		_w22579_
	);
	LUT2 #(
		.INIT('h2)
	) name16753 (
		_w22364_,
		_w22376_,
		_w22580_
	);
	LUT4 #(
		.INIT('h00fd)
	) name16754 (
		_w22350_,
		_w22349_,
		_w22354_,
		_w22363_,
		_w22581_
	);
	LUT3 #(
		.INIT('h10)
	) name16755 (
		_w22374_,
		_w22375_,
		_w22581_,
		_w22582_
	);
	LUT4 #(
		.INIT('h7077)
	) name16756 (
		_w22575_,
		_w22579_,
		_w22580_,
		_w22582_,
		_w22583_
	);
	LUT3 #(
		.INIT('h56)
	) name16757 (
		\u1_L2_reg[26]/NET0131 ,
		_w22572_,
		_w22583_,
		_w22584_
	);
	LUT4 #(
		.INIT('h779a)
	) name16758 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22585_
	);
	LUT4 #(
		.INIT('h0e02)
	) name16759 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22586_
	);
	LUT4 #(
		.INIT('hf17d)
	) name16760 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22587_
	);
	LUT4 #(
		.INIT('h1000)
	) name16761 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22588_
	);
	LUT4 #(
		.INIT('h00e4)
	) name16762 (
		_w22316_,
		_w22587_,
		_w22585_,
		_w22588_,
		_w22589_
	);
	LUT2 #(
		.INIT('h1)
	) name16763 (
		_w22315_,
		_w22589_,
		_w22590_
	);
	LUT4 #(
		.INIT('hdd7d)
	) name16764 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22591_
	);
	LUT2 #(
		.INIT('h2)
	) name16765 (
		_w22316_,
		_w22591_,
		_w22592_
	);
	LUT3 #(
		.INIT('h48)
	) name16766 (
		_w22318_,
		_w22319_,
		_w22320_,
		_w22593_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name16767 (
		_w22317_,
		_w22319_,
		_w22316_,
		_w22320_,
		_w22594_
	);
	LUT3 #(
		.INIT('h01)
	) name16768 (
		_w22586_,
		_w22594_,
		_w22593_,
		_w22595_
	);
	LUT4 #(
		.INIT('h0004)
	) name16769 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22596_
	);
	LUT4 #(
		.INIT('h2000)
	) name16770 (
		_w22317_,
		_w22319_,
		_w22316_,
		_w22320_,
		_w22597_
	);
	LUT2 #(
		.INIT('h1)
	) name16771 (
		_w22596_,
		_w22597_,
		_w22598_
	);
	LUT4 #(
		.INIT('h5700)
	) name16772 (
		_w22315_,
		_w22592_,
		_w22595_,
		_w22598_,
		_w22599_
	);
	LUT3 #(
		.INIT('h9a)
	) name16773 (
		\u1_L2_reg[29]/NET0131 ,
		_w22590_,
		_w22599_,
		_w22600_
	);
	LUT4 #(
		.INIT('hc693)
	) name16774 (
		decrypt_pad,
		\u1_R2_reg[8]/NET0131 ,
		\u1_uk_K_r2_reg[17]/NET0131 ,
		\u1_uk_K_r2_reg[54]/NET0131 ,
		_w22601_
	);
	LUT4 #(
		.INIT('hc693)
	) name16775 (
		decrypt_pad,
		\u1_R2_reg[7]/NET0131 ,
		\u1_uk_K_r2_reg[26]/NET0131 ,
		\u1_uk_K_r2_reg[6]/NET0131 ,
		_w22602_
	);
	LUT4 #(
		.INIT('hc693)
	) name16776 (
		decrypt_pad,
		\u1_R2_reg[5]/NET0131 ,
		\u1_uk_K_r2_reg[41]/NET0131 ,
		\u1_uk_K_r2_reg[46]/NET0131 ,
		_w22603_
	);
	LUT4 #(
		.INIT('hc963)
	) name16777 (
		decrypt_pad,
		\u1_R2_reg[4]/NET0131 ,
		\u1_uk_K_r2_reg[10]/NET0131 ,
		\u1_uk_K_r2_reg[5]/NET0131 ,
		_w22604_
	);
	LUT4 #(
		.INIT('hc963)
	) name16778 (
		decrypt_pad,
		\u1_R2_reg[9]/NET0131 ,
		\u1_uk_K_r2_reg[34]/NET0131 ,
		\u1_uk_K_r2_reg[54]/NET0131 ,
		_w22605_
	);
	LUT4 #(
		.INIT('hc963)
	) name16779 (
		decrypt_pad,
		\u1_R2_reg[6]/NET0131 ,
		\u1_uk_K_r2_reg[12]/NET0131 ,
		\u1_uk_K_r2_reg[32]/NET0131 ,
		_w22606_
	);
	LUT4 #(
		.INIT('h59fb)
	) name16780 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22607_
	);
	LUT2 #(
		.INIT('h1)
	) name16781 (
		_w22602_,
		_w22607_,
		_w22608_
	);
	LUT4 #(
		.INIT('h0034)
	) name16782 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22609_
	);
	LUT4 #(
		.INIT('h0800)
	) name16783 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22610_
	);
	LUT4 #(
		.INIT('h0004)
	) name16784 (
		_w22602_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22611_
	);
	LUT4 #(
		.INIT('h4000)
	) name16785 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22612_
	);
	LUT4 #(
		.INIT('h0007)
	) name16786 (
		_w22602_,
		_w22610_,
		_w22611_,
		_w22612_,
		_w22613_
	);
	LUT4 #(
		.INIT('h5455)
	) name16787 (
		_w22601_,
		_w22608_,
		_w22609_,
		_w22613_,
		_w22614_
	);
	LUT4 #(
		.INIT('he6ee)
	) name16788 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22615_
	);
	LUT4 #(
		.INIT('h4044)
	) name16789 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22616_
	);
	LUT3 #(
		.INIT('h51)
	) name16790 (
		_w22602_,
		_w22603_,
		_w22606_,
		_w22617_
	);
	LUT4 #(
		.INIT('hf200)
	) name16791 (
		_w22601_,
		_w22615_,
		_w22616_,
		_w22617_,
		_w22618_
	);
	LUT4 #(
		.INIT('h0002)
	) name16792 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22619_
	);
	LUT4 #(
		.INIT('h80a0)
	) name16793 (
		_w22602_,
		_w22604_,
		_w22603_,
		_w22606_,
		_w22620_
	);
	LUT4 #(
		.INIT('h0080)
	) name16794 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22621_
	);
	LUT4 #(
		.INIT('haaa8)
	) name16795 (
		_w22601_,
		_w22619_,
		_w22620_,
		_w22621_,
		_w22622_
	);
	LUT3 #(
		.INIT('ha2)
	) name16796 (
		_w22604_,
		_w22603_,
		_w22606_,
		_w22623_
	);
	LUT3 #(
		.INIT('h45)
	) name16797 (
		_w22604_,
		_w22603_,
		_w22606_,
		_w22624_
	);
	LUT3 #(
		.INIT('h8a)
	) name16798 (
		_w22602_,
		_w22604_,
		_w22605_,
		_w22625_
	);
	LUT3 #(
		.INIT('h10)
	) name16799 (
		_w22624_,
		_w22623_,
		_w22625_,
		_w22626_
	);
	LUT3 #(
		.INIT('h01)
	) name16800 (
		_w22622_,
		_w22626_,
		_w22618_,
		_w22627_
	);
	LUT3 #(
		.INIT('h65)
	) name16801 (
		\u1_L2_reg[2]/NET0131 ,
		_w22614_,
		_w22627_,
		_w22628_
	);
	LUT2 #(
		.INIT('h1)
	) name16802 (
		_w22604_,
		_w22606_,
		_w22629_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name16803 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22630_
	);
	LUT2 #(
		.INIT('h2)
	) name16804 (
		_w22602_,
		_w22630_,
		_w22631_
	);
	LUT4 #(
		.INIT('hbfae)
	) name16805 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22632_
	);
	LUT2 #(
		.INIT('h1)
	) name16806 (
		_w22602_,
		_w22632_,
		_w22633_
	);
	LUT2 #(
		.INIT('h8)
	) name16807 (
		_w22602_,
		_w22604_,
		_w22634_
	);
	LUT4 #(
		.INIT('h7737)
	) name16808 (
		_w22602_,
		_w22604_,
		_w22605_,
		_w22603_,
		_w22635_
	);
	LUT4 #(
		.INIT('h0400)
	) name16809 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22636_
	);
	LUT3 #(
		.INIT('h0e)
	) name16810 (
		_w22606_,
		_w22635_,
		_w22636_,
		_w22637_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name16811 (
		_w22601_,
		_w22633_,
		_w22631_,
		_w22637_,
		_w22638_
	);
	LUT4 #(
		.INIT('hdaff)
	) name16812 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22639_
	);
	LUT2 #(
		.INIT('h1)
	) name16813 (
		_w22602_,
		_w22639_,
		_w22640_
	);
	LUT3 #(
		.INIT('h02)
	) name16814 (
		_w22604_,
		_w22605_,
		_w22606_,
		_w22641_
	);
	LUT4 #(
		.INIT('h1145)
	) name16815 (
		_w22602_,
		_w22604_,
		_w22605_,
		_w22603_,
		_w22642_
	);
	LUT4 #(
		.INIT('h7077)
	) name16816 (
		_w22602_,
		_w22632_,
		_w22641_,
		_w22642_,
		_w22643_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name16817 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22644_
	);
	LUT4 #(
		.INIT('h2322)
	) name16818 (
		_w22601_,
		_w22640_,
		_w22643_,
		_w22644_,
		_w22645_
	);
	LUT3 #(
		.INIT('h65)
	) name16819 (
		\u1_L2_reg[28]/NET0131 ,
		_w22638_,
		_w22645_,
		_w22646_
	);
	LUT4 #(
		.INIT('h2000)
	) name16820 (
		_w22318_,
		_w22319_,
		_w22316_,
		_w22320_,
		_w22647_
	);
	LUT4 #(
		.INIT('h7f00)
	) name16821 (
		_w22317_,
		_w22319_,
		_w22320_,
		_w22315_,
		_w22648_
	);
	LUT2 #(
		.INIT('h4)
	) name16822 (
		_w22647_,
		_w22648_,
		_w22649_
	);
	LUT3 #(
		.INIT('h51)
	) name16823 (
		_w22343_,
		_w22327_,
		_w22321_,
		_w22650_
	);
	LUT4 #(
		.INIT('hf070)
	) name16824 (
		_w22317_,
		_w22318_,
		_w22316_,
		_w22320_,
		_w22651_
	);
	LUT4 #(
		.INIT('hbcff)
	) name16825 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22652_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name16826 (
		_w22317_,
		_w22318_,
		_w22316_,
		_w22320_,
		_w22653_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name16827 (
		_w22588_,
		_w22651_,
		_w22652_,
		_w22653_,
		_w22654_
	);
	LUT3 #(
		.INIT('h01)
	) name16828 (
		_w22315_,
		_w22328_,
		_w22596_,
		_w22655_
	);
	LUT4 #(
		.INIT('h7077)
	) name16829 (
		_w22649_,
		_w22650_,
		_w22654_,
		_w22655_,
		_w22656_
	);
	LUT3 #(
		.INIT('h31)
	) name16830 (
		_w22317_,
		_w22318_,
		_w22320_,
		_w22657_
	);
	LUT4 #(
		.INIT('hd060)
	) name16831 (
		_w22317_,
		_w22318_,
		_w22316_,
		_w22320_,
		_w22658_
	);
	LUT4 #(
		.INIT('h070b)
	) name16832 (
		_w22317_,
		_w22318_,
		_w22316_,
		_w22320_,
		_w22659_
	);
	LUT4 #(
		.INIT('h3331)
	) name16833 (
		_w22319_,
		_w22345_,
		_w22659_,
		_w22658_,
		_w22660_
	);
	LUT3 #(
		.INIT('h65)
	) name16834 (
		\u1_L2_reg[4]/NET0131 ,
		_w22656_,
		_w22660_,
		_w22661_
	);
	LUT3 #(
		.INIT('h10)
	) name16835 (
		_w22605_,
		_w22603_,
		_w22606_,
		_w22662_
	);
	LUT4 #(
		.INIT('h5515)
	) name16836 (
		_w22602_,
		_w22604_,
		_w22605_,
		_w22603_,
		_w22663_
	);
	LUT3 #(
		.INIT('h40)
	) name16837 (
		_w22604_,
		_w22605_,
		_w22606_,
		_w22664_
	);
	LUT4 #(
		.INIT('haaa8)
	) name16838 (
		_w22602_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22665_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16839 (
		_w22662_,
		_w22663_,
		_w22664_,
		_w22665_,
		_w22666_
	);
	LUT4 #(
		.INIT('h0010)
	) name16840 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22667_
	);
	LUT4 #(
		.INIT('h0002)
	) name16841 (
		_w22601_,
		_w22611_,
		_w22612_,
		_w22667_,
		_w22668_
	);
	LUT2 #(
		.INIT('h4)
	) name16842 (
		_w22666_,
		_w22668_,
		_w22669_
	);
	LUT3 #(
		.INIT('hc8)
	) name16843 (
		_w22602_,
		_w22605_,
		_w22603_,
		_w22670_
	);
	LUT2 #(
		.INIT('h8)
	) name16844 (
		_w22629_,
		_w22670_,
		_w22671_
	);
	LUT3 #(
		.INIT('hb0)
	) name16845 (
		_w22605_,
		_w22603_,
		_w22606_,
		_w22672_
	);
	LUT3 #(
		.INIT('h15)
	) name16846 (
		_w22601_,
		_w22634_,
		_w22672_,
		_w22673_
	);
	LUT3 #(
		.INIT('h10)
	) name16847 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22674_
	);
	LUT4 #(
		.INIT('h0001)
	) name16848 (
		_w22602_,
		_w22619_,
		_w22636_,
		_w22674_,
		_w22675_
	);
	LUT3 #(
		.INIT('h40)
	) name16849 (
		_w22671_,
		_w22673_,
		_w22675_,
		_w22676_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name16850 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22677_
	);
	LUT4 #(
		.INIT('h0929)
	) name16851 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22678_
	);
	LUT2 #(
		.INIT('h2)
	) name16852 (
		_w22602_,
		_w22678_,
		_w22679_
	);
	LUT3 #(
		.INIT('h40)
	) name16853 (
		_w22671_,
		_w22673_,
		_w22679_,
		_w22680_
	);
	LUT4 #(
		.INIT('h001f)
	) name16854 (
		_w22669_,
		_w22676_,
		_w22677_,
		_w22680_,
		_w22681_
	);
	LUT2 #(
		.INIT('h9)
	) name16855 (
		\u1_L2_reg[13]/NET0131 ,
		_w22681_,
		_w22682_
	);
	LUT4 #(
		.INIT('h0201)
	) name16856 (
		_w22317_,
		_w22318_,
		_w22316_,
		_w22320_,
		_w22683_
	);
	LUT4 #(
		.INIT('hf700)
	) name16857 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22316_,
		_w22684_
	);
	LUT4 #(
		.INIT('h8000)
	) name16858 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22685_
	);
	LUT4 #(
		.INIT('h0045)
	) name16859 (
		_w22315_,
		_w22657_,
		_w22684_,
		_w22685_,
		_w22686_
	);
	LUT4 #(
		.INIT('h2010)
	) name16860 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22687_
	);
	LUT3 #(
		.INIT('h04)
	) name16861 (
		_w22332_,
		_w22315_,
		_w22687_,
		_w22688_
	);
	LUT4 #(
		.INIT('h010a)
	) name16862 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22320_,
		_w22689_
	);
	LUT4 #(
		.INIT('h0844)
	) name16863 (
		_w22317_,
		_w22318_,
		_w22319_,
		_w22316_,
		_w22690_
	);
	LUT2 #(
		.INIT('h1)
	) name16864 (
		_w22689_,
		_w22690_,
		_w22691_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name16865 (
		_w22683_,
		_w22686_,
		_w22688_,
		_w22691_,
		_w22692_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name16866 (
		_w22317_,
		_w22319_,
		_w22341_,
		_w22328_,
		_w22693_
	);
	LUT3 #(
		.INIT('h65)
	) name16867 (
		\u1_L2_reg[19]/NET0131 ,
		_w22692_,
		_w22693_,
		_w22694_
	);
	LUT4 #(
		.INIT('hfcd3)
	) name16868 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22695_
	);
	LUT4 #(
		.INIT('heffb)
	) name16869 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22696_
	);
	LUT4 #(
		.INIT('h0233)
	) name16870 (
		_w22284_,
		_w22291_,
		_w22695_,
		_w22696_,
		_w22697_
	);
	LUT4 #(
		.INIT('h02a0)
	) name16871 (
		_w22291_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22698_
	);
	LUT3 #(
		.INIT('h54)
	) name16872 (
		_w22303_,
		_w22309_,
		_w22698_,
		_w22699_
	);
	LUT3 #(
		.INIT('h8c)
	) name16873 (
		_w22287_,
		_w22291_,
		_w22285_,
		_w22700_
	);
	LUT2 #(
		.INIT('h8)
	) name16874 (
		_w22304_,
		_w22700_,
		_w22701_
	);
	LUT4 #(
		.INIT('h002a)
	) name16875 (
		_w22284_,
		_w22295_,
		_w22307_,
		_w22486_,
		_w22702_
	);
	LUT4 #(
		.INIT('h1554)
	) name16876 (
		_w22284_,
		_w22287_,
		_w22288_,
		_w22286_,
		_w22703_
	);
	LUT3 #(
		.INIT('h47)
	) name16877 (
		_w22287_,
		_w22288_,
		_w22286_,
		_w22704_
	);
	LUT3 #(
		.INIT('h07)
	) name16878 (
		_w22287_,
		_w22288_,
		_w22286_,
		_w22705_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name16879 (
		_w22291_,
		_w22285_,
		_w22704_,
		_w22705_,
		_w22706_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name16880 (
		_w22701_,
		_w22702_,
		_w22703_,
		_w22706_,
		_w22707_
	);
	LUT4 #(
		.INIT('haaa9)
	) name16881 (
		\u1_L2_reg[23]/NET0131 ,
		_w22699_,
		_w22707_,
		_w22697_,
		_w22708_
	);
	LUT4 #(
		.INIT('hb7b4)
	) name16882 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22709_
	);
	LUT2 #(
		.INIT('h1)
	) name16883 (
		_w22391_,
		_w22709_,
		_w22710_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name16884 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22711_
	);
	LUT4 #(
		.INIT('h80aa)
	) name16885 (
		_w22391_,
		_w22388_,
		_w22389_,
		_w22387_,
		_w22712_
	);
	LUT4 #(
		.INIT('he7dd)
	) name16886 (
		_w22388_,
		_w22389_,
		_w22387_,
		_w22386_,
		_w22713_
	);
	LUT3 #(
		.INIT('hb0)
	) name16887 (
		_w22711_,
		_w22712_,
		_w22713_,
		_w22714_
	);
	LUT3 #(
		.INIT('h8a)
	) name16888 (
		_w22385_,
		_w22710_,
		_w22714_,
		_w22715_
	);
	LUT4 #(
		.INIT('haa8a)
	) name16889 (
		_w22391_,
		_w22388_,
		_w22389_,
		_w22386_,
		_w22716_
	);
	LUT4 #(
		.INIT('h4544)
	) name16890 (
		_w22385_,
		_w22410_,
		_w22408_,
		_w22716_,
		_w22717_
	);
	LUT2 #(
		.INIT('h4)
	) name16891 (
		_w22391_,
		_w22409_,
		_w22718_
	);
	LUT3 #(
		.INIT('h10)
	) name16892 (
		_w22404_,
		_w22407_,
		_w22529_,
		_w22719_
	);
	LUT4 #(
		.INIT('h0200)
	) name16893 (
		_w22391_,
		_w22388_,
		_w22389_,
		_w22386_,
		_w22720_
	);
	LUT3 #(
		.INIT('h07)
	) name16894 (
		_w22403_,
		_w22395_,
		_w22720_,
		_w22721_
	);
	LUT4 #(
		.INIT('h0100)
	) name16895 (
		_w22717_,
		_w22719_,
		_w22718_,
		_w22721_,
		_w22722_
	);
	LUT3 #(
		.INIT('h65)
	) name16896 (
		\u1_L2_reg[27]/NET0131 ,
		_w22715_,
		_w22722_,
		_w22723_
	);
	LUT2 #(
		.INIT('h9)
	) name16897 (
		_w22256_,
		_w22258_,
		_w22724_
	);
	LUT4 #(
		.INIT('hd003)
	) name16898 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22725_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name16899 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22726_
	);
	LUT3 #(
		.INIT('h01)
	) name16900 (
		_w22259_,
		_w22726_,
		_w22725_,
		_w22727_
	);
	LUT4 #(
		.INIT('h0800)
	) name16901 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22728_
	);
	LUT4 #(
		.INIT('hb5bc)
	) name16902 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22729_
	);
	LUT3 #(
		.INIT('h31)
	) name16903 (
		_w22259_,
		_w22728_,
		_w22729_,
		_w22730_
	);
	LUT3 #(
		.INIT('h8a)
	) name16904 (
		_w22253_,
		_w22727_,
		_w22730_,
		_w22731_
	);
	LUT3 #(
		.INIT('h40)
	) name16905 (
		_w22255_,
		_w22256_,
		_w22258_,
		_w22732_
	);
	LUT4 #(
		.INIT('hab89)
	) name16906 (
		_w22259_,
		_w22436_,
		_w22438_,
		_w22732_,
		_w22733_
	);
	LUT4 #(
		.INIT('h7bd7)
	) name16907 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22734_
	);
	LUT4 #(
		.INIT('h00c8)
	) name16908 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22259_,
		_w22735_
	);
	LUT4 #(
		.INIT('h135f)
	) name16909 (
		_w22259_,
		_w22274_,
		_w22266_,
		_w22735_,
		_w22736_
	);
	LUT4 #(
		.INIT('hba00)
	) name16910 (
		_w22253_,
		_w22733_,
		_w22734_,
		_w22736_,
		_w22737_
	);
	LUT3 #(
		.INIT('h65)
	) name16911 (
		\u1_L2_reg[32]/NET0131 ,
		_w22731_,
		_w22737_,
		_w22738_
	);
	LUT4 #(
		.INIT('hc693)
	) name16912 (
		decrypt_pad,
		\u1_R2_reg[11]/NET0131 ,
		\u1_uk_K_r2_reg[12]/NET0131 ,
		\u1_uk_K_r2_reg[17]/NET0131 ,
		_w22739_
	);
	LUT4 #(
		.INIT('hc693)
	) name16913 (
		decrypt_pad,
		\u1_R2_reg[12]/NET0131 ,
		\u1_uk_K_r2_reg[27]/NET0131 ,
		\u1_uk_K_r2_reg[32]/NET0131 ,
		_w22740_
	);
	LUT4 #(
		.INIT('hc693)
	) name16914 (
		decrypt_pad,
		\u1_R2_reg[9]/NET0131 ,
		\u1_uk_K_r2_reg[3]/NET0131 ,
		\u1_uk_K_r2_reg[40]/NET0131 ,
		_w22741_
	);
	LUT4 #(
		.INIT('hc963)
	) name16915 (
		decrypt_pad,
		\u1_R2_reg[13]/NET0131 ,
		\u1_uk_K_r2_reg[20]/NET0131 ,
		\u1_uk_K_r2_reg[40]/NET0131 ,
		_w22742_
	);
	LUT4 #(
		.INIT('hc693)
	) name16916 (
		decrypt_pad,
		\u1_R2_reg[10]/NET0131 ,
		\u1_uk_K_r2_reg[11]/NET0131 ,
		\u1_uk_K_r2_reg[48]/NET0131 ,
		_w22743_
	);
	LUT4 #(
		.INIT('hc963)
	) name16917 (
		decrypt_pad,
		\u1_R2_reg[8]/NET0131 ,
		\u1_uk_K_r2_reg[11]/NET0131 ,
		\u1_uk_K_r2_reg[6]/NET0131 ,
		_w22744_
	);
	LUT4 #(
		.INIT('hf35f)
	) name16918 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22745_
	);
	LUT4 #(
		.INIT('ha25f)
	) name16919 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22746_
	);
	LUT2 #(
		.INIT('h1)
	) name16920 (
		_w22744_,
		_w22742_,
		_w22747_
	);
	LUT4 #(
		.INIT('h0001)
	) name16921 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22748_
	);
	LUT4 #(
		.INIT('hbbfe)
	) name16922 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22749_
	);
	LUT4 #(
		.INIT('h08cc)
	) name16923 (
		_w22740_,
		_w22739_,
		_w22746_,
		_w22749_,
		_w22750_
	);
	LUT2 #(
		.INIT('h6)
	) name16924 (
		_w22744_,
		_w22742_,
		_w22751_
	);
	LUT4 #(
		.INIT('he00e)
	) name16925 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22752_
	);
	LUT4 #(
		.INIT('h6006)
	) name16926 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22753_
	);
	LUT4 #(
		.INIT('h0800)
	) name16927 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22754_
	);
	LUT2 #(
		.INIT('h4)
	) name16928 (
		_w22739_,
		_w22754_,
		_w22755_
	);
	LUT4 #(
		.INIT('h1101)
	) name16929 (
		_w22741_,
		_w22743_,
		_w22739_,
		_w22744_,
		_w22756_
	);
	LUT4 #(
		.INIT('h0020)
	) name16930 (
		_w22741_,
		_w22743_,
		_w22739_,
		_w22744_,
		_w22757_
	);
	LUT4 #(
		.INIT('h0080)
	) name16931 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22758_
	);
	LUT4 #(
		.INIT('h0111)
	) name16932 (
		_w22757_,
		_w22758_,
		_w22751_,
		_w22756_,
		_w22759_
	);
	LUT4 #(
		.INIT('h5455)
	) name16933 (
		_w22740_,
		_w22755_,
		_w22753_,
		_w22759_,
		_w22760_
	);
	LUT3 #(
		.INIT('h80)
	) name16934 (
		_w22740_,
		_w22741_,
		_w22743_,
		_w22761_
	);
	LUT3 #(
		.INIT('h0d)
	) name16935 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22762_
	);
	LUT4 #(
		.INIT('h0802)
	) name16936 (
		_w22740_,
		_w22741_,
		_w22739_,
		_w22742_,
		_w22763_
	);
	LUT4 #(
		.INIT('h7077)
	) name16937 (
		_w22747_,
		_w22761_,
		_w22762_,
		_w22763_,
		_w22764_
	);
	LUT4 #(
		.INIT('h5655)
	) name16938 (
		\u1_L2_reg[6]/NET0131 ,
		_w22760_,
		_w22750_,
		_w22764_,
		_w22765_
	);
	LUT4 #(
		.INIT('hf126)
	) name16939 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22766_
	);
	LUT4 #(
		.INIT('h2880)
	) name16940 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22767_
	);
	LUT4 #(
		.INIT('h5004)
	) name16941 (
		_w22254_,
		_w22255_,
		_w22256_,
		_w22258_,
		_w22768_
	);
	LUT4 #(
		.INIT('h1302)
	) name16942 (
		_w22259_,
		_w22767_,
		_w22768_,
		_w22766_,
		_w22769_
	);
	LUT2 #(
		.INIT('h2)
	) name16943 (
		_w22253_,
		_w22769_,
		_w22770_
	);
	LUT2 #(
		.INIT('h4)
	) name16944 (
		_w22259_,
		_w22767_,
		_w22771_
	);
	LUT2 #(
		.INIT('h2)
	) name16945 (
		_w22253_,
		_w22259_,
		_w22772_
	);
	LUT3 #(
		.INIT('h4c)
	) name16946 (
		_w22255_,
		_w22256_,
		_w22258_,
		_w22773_
	);
	LUT4 #(
		.INIT('h8a00)
	) name16947 (
		_w22254_,
		_w22256_,
		_w22258_,
		_w22259_,
		_w22774_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name16948 (
		_w22260_,
		_w22724_,
		_w22773_,
		_w22774_,
		_w22775_
	);
	LUT3 #(
		.INIT('h45)
	) name16949 (
		_w22273_,
		_w22259_,
		_w22768_,
		_w22776_
	);
	LUT4 #(
		.INIT('h0133)
	) name16950 (
		_w22253_,
		_w22772_,
		_w22775_,
		_w22776_,
		_w22777_
	);
	LUT4 #(
		.INIT('h5556)
	) name16951 (
		\u1_L2_reg[7]/NET0131 ,
		_w22771_,
		_w22777_,
		_w22770_,
		_w22778_
	);
	LUT4 #(
		.INIT('hff76)
	) name16952 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22779_
	);
	LUT3 #(
		.INIT('h02)
	) name16953 (
		_w22452_,
		_w22451_,
		_w22450_,
		_w22780_
	);
	LUT4 #(
		.INIT('h0031)
	) name16954 (
		_w22450_,
		_w22478_,
		_w22779_,
		_w22780_,
		_w22781_
	);
	LUT2 #(
		.INIT('h2)
	) name16955 (
		_w22449_,
		_w22781_,
		_w22782_
	);
	LUT4 #(
		.INIT('h8000)
	) name16956 (
		_w22452_,
		_w22453_,
		_w22454_,
		_w22450_,
		_w22783_
	);
	LUT3 #(
		.INIT('h04)
	) name16957 (
		_w22460_,
		_w22562_,
		_w22783_,
		_w22784_
	);
	LUT4 #(
		.INIT('hbb73)
	) name16958 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22785_
	);
	LUT3 #(
		.INIT('h72)
	) name16959 (
		_w22450_,
		_w22456_,
		_w22785_,
		_w22786_
	);
	LUT4 #(
		.INIT('hcbbf)
	) name16960 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22787_
	);
	LUT4 #(
		.INIT('haf23)
	) name16961 (
		_w22453_,
		_w22450_,
		_w22564_,
		_w22787_,
		_w22788_
	);
	LUT4 #(
		.INIT('hea00)
	) name16962 (
		_w22449_,
		_w22784_,
		_w22786_,
		_w22788_,
		_w22789_
	);
	LUT3 #(
		.INIT('h65)
	) name16963 (
		\u1_L2_reg[8]/NET0131 ,
		_w22782_,
		_w22789_,
		_w22790_
	);
	LUT3 #(
		.INIT('h80)
	) name16964 (
		_w22741_,
		_w22744_,
		_w22742_,
		_w22791_
	);
	LUT4 #(
		.INIT('h5aa7)
	) name16965 (
		_w22741_,
		_w22739_,
		_w22744_,
		_w22742_,
		_w22792_
	);
	LUT2 #(
		.INIT('h1)
	) name16966 (
		_w22743_,
		_w22792_,
		_w22793_
	);
	LUT4 #(
		.INIT('h0012)
	) name16967 (
		_w22743_,
		_w22739_,
		_w22744_,
		_w22742_,
		_w22794_
	);
	LUT3 #(
		.INIT('h02)
	) name16968 (
		_w22740_,
		_w22754_,
		_w22794_,
		_w22795_
	);
	LUT4 #(
		.INIT('h5afc)
	) name16969 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22796_
	);
	LUT2 #(
		.INIT('h1)
	) name16970 (
		_w22739_,
		_w22796_,
		_w22797_
	);
	LUT4 #(
		.INIT('h4880)
	) name16971 (
		_w22741_,
		_w22739_,
		_w22744_,
		_w22742_,
		_w22798_
	);
	LUT3 #(
		.INIT('h01)
	) name16972 (
		_w22740_,
		_w22748_,
		_w22798_,
		_w22799_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name16973 (
		_w22793_,
		_w22795_,
		_w22797_,
		_w22799_,
		_w22800_
	);
	LUT4 #(
		.INIT('h0400)
	) name16974 (
		_w22741_,
		_w22743_,
		_w22739_,
		_w22744_,
		_w22801_
	);
	LUT4 #(
		.INIT('hff7b)
	) name16975 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22802_
	);
	LUT3 #(
		.INIT('h31)
	) name16976 (
		_w22739_,
		_w22801_,
		_w22802_,
		_w22803_
	);
	LUT3 #(
		.INIT('h65)
	) name16977 (
		\u1_L2_reg[16]/NET0131 ,
		_w22800_,
		_w22803_,
		_w22804_
	);
	LUT4 #(
		.INIT('hefbe)
	) name16978 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22805_
	);
	LUT3 #(
		.INIT('h40)
	) name16979 (
		_w22739_,
		_w22745_,
		_w22805_,
		_w22806_
	);
	LUT3 #(
		.INIT('hed)
	) name16980 (
		_w22743_,
		_w22744_,
		_w22742_,
		_w22807_
	);
	LUT3 #(
		.INIT('h02)
	) name16981 (
		_w22741_,
		_w22744_,
		_w22742_,
		_w22808_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name16982 (
		_w22741_,
		_w22743_,
		_w22739_,
		_w22744_,
		_w22809_
	);
	LUT3 #(
		.INIT('h20)
	) name16983 (
		_w22807_,
		_w22808_,
		_w22809_,
		_w22810_
	);
	LUT3 #(
		.INIT('h54)
	) name16984 (
		_w22740_,
		_w22806_,
		_w22810_,
		_w22811_
	);
	LUT2 #(
		.INIT('h4)
	) name16985 (
		_w22743_,
		_w22739_,
		_w22812_
	);
	LUT3 #(
		.INIT('h45)
	) name16986 (
		_w22741_,
		_w22744_,
		_w22742_,
		_w22813_
	);
	LUT2 #(
		.INIT('h8)
	) name16987 (
		_w22812_,
		_w22813_,
		_w22814_
	);
	LUT3 #(
		.INIT('h2a)
	) name16988 (
		_w22740_,
		_w22751_,
		_w22756_,
		_w22815_
	);
	LUT4 #(
		.INIT('h737f)
	) name16989 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22816_
	);
	LUT3 #(
		.INIT('hb1)
	) name16990 (
		_w22739_,
		_w22752_,
		_w22816_,
		_w22817_
	);
	LUT3 #(
		.INIT('h40)
	) name16991 (
		_w22814_,
		_w22815_,
		_w22817_,
		_w22818_
	);
	LUT2 #(
		.INIT('h2)
	) name16992 (
		_w22743_,
		_w22739_,
		_w22819_
	);
	LUT3 #(
		.INIT('he4)
	) name16993 (
		_w22741_,
		_w22744_,
		_w22742_,
		_w22820_
	);
	LUT4 #(
		.INIT('h0444)
	) name16994 (
		_w22743_,
		_w22739_,
		_w22744_,
		_w22742_,
		_w22821_
	);
	LUT4 #(
		.INIT('h0777)
	) name16995 (
		_w22791_,
		_w22819_,
		_w22820_,
		_w22821_,
		_w22822_
	);
	LUT4 #(
		.INIT('ha955)
	) name16996 (
		\u1_L2_reg[24]/NET0131 ,
		_w22811_,
		_w22818_,
		_w22822_,
		_w22823_
	);
	LUT4 #(
		.INIT('hfce3)
	) name16997 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22824_
	);
	LUT4 #(
		.INIT('h0888)
	) name16998 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22825_
	);
	LUT4 #(
		.INIT('h3f35)
	) name16999 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22826_
	);
	LUT4 #(
		.INIT('h3210)
	) name17000 (
		_w22739_,
		_w22825_,
		_w22826_,
		_w22824_,
		_w22827_
	);
	LUT2 #(
		.INIT('h2)
	) name17001 (
		_w22740_,
		_w22827_,
		_w22828_
	);
	LUT3 #(
		.INIT('h13)
	) name17002 (
		_w22743_,
		_w22739_,
		_w22744_,
		_w22829_
	);
	LUT4 #(
		.INIT('hebfe)
	) name17003 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22830_
	);
	LUT4 #(
		.INIT('h4055)
	) name17004 (
		_w22740_,
		_w22820_,
		_w22829_,
		_w22830_,
		_w22831_
	);
	LUT4 #(
		.INIT('h0008)
	) name17005 (
		_w22741_,
		_w22743_,
		_w22739_,
		_w22742_,
		_w22832_
	);
	LUT4 #(
		.INIT('h3f9d)
	) name17006 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22833_
	);
	LUT4 #(
		.INIT('h4000)
	) name17007 (
		_w22741_,
		_w22743_,
		_w22744_,
		_w22742_,
		_w22834_
	);
	LUT4 #(
		.INIT('hcc04)
	) name17008 (
		_w22740_,
		_w22739_,
		_w22833_,
		_w22834_,
		_w22835_
	);
	LUT3 #(
		.INIT('h01)
	) name17009 (
		_w22832_,
		_w22835_,
		_w22831_,
		_w22836_
	);
	LUT3 #(
		.INIT('h9a)
	) name17010 (
		\u1_L2_reg[30]/NET0131 ,
		_w22828_,
		_w22836_,
		_w22837_
	);
	LUT4 #(
		.INIT('he6f7)
	) name17011 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22838_
	);
	LUT4 #(
		.INIT('hf7df)
	) name17012 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22839_
	);
	LUT4 #(
		.INIT('hb100)
	) name17013 (
		_w22450_,
		_w22475_,
		_w22838_,
		_w22839_,
		_w22840_
	);
	LUT2 #(
		.INIT('h2)
	) name17014 (
		_w22449_,
		_w22840_,
		_w22841_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name17015 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22842_
	);
	LUT4 #(
		.INIT('h00d0)
	) name17016 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22843_
	);
	LUT4 #(
		.INIT('h2e26)
	) name17017 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22844_
	);
	LUT4 #(
		.INIT('h3210)
	) name17018 (
		_w22450_,
		_w22843_,
		_w22844_,
		_w22842_,
		_w22845_
	);
	LUT4 #(
		.INIT('hfd7e)
	) name17019 (
		_w22452_,
		_w22453_,
		_w22451_,
		_w22454_,
		_w22846_
	);
	LUT2 #(
		.INIT('h1)
	) name17020 (
		_w22450_,
		_w22846_,
		_w22847_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name17021 (
		_w22451_,
		_w22450_,
		_w22458_,
		_w22455_,
		_w22848_
	);
	LUT4 #(
		.INIT('h0e00)
	) name17022 (
		_w22449_,
		_w22845_,
		_w22847_,
		_w22848_,
		_w22849_
	);
	LUT3 #(
		.INIT('h65)
	) name17023 (
		\u1_L2_reg[3]/NET0131 ,
		_w22841_,
		_w22849_,
		_w22850_
	);
	LUT4 #(
		.INIT('hdc33)
	) name17024 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22851_
	);
	LUT2 #(
		.INIT('h2)
	) name17025 (
		_w22291_,
		_w22851_,
		_w22852_
	);
	LUT4 #(
		.INIT('h0082)
	) name17026 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22853_
	);
	LUT3 #(
		.INIT('h25)
	) name17027 (
		_w22288_,
		_w22285_,
		_w22286_,
		_w22854_
	);
	LUT4 #(
		.INIT('h0411)
	) name17028 (
		_w22291_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22855_
	);
	LUT4 #(
		.INIT('h4000)
	) name17029 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22856_
	);
	LUT3 #(
		.INIT('h01)
	) name17030 (
		_w22855_,
		_w22853_,
		_w22856_,
		_w22857_
	);
	LUT3 #(
		.INIT('h45)
	) name17031 (
		_w22284_,
		_w22852_,
		_w22857_,
		_w22858_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name17032 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22859_
	);
	LUT2 #(
		.INIT('h1)
	) name17033 (
		_w22291_,
		_w22859_,
		_w22860_
	);
	LUT4 #(
		.INIT('h8228)
	) name17034 (
		_w22287_,
		_w22288_,
		_w22285_,
		_w22286_,
		_w22861_
	);
	LUT4 #(
		.INIT('h0013)
	) name17035 (
		_w22292_,
		_w22489_,
		_w22854_,
		_w22861_,
		_w22862_
	);
	LUT3 #(
		.INIT('h31)
	) name17036 (
		_w22284_,
		_w22860_,
		_w22862_,
		_w22863_
	);
	LUT3 #(
		.INIT('h65)
	) name17037 (
		\u1_L2_reg[9]/NET0131 ,
		_w22858_,
		_w22863_,
		_w22864_
	);
	LUT4 #(
		.INIT('h0a20)
	) name17038 (
		_w22602_,
		_w22604_,
		_w22605_,
		_w22603_,
		_w22865_
	);
	LUT3 #(
		.INIT('he4)
	) name17039 (
		_w22605_,
		_w22603_,
		_w22606_,
		_w22866_
	);
	LUT3 #(
		.INIT('h74)
	) name17040 (
		_w22602_,
		_w22604_,
		_w22606_,
		_w22867_
	);
	LUT4 #(
		.INIT('h8a88)
	) name17041 (
		_w22601_,
		_w22865_,
		_w22866_,
		_w22867_,
		_w22868_
	);
	LUT4 #(
		.INIT('h8000)
	) name17042 (
		_w22602_,
		_w22604_,
		_w22605_,
		_w22603_,
		_w22869_
	);
	LUT4 #(
		.INIT('hdffc)
	) name17043 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22870_
	);
	LUT4 #(
		.INIT('h1003)
	) name17044 (
		_w22602_,
		_w22604_,
		_w22603_,
		_w22606_,
		_w22871_
	);
	LUT4 #(
		.INIT('h0100)
	) name17045 (
		_w22610_,
		_w22869_,
		_w22871_,
		_w22870_,
		_w22872_
	);
	LUT4 #(
		.INIT('h1000)
	) name17046 (
		_w22602_,
		_w22604_,
		_w22605_,
		_w22603_,
		_w22873_
	);
	LUT4 #(
		.INIT('h77ef)
	) name17047 (
		_w22604_,
		_w22605_,
		_w22603_,
		_w22606_,
		_w22874_
	);
	LUT3 #(
		.INIT('h31)
	) name17048 (
		_w22602_,
		_w22873_,
		_w22874_,
		_w22875_
	);
	LUT4 #(
		.INIT('h0e00)
	) name17049 (
		_w22601_,
		_w22872_,
		_w22868_,
		_w22875_,
		_w22876_
	);
	LUT2 #(
		.INIT('h9)
	) name17050 (
		\u1_L2_reg[18]/NET0131 ,
		_w22876_,
		_w22877_
	);
	LUT4 #(
		.INIT('hc963)
	) name17051 (
		decrypt_pad,
		\u1_R1_reg[4]/NET0131 ,
		\u1_uk_K_r1_reg[10]/P0001 ,
		\u1_uk_K_r1_reg[34]/NET0131 ,
		_w22878_
	);
	LUT4 #(
		.INIT('hc693)
	) name17052 (
		decrypt_pad,
		\u1_R1_reg[32]/NET0131 ,
		\u1_uk_K_r1_reg[11]/NET0131 ,
		\u1_uk_K_r1_reg[19]/NET0131 ,
		_w22879_
	);
	LUT4 #(
		.INIT('hc693)
	) name17053 (
		decrypt_pad,
		\u1_R1_reg[1]/NET0131 ,
		\u1_uk_K_r1_reg[32]/NET0131 ,
		\u1_uk_K_r1_reg[40]/NET0131 ,
		_w22880_
	);
	LUT4 #(
		.INIT('hc693)
	) name17054 (
		decrypt_pad,
		\u1_R1_reg[2]/NET0131 ,
		\u1_uk_K_r1_reg[47]/NET0131 ,
		\u1_uk_K_r1_reg[55]/NET0131 ,
		_w22881_
	);
	LUT4 #(
		.INIT('hc963)
	) name17055 (
		decrypt_pad,
		\u1_R1_reg[5]/NET0131 ,
		\u1_uk_K_r1_reg[13]/NET0131 ,
		\u1_uk_K_r1_reg[5]/NET0131 ,
		_w22882_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name17056 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22883_
	);
	LUT2 #(
		.INIT('h1)
	) name17057 (
		_w22882_,
		_w22879_,
		_w22884_
	);
	LUT4 #(
		.INIT('hc693)
	) name17058 (
		decrypt_pad,
		\u1_R1_reg[3]/NET0131 ,
		\u1_uk_K_r1_reg[24]/NET0131 ,
		\u1_uk_K_r1_reg[32]/NET0131 ,
		_w22885_
	);
	LUT2 #(
		.INIT('h4)
	) name17059 (
		_w22881_,
		_w22885_,
		_w22886_
	);
	LUT3 #(
		.INIT('hb0)
	) name17060 (
		_w22881_,
		_w22885_,
		_w22880_,
		_w22887_
	);
	LUT3 #(
		.INIT('h01)
	) name17061 (
		_w22884_,
		_w22887_,
		_w22883_,
		_w22888_
	);
	LUT3 #(
		.INIT('h02)
	) name17062 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22889_
	);
	LUT4 #(
		.INIT('hfd31)
	) name17063 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22890_
	);
	LUT4 #(
		.INIT('h300a)
	) name17064 (
		_w22881_,
		_w22885_,
		_w22879_,
		_w22880_,
		_w22891_
	);
	LUT3 #(
		.INIT('h0d)
	) name17065 (
		_w22885_,
		_w22890_,
		_w22891_,
		_w22892_
	);
	LUT3 #(
		.INIT('h8a)
	) name17066 (
		_w22878_,
		_w22888_,
		_w22892_,
		_w22893_
	);
	LUT3 #(
		.INIT('he6)
	) name17067 (
		_w22881_,
		_w22879_,
		_w22880_,
		_w22894_
	);
	LUT3 #(
		.INIT('h51)
	) name17068 (
		_w22885_,
		_w22882_,
		_w22880_,
		_w22895_
	);
	LUT2 #(
		.INIT('h4)
	) name17069 (
		_w22894_,
		_w22895_,
		_w22896_
	);
	LUT2 #(
		.INIT('h8)
	) name17070 (
		_w22881_,
		_w22885_,
		_w22897_
	);
	LUT3 #(
		.INIT('h60)
	) name17071 (
		_w22882_,
		_w22879_,
		_w22880_,
		_w22898_
	);
	LUT4 #(
		.INIT('h7c3f)
	) name17072 (
		_w22885_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22899_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name17073 (
		_w22881_,
		_w22885_,
		_w22898_,
		_w22899_,
		_w22900_
	);
	LUT2 #(
		.INIT('h2)
	) name17074 (
		_w22885_,
		_w22880_,
		_w22901_
	);
	LUT3 #(
		.INIT('had)
	) name17075 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22902_
	);
	LUT4 #(
		.INIT('h8000)
	) name17076 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22903_
	);
	LUT4 #(
		.INIT('h0008)
	) name17077 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22904_
	);
	LUT4 #(
		.INIT('h6ef7)
	) name17078 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22905_
	);
	LUT4 #(
		.INIT('hfda8)
	) name17079 (
		_w22885_,
		_w22880_,
		_w22902_,
		_w22905_,
		_w22906_
	);
	LUT4 #(
		.INIT('hba00)
	) name17080 (
		_w22878_,
		_w22896_,
		_w22900_,
		_w22906_,
		_w22907_
	);
	LUT3 #(
		.INIT('h65)
	) name17081 (
		\u1_L1_reg[31]/NET0131 ,
		_w22893_,
		_w22907_,
		_w22908_
	);
	LUT4 #(
		.INIT('hc693)
	) name17082 (
		decrypt_pad,
		\u1_R1_reg[24]/NET0131 ,
		\u1_uk_K_r1_reg[1]/NET0131 ,
		\u1_uk_K_r1_reg[7]/P0001 ,
		_w22909_
	);
	LUT4 #(
		.INIT('hc693)
	) name17083 (
		decrypt_pad,
		\u1_R1_reg[20]/NET0131 ,
		\u1_uk_K_r1_reg[35]/NET0131 ,
		\u1_uk_K_r1_reg[45]/NET0131 ,
		_w22910_
	);
	LUT4 #(
		.INIT('hc963)
	) name17084 (
		decrypt_pad,
		\u1_R1_reg[21]/NET0131 ,
		\u1_uk_K_r1_reg[1]/NET0131 ,
		\u1_uk_K_r1_reg[50]/NET0131 ,
		_w22911_
	);
	LUT4 #(
		.INIT('hc963)
	) name17085 (
		decrypt_pad,
		\u1_R1_reg[25]/NET0131 ,
		\u1_uk_K_r1_reg[2]/NET0131 ,
		\u1_uk_K_r1_reg[51]/NET0131 ,
		_w22912_
	);
	LUT4 #(
		.INIT('hc963)
	) name17086 (
		decrypt_pad,
		\u1_R1_reg[22]/NET0131 ,
		\u1_uk_K_r1_reg[23]/NET0131 ,
		\u1_uk_K_r1_reg[45]/NET0131 ,
		_w22913_
	);
	LUT4 #(
		.INIT('h4155)
	) name17087 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22914_
	);
	LUT3 #(
		.INIT('h80)
	) name17088 (
		_w22913_,
		_w22910_,
		_w22912_,
		_w22915_
	);
	LUT4 #(
		.INIT('hc693)
	) name17089 (
		decrypt_pad,
		\u1_R1_reg[23]/NET0131 ,
		\u1_uk_K_r1_reg[30]/NET0131 ,
		\u1_uk_K_r1_reg[36]/NET0131 ,
		_w22916_
	);
	LUT4 #(
		.INIT('h00df)
	) name17090 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22916_,
		_w22917_
	);
	LUT3 #(
		.INIT('h10)
	) name17091 (
		_w22915_,
		_w22914_,
		_w22917_,
		_w22918_
	);
	LUT4 #(
		.INIT('h0004)
	) name17092 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22919_
	);
	LUT4 #(
		.INIT('h1fdb)
	) name17093 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22920_
	);
	LUT2 #(
		.INIT('h2)
	) name17094 (
		_w22916_,
		_w22920_,
		_w22921_
	);
	LUT3 #(
		.INIT('ha8)
	) name17095 (
		_w22909_,
		_w22918_,
		_w22921_,
		_w22922_
	);
	LUT4 #(
		.INIT('h1900)
	) name17096 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22916_,
		_w22923_
	);
	LUT4 #(
		.INIT('h0040)
	) name17097 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22924_
	);
	LUT3 #(
		.INIT('h10)
	) name17098 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w22925_
	);
	LUT4 #(
		.INIT('h1000)
	) name17099 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w22916_,
		_w22926_
	);
	LUT3 #(
		.INIT('h01)
	) name17100 (
		_w22924_,
		_w22926_,
		_w22923_,
		_w22927_
	);
	LUT2 #(
		.INIT('h1)
	) name17101 (
		_w22913_,
		_w22916_,
		_w22928_
	);
	LUT4 #(
		.INIT('h0004)
	) name17102 (
		_w22913_,
		_w22910_,
		_w22912_,
		_w22916_,
		_w22929_
	);
	LUT4 #(
		.INIT('h0800)
	) name17103 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22930_
	);
	LUT4 #(
		.INIT('h0060)
	) name17104 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22916_,
		_w22931_
	);
	LUT3 #(
		.INIT('h01)
	) name17105 (
		_w22929_,
		_w22930_,
		_w22931_,
		_w22932_
	);
	LUT3 #(
		.INIT('h15)
	) name17106 (
		_w22909_,
		_w22927_,
		_w22932_,
		_w22933_
	);
	LUT4 #(
		.INIT('h77ef)
	) name17107 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22934_
	);
	LUT2 #(
		.INIT('h2)
	) name17108 (
		_w22916_,
		_w22934_,
		_w22935_
	);
	LUT3 #(
		.INIT('hf6)
	) name17109 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w22936_
	);
	LUT4 #(
		.INIT('hbfae)
	) name17110 (
		_w22913_,
		_w22916_,
		_w22925_,
		_w22936_,
		_w22937_
	);
	LUT2 #(
		.INIT('h4)
	) name17111 (
		_w22935_,
		_w22937_,
		_w22938_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name17112 (
		\u1_L1_reg[11]/NET0131 ,
		_w22933_,
		_w22922_,
		_w22938_,
		_w22939_
	);
	LUT4 #(
		.INIT('hc963)
	) name17113 (
		decrypt_pad,
		\u1_R1_reg[28]/NET0131 ,
		\u1_uk_K_r1_reg[14]/NET0131 ,
		\u1_uk_K_r1_reg[8]/NET0131 ,
		_w22940_
	);
	LUT4 #(
		.INIT('hc693)
	) name17114 (
		decrypt_pad,
		\u1_R1_reg[24]/NET0131 ,
		\u1_uk_K_r1_reg[23]/NET0131 ,
		\u1_uk_K_r1_reg[29]/NET0131 ,
		_w22941_
	);
	LUT4 #(
		.INIT('hc693)
	) name17115 (
		decrypt_pad,
		\u1_R1_reg[26]/NET0131 ,
		\u1_uk_K_r1_reg[43]/NET0131 ,
		\u1_uk_K_r1_reg[49]/NET0131 ,
		_w22942_
	);
	LUT4 #(
		.INIT('hc693)
	) name17116 (
		decrypt_pad,
		\u1_R1_reg[25]/NET0131 ,
		\u1_uk_K_r1_reg[31]/NET0131 ,
		\u1_uk_K_r1_reg[9]/NET0131 ,
		_w22943_
	);
	LUT4 #(
		.INIT('hc693)
	) name17117 (
		decrypt_pad,
		\u1_R1_reg[27]/NET0131 ,
		\u1_uk_K_r1_reg[21]/NET0131 ,
		\u1_uk_K_r1_reg[31]/NET0131 ,
		_w22944_
	);
	LUT4 #(
		.INIT('hc693)
	) name17118 (
		decrypt_pad,
		\u1_R1_reg[29]/NET0131 ,
		\u1_uk_K_r1_reg[0]/NET0131 ,
		\u1_uk_K_r1_reg[37]/NET0131 ,
		_w22945_
	);
	LUT4 #(
		.INIT('hfc3a)
	) name17119 (
		_w22945_,
		_w22943_,
		_w22942_,
		_w22944_,
		_w22946_
	);
	LUT2 #(
		.INIT('h2)
	) name17120 (
		_w22941_,
		_w22946_,
		_w22947_
	);
	LUT4 #(
		.INIT('h0100)
	) name17121 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w22948_
	);
	LUT2 #(
		.INIT('h6)
	) name17122 (
		_w22941_,
		_w22942_,
		_w22949_
	);
	LUT3 #(
		.INIT('h8a)
	) name17123 (
		_w22945_,
		_w22943_,
		_w22944_,
		_w22950_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name17124 (
		_w22948_,
		_w22944_,
		_w22949_,
		_w22950_,
		_w22951_
	);
	LUT4 #(
		.INIT('h0100)
	) name17125 (
		_w22945_,
		_w22943_,
		_w22942_,
		_w22944_,
		_w22952_
	);
	LUT4 #(
		.INIT('h0082)
	) name17126 (
		_w22943_,
		_w22941_,
		_w22942_,
		_w22944_,
		_w22953_
	);
	LUT2 #(
		.INIT('h1)
	) name17127 (
		_w22952_,
		_w22953_,
		_w22954_
	);
	LUT4 #(
		.INIT('hba00)
	) name17128 (
		_w22940_,
		_w22947_,
		_w22951_,
		_w22954_,
		_w22955_
	);
	LUT4 #(
		.INIT('hf47c)
	) name17129 (
		_w22940_,
		_w22945_,
		_w22943_,
		_w22942_,
		_w22956_
	);
	LUT4 #(
		.INIT('h0600)
	) name17130 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w22957_
	);
	LUT4 #(
		.INIT('hcc08)
	) name17131 (
		_w22941_,
		_w22944_,
		_w22956_,
		_w22957_,
		_w22958_
	);
	LUT2 #(
		.INIT('h2)
	) name17132 (
		_w22945_,
		_w22941_,
		_w22959_
	);
	LUT4 #(
		.INIT('hf700)
	) name17133 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w22960_
	);
	LUT3 #(
		.INIT('h20)
	) name17134 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22961_
	);
	LUT4 #(
		.INIT('h0028)
	) name17135 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22944_,
		_w22962_
	);
	LUT4 #(
		.INIT('h0200)
	) name17136 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w22963_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name17137 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w22964_
	);
	LUT4 #(
		.INIT('h20aa)
	) name17138 (
		_w22940_,
		_w22960_,
		_w22962_,
		_w22964_,
		_w22965_
	);
	LUT2 #(
		.INIT('h1)
	) name17139 (
		_w22958_,
		_w22965_,
		_w22966_
	);
	LUT3 #(
		.INIT('h95)
	) name17140 (
		\u1_L1_reg[22]/NET0131 ,
		_w22955_,
		_w22966_,
		_w22967_
	);
	LUT4 #(
		.INIT('hfe3c)
	) name17141 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22968_
	);
	LUT2 #(
		.INIT('h1)
	) name17142 (
		_w22885_,
		_w22968_,
		_w22969_
	);
	LUT4 #(
		.INIT('h35f3)
	) name17143 (
		_w22881_,
		_w22885_,
		_w22882_,
		_w22880_,
		_w22970_
	);
	LUT4 #(
		.INIT('h0501)
	) name17144 (
		_w22878_,
		_w22879_,
		_w22904_,
		_w22970_,
		_w22971_
	);
	LUT4 #(
		.INIT('h0040)
	) name17145 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22972_
	);
	LUT4 #(
		.INIT('hf0b5)
	) name17146 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22973_
	);
	LUT2 #(
		.INIT('h2)
	) name17147 (
		_w22885_,
		_w22973_,
		_w22974_
	);
	LUT4 #(
		.INIT('h1000)
	) name17148 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w22975_
	);
	LUT4 #(
		.INIT('h2021)
	) name17149 (
		_w22881_,
		_w22885_,
		_w22879_,
		_w22880_,
		_w22976_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name17150 (
		_w22878_,
		_w22881_,
		_w22882_,
		_w22880_,
		_w22977_
	);
	LUT3 #(
		.INIT('h10)
	) name17151 (
		_w22976_,
		_w22975_,
		_w22977_,
		_w22978_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17152 (
		_w22969_,
		_w22971_,
		_w22974_,
		_w22978_,
		_w22979_
	);
	LUT3 #(
		.INIT('he0)
	) name17153 (
		_w22881_,
		_w22882_,
		_w22880_,
		_w22980_
	);
	LUT4 #(
		.INIT('h004c)
	) name17154 (
		_w22881_,
		_w22885_,
		_w22882_,
		_w22879_,
		_w22981_
	);
	LUT2 #(
		.INIT('h8)
	) name17155 (
		_w22980_,
		_w22981_,
		_w22982_
	);
	LUT3 #(
		.INIT('h56)
	) name17156 (
		\u1_L1_reg[17]/NET0131 ,
		_w22979_,
		_w22982_,
		_w22983_
	);
	LUT4 #(
		.INIT('h3fd2)
	) name17157 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22984_
	);
	LUT4 #(
		.INIT('h0200)
	) name17158 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22985_
	);
	LUT4 #(
		.INIT('hab6f)
	) name17159 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22986_
	);
	LUT4 #(
		.INIT('h3120)
	) name17160 (
		_w22916_,
		_w22985_,
		_w22984_,
		_w22986_,
		_w22987_
	);
	LUT2 #(
		.INIT('h1)
	) name17161 (
		_w22909_,
		_w22987_,
		_w22988_
	);
	LUT4 #(
		.INIT('hcf6f)
	) name17162 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22989_
	);
	LUT2 #(
		.INIT('h2)
	) name17163 (
		_w22916_,
		_w22989_,
		_w22990_
	);
	LUT4 #(
		.INIT('h77dc)
	) name17164 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22991_
	);
	LUT2 #(
		.INIT('h1)
	) name17165 (
		_w22916_,
		_w22991_,
		_w22992_
	);
	LUT4 #(
		.INIT('h0102)
	) name17166 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w22993_
	);
	LUT3 #(
		.INIT('h01)
	) name17167 (
		_w22929_,
		_w22930_,
		_w22993_,
		_w22994_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name17168 (
		_w22909_,
		_w22992_,
		_w22990_,
		_w22994_,
		_w22995_
	);
	LUT4 #(
		.INIT('h4000)
	) name17169 (
		_w22913_,
		_w22911_,
		_w22912_,
		_w22916_,
		_w22996_
	);
	LUT2 #(
		.INIT('h1)
	) name17170 (
		_w22919_,
		_w22996_,
		_w22997_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name17171 (
		\u1_L1_reg[29]/NET0131 ,
		_w22995_,
		_w22988_,
		_w22997_,
		_w22998_
	);
	LUT4 #(
		.INIT('hc693)
	) name17172 (
		decrypt_pad,
		\u1_R1_reg[7]/NET0131 ,
		\u1_uk_K_r1_reg[12]/NET0131 ,
		\u1_uk_K_r1_reg[20]/NET0131 ,
		_w22999_
	);
	LUT4 #(
		.INIT('hc693)
	) name17173 (
		decrypt_pad,
		\u1_R1_reg[5]/NET0131 ,
		\u1_uk_K_r1_reg[27]/NET0131 ,
		\u1_uk_K_r1_reg[3]/NET0131 ,
		_w23000_
	);
	LUT4 #(
		.INIT('hc693)
	) name17174 (
		decrypt_pad,
		\u1_R1_reg[6]/NET0131 ,
		\u1_uk_K_r1_reg[18]/NET0131 ,
		\u1_uk_K_r1_reg[26]/NET0131 ,
		_w23001_
	);
	LUT2 #(
		.INIT('h2)
	) name17175 (
		_w23000_,
		_w23001_,
		_w23002_
	);
	LUT4 #(
		.INIT('hc963)
	) name17176 (
		decrypt_pad,
		\u1_R1_reg[8]/NET0131 ,
		\u1_uk_K_r1_reg[11]/NET0131 ,
		\u1_uk_K_r1_reg[3]/NET0131 ,
		_w23003_
	);
	LUT4 #(
		.INIT('hc963)
	) name17177 (
		decrypt_pad,
		\u1_R1_reg[4]/NET0131 ,
		\u1_uk_K_r1_reg[24]/NET0131 ,
		\u1_uk_K_r1_reg[48]/NET0131 ,
		_w23004_
	);
	LUT4 #(
		.INIT('hc693)
	) name17178 (
		decrypt_pad,
		\u1_R1_reg[9]/NET0131 ,
		\u1_uk_K_r1_reg[40]/NET0131 ,
		\u1_uk_K_r1_reg[48]/NET0131 ,
		_w23005_
	);
	LUT4 #(
		.INIT('h0800)
	) name17179 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23006_
	);
	LUT4 #(
		.INIT('he6ee)
	) name17180 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23007_
	);
	LUT4 #(
		.INIT('h4044)
	) name17181 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23008_
	);
	LUT4 #(
		.INIT('h3302)
	) name17182 (
		_w23003_,
		_w23002_,
		_w23007_,
		_w23008_,
		_w23009_
	);
	LUT4 #(
		.INIT('h0100)
	) name17183 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23010_
	);
	LUT4 #(
		.INIT('hf700)
	) name17184 (
		_w23004_,
		_w23000_,
		_w23001_,
		_w22999_,
		_w23011_
	);
	LUT2 #(
		.INIT('h4)
	) name17185 (
		_w23010_,
		_w23011_,
		_w23012_
	);
	LUT3 #(
		.INIT('h0e)
	) name17186 (
		_w22999_,
		_w23009_,
		_w23012_,
		_w23013_
	);
	LUT4 #(
		.INIT('h59fb)
	) name17187 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23014_
	);
	LUT2 #(
		.INIT('h1)
	) name17188 (
		_w22999_,
		_w23014_,
		_w23015_
	);
	LUT4 #(
		.INIT('h0034)
	) name17189 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23016_
	);
	LUT2 #(
		.INIT('h2)
	) name17190 (
		_w23005_,
		_w23001_,
		_w23017_
	);
	LUT4 #(
		.INIT('h0002)
	) name17191 (
		_w23005_,
		_w23000_,
		_w23001_,
		_w22999_,
		_w23018_
	);
	LUT4 #(
		.INIT('h4000)
	) name17192 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23019_
	);
	LUT4 #(
		.INIT('h0007)
	) name17193 (
		_w23006_,
		_w22999_,
		_w23018_,
		_w23019_,
		_w23020_
	);
	LUT4 #(
		.INIT('h5455)
	) name17194 (
		_w23003_,
		_w23015_,
		_w23016_,
		_w23020_,
		_w23021_
	);
	LUT4 #(
		.INIT('h0082)
	) name17195 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23022_
	);
	LUT4 #(
		.INIT('h8c00)
	) name17196 (
		_w23004_,
		_w23000_,
		_w23001_,
		_w22999_,
		_w23023_
	);
	LUT3 #(
		.INIT('ha8)
	) name17197 (
		_w23003_,
		_w23022_,
		_w23023_,
		_w23024_
	);
	LUT4 #(
		.INIT('h5556)
	) name17198 (
		\u1_L1_reg[2]/NET0131 ,
		_w23021_,
		_w23024_,
		_w23013_,
		_w23025_
	);
	LUT4 #(
		.INIT('hb9cf)
	) name17199 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w23026_
	);
	LUT4 #(
		.INIT('he63f)
	) name17200 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w23027_
	);
	LUT4 #(
		.INIT('h3120)
	) name17201 (
		_w22916_,
		_w22919_,
		_w23027_,
		_w23026_,
		_w23028_
	);
	LUT4 #(
		.INIT('h5fef)
	) name17202 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w23029_
	);
	LUT3 #(
		.INIT('ha2)
	) name17203 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w23030_
	);
	LUT4 #(
		.INIT('h4000)
	) name17204 (
		_w22913_,
		_w22910_,
		_w22912_,
		_w22916_,
		_w23031_
	);
	LUT4 #(
		.INIT('h0d00)
	) name17205 (
		_w22928_,
		_w23030_,
		_w23031_,
		_w23029_,
		_w23032_
	);
	LUT4 #(
		.INIT('hb600)
	) name17206 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w22916_,
		_w23033_
	);
	LUT4 #(
		.INIT('h007d)
	) name17207 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w22916_,
		_w23034_
	);
	LUT4 #(
		.INIT('h0001)
	) name17208 (
		_w22913_,
		_w22910_,
		_w22912_,
		_w22916_,
		_w23035_
	);
	LUT4 #(
		.INIT('h00fd)
	) name17209 (
		_w22913_,
		_w23034_,
		_w23033_,
		_w23035_,
		_w23036_
	);
	LUT4 #(
		.INIT('he400)
	) name17210 (
		_w22909_,
		_w23028_,
		_w23032_,
		_w23036_,
		_w23037_
	);
	LUT2 #(
		.INIT('h9)
	) name17211 (
		\u1_L1_reg[4]/NET0131 ,
		_w23037_,
		_w23038_
	);
	LUT4 #(
		.INIT('hc693)
	) name17212 (
		decrypt_pad,
		\u1_R1_reg[32]/NET0131 ,
		\u1_uk_K_r1_reg[28]/NET0131 ,
		\u1_uk_K_r1_reg[38]/NET0131 ,
		_w23039_
	);
	LUT4 #(
		.INIT('hc693)
	) name17213 (
		decrypt_pad,
		\u1_R1_reg[28]/NET0131 ,
		\u1_uk_K_r1_reg[37]/NET0131 ,
		\u1_uk_K_r1_reg[43]/NET0131 ,
		_w23040_
	);
	LUT4 #(
		.INIT('hc963)
	) name17214 (
		decrypt_pad,
		\u1_R1_reg[29]/NET0131 ,
		\u1_uk_K_r1_reg[15]/NET0131 ,
		\u1_uk_K_r1_reg[9]/NET0131 ,
		_w23041_
	);
	LUT4 #(
		.INIT('hc963)
	) name17215 (
		decrypt_pad,
		\u1_R1_reg[30]/NET0131 ,
		\u1_uk_K_r1_reg[16]/NET0131 ,
		\u1_uk_K_r1_reg[38]/NET0131 ,
		_w23042_
	);
	LUT4 #(
		.INIT('hc963)
	) name17216 (
		decrypt_pad,
		\u1_R1_reg[1]/NET0131 ,
		\u1_uk_K_r1_reg[0]/NET0131 ,
		\u1_uk_K_r1_reg[49]/NET0131 ,
		_w23043_
	);
	LUT4 #(
		.INIT('h0020)
	) name17217 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23044_
	);
	LUT4 #(
		.INIT('hc693)
	) name17218 (
		decrypt_pad,
		\u1_R1_reg[31]/P0001 ,
		\u1_uk_K_r1_reg[22]/NET0131 ,
		\u1_uk_K_r1_reg[28]/NET0131 ,
		_w23045_
	);
	LUT4 #(
		.INIT('hef00)
	) name17219 (
		_w23040_,
		_w23041_,
		_w23043_,
		_w23045_,
		_w23046_
	);
	LUT2 #(
		.INIT('h8)
	) name17220 (
		_w23041_,
		_w23043_,
		_w23047_
	);
	LUT3 #(
		.INIT('h0d)
	) name17221 (
		_w23040_,
		_w23042_,
		_w23045_,
		_w23048_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17222 (
		_w23044_,
		_w23046_,
		_w23047_,
		_w23048_,
		_w23049_
	);
	LUT4 #(
		.INIT('h0008)
	) name17223 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23050_
	);
	LUT4 #(
		.INIT('h7f7a)
	) name17224 (
		_w23040_,
		_w23041_,
		_w23043_,
		_w23045_,
		_w23051_
	);
	LUT3 #(
		.INIT('h31)
	) name17225 (
		_w23042_,
		_w23050_,
		_w23051_,
		_w23052_
	);
	LUT3 #(
		.INIT('h45)
	) name17226 (
		_w23039_,
		_w23049_,
		_w23052_,
		_w23053_
	);
	LUT4 #(
		.INIT('hf531)
	) name17227 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23054_
	);
	LUT3 #(
		.INIT('h02)
	) name17228 (
		_w23045_,
		_w23054_,
		_w23050_,
		_w23055_
	);
	LUT4 #(
		.INIT('h4000)
	) name17229 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23056_
	);
	LUT4 #(
		.INIT('h0001)
	) name17230 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23045_,
		_w23057_
	);
	LUT2 #(
		.INIT('h1)
	) name17231 (
		_w23056_,
		_w23057_,
		_w23058_
	);
	LUT3 #(
		.INIT('h8a)
	) name17232 (
		_w23039_,
		_w23055_,
		_w23058_,
		_w23059_
	);
	LUT4 #(
		.INIT('h0041)
	) name17233 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23060_
	);
	LUT4 #(
		.INIT('h1000)
	) name17234 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23061_
	);
	LUT4 #(
		.INIT('h0200)
	) name17235 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23062_
	);
	LUT4 #(
		.INIT('h0002)
	) name17236 (
		_w23045_,
		_w23061_,
		_w23060_,
		_w23062_,
		_w23063_
	);
	LUT4 #(
		.INIT('h0800)
	) name17237 (
		_w23039_,
		_w23040_,
		_w23041_,
		_w23042_,
		_w23064_
	);
	LUT3 #(
		.INIT('h01)
	) name17238 (
		_w23045_,
		_w23050_,
		_w23064_,
		_w23065_
	);
	LUT2 #(
		.INIT('h1)
	) name17239 (
		_w23063_,
		_w23065_,
		_w23066_
	);
	LUT4 #(
		.INIT('haaa9)
	) name17240 (
		\u1_L1_reg[5]/NET0131 ,
		_w23059_,
		_w23066_,
		_w23053_,
		_w23067_
	);
	LUT4 #(
		.INIT('hc963)
	) name17241 (
		decrypt_pad,
		\u1_R1_reg[16]/NET0131 ,
		\u1_uk_K_r1_reg[12]/NET0131 ,
		\u1_uk_K_r1_reg[4]/NET0131 ,
		_w23068_
	);
	LUT4 #(
		.INIT('hc963)
	) name17242 (
		decrypt_pad,
		\u1_R1_reg[15]/NET0131 ,
		\u1_uk_K_r1_reg[4]/NET0131 ,
		\u1_uk_K_r1_reg[53]/NET0131 ,
		_w23069_
	);
	LUT4 #(
		.INIT('hc693)
	) name17243 (
		decrypt_pad,
		\u1_R1_reg[13]/NET0131 ,
		\u1_uk_K_r1_reg[19]/NET0131 ,
		\u1_uk_K_r1_reg[27]/NET0131 ,
		_w23070_
	);
	LUT4 #(
		.INIT('hc693)
	) name17244 (
		decrypt_pad,
		\u1_R1_reg[12]/NET0131 ,
		\u1_uk_K_r1_reg[25]/NET0131 ,
		\u1_uk_K_r1_reg[33]/NET0131 ,
		_w23071_
	);
	LUT4 #(
		.INIT('hc963)
	) name17245 (
		decrypt_pad,
		\u1_R1_reg[17]/NET0131 ,
		\u1_uk_K_r1_reg[17]/NET0131 ,
		\u1_uk_K_r1_reg[41]/NET0131 ,
		_w23072_
	);
	LUT4 #(
		.INIT('hc693)
	) name17246 (
		decrypt_pad,
		\u1_R1_reg[14]/NET0131 ,
		\u1_uk_K_r1_reg[20]/NET0131 ,
		\u1_uk_K_r1_reg[53]/NET0131 ,
		_w23073_
	);
	LUT4 #(
		.INIT('h1000)
	) name17247 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23074_
	);
	LUT4 #(
		.INIT('heff3)
	) name17248 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23075_
	);
	LUT2 #(
		.INIT('h2)
	) name17249 (
		_w23069_,
		_w23075_,
		_w23076_
	);
	LUT4 #(
		.INIT('h8200)
	) name17250 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23077_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name17251 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23078_
	);
	LUT4 #(
		.INIT('h4044)
	) name17252 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23079_
	);
	LUT4 #(
		.INIT('h3332)
	) name17253 (
		_w23069_,
		_w23077_,
		_w23079_,
		_w23078_,
		_w23080_
	);
	LUT3 #(
		.INIT('h8a)
	) name17254 (
		_w23068_,
		_w23076_,
		_w23080_,
		_w23081_
	);
	LUT4 #(
		.INIT('hdacf)
	) name17255 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23082_
	);
	LUT2 #(
		.INIT('h4)
	) name17256 (
		_w23082_,
		_w23069_,
		_w23083_
	);
	LUT4 #(
		.INIT('h0009)
	) name17257 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23084_
	);
	LUT4 #(
		.INIT('h0040)
	) name17258 (
		_w23073_,
		_w23071_,
		_w23072_,
		_w23069_,
		_w23085_
	);
	LUT3 #(
		.INIT('h40)
	) name17259 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23086_
	);
	LUT2 #(
		.INIT('h1)
	) name17260 (
		_w23070_,
		_w23069_,
		_w23087_
	);
	LUT4 #(
		.INIT('h0001)
	) name17261 (
		_w23070_,
		_w23071_,
		_w23072_,
		_w23069_,
		_w23088_
	);
	LUT4 #(
		.INIT('h0001)
	) name17262 (
		_w23086_,
		_w23084_,
		_w23088_,
		_w23085_,
		_w23089_
	);
	LUT3 #(
		.INIT('h45)
	) name17263 (
		_w23068_,
		_w23083_,
		_w23089_,
		_w23090_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name17264 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23091_
	);
	LUT2 #(
		.INIT('h1)
	) name17265 (
		_w23069_,
		_w23091_,
		_w23092_
	);
	LUT2 #(
		.INIT('h8)
	) name17266 (
		_w23070_,
		_w23069_,
		_w23093_
	);
	LUT4 #(
		.INIT('h0800)
	) name17267 (
		_w23070_,
		_w23071_,
		_w23072_,
		_w23069_,
		_w23094_
	);
	LUT2 #(
		.INIT('h8)
	) name17268 (
		_w23073_,
		_w23069_,
		_w23095_
	);
	LUT4 #(
		.INIT('h0800)
	) name17269 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23069_,
		_w23096_
	);
	LUT3 #(
		.INIT('h0b)
	) name17270 (
		_w23073_,
		_w23094_,
		_w23096_,
		_w23097_
	);
	LUT2 #(
		.INIT('h4)
	) name17271 (
		_w23092_,
		_w23097_,
		_w23098_
	);
	LUT4 #(
		.INIT('h5655)
	) name17272 (
		\u1_L1_reg[10]/NET0131 ,
		_w23090_,
		_w23081_,
		_w23098_,
		_w23099_
	);
	LUT3 #(
		.INIT('h09)
	) name17273 (
		_w22945_,
		_w22943_,
		_w22944_,
		_w23100_
	);
	LUT4 #(
		.INIT('h0004)
	) name17274 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23101_
	);
	LUT3 #(
		.INIT('h27)
	) name17275 (
		_w22943_,
		_w22942_,
		_w22944_,
		_w23102_
	);
	LUT4 #(
		.INIT('h0031)
	) name17276 (
		_w22959_,
		_w23101_,
		_w23102_,
		_w23100_,
		_w23103_
	);
	LUT3 #(
		.INIT('h04)
	) name17277 (
		_w22945_,
		_w22941_,
		_w22942_,
		_w23104_
	);
	LUT4 #(
		.INIT('h2010)
	) name17278 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23105_
	);
	LUT3 #(
		.INIT('h08)
	) name17279 (
		_w22941_,
		_w22942_,
		_w22944_,
		_w23106_
	);
	LUT4 #(
		.INIT('h0001)
	) name17280 (
		_w22940_,
		_w22948_,
		_w23105_,
		_w23106_,
		_w23107_
	);
	LUT2 #(
		.INIT('h9)
	) name17281 (
		_w22945_,
		_w22941_,
		_w23108_
	);
	LUT4 #(
		.INIT('h4050)
	) name17282 (
		_w22943_,
		_w22941_,
		_w22942_,
		_w22944_,
		_w23109_
	);
	LUT4 #(
		.INIT('h0400)
	) name17283 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23110_
	);
	LUT4 #(
		.INIT('h2022)
	) name17284 (
		_w22940_,
		_w23110_,
		_w23108_,
		_w23109_,
		_w23111_
	);
	LUT4 #(
		.INIT('h0028)
	) name17285 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23112_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name17286 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23113_
	);
	LUT3 #(
		.INIT('h31)
	) name17287 (
		_w22944_,
		_w23112_,
		_w23113_,
		_w23114_
	);
	LUT4 #(
		.INIT('h0777)
	) name17288 (
		_w23103_,
		_w23107_,
		_w23111_,
		_w23114_,
		_w23115_
	);
	LUT2 #(
		.INIT('h6)
	) name17289 (
		\u1_L1_reg[12]/NET0131 ,
		_w23115_,
		_w23116_
	);
	LUT3 #(
		.INIT('h08)
	) name17290 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23117_
	);
	LUT4 #(
		.INIT('h00ef)
	) name17291 (
		_w23005_,
		_w23000_,
		_w23001_,
		_w22999_,
		_w23118_
	);
	LUT3 #(
		.INIT('h40)
	) name17292 (
		_w23004_,
		_w23005_,
		_w23001_,
		_w23119_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17293 (
		_w23005_,
		_w23000_,
		_w23001_,
		_w22999_,
		_w23120_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17294 (
		_w23117_,
		_w23118_,
		_w23119_,
		_w23120_,
		_w23121_
	);
	LUT4 #(
		.INIT('h0010)
	) name17295 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23122_
	);
	LUT4 #(
		.INIT('h0002)
	) name17296 (
		_w23003_,
		_w23018_,
		_w23019_,
		_w23122_,
		_w23123_
	);
	LUT2 #(
		.INIT('h4)
	) name17297 (
		_w23121_,
		_w23123_,
		_w23124_
	);
	LUT3 #(
		.INIT('h54)
	) name17298 (
		_w23004_,
		_w23000_,
		_w22999_,
		_w23125_
	);
	LUT2 #(
		.INIT('h8)
	) name17299 (
		_w23017_,
		_w23125_,
		_w23126_
	);
	LUT2 #(
		.INIT('h8)
	) name17300 (
		_w23004_,
		_w22999_,
		_w23127_
	);
	LUT3 #(
		.INIT('hb0)
	) name17301 (
		_w23005_,
		_w23000_,
		_w23001_,
		_w23128_
	);
	LUT3 #(
		.INIT('h15)
	) name17302 (
		_w23003_,
		_w23127_,
		_w23128_,
		_w23129_
	);
	LUT4 #(
		.INIT('h0400)
	) name17303 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23130_
	);
	LUT4 #(
		.INIT('h0002)
	) name17304 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23131_
	);
	LUT4 #(
		.INIT('h00ef)
	) name17305 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w22999_,
		_w23132_
	);
	LUT3 #(
		.INIT('h10)
	) name17306 (
		_w23131_,
		_w23130_,
		_w23132_,
		_w23133_
	);
	LUT3 #(
		.INIT('h40)
	) name17307 (
		_w23126_,
		_w23129_,
		_w23133_,
		_w23134_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name17308 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23135_
	);
	LUT3 #(
		.INIT('h09)
	) name17309 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23136_
	);
	LUT3 #(
		.INIT('h02)
	) name17310 (
		_w23004_,
		_w23005_,
		_w23001_,
		_w23137_
	);
	LUT4 #(
		.INIT('h0020)
	) name17311 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23138_
	);
	LUT3 #(
		.INIT('h02)
	) name17312 (
		_w22999_,
		_w23138_,
		_w23136_,
		_w23139_
	);
	LUT3 #(
		.INIT('h40)
	) name17313 (
		_w23126_,
		_w23129_,
		_w23139_,
		_w23140_
	);
	LUT4 #(
		.INIT('h001f)
	) name17314 (
		_w23124_,
		_w23134_,
		_w23135_,
		_w23140_,
		_w23141_
	);
	LUT2 #(
		.INIT('h9)
	) name17315 (
		\u1_L1_reg[13]/NET0131 ,
		_w23141_,
		_w23142_
	);
	LUT4 #(
		.INIT('h8b73)
	) name17316 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23143_
	);
	LUT2 #(
		.INIT('h2)
	) name17317 (
		_w14634_,
		_w23143_,
		_w23144_
	);
	LUT2 #(
		.INIT('h1)
	) name17318 (
		_w14635_,
		_w14634_,
		_w23145_
	);
	LUT3 #(
		.INIT('hf6)
	) name17319 (
		_w14637_,
		_w14638_,
		_w14636_,
		_w23146_
	);
	LUT2 #(
		.INIT('h2)
	) name17320 (
		_w23145_,
		_w23146_,
		_w23147_
	);
	LUT4 #(
		.INIT('h0200)
	) name17321 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23148_
	);
	LUT4 #(
		.INIT('h1000)
	) name17322 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23149_
	);
	LUT3 #(
		.INIT('hc4)
	) name17323 (
		_w14635_,
		_w14638_,
		_w14634_,
		_w23150_
	);
	LUT4 #(
		.INIT('hc400)
	) name17324 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23151_
	);
	LUT4 #(
		.INIT('h0045)
	) name17325 (
		_w23149_,
		_w23150_,
		_w23151_,
		_w23148_,
		_w23152_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name17326 (
		_w14633_,
		_w23147_,
		_w23144_,
		_w23152_,
		_w23153_
	);
	LUT4 #(
		.INIT('h0100)
	) name17327 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23154_
	);
	LUT4 #(
		.INIT('h9ed3)
	) name17328 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23155_
	);
	LUT4 #(
		.INIT('h77ac)
	) name17329 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23156_
	);
	LUT4 #(
		.INIT('h0810)
	) name17330 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23157_
	);
	LUT4 #(
		.INIT('h00d8)
	) name17331 (
		_w14634_,
		_w23156_,
		_w23155_,
		_w23157_,
		_w23158_
	);
	LUT4 #(
		.INIT('heffd)
	) name17332 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23159_
	);
	LUT4 #(
		.INIT('h0008)
	) name17333 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23160_
	);
	LUT4 #(
		.INIT('hffd7)
	) name17334 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23161_
	);
	LUT3 #(
		.INIT('hd8)
	) name17335 (
		_w14634_,
		_w23159_,
		_w23161_,
		_w23162_
	);
	LUT3 #(
		.INIT('he0)
	) name17336 (
		_w14633_,
		_w23158_,
		_w23162_,
		_w23163_
	);
	LUT3 #(
		.INIT('h65)
	) name17337 (
		\u1_L1_reg[14]/NET0131 ,
		_w23153_,
		_w23163_,
		_w23164_
	);
	LUT3 #(
		.INIT('h71)
	) name17338 (
		_w23073_,
		_w23071_,
		_w23072_,
		_w23165_
	);
	LUT4 #(
		.INIT('h008e)
	) name17339 (
		_w23073_,
		_w23071_,
		_w23072_,
		_w23069_,
		_w23166_
	);
	LUT3 #(
		.INIT('h10)
	) name17340 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23167_
	);
	LUT3 #(
		.INIT('hb0)
	) name17341 (
		_w23070_,
		_w23072_,
		_w23069_,
		_w23168_
	);
	LUT4 #(
		.INIT('h1011)
	) name17342 (
		_w23087_,
		_w23166_,
		_w23167_,
		_w23168_,
		_w23169_
	);
	LUT3 #(
		.INIT('h08)
	) name17343 (
		_w23073_,
		_w23071_,
		_w23072_,
		_w23170_
	);
	LUT4 #(
		.INIT('h0080)
	) name17344 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23171_
	);
	LUT4 #(
		.INIT('haaa2)
	) name17345 (
		_w23068_,
		_w23073_,
		_w23070_,
		_w23071_,
		_w23172_
	);
	LUT2 #(
		.INIT('h4)
	) name17346 (
		_w23171_,
		_w23172_,
		_w23173_
	);
	LUT3 #(
		.INIT('h04)
	) name17347 (
		_w23073_,
		_w23071_,
		_w23072_,
		_w23174_
	);
	LUT4 #(
		.INIT('h00bf)
	) name17348 (
		_w23070_,
		_w23071_,
		_w23072_,
		_w23069_,
		_w23175_
	);
	LUT4 #(
		.INIT('h0020)
	) name17349 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23176_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17350 (
		_w23073_,
		_w23071_,
		_w23072_,
		_w23069_,
		_w23177_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17351 (
		_w23174_,
		_w23175_,
		_w23176_,
		_w23177_,
		_w23178_
	);
	LUT4 #(
		.INIT('h8400)
	) name17352 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23179_
	);
	LUT4 #(
		.INIT('h0040)
	) name17353 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23180_
	);
	LUT3 #(
		.INIT('h01)
	) name17354 (
		_w23068_,
		_w23179_,
		_w23180_,
		_w23181_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17355 (
		_w23169_,
		_w23173_,
		_w23178_,
		_w23181_,
		_w23182_
	);
	LUT3 #(
		.INIT('h6d)
	) name17356 (
		_w23070_,
		_w23071_,
		_w23072_,
		_w23183_
	);
	LUT2 #(
		.INIT('h2)
	) name17357 (
		_w23095_,
		_w23183_,
		_w23184_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name17358 (
		_w23073_,
		_w23069_,
		_w23088_,
		_w23171_,
		_w23185_
	);
	LUT2 #(
		.INIT('h4)
	) name17359 (
		_w23184_,
		_w23185_,
		_w23186_
	);
	LUT3 #(
		.INIT('h65)
	) name17360 (
		\u1_L1_reg[1]/NET0131 ,
		_w23182_,
		_w23186_,
		_w23187_
	);
	LUT4 #(
		.INIT('hfcd3)
	) name17361 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w23188_
	);
	LUT4 #(
		.INIT('heffb)
	) name17362 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w23189_
	);
	LUT4 #(
		.INIT('h0233)
	) name17363 (
		_w22878_,
		_w22885_,
		_w23188_,
		_w23189_,
		_w23190_
	);
	LUT4 #(
		.INIT('h02a0)
	) name17364 (
		_w22885_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w23191_
	);
	LUT3 #(
		.INIT('h54)
	) name17365 (
		_w22897_,
		_w22903_,
		_w23191_,
		_w23192_
	);
	LUT3 #(
		.INIT('h8c)
	) name17366 (
		_w22881_,
		_w22885_,
		_w22879_,
		_w23193_
	);
	LUT2 #(
		.INIT('h8)
	) name17367 (
		_w22898_,
		_w23193_,
		_w23194_
	);
	LUT4 #(
		.INIT('h002a)
	) name17368 (
		_w22878_,
		_w22889_,
		_w22901_,
		_w22972_,
		_w23195_
	);
	LUT4 #(
		.INIT('h1554)
	) name17369 (
		_w22878_,
		_w22881_,
		_w22882_,
		_w22880_,
		_w23196_
	);
	LUT3 #(
		.INIT('h47)
	) name17370 (
		_w22881_,
		_w22882_,
		_w22880_,
		_w23197_
	);
	LUT3 #(
		.INIT('h07)
	) name17371 (
		_w22881_,
		_w22882_,
		_w22880_,
		_w23198_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name17372 (
		_w22885_,
		_w22879_,
		_w23197_,
		_w23198_,
		_w23199_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name17373 (
		_w23194_,
		_w23195_,
		_w23196_,
		_w23199_,
		_w23200_
	);
	LUT4 #(
		.INIT('haaa9)
	) name17374 (
		\u1_L1_reg[23]/NET0131 ,
		_w23192_,
		_w23200_,
		_w23190_,
		_w23201_
	);
	LUT4 #(
		.INIT('h5eff)
	) name17375 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23202_
	);
	LUT3 #(
		.INIT('hf6)
	) name17376 (
		_w23073_,
		_w23071_,
		_w23072_,
		_w23203_
	);
	LUT4 #(
		.INIT('hf578)
	) name17377 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23204_
	);
	LUT4 #(
		.INIT('hfc10)
	) name17378 (
		_w23070_,
		_w23069_,
		_w23202_,
		_w23204_,
		_w23205_
	);
	LUT2 #(
		.INIT('h2)
	) name17379 (
		_w23068_,
		_w23205_,
		_w23206_
	);
	LUT4 #(
		.INIT('h0400)
	) name17380 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23207_
	);
	LUT4 #(
		.INIT('hebef)
	) name17381 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23208_
	);
	LUT4 #(
		.INIT('h0455)
	) name17382 (
		_w23068_,
		_w23093_,
		_w23165_,
		_w23208_,
		_w23209_
	);
	LUT4 #(
		.INIT('hfdcc)
	) name17383 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23210_
	);
	LUT4 #(
		.INIT('h4004)
	) name17384 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23072_,
		_w23211_
	);
	LUT4 #(
		.INIT('h3301)
	) name17385 (
		_w23068_,
		_w23069_,
		_w23210_,
		_w23211_,
		_w23212_
	);
	LUT3 #(
		.INIT('heb)
	) name17386 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23213_
	);
	LUT2 #(
		.INIT('h8)
	) name17387 (
		_w23072_,
		_w23069_,
		_w23214_
	);
	LUT4 #(
		.INIT('h7077)
	) name17388 (
		_w23087_,
		_w23174_,
		_w23213_,
		_w23214_,
		_w23215_
	);
	LUT3 #(
		.INIT('h10)
	) name17389 (
		_w23212_,
		_w23209_,
		_w23215_,
		_w23216_
	);
	LUT3 #(
		.INIT('h65)
	) name17390 (
		\u1_L1_reg[26]/NET0131 ,
		_w23206_,
		_w23216_,
		_w23217_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name17391 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23218_
	);
	LUT2 #(
		.INIT('h2)
	) name17392 (
		_w22999_,
		_w23218_,
		_w23219_
	);
	LUT4 #(
		.INIT('h55f7)
	) name17393 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w22999_,
		_w23220_
	);
	LUT2 #(
		.INIT('h1)
	) name17394 (
		_w23001_,
		_w23220_,
		_w23221_
	);
	LUT4 #(
		.INIT('hbfae)
	) name17395 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23222_
	);
	LUT3 #(
		.INIT('h32)
	) name17396 (
		_w22999_,
		_w23130_,
		_w23222_,
		_w23223_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name17397 (
		_w23003_,
		_w23221_,
		_w23219_,
		_w23223_,
		_w23224_
	);
	LUT4 #(
		.INIT('hdaff)
	) name17398 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23225_
	);
	LUT2 #(
		.INIT('h1)
	) name17399 (
		_w22999_,
		_w23225_,
		_w23226_
	);
	LUT4 #(
		.INIT('h005b)
	) name17400 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w22999_,
		_w23227_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name17401 (
		_w22999_,
		_w23137_,
		_w23222_,
		_w23227_,
		_w23228_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name17402 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23229_
	);
	LUT4 #(
		.INIT('h2322)
	) name17403 (
		_w23003_,
		_w23226_,
		_w23228_,
		_w23229_,
		_w23230_
	);
	LUT3 #(
		.INIT('h65)
	) name17404 (
		\u1_L1_reg[28]/NET0131 ,
		_w23224_,
		_w23230_,
		_w23231_
	);
	LUT4 #(
		.INIT('h3eff)
	) name17405 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23232_
	);
	LUT4 #(
		.INIT('hf33b)
	) name17406 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23233_
	);
	LUT4 #(
		.INIT('hdfad)
	) name17407 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23234_
	);
	LUT4 #(
		.INIT('hd800)
	) name17408 (
		_w14634_,
		_w23232_,
		_w23233_,
		_w23234_,
		_w23235_
	);
	LUT4 #(
		.INIT('h0001)
	) name17409 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23236_
	);
	LUT4 #(
		.INIT('hf3fe)
	) name17410 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23237_
	);
	LUT3 #(
		.INIT('h10)
	) name17411 (
		_w14635_,
		_w14634_,
		_w14636_,
		_w23238_
	);
	LUT4 #(
		.INIT('h00c4)
	) name17412 (
		_w14634_,
		_w23161_,
		_w23237_,
		_w23238_,
		_w23239_
	);
	LUT4 #(
		.INIT('hdf9f)
	) name17413 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23240_
	);
	LUT4 #(
		.INIT('he4ee)
	) name17414 (
		_w14634_,
		_w23148_,
		_w23160_,
		_w23240_,
		_w23241_
	);
	LUT4 #(
		.INIT('h0d08)
	) name17415 (
		_w14633_,
		_w23239_,
		_w23241_,
		_w23235_,
		_w23242_
	);
	LUT2 #(
		.INIT('h9)
	) name17416 (
		\u1_L1_reg[8]/NET0131 ,
		_w23242_,
		_w23243_
	);
	LUT4 #(
		.INIT('h0002)
	) name17417 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23244_
	);
	LUT4 #(
		.INIT('h6673)
	) name17418 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23245_
	);
	LUT4 #(
		.INIT('h5054)
	) name17419 (
		_w23039_,
		_w23045_,
		_w23244_,
		_w23245_,
		_w23246_
	);
	LUT4 #(
		.INIT('h0040)
	) name17420 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23247_
	);
	LUT4 #(
		.INIT('h0040)
	) name17421 (
		_w23041_,
		_w23042_,
		_w23043_,
		_w23045_,
		_w23248_
	);
	LUT4 #(
		.INIT('h2000)
	) name17422 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23249_
	);
	LUT2 #(
		.INIT('h4)
	) name17423 (
		_w23041_,
		_w23045_,
		_w23250_
	);
	LUT4 #(
		.INIT('h0100)
	) name17424 (
		_w23040_,
		_w23041_,
		_w23043_,
		_w23045_,
		_w23251_
	);
	LUT3 #(
		.INIT('h08)
	) name17425 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23252_
	);
	LUT4 #(
		.INIT('h0001)
	) name17426 (
		_w23248_,
		_w23249_,
		_w23251_,
		_w23252_,
		_w23253_
	);
	LUT3 #(
		.INIT('h8a)
	) name17427 (
		_w23039_,
		_w23247_,
		_w23253_,
		_w23254_
	);
	LUT4 #(
		.INIT('h4100)
	) name17428 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23255_
	);
	LUT2 #(
		.INIT('h2)
	) name17429 (
		_w23045_,
		_w23255_,
		_w23256_
	);
	LUT4 #(
		.INIT('h0c04)
	) name17430 (
		_w23039_,
		_w23040_,
		_w23041_,
		_w23042_,
		_w23257_
	);
	LUT4 #(
		.INIT('h0400)
	) name17431 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23258_
	);
	LUT4 #(
		.INIT('h0001)
	) name17432 (
		_w23045_,
		_w23060_,
		_w23258_,
		_w23257_,
		_w23259_
	);
	LUT2 #(
		.INIT('h1)
	) name17433 (
		_w23256_,
		_w23259_,
		_w23260_
	);
	LUT4 #(
		.INIT('h5556)
	) name17434 (
		\u1_L1_reg[15]/P0001 ,
		_w23246_,
		_w23254_,
		_w23260_,
		_w23261_
	);
	LUT4 #(
		.INIT('h0040)
	) name17435 (
		_w23040_,
		_w23042_,
		_w23043_,
		_w23045_,
		_w23262_
	);
	LUT4 #(
		.INIT('hffde)
	) name17436 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23263_
	);
	LUT2 #(
		.INIT('h4)
	) name17437 (
		_w23262_,
		_w23263_,
		_w23264_
	);
	LUT4 #(
		.INIT('h0004)
	) name17438 (
		_w23040_,
		_w23041_,
		_w23043_,
		_w23045_,
		_w23265_
	);
	LUT4 #(
		.INIT('h4555)
	) name17439 (
		_w23039_,
		_w23040_,
		_w23041_,
		_w23042_,
		_w23266_
	);
	LUT2 #(
		.INIT('h4)
	) name17440 (
		_w23265_,
		_w23266_,
		_w23267_
	);
	LUT3 #(
		.INIT('h20)
	) name17441 (
		_w23040_,
		_w23042_,
		_w23043_,
		_w23268_
	);
	LUT3 #(
		.INIT('h4e)
	) name17442 (
		_w23041_,
		_w23042_,
		_w23043_,
		_w23269_
	);
	LUT2 #(
		.INIT('h8)
	) name17443 (
		_w23040_,
		_w23045_,
		_w23270_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name17444 (
		_w23250_,
		_w23268_,
		_w23269_,
		_w23270_,
		_w23271_
	);
	LUT3 #(
		.INIT('h80)
	) name17445 (
		_w23264_,
		_w23267_,
		_w23271_,
		_w23272_
	);
	LUT4 #(
		.INIT('hc480)
	) name17446 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23273_
	);
	LUT4 #(
		.INIT('hef00)
	) name17447 (
		_w23041_,
		_w23042_,
		_w23043_,
		_w23045_,
		_w23274_
	);
	LUT4 #(
		.INIT('h00fd)
	) name17448 (
		_w23040_,
		_w23042_,
		_w23043_,
		_w23045_,
		_w23275_
	);
	LUT4 #(
		.INIT('h8acf)
	) name17449 (
		_w23249_,
		_w23273_,
		_w23274_,
		_w23275_,
		_w23276_
	);
	LUT4 #(
		.INIT('h0190)
	) name17450 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23277_
	);
	LUT2 #(
		.INIT('h2)
	) name17451 (
		_w23039_,
		_w23277_,
		_w23278_
	);
	LUT2 #(
		.INIT('h4)
	) name17452 (
		_w23276_,
		_w23278_,
		_w23279_
	);
	LUT3 #(
		.INIT('h02)
	) name17453 (
		_w23040_,
		_w23042_,
		_w23045_,
		_w23280_
	);
	LUT4 #(
		.INIT('h0100)
	) name17454 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23045_,
		_w23281_
	);
	LUT3 #(
		.INIT('h07)
	) name17455 (
		_w23047_,
		_w23280_,
		_w23281_,
		_w23282_
	);
	LUT4 #(
		.INIT('ha955)
	) name17456 (
		\u1_L1_reg[21]/NET0131 ,
		_w23272_,
		_w23279_,
		_w23282_,
		_w23283_
	);
	LUT4 #(
		.INIT('h77fb)
	) name17457 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23284_
	);
	LUT2 #(
		.INIT('h2)
	) name17458 (
		_w23045_,
		_w23284_,
		_w23285_
	);
	LUT4 #(
		.INIT('h1054)
	) name17459 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23286_
	);
	LUT4 #(
		.INIT('h005d)
	) name17460 (
		_w23040_,
		_w23041_,
		_w23043_,
		_w23045_,
		_w23287_
	);
	LUT4 #(
		.INIT('hbcdf)
	) name17461 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23288_
	);
	LUT3 #(
		.INIT('hb0)
	) name17462 (
		_w23286_,
		_w23287_,
		_w23288_,
		_w23289_
	);
	LUT3 #(
		.INIT('h8a)
	) name17463 (
		_w23039_,
		_w23285_,
		_w23289_,
		_w23290_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17464 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23045_,
		_w23291_
	);
	LUT3 #(
		.INIT('h2d)
	) name17465 (
		_w23041_,
		_w23042_,
		_w23043_,
		_w23292_
	);
	LUT2 #(
		.INIT('h8)
	) name17466 (
		_w23291_,
		_w23292_,
		_w23293_
	);
	LUT4 #(
		.INIT('h0080)
	) name17467 (
		_w23040_,
		_w23042_,
		_w23043_,
		_w23045_,
		_w23294_
	);
	LUT3 #(
		.INIT('h01)
	) name17468 (
		_w23061_,
		_w23265_,
		_w23294_,
		_w23295_
	);
	LUT4 #(
		.INIT('h0400)
	) name17469 (
		_w23041_,
		_w23042_,
		_w23043_,
		_w23045_,
		_w23296_
	);
	LUT4 #(
		.INIT('hfdb7)
	) name17470 (
		_w23040_,
		_w23041_,
		_w23042_,
		_w23043_,
		_w23297_
	);
	LUT3 #(
		.INIT('h32)
	) name17471 (
		_w23045_,
		_w23296_,
		_w23297_,
		_w23298_
	);
	LUT4 #(
		.INIT('hba00)
	) name17472 (
		_w23039_,
		_w23293_,
		_w23295_,
		_w23298_,
		_w23299_
	);
	LUT3 #(
		.INIT('h65)
	) name17473 (
		\u1_L1_reg[27]/NET0131 ,
		_w23290_,
		_w23299_,
		_w23300_
	);
	LUT4 #(
		.INIT('h4000)
	) name17474 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23301_
	);
	LUT3 #(
		.INIT('h09)
	) name17475 (
		_w22945_,
		_w22941_,
		_w22942_,
		_w23302_
	);
	LUT4 #(
		.INIT('h2012)
	) name17476 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23303_
	);
	LUT4 #(
		.INIT('h00fb)
	) name17477 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22944_,
		_w23304_
	);
	LUT4 #(
		.INIT('h0189)
	) name17478 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23305_
	);
	LUT4 #(
		.INIT('hbf00)
	) name17479 (
		_w22945_,
		_w22941_,
		_w22942_,
		_w22944_,
		_w23306_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17480 (
		_w23303_,
		_w23304_,
		_w23305_,
		_w23306_,
		_w23307_
	);
	LUT3 #(
		.INIT('ha8)
	) name17481 (
		_w22940_,
		_w23301_,
		_w23307_,
		_w23308_
	);
	LUT4 #(
		.INIT('h79bf)
	) name17482 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23309_
	);
	LUT4 #(
		.INIT('h5057)
	) name17483 (
		_w22944_,
		_w22961_,
		_w23104_,
		_w23100_,
		_w23310_
	);
	LUT4 #(
		.INIT('h008c)
	) name17484 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22944_,
		_w23311_
	);
	LUT4 #(
		.INIT('h135f)
	) name17485 (
		_w22944_,
		_w22949_,
		_w22963_,
		_w23311_,
		_w23312_
	);
	LUT4 #(
		.INIT('hea00)
	) name17486 (
		_w22940_,
		_w23309_,
		_w23310_,
		_w23312_,
		_w23313_
	);
	LUT3 #(
		.INIT('h65)
	) name17487 (
		\u1_L1_reg[32]/NET0131 ,
		_w23308_,
		_w23313_,
		_w23314_
	);
	LUT3 #(
		.INIT('hb0)
	) name17488 (
		_w14635_,
		_w14637_,
		_w14636_,
		_w23315_
	);
	LUT4 #(
		.INIT('hf040)
	) name17489 (
		_w14637_,
		_w14638_,
		_w14634_,
		_w14636_,
		_w23316_
	);
	LUT4 #(
		.INIT('h0008)
	) name17490 (
		_w14637_,
		_w14638_,
		_w14634_,
		_w14636_,
		_w23317_
	);
	LUT4 #(
		.INIT('hbdff)
	) name17491 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23318_
	);
	LUT4 #(
		.INIT('h4500)
	) name17492 (
		_w23317_,
		_w23315_,
		_w23316_,
		_w23318_,
		_w23319_
	);
	LUT2 #(
		.INIT('h2)
	) name17493 (
		_w14633_,
		_w23319_,
		_w23320_
	);
	LUT4 #(
		.INIT('h7344)
	) name17494 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23321_
	);
	LUT4 #(
		.INIT('h080a)
	) name17495 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23322_
	);
	LUT4 #(
		.INIT('hcfbb)
	) name17496 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23323_
	);
	LUT4 #(
		.INIT('h3120)
	) name17497 (
		_w14634_,
		_w23322_,
		_w23323_,
		_w23321_,
		_w23324_
	);
	LUT3 #(
		.INIT('h02)
	) name17498 (
		_w14634_,
		_w23154_,
		_w23160_,
		_w23325_
	);
	LUT4 #(
		.INIT('h0800)
	) name17499 (
		_w14635_,
		_w14637_,
		_w14638_,
		_w14636_,
		_w23326_
	);
	LUT4 #(
		.INIT('h0001)
	) name17500 (
		_w14634_,
		_w23149_,
		_w23236_,
		_w23326_,
		_w23327_
	);
	LUT4 #(
		.INIT('heee0)
	) name17501 (
		_w14633_,
		_w23324_,
		_w23325_,
		_w23327_,
		_w23328_
	);
	LUT3 #(
		.INIT('h65)
	) name17502 (
		\u1_L1_reg[3]/NET0131 ,
		_w23320_,
		_w23328_,
		_w23329_
	);
	LUT4 #(
		.INIT('hc693)
	) name17503 (
		decrypt_pad,
		\u1_R1_reg[11]/NET0131 ,
		\u1_uk_K_r1_reg[55]/NET0131 ,
		\u1_uk_K_r1_reg[6]/NET0131 ,
		_w23330_
	);
	LUT4 #(
		.INIT('hc693)
	) name17504 (
		decrypt_pad,
		\u1_R1_reg[12]/NET0131 ,
		\u1_uk_K_r1_reg[13]/NET0131 ,
		\u1_uk_K_r1_reg[46]/NET0131 ,
		_w23331_
	);
	LUT4 #(
		.INIT('hc693)
	) name17505 (
		decrypt_pad,
		\u1_R1_reg[13]/NET0131 ,
		\u1_uk_K_r1_reg[26]/NET0131 ,
		\u1_uk_K_r1_reg[34]/NET0131 ,
		_w23332_
	);
	LUT4 #(
		.INIT('hc693)
	) name17506 (
		decrypt_pad,
		\u1_R1_reg[9]/NET0131 ,
		\u1_uk_K_r1_reg[46]/NET0131 ,
		\u1_uk_K_r1_reg[54]/NET0131 ,
		_w23333_
	);
	LUT4 #(
		.INIT('hc693)
	) name17507 (
		decrypt_pad,
		\u1_R1_reg[8]/NET0131 ,
		\u1_uk_K_r1_reg[17]/NET0131 ,
		\u1_uk_K_r1_reg[25]/NET0131 ,
		_w23334_
	);
	LUT4 #(
		.INIT('hc693)
	) name17508 (
		decrypt_pad,
		\u1_R1_reg[10]/NET0131 ,
		\u1_uk_K_r1_reg[54]/NET0131 ,
		\u1_uk_K_r1_reg[5]/NET0131 ,
		_w23335_
	);
	LUT4 #(
		.INIT('h95b5)
	) name17509 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23336_
	);
	LUT2 #(
		.INIT('h1)
	) name17510 (
		_w23332_,
		_w23334_,
		_w23337_
	);
	LUT4 #(
		.INIT('h0001)
	) name17511 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23338_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name17512 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23339_
	);
	LUT4 #(
		.INIT('h08cc)
	) name17513 (
		_w23331_,
		_w23330_,
		_w23336_,
		_w23339_,
		_w23340_
	);
	LUT2 #(
		.INIT('h8)
	) name17514 (
		_w23332_,
		_w23334_,
		_w23341_
	);
	LUT2 #(
		.INIT('h6)
	) name17515 (
		_w23332_,
		_w23334_,
		_w23342_
	);
	LUT4 #(
		.INIT('h000d)
	) name17516 (
		_w23330_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23343_
	);
	LUT4 #(
		.INIT('h0020)
	) name17517 (
		_w23330_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23344_
	);
	LUT4 #(
		.INIT('h4000)
	) name17518 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23345_
	);
	LUT4 #(
		.INIT('h0103)
	) name17519 (
		_w23342_,
		_w23344_,
		_w23345_,
		_w23343_,
		_w23346_
	);
	LUT3 #(
		.INIT('h20)
	) name17520 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23347_
	);
	LUT4 #(
		.INIT('h2000)
	) name17521 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23348_
	);
	LUT4 #(
		.INIT('h9990)
	) name17522 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23349_
	);
	LUT4 #(
		.INIT('h0990)
	) name17523 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23350_
	);
	LUT3 #(
		.INIT('h0b)
	) name17524 (
		_w23330_,
		_w23348_,
		_w23350_,
		_w23351_
	);
	LUT3 #(
		.INIT('h80)
	) name17525 (
		_w23331_,
		_w23333_,
		_w23335_,
		_w23352_
	);
	LUT3 #(
		.INIT('h80)
	) name17526 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23353_
	);
	LUT4 #(
		.INIT('h7b5b)
	) name17527 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23354_
	);
	LUT2 #(
		.INIT('h2)
	) name17528 (
		_w23331_,
		_w23330_,
		_w23355_
	);
	LUT4 #(
		.INIT('h7077)
	) name17529 (
		_w23337_,
		_w23352_,
		_w23354_,
		_w23355_,
		_w23356_
	);
	LUT4 #(
		.INIT('hea00)
	) name17530 (
		_w23331_,
		_w23346_,
		_w23351_,
		_w23356_,
		_w23357_
	);
	LUT3 #(
		.INIT('h65)
	) name17531 (
		\u1_L1_reg[6]/NET0131 ,
		_w23340_,
		_w23357_,
		_w23358_
	);
	LUT4 #(
		.INIT('h00a4)
	) name17532 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23359_
	);
	LUT2 #(
		.INIT('h2)
	) name17533 (
		_w22944_,
		_w23359_,
		_w23360_
	);
	LUT3 #(
		.INIT('h21)
	) name17534 (
		_w22943_,
		_w22941_,
		_w22942_,
		_w23361_
	);
	LUT3 #(
		.INIT('h48)
	) name17535 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w23362_
	);
	LUT4 #(
		.INIT('h00bf)
	) name17536 (
		_w22945_,
		_w22941_,
		_w22942_,
		_w22944_,
		_w23363_
	);
	LUT3 #(
		.INIT('h10)
	) name17537 (
		_w23362_,
		_w23361_,
		_w23363_,
		_w23364_
	);
	LUT4 #(
		.INIT('h6800)
	) name17538 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23365_
	);
	LUT2 #(
		.INIT('h2)
	) name17539 (
		_w22940_,
		_w23365_,
		_w23366_
	);
	LUT4 #(
		.INIT('h4800)
	) name17540 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22942_,
		_w23367_
	);
	LUT4 #(
		.INIT('hdf00)
	) name17541 (
		_w22945_,
		_w22943_,
		_w22941_,
		_w22944_,
		_w23368_
	);
	LUT4 #(
		.INIT('h5455)
	) name17542 (
		_w22940_,
		_w23302_,
		_w23367_,
		_w23368_,
		_w23369_
	);
	LUT4 #(
		.INIT('h001f)
	) name17543 (
		_w23360_,
		_w23364_,
		_w23366_,
		_w23369_,
		_w23370_
	);
	LUT2 #(
		.INIT('h4)
	) name17544 (
		_w22944_,
		_w23365_,
		_w23371_
	);
	LUT2 #(
		.INIT('h2)
	) name17545 (
		_w22940_,
		_w22944_,
		_w23372_
	);
	LUT4 #(
		.INIT('h00ba)
	) name17546 (
		_w22948_,
		_w22944_,
		_w23359_,
		_w23372_,
		_w23373_
	);
	LUT2 #(
		.INIT('h1)
	) name17547 (
		_w23371_,
		_w23373_,
		_w23374_
	);
	LUT3 #(
		.INIT('h65)
	) name17548 (
		\u1_L1_reg[7]/NET0131 ,
		_w23370_,
		_w23374_,
		_w23375_
	);
	LUT4 #(
		.INIT('hdc33)
	) name17549 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w23376_
	);
	LUT2 #(
		.INIT('h2)
	) name17550 (
		_w22885_,
		_w23376_,
		_w23377_
	);
	LUT4 #(
		.INIT('h0082)
	) name17551 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w23378_
	);
	LUT3 #(
		.INIT('h25)
	) name17552 (
		_w22882_,
		_w22879_,
		_w22880_,
		_w23379_
	);
	LUT4 #(
		.INIT('h0411)
	) name17553 (
		_w22885_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w23380_
	);
	LUT4 #(
		.INIT('h4000)
	) name17554 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w23381_
	);
	LUT3 #(
		.INIT('h01)
	) name17555 (
		_w23380_,
		_w23378_,
		_w23381_,
		_w23382_
	);
	LUT3 #(
		.INIT('h45)
	) name17556 (
		_w22878_,
		_w23377_,
		_w23382_,
		_w23383_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name17557 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w23384_
	);
	LUT2 #(
		.INIT('h1)
	) name17558 (
		_w22885_,
		_w23384_,
		_w23385_
	);
	LUT4 #(
		.INIT('h8228)
	) name17559 (
		_w22881_,
		_w22882_,
		_w22879_,
		_w22880_,
		_w23386_
	);
	LUT4 #(
		.INIT('h0013)
	) name17560 (
		_w22886_,
		_w22975_,
		_w23379_,
		_w23386_,
		_w23387_
	);
	LUT3 #(
		.INIT('h31)
	) name17561 (
		_w22878_,
		_w23385_,
		_w23387_,
		_w23388_
	);
	LUT3 #(
		.INIT('h65)
	) name17562 (
		\u1_L1_reg[9]/NET0131 ,
		_w23383_,
		_w23388_,
		_w23389_
	);
	LUT4 #(
		.INIT('h3dc3)
	) name17563 (
		_w23330_,
		_w23332_,
		_w23334_,
		_w23333_,
		_w23390_
	);
	LUT4 #(
		.INIT('h0110)
	) name17564 (
		_w23330_,
		_w23332_,
		_w23334_,
		_w23335_,
		_w23391_
	);
	LUT4 #(
		.INIT('h0074)
	) name17565 (
		_w23347_,
		_w23335_,
		_w23390_,
		_w23391_,
		_w23392_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name17566 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23393_
	);
	LUT4 #(
		.INIT('h2880)
	) name17567 (
		_w23330_,
		_w23332_,
		_w23334_,
		_w23333_,
		_w23394_
	);
	LUT4 #(
		.INIT('h0032)
	) name17568 (
		_w23330_,
		_w23338_,
		_w23393_,
		_w23394_,
		_w23395_
	);
	LUT4 #(
		.INIT('hbeff)
	) name17569 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23396_
	);
	LUT4 #(
		.INIT('h0400)
	) name17570 (
		_w23330_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23397_
	);
	LUT3 #(
		.INIT('h0d)
	) name17571 (
		_w23330_,
		_w23396_,
		_w23397_,
		_w23398_
	);
	LUT4 #(
		.INIT('he400)
	) name17572 (
		_w23331_,
		_w23395_,
		_w23392_,
		_w23398_,
		_w23399_
	);
	LUT2 #(
		.INIT('h9)
	) name17573 (
		\u1_L1_reg[16]/NET0131 ,
		_w23399_,
		_w23400_
	);
	LUT4 #(
		.INIT('h3400)
	) name17574 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w22999_,
		_w23401_
	);
	LUT4 #(
		.INIT('hfd75)
	) name17575 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23402_
	);
	LUT4 #(
		.INIT('h0a08)
	) name17576 (
		_w23003_,
		_w22999_,
		_w23010_,
		_w23402_,
		_w23403_
	);
	LUT4 #(
		.INIT('h0141)
	) name17577 (
		_w23004_,
		_w23000_,
		_w23001_,
		_w22999_,
		_w23404_
	);
	LUT4 #(
		.INIT('h8000)
	) name17578 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w22999_,
		_w23405_
	);
	LUT4 #(
		.INIT('hdffc)
	) name17579 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23406_
	);
	LUT4 #(
		.INIT('h0100)
	) name17580 (
		_w23003_,
		_w23006_,
		_w23405_,
		_w23406_,
		_w23407_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17581 (
		_w23401_,
		_w23403_,
		_w23404_,
		_w23407_,
		_w23408_
	);
	LUT4 #(
		.INIT('h0040)
	) name17582 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w22999_,
		_w23409_
	);
	LUT4 #(
		.INIT('h77ef)
	) name17583 (
		_w23004_,
		_w23005_,
		_w23000_,
		_w23001_,
		_w23410_
	);
	LUT3 #(
		.INIT('h31)
	) name17584 (
		_w22999_,
		_w23409_,
		_w23410_,
		_w23411_
	);
	LUT3 #(
		.INIT('h65)
	) name17585 (
		\u1_L1_reg[18]/NET0131 ,
		_w23408_,
		_w23411_,
		_w23412_
	);
	LUT2 #(
		.INIT('h4)
	) name17586 (
		_w23330_,
		_w23349_,
		_w23413_
	);
	LUT4 #(
		.INIT('h1dff)
	) name17587 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23414_
	);
	LUT2 #(
		.INIT('h2)
	) name17588 (
		_w23330_,
		_w23414_,
		_w23415_
	);
	LUT2 #(
		.INIT('h2)
	) name17589 (
		_w23330_,
		_w23335_,
		_w23416_
	);
	LUT3 #(
		.INIT('h0d)
	) name17590 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23417_
	);
	LUT4 #(
		.INIT('h0777)
	) name17591 (
		_w23342_,
		_w23343_,
		_w23416_,
		_w23417_,
		_w23418_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name17592 (
		_w23331_,
		_w23415_,
		_w23413_,
		_w23418_,
		_w23419_
	);
	LUT4 #(
		.INIT('he2cd)
	) name17593 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23420_
	);
	LUT4 #(
		.INIT('h0400)
	) name17594 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23421_
	);
	LUT4 #(
		.INIT('h5504)
	) name17595 (
		_w23331_,
		_w23330_,
		_w23420_,
		_w23421_,
		_w23422_
	);
	LUT4 #(
		.INIT('h0009)
	) name17596 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23423_
	);
	LUT4 #(
		.INIT('h9db6)
	) name17597 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23424_
	);
	LUT2 #(
		.INIT('h1)
	) name17598 (
		_w23331_,
		_w23330_,
		_w23425_
	);
	LUT2 #(
		.INIT('h4)
	) name17599 (
		_w23424_,
		_w23425_,
		_w23426_
	);
	LUT3 #(
		.INIT('hdb)
	) name17600 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23427_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name17601 (
		_w23330_,
		_w23335_,
		_w23353_,
		_w23427_,
		_w23428_
	);
	LUT3 #(
		.INIT('h10)
	) name17602 (
		_w23422_,
		_w23426_,
		_w23428_,
		_w23429_
	);
	LUT3 #(
		.INIT('h65)
	) name17603 (
		\u1_L1_reg[24]/NET0131 ,
		_w23419_,
		_w23429_,
		_w23430_
	);
	LUT4 #(
		.INIT('h0200)
	) name17604 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23431_
	);
	LUT3 #(
		.INIT('h01)
	) name17605 (
		_w23331_,
		_w23423_,
		_w23431_,
		_w23432_
	);
	LUT2 #(
		.INIT('h8)
	) name17606 (
		_w23334_,
		_w23335_,
		_w23433_
	);
	LUT4 #(
		.INIT('h73af)
	) name17607 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23434_
	);
	LUT4 #(
		.INIT('hdf53)
	) name17608 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23435_
	);
	LUT3 #(
		.INIT('hd8)
	) name17609 (
		_w23330_,
		_w23434_,
		_w23435_,
		_w23436_
	);
	LUT4 #(
		.INIT('heed9)
	) name17610 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23437_
	);
	LUT4 #(
		.INIT('h23ef)
	) name17611 (
		_w23332_,
		_w23334_,
		_w23333_,
		_w23335_,
		_w23438_
	);
	LUT4 #(
		.INIT('ha820)
	) name17612 (
		_w23331_,
		_w23330_,
		_w23438_,
		_w23437_,
		_w23439_
	);
	LUT3 #(
		.INIT('h07)
	) name17613 (
		_w23432_,
		_w23436_,
		_w23439_,
		_w23440_
	);
	LUT3 #(
		.INIT('h08)
	) name17614 (
		_w23330_,
		_w23332_,
		_w23333_,
		_w23441_
	);
	LUT2 #(
		.INIT('h8)
	) name17615 (
		_w23433_,
		_w23441_,
		_w23442_
	);
	LUT4 #(
		.INIT('h1000)
	) name17616 (
		_w23330_,
		_w23332_,
		_w23333_,
		_w23335_,
		_w23443_
	);
	LUT3 #(
		.INIT('h0b)
	) name17617 (
		_w23341_,
		_w23352_,
		_w23443_,
		_w23444_
	);
	LUT2 #(
		.INIT('h4)
	) name17618 (
		_w23442_,
		_w23444_,
		_w23445_
	);
	LUT3 #(
		.INIT('h9a)
	) name17619 (
		\u1_L1_reg[30]/NET0131 ,
		_w23440_,
		_w23445_,
		_w23446_
	);
	LUT4 #(
		.INIT('hc963)
	) name17620 (
		decrypt_pad,
		\u1_R0_reg[27]/NET0131 ,
		\u1_uk_K_r0_reg[45]/NET0131 ,
		\u1_uk_K_r0_reg[7]/NET0131 ,
		_w23447_
	);
	LUT4 #(
		.INIT('hc963)
	) name17621 (
		decrypt_pad,
		\u1_R0_reg[24]/NET0131 ,
		\u1_uk_K_r0_reg[43]/NET0131 ,
		\u1_uk_K_r0_reg[9]/NET0131 ,
		_w23448_
	);
	LUT4 #(
		.INIT('hc693)
	) name17622 (
		decrypt_pad,
		\u1_R0_reg[29]/NET0131 ,
		\u1_uk_K_r0_reg[45]/NET0131 ,
		\u1_uk_K_r0_reg[51]/NET0131 ,
		_w23449_
	);
	LUT4 #(
		.INIT('hc963)
	) name17623 (
		decrypt_pad,
		\u1_R0_reg[25]/NET0131 ,
		\u1_uk_K_r0_reg[23]/NET0131 ,
		\u1_uk_K_r0_reg[44]/NET0131 ,
		_w23450_
	);
	LUT4 #(
		.INIT('hc963)
	) name17624 (
		decrypt_pad,
		\u1_R0_reg[28]/NET0131 ,
		\u1_uk_K_r0_reg[28]/NET0131 ,
		\u1_uk_K_r0_reg[49]/NET0131 ,
		_w23451_
	);
	LUT4 #(
		.INIT('hc693)
	) name17625 (
		decrypt_pad,
		\u1_R0_reg[26]/NET0131 ,
		\u1_uk_K_r0_reg[29]/NET0131 ,
		\u1_uk_K_r0_reg[8]/NET0131 ,
		_w23452_
	);
	LUT2 #(
		.INIT('h4)
	) name17626 (
		_w23450_,
		_w23452_,
		_w23453_
	);
	LUT4 #(
		.INIT('hf47c)
	) name17627 (
		_w23451_,
		_w23449_,
		_w23450_,
		_w23452_,
		_w23454_
	);
	LUT4 #(
		.INIT('h0400)
	) name17628 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23455_
	);
	LUT4 #(
		.INIT('hf9ee)
	) name17629 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23456_
	);
	LUT4 #(
		.INIT('h08cc)
	) name17630 (
		_w23448_,
		_w23447_,
		_w23454_,
		_w23456_,
		_w23457_
	);
	LUT4 #(
		.INIT('h0100)
	) name17631 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23458_
	);
	LUT4 #(
		.INIT('h1ebf)
	) name17632 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23459_
	);
	LUT2 #(
		.INIT('h1)
	) name17633 (
		_w23447_,
		_w23459_,
		_w23460_
	);
	LUT2 #(
		.INIT('h6)
	) name17634 (
		_w23448_,
		_w23452_,
		_w23461_
	);
	LUT4 #(
		.INIT('h8008)
	) name17635 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23462_
	);
	LUT4 #(
		.INIT('hcfe5)
	) name17636 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23447_,
		_w23463_
	);
	LUT3 #(
		.INIT('h32)
	) name17637 (
		_w23452_,
		_w23462_,
		_w23463_,
		_w23464_
	);
	LUT3 #(
		.INIT('h45)
	) name17638 (
		_w23451_,
		_w23460_,
		_w23464_,
		_w23465_
	);
	LUT4 #(
		.INIT('h0082)
	) name17639 (
		_w23450_,
		_w23448_,
		_w23452_,
		_w23447_,
		_w23466_
	);
	LUT3 #(
		.INIT('h20)
	) name17640 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23467_
	);
	LUT4 #(
		.INIT('h0020)
	) name17641 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23468_
	);
	LUT4 #(
		.INIT('hf7d7)
	) name17642 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23469_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name17643 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23470_
	);
	LUT4 #(
		.INIT('h02aa)
	) name17644 (
		_w23451_,
		_w23447_,
		_w23469_,
		_w23470_,
		_w23471_
	);
	LUT2 #(
		.INIT('h1)
	) name17645 (
		_w23466_,
		_w23471_,
		_w23472_
	);
	LUT4 #(
		.INIT('h5655)
	) name17646 (
		\u1_L0_reg[22]/NET0131 ,
		_w23465_,
		_w23457_,
		_w23472_,
		_w23473_
	);
	LUT4 #(
		.INIT('hc963)
	) name17647 (
		decrypt_pad,
		\u1_R0_reg[24]/NET0131 ,
		\u1_uk_K_r0_reg[21]/NET0131 ,
		\u1_uk_K_r0_reg[42]/NET0131 ,
		_w23474_
	);
	LUT4 #(
		.INIT('hc693)
	) name17648 (
		decrypt_pad,
		\u1_R0_reg[22]/NET0131 ,
		\u1_uk_K_r0_reg[31]/NET0131 ,
		\u1_uk_K_r0_reg[37]/NET0131 ,
		_w23475_
	);
	LUT4 #(
		.INIT('hc963)
	) name17649 (
		decrypt_pad,
		\u1_R0_reg[20]/NET0131 ,
		\u1_uk_K_r0_reg[0]/NET0131 ,
		\u1_uk_K_r0_reg[21]/NET0131 ,
		_w23476_
	);
	LUT4 #(
		.INIT('hc963)
	) name17650 (
		decrypt_pad,
		\u1_R0_reg[21]/NET0131 ,
		\u1_uk_K_r0_reg[15]/NET0131 ,
		\u1_uk_K_r0_reg[36]/NET0131 ,
		_w23477_
	);
	LUT4 #(
		.INIT('hc963)
	) name17651 (
		decrypt_pad,
		\u1_R0_reg[25]/NET0131 ,
		\u1_uk_K_r0_reg[16]/NET0131 ,
		\u1_uk_K_r0_reg[37]/NET0131 ,
		_w23478_
	);
	LUT4 #(
		.INIT('ha280)
	) name17652 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23479_
	);
	LUT4 #(
		.INIT('hc693)
	) name17653 (
		decrypt_pad,
		\u1_R0_reg[23]/NET0131 ,
		\u1_uk_K_r0_reg[16]/NET0131 ,
		\u1_uk_K_r0_reg[50]/NET0131 ,
		_w23480_
	);
	LUT4 #(
		.INIT('h4555)
	) name17654 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23481_
	);
	LUT3 #(
		.INIT('h01)
	) name17655 (
		_w23480_,
		_w23481_,
		_w23479_,
		_w23482_
	);
	LUT4 #(
		.INIT('h0004)
	) name17656 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23483_
	);
	LUT4 #(
		.INIT('h1dfb)
	) name17657 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23484_
	);
	LUT2 #(
		.INIT('h1)
	) name17658 (
		_w23475_,
		_w23480_,
		_w23485_
	);
	LUT4 #(
		.INIT('h1000)
	) name17659 (
		_w23475_,
		_w23480_,
		_w23476_,
		_w23478_,
		_w23486_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name17660 (
		_w23480_,
		_w23477_,
		_w23484_,
		_w23486_,
		_w23487_
	);
	LUT3 #(
		.INIT('h8a)
	) name17661 (
		_w23474_,
		_w23482_,
		_w23487_,
		_w23488_
	);
	LUT3 #(
		.INIT('h8a)
	) name17662 (
		_w23476_,
		_w23478_,
		_w23477_,
		_w23489_
	);
	LUT3 #(
		.INIT('h54)
	) name17663 (
		_w23475_,
		_w23480_,
		_w23476_,
		_w23490_
	);
	LUT4 #(
		.INIT('h0020)
	) name17664 (
		_w23480_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23491_
	);
	LUT2 #(
		.INIT('h8)
	) name17665 (
		_w23475_,
		_w23480_,
		_w23492_
	);
	LUT4 #(
		.INIT('h0080)
	) name17666 (
		_w23475_,
		_w23480_,
		_w23476_,
		_w23477_,
		_w23493_
	);
	LUT4 #(
		.INIT('h1011)
	) name17667 (
		_w23491_,
		_w23493_,
		_w23489_,
		_w23490_,
		_w23494_
	);
	LUT4 #(
		.INIT('h0080)
	) name17668 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23495_
	);
	LUT4 #(
		.INIT('h0010)
	) name17669 (
		_w23475_,
		_w23480_,
		_w23476_,
		_w23478_,
		_w23496_
	);
	LUT4 #(
		.INIT('h1200)
	) name17670 (
		_w23475_,
		_w23480_,
		_w23476_,
		_w23477_,
		_w23497_
	);
	LUT3 #(
		.INIT('h01)
	) name17671 (
		_w23495_,
		_w23496_,
		_w23497_,
		_w23498_
	);
	LUT3 #(
		.INIT('h15)
	) name17672 (
		_w23474_,
		_w23494_,
		_w23498_,
		_w23499_
	);
	LUT4 #(
		.INIT('hfbdf)
	) name17673 (
		_w23480_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23500_
	);
	LUT2 #(
		.INIT('h1)
	) name17674 (
		_w23475_,
		_w23500_,
		_w23501_
	);
	LUT3 #(
		.INIT('h01)
	) name17675 (
		_w23476_,
		_w23478_,
		_w23477_,
		_w23502_
	);
	LUT4 #(
		.INIT('h7e7f)
	) name17676 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23503_
	);
	LUT4 #(
		.INIT('hef23)
	) name17677 (
		_w23475_,
		_w23480_,
		_w23502_,
		_w23503_,
		_w23504_
	);
	LUT2 #(
		.INIT('h4)
	) name17678 (
		_w23501_,
		_w23504_,
		_w23505_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name17679 (
		\u1_L0_reg[11]/NET0131 ,
		_w23488_,
		_w23499_,
		_w23505_,
		_w23506_
	);
	LUT4 #(
		.INIT('hc963)
	) name17680 (
		decrypt_pad,
		\u1_R0_reg[15]/NET0131 ,
		\u1_uk_K_r0_reg[18]/NET0131 ,
		\u1_uk_K_r0_reg[39]/NET0131 ,
		_w23507_
	);
	LUT4 #(
		.INIT('hc963)
	) name17681 (
		decrypt_pad,
		\u1_R0_reg[13]/NET0131 ,
		\u1_uk_K_r0_reg[41]/NET0131 ,
		\u1_uk_K_r0_reg[5]/NET0131 ,
		_w23508_
	);
	LUT4 #(
		.INIT('hc693)
	) name17682 (
		decrypt_pad,
		\u1_R0_reg[12]/NET0131 ,
		\u1_uk_K_r0_reg[11]/NET0131 ,
		\u1_uk_K_r0_reg[47]/NET0131 ,
		_w23509_
	);
	LUT4 #(
		.INIT('hc963)
	) name17683 (
		decrypt_pad,
		\u1_R0_reg[14]/NET0131 ,
		\u1_uk_K_r0_reg[10]/NET0131 ,
		\u1_uk_K_r0_reg[6]/NET0131 ,
		_w23510_
	);
	LUT4 #(
		.INIT('hc693)
	) name17684 (
		decrypt_pad,
		\u1_R0_reg[17]/NET0131 ,
		\u1_uk_K_r0_reg[27]/NET0131 ,
		\u1_uk_K_r0_reg[6]/NET0131 ,
		_w23511_
	);
	LUT4 #(
		.INIT('h0200)
	) name17685 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23512_
	);
	LUT2 #(
		.INIT('h1)
	) name17686 (
		_w23507_,
		_w23512_,
		_w23513_
	);
	LUT3 #(
		.INIT('h01)
	) name17687 (
		_w23508_,
		_w23509_,
		_w23511_,
		_w23514_
	);
	LUT4 #(
		.INIT('h0001)
	) name17688 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23515_
	);
	LUT4 #(
		.INIT('h0040)
	) name17689 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23516_
	);
	LUT4 #(
		.INIT('h0008)
	) name17690 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23517_
	);
	LUT4 #(
		.INIT('h0002)
	) name17691 (
		_w23507_,
		_w23516_,
		_w23517_,
		_w23515_,
		_w23518_
	);
	LUT2 #(
		.INIT('h1)
	) name17692 (
		_w23513_,
		_w23518_,
		_w23519_
	);
	LUT3 #(
		.INIT('h10)
	) name17693 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23520_
	);
	LUT2 #(
		.INIT('h1)
	) name17694 (
		_w23507_,
		_w23511_,
		_w23521_
	);
	LUT4 #(
		.INIT('hc963)
	) name17695 (
		decrypt_pad,
		\u1_R0_reg[16]/NET0131 ,
		\u1_uk_K_r0_reg[26]/NET0131 ,
		\u1_uk_K_r0_reg[47]/NET0131 ,
		_w23522_
	);
	LUT2 #(
		.INIT('h9)
	) name17696 (
		_w23508_,
		_w23509_,
		_w23523_
	);
	LUT2 #(
		.INIT('h1)
	) name17697 (
		_w23507_,
		_w23510_,
		_w23524_
	);
	LUT4 #(
		.INIT('h0014)
	) name17698 (
		_w23507_,
		_w23508_,
		_w23509_,
		_w23510_,
		_w23525_
	);
	LUT4 #(
		.INIT('h0222)
	) name17699 (
		_w23522_,
		_w23525_,
		_w23520_,
		_w23521_,
		_w23526_
	);
	LUT4 #(
		.INIT('h7dff)
	) name17700 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23527_
	);
	LUT4 #(
		.INIT('h0280)
	) name17701 (
		_w23507_,
		_w23508_,
		_w23509_,
		_w23511_,
		_w23528_
	);
	LUT2 #(
		.INIT('h2)
	) name17702 (
		_w23527_,
		_w23528_,
		_w23529_
	);
	LUT4 #(
		.INIT('h2aa8)
	) name17703 (
		_w23507_,
		_w23508_,
		_w23509_,
		_w23511_,
		_w23530_
	);
	LUT3 #(
		.INIT('h08)
	) name17704 (
		_w23509_,
		_w23510_,
		_w23511_,
		_w23531_
	);
	LUT3 #(
		.INIT('h45)
	) name17705 (
		_w23507_,
		_w23508_,
		_w23511_,
		_w23532_
	);
	LUT3 #(
		.INIT('h45)
	) name17706 (
		_w23530_,
		_w23531_,
		_w23532_,
		_w23533_
	);
	LUT4 #(
		.INIT('hffde)
	) name17707 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23534_
	);
	LUT4 #(
		.INIT('h0800)
	) name17708 (
		_w23507_,
		_w23508_,
		_w23509_,
		_w23510_,
		_w23535_
	);
	LUT4 #(
		.INIT('h0400)
	) name17709 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23536_
	);
	LUT4 #(
		.INIT('h0004)
	) name17710 (
		_w23522_,
		_w23534_,
		_w23536_,
		_w23535_,
		_w23537_
	);
	LUT4 #(
		.INIT('h7077)
	) name17711 (
		_w23526_,
		_w23529_,
		_w23533_,
		_w23537_,
		_w23538_
	);
	LUT3 #(
		.INIT('h56)
	) name17712 (
		\u1_L0_reg[20]/NET0131 ,
		_w23519_,
		_w23538_,
		_w23539_
	);
	LUT4 #(
		.INIT('hc693)
	) name17713 (
		decrypt_pad,
		\u1_R0_reg[32]/NET0131 ,
		\u1_uk_K_r0_reg[14]/NET0131 ,
		\u1_uk_K_r0_reg[52]/P0001 ,
		_w23540_
	);
	LUT4 #(
		.INIT('hc963)
	) name17714 (
		decrypt_pad,
		\u1_R0_reg[30]/NET0131 ,
		\u1_uk_K_r0_reg[30]/NET0131 ,
		\u1_uk_K_r0_reg[51]/NET0131 ,
		_w23541_
	);
	LUT4 #(
		.INIT('hc693)
	) name17715 (
		decrypt_pad,
		\u1_R0_reg[28]/NET0131 ,
		\u1_uk_K_r0_reg[23]/NET0131 ,
		\u1_uk_K_r0_reg[2]/NET0131 ,
		_w23542_
	);
	LUT4 #(
		.INIT('hc963)
	) name17716 (
		decrypt_pad,
		\u1_R0_reg[1]/NET0131 ,
		\u1_uk_K_r0_reg[14]/NET0131 ,
		\u1_uk_K_r0_reg[35]/NET0131 ,
		_w23543_
	);
	LUT4 #(
		.INIT('hc963)
	) name17717 (
		decrypt_pad,
		\u1_R0_reg[29]/NET0131 ,
		\u1_uk_K_r0_reg[29]/NET0131 ,
		\u1_uk_K_r0_reg[50]/NET0131 ,
		_w23544_
	);
	LUT4 #(
		.INIT('h0800)
	) name17718 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23545_
	);
	LUT4 #(
		.INIT('hc963)
	) name17719 (
		decrypt_pad,
		\u1_R0_reg[31]/P0001 ,
		\u1_uk_K_r0_reg[42]/NET0131 ,
		\u1_uk_K_r0_reg[8]/NET0131 ,
		_w23546_
	);
	LUT4 #(
		.INIT('h4555)
	) name17720 (
		_w23546_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23547_
	);
	LUT4 #(
		.INIT('h4554)
	) name17721 (
		_w23546_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23548_
	);
	LUT2 #(
		.INIT('h2)
	) name17722 (
		_w23542_,
		_w23541_,
		_w23549_
	);
	LUT2 #(
		.INIT('h4)
	) name17723 (
		_w23543_,
		_w23544_,
		_w23550_
	);
	LUT4 #(
		.INIT('h070d)
	) name17724 (
		_w23546_,
		_w23549_,
		_w23548_,
		_w23550_,
		_w23551_
	);
	LUT3 #(
		.INIT('ha8)
	) name17725 (
		_w23540_,
		_w23545_,
		_w23551_,
		_w23552_
	);
	LUT4 #(
		.INIT('h1000)
	) name17726 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23553_
	);
	LUT4 #(
		.INIT('haaa2)
	) name17727 (
		_w23546_,
		_w23543_,
		_w23544_,
		_w23542_,
		_w23554_
	);
	LUT3 #(
		.INIT('h10)
	) name17728 (
		_w23543_,
		_w23542_,
		_w23541_,
		_w23555_
	);
	LUT3 #(
		.INIT('h15)
	) name17729 (
		_w23546_,
		_w23543_,
		_w23544_,
		_w23556_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17730 (
		_w23553_,
		_w23554_,
		_w23555_,
		_w23556_,
		_w23557_
	);
	LUT3 #(
		.INIT('h04)
	) name17731 (
		_w23546_,
		_w23542_,
		_w23541_,
		_w23558_
	);
	LUT3 #(
		.INIT('h2a)
	) name17732 (
		_w23543_,
		_w23542_,
		_w23541_,
		_w23559_
	);
	LUT4 #(
		.INIT('h8040)
	) name17733 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23560_
	);
	LUT2 #(
		.INIT('h1)
	) name17734 (
		_w23558_,
		_w23560_,
		_w23561_
	);
	LUT3 #(
		.INIT('h51)
	) name17735 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23562_
	);
	LUT4 #(
		.INIT('hae22)
	) name17736 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23563_
	);
	LUT4 #(
		.INIT('h0420)
	) name17737 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23564_
	);
	LUT4 #(
		.INIT('h0200)
	) name17738 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23565_
	);
	LUT4 #(
		.INIT('h0001)
	) name17739 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23566_
	);
	LUT4 #(
		.INIT('hf9de)
	) name17740 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23567_
	);
	LUT4 #(
		.INIT('h31f5)
	) name17741 (
		_w23546_,
		_w23558_,
		_w23567_,
		_w23550_,
		_w23568_
	);
	LUT4 #(
		.INIT('hba00)
	) name17742 (
		_w23540_,
		_w23557_,
		_w23561_,
		_w23568_,
		_w23569_
	);
	LUT3 #(
		.INIT('h9a)
	) name17743 (
		\u1_L0_reg[5]/NET0131 ,
		_w23552_,
		_w23569_,
		_w23570_
	);
	LUT4 #(
		.INIT('hc693)
	) name17744 (
		decrypt_pad,
		\u1_R0_reg[4]/NET0131 ,
		\u1_uk_K_r0_reg[20]/NET0131 ,
		\u1_uk_K_r0_reg[24]/NET0131 ,
		_w23571_
	);
	LUT4 #(
		.INIT('hc693)
	) name17745 (
		decrypt_pad,
		\u1_R0_reg[3]/NET0131 ,
		\u1_uk_K_r0_reg[10]/NET0131 ,
		\u1_uk_K_r0_reg[46]/NET0131 ,
		_w23572_
	);
	LUT4 #(
		.INIT('hc693)
	) name17746 (
		decrypt_pad,
		\u1_R0_reg[1]/NET0131 ,
		\u1_uk_K_r0_reg[18]/NET0131 ,
		\u1_uk_K_r0_reg[54]/NET0131 ,
		_w23573_
	);
	LUT4 #(
		.INIT('hc963)
	) name17747 (
		decrypt_pad,
		\u1_R0_reg[5]/NET0131 ,
		\u1_uk_K_r0_reg[27]/NET0131 ,
		\u1_uk_K_r0_reg[48]/NET0131 ,
		_w23574_
	);
	LUT4 #(
		.INIT('hc963)
	) name17748 (
		decrypt_pad,
		\u1_R0_reg[2]/NET0131 ,
		\u1_uk_K_r0_reg[12]/NET0131 ,
		\u1_uk_K_r0_reg[33]/NET0131 ,
		_w23575_
	);
	LUT4 #(
		.INIT('hc963)
	) name17749 (
		decrypt_pad,
		\u1_R0_reg[32]/NET0131 ,
		\u1_uk_K_r0_reg[33]/NET0131 ,
		\u1_uk_K_r0_reg[54]/NET0131 ,
		_w23576_
	);
	LUT4 #(
		.INIT('hf0dd)
	) name17750 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23577_
	);
	LUT2 #(
		.INIT('h2)
	) name17751 (
		_w23572_,
		_w23577_,
		_w23578_
	);
	LUT4 #(
		.INIT('hafac)
	) name17752 (
		_w23572_,
		_w23575_,
		_w23573_,
		_w23574_,
		_w23579_
	);
	LUT2 #(
		.INIT('h2)
	) name17753 (
		_w23572_,
		_w23575_,
		_w23580_
	);
	LUT3 #(
		.INIT('hd0)
	) name17754 (
		_w23572_,
		_w23575_,
		_w23573_,
		_w23581_
	);
	LUT3 #(
		.INIT('h32)
	) name17755 (
		_w23575_,
		_w23576_,
		_w23574_,
		_w23582_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name17756 (
		_w23576_,
		_w23579_,
		_w23581_,
		_w23582_,
		_w23583_
	);
	LUT3 #(
		.INIT('h8a)
	) name17757 (
		_w23571_,
		_w23578_,
		_w23583_,
		_w23584_
	);
	LUT4 #(
		.INIT('hefe6)
	) name17758 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23585_
	);
	LUT2 #(
		.INIT('h1)
	) name17759 (
		_w23572_,
		_w23585_,
		_w23586_
	);
	LUT2 #(
		.INIT('h1)
	) name17760 (
		_w23576_,
		_w23574_,
		_w23587_
	);
	LUT3 #(
		.INIT('h48)
	) name17761 (
		_w23576_,
		_w23573_,
		_w23574_,
		_w23588_
	);
	LUT4 #(
		.INIT('h73cf)
	) name17762 (
		_w23572_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23589_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name17763 (
		_w23572_,
		_w23575_,
		_w23588_,
		_w23589_,
		_w23590_
	);
	LUT3 #(
		.INIT('h45)
	) name17764 (
		_w23571_,
		_w23586_,
		_w23590_,
		_w23591_
	);
	LUT4 #(
		.INIT('h7daf)
	) name17765 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23592_
	);
	LUT2 #(
		.INIT('h1)
	) name17766 (
		_w23572_,
		_w23592_,
		_w23593_
	);
	LUT4 #(
		.INIT('h0020)
	) name17767 (
		_w23572_,
		_w23575_,
		_w23576_,
		_w23573_,
		_w23594_
	);
	LUT3 #(
		.INIT('h08)
	) name17768 (
		_w23572_,
		_w23575_,
		_w23573_,
		_w23595_
	);
	LUT3 #(
		.INIT('h15)
	) name17769 (
		_w23594_,
		_w23587_,
		_w23595_,
		_w23596_
	);
	LUT2 #(
		.INIT('h4)
	) name17770 (
		_w23593_,
		_w23596_,
		_w23597_
	);
	LUT4 #(
		.INIT('h5655)
	) name17771 (
		\u1_L0_reg[31]/NET0131 ,
		_w23591_,
		_w23584_,
		_w23597_,
		_w23598_
	);
	LUT4 #(
		.INIT('hf7d6)
	) name17772 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23599_
	);
	LUT3 #(
		.INIT('h20)
	) name17773 (
		_w23509_,
		_w23510_,
		_w23511_,
		_w23600_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17774 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23601_
	);
	LUT4 #(
		.INIT('haba1)
	) name17775 (
		_w23507_,
		_w23514_,
		_w23600_,
		_w23601_,
		_w23602_
	);
	LUT3 #(
		.INIT('h15)
	) name17776 (
		_w23522_,
		_w23599_,
		_w23602_,
		_w23603_
	);
	LUT4 #(
		.INIT('hfd3b)
	) name17777 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23604_
	);
	LUT4 #(
		.INIT('h9000)
	) name17778 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23605_
	);
	LUT4 #(
		.INIT('hfbdd)
	) name17779 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23606_
	);
	LUT4 #(
		.INIT('h3120)
	) name17780 (
		_w23507_,
		_w23605_,
		_w23606_,
		_w23604_,
		_w23607_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name17781 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23608_
	);
	LUT4 #(
		.INIT('h0702)
	) name17782 (
		_w23507_,
		_w23517_,
		_w23535_,
		_w23608_,
		_w23609_
	);
	LUT3 #(
		.INIT('hd0)
	) name17783 (
		_w23522_,
		_w23607_,
		_w23609_,
		_w23610_
	);
	LUT3 #(
		.INIT('h65)
	) name17784 (
		\u1_L0_reg[10]/NET0131 ,
		_w23603_,
		_w23610_,
		_w23611_
	);
	LUT3 #(
		.INIT('h07)
	) name17785 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23612_
	);
	LUT3 #(
		.INIT('h4c)
	) name17786 (
		_w23448_,
		_w23452_,
		_w23447_,
		_w23613_
	);
	LUT3 #(
		.INIT('h09)
	) name17787 (
		_w23449_,
		_w23450_,
		_w23447_,
		_w23614_
	);
	LUT4 #(
		.INIT('h5514)
	) name17788 (
		_w23451_,
		_w23449_,
		_w23450_,
		_w23447_,
		_w23615_
	);
	LUT3 #(
		.INIT('hb0)
	) name17789 (
		_w23612_,
		_w23613_,
		_w23615_,
		_w23616_
	);
	LUT4 #(
		.INIT('h2104)
	) name17790 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23617_
	);
	LUT3 #(
		.INIT('h04)
	) name17791 (
		_w23449_,
		_w23448_,
		_w23452_,
		_w23618_
	);
	LUT3 #(
		.INIT('h20)
	) name17792 (
		_w23449_,
		_w23448_,
		_w23447_,
		_w23619_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name17793 (
		_w23449_,
		_w23448_,
		_w23452_,
		_w23447_,
		_w23620_
	);
	LUT3 #(
		.INIT('h32)
	) name17794 (
		_w23450_,
		_w23617_,
		_w23620_,
		_w23621_
	);
	LUT4 #(
		.INIT('h0008)
	) name17795 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23622_
	);
	LUT4 #(
		.INIT('h0002)
	) name17796 (
		_w23451_,
		_w23468_,
		_w23455_,
		_w23622_,
		_w23623_
	);
	LUT3 #(
		.INIT('hb9)
	) name17797 (
		_w23449_,
		_w23448_,
		_w23447_,
		_w23624_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name17798 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23625_
	);
	LUT4 #(
		.INIT('hf351)
	) name17799 (
		_w23447_,
		_w23453_,
		_w23624_,
		_w23625_,
		_w23626_
	);
	LUT4 #(
		.INIT('h0777)
	) name17800 (
		_w23616_,
		_w23621_,
		_w23623_,
		_w23626_,
		_w23627_
	);
	LUT2 #(
		.INIT('h6)
	) name17801 (
		\u1_L0_reg[12]/NET0131 ,
		_w23627_,
		_w23628_
	);
	LUT4 #(
		.INIT('hc693)
	) name17802 (
		decrypt_pad,
		\u1_R0_reg[20]/NET0131 ,
		\u1_uk_K_r0_reg[30]/NET0131 ,
		\u1_uk_K_r0_reg[9]/NET0131 ,
		_w23629_
	);
	LUT4 #(
		.INIT('hc693)
	) name17803 (
		decrypt_pad,
		\u1_R0_reg[19]/NET0131 ,
		\u1_uk_K_r0_reg[15]/NET0131 ,
		\u1_uk_K_r0_reg[49]/NET0131 ,
		_w23630_
	);
	LUT4 #(
		.INIT('hc693)
	) name17804 (
		decrypt_pad,
		\u1_R0_reg[21]/NET0131 ,
		\u1_uk_K_r0_reg[0]/NET0131 ,
		\u1_uk_K_r0_reg[38]/NET0131 ,
		_w23631_
	);
	LUT4 #(
		.INIT('hc693)
	) name17805 (
		decrypt_pad,
		\u1_R0_reg[17]/NET0131 ,
		\u1_uk_K_r0_reg[38]/NET0131 ,
		\u1_uk_K_r0_reg[44]/NET0131 ,
		_w23632_
	);
	LUT4 #(
		.INIT('hc963)
	) name17806 (
		decrypt_pad,
		\u1_R0_reg[16]/NET0131 ,
		\u1_uk_K_r0_reg[22]/NET0131 ,
		\u1_uk_K_r0_reg[43]/NET0131 ,
		_w23633_
	);
	LUT4 #(
		.INIT('hc693)
	) name17807 (
		decrypt_pad,
		\u1_R0_reg[18]/NET0131 ,
		\u1_uk_K_r0_reg[28]/NET0131 ,
		\u1_uk_K_r0_reg[7]/NET0131 ,
		_w23634_
	);
	LUT4 #(
		.INIT('h8d75)
	) name17808 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23635_
	);
	LUT2 #(
		.INIT('h2)
	) name17809 (
		_w23630_,
		_w23635_,
		_w23636_
	);
	LUT2 #(
		.INIT('h1)
	) name17810 (
		_w23634_,
		_w23630_,
		_w23637_
	);
	LUT3 #(
		.INIT('h08)
	) name17811 (
		_w23631_,
		_w23632_,
		_w23633_,
		_w23638_
	);
	LUT3 #(
		.INIT('hf6)
	) name17812 (
		_w23631_,
		_w23632_,
		_w23633_,
		_w23639_
	);
	LUT2 #(
		.INIT('h2)
	) name17813 (
		_w23637_,
		_w23639_,
		_w23640_
	);
	LUT4 #(
		.INIT('h0400)
	) name17814 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23641_
	);
	LUT2 #(
		.INIT('h2)
	) name17815 (
		_w23634_,
		_w23630_,
		_w23642_
	);
	LUT3 #(
		.INIT('h80)
	) name17816 (
		_w23631_,
		_w23632_,
		_w23633_,
		_w23643_
	);
	LUT4 #(
		.INIT('h1000)
	) name17817 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23644_
	);
	LUT4 #(
		.INIT('hedff)
	) name17818 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23645_
	);
	LUT4 #(
		.INIT('h1500)
	) name17819 (
		_w23641_,
		_w23642_,
		_w23643_,
		_w23645_,
		_w23646_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name17820 (
		_w23629_,
		_w23636_,
		_w23640_,
		_w23646_,
		_w23647_
	);
	LUT4 #(
		.INIT('hf5cf)
	) name17821 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23648_
	);
	LUT4 #(
		.INIT('h0810)
	) name17822 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23649_
	);
	LUT4 #(
		.INIT('h2000)
	) name17823 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23650_
	);
	LUT4 #(
		.INIT('h00fd)
	) name17824 (
		_w23631_,
		_w23632_,
		_w23633_,
		_w23630_,
		_w23651_
	);
	LUT4 #(
		.INIT('h0100)
	) name17825 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23652_
	);
	LUT4 #(
		.INIT('hbebf)
	) name17826 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23653_
	);
	LUT3 #(
		.INIT('h40)
	) name17827 (
		_w23650_,
		_w23651_,
		_w23653_,
		_w23654_
	);
	LUT4 #(
		.INIT('h8830)
	) name17828 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23655_
	);
	LUT4 #(
		.INIT('hfe00)
	) name17829 (
		_w23631_,
		_w23632_,
		_w23633_,
		_w23630_,
		_w23656_
	);
	LUT2 #(
		.INIT('h4)
	) name17830 (
		_w23655_,
		_w23656_,
		_w23657_
	);
	LUT4 #(
		.INIT('h00ab)
	) name17831 (
		_w23649_,
		_w23654_,
		_w23657_,
		_w23629_,
		_w23658_
	);
	LUT4 #(
		.INIT('h0008)
	) name17832 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23659_
	);
	LUT4 #(
		.INIT('h0048)
	) name17833 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23660_
	);
	LUT4 #(
		.INIT('heffb)
	) name17834 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23661_
	);
	LUT3 #(
		.INIT('hb1)
	) name17835 (
		_w23630_,
		_w23660_,
		_w23661_,
		_w23662_
	);
	LUT4 #(
		.INIT('h5655)
	) name17836 (
		\u1_L0_reg[14]/NET0131 ,
		_w23658_,
		_w23647_,
		_w23662_,
		_w23663_
	);
	LUT2 #(
		.INIT('h4)
	) name17837 (
		_w23546_,
		_w23543_,
		_w23664_
	);
	LUT4 #(
		.INIT('h0400)
	) name17838 (
		_w23546_,
		_w23543_,
		_w23544_,
		_w23541_,
		_w23665_
	);
	LUT3 #(
		.INIT('h08)
	) name17839 (
		_w23544_,
		_w23542_,
		_w23541_,
		_w23666_
	);
	LUT4 #(
		.INIT('h0002)
	) name17840 (
		_w23546_,
		_w23543_,
		_w23544_,
		_w23542_,
		_w23667_
	);
	LUT4 #(
		.INIT('h0002)
	) name17841 (
		_w23540_,
		_w23665_,
		_w23666_,
		_w23667_,
		_w23668_
	);
	LUT4 #(
		.INIT('h0400)
	) name17842 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23669_
	);
	LUT4 #(
		.INIT('h2000)
	) name17843 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23670_
	);
	LUT4 #(
		.INIT('hdbff)
	) name17844 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23671_
	);
	LUT4 #(
		.INIT('h3d39)
	) name17845 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23672_
	);
	LUT4 #(
		.INIT('h0010)
	) name17846 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23673_
	);
	LUT4 #(
		.INIT('h0051)
	) name17847 (
		_w23540_,
		_w23546_,
		_w23672_,
		_w23673_,
		_w23674_
	);
	LUT3 #(
		.INIT('h07)
	) name17848 (
		_w23668_,
		_w23671_,
		_w23674_,
		_w23675_
	);
	LUT4 #(
		.INIT('hfff6)
	) name17849 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23676_
	);
	LUT3 #(
		.INIT('h20)
	) name17850 (
		_w23547_,
		_w23669_,
		_w23676_,
		_w23677_
	);
	LUT4 #(
		.INIT('h0002)
	) name17851 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23678_
	);
	LUT3 #(
		.INIT('h02)
	) name17852 (
		_w23546_,
		_w23545_,
		_w23678_,
		_w23679_
	);
	LUT2 #(
		.INIT('h1)
	) name17853 (
		_w23540_,
		_w23546_,
		_w23680_
	);
	LUT4 #(
		.INIT('h0100)
	) name17854 (
		_w23540_,
		_w23546_,
		_w23544_,
		_w23542_,
		_w23681_
	);
	LUT3 #(
		.INIT('h0e)
	) name17855 (
		_w23677_,
		_w23679_,
		_w23681_,
		_w23682_
	);
	LUT3 #(
		.INIT('h65)
	) name17856 (
		\u1_L0_reg[15]/P0001 ,
		_w23675_,
		_w23682_,
		_w23683_
	);
	LUT4 #(
		.INIT('h32ff)
	) name17857 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23684_
	);
	LUT3 #(
		.INIT('h51)
	) name17858 (
		_w23507_,
		_w23509_,
		_w23510_,
		_w23685_
	);
	LUT2 #(
		.INIT('h4)
	) name17859 (
		_w23684_,
		_w23685_,
		_w23686_
	);
	LUT4 #(
		.INIT('h0002)
	) name17860 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23687_
	);
	LUT4 #(
		.INIT('h2000)
	) name17861 (
		_w23507_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23688_
	);
	LUT3 #(
		.INIT('h02)
	) name17862 (
		_w23522_,
		_w23688_,
		_w23687_,
		_w23689_
	);
	LUT4 #(
		.INIT('h2080)
	) name17863 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23690_
	);
	LUT4 #(
		.INIT('h0002)
	) name17864 (
		_w23507_,
		_w23508_,
		_w23509_,
		_w23511_,
		_w23691_
	);
	LUT2 #(
		.INIT('h1)
	) name17865 (
		_w23690_,
		_w23691_,
		_w23692_
	);
	LUT3 #(
		.INIT('h40)
	) name17866 (
		_w23686_,
		_w23689_,
		_w23692_,
		_w23693_
	);
	LUT3 #(
		.INIT('h71)
	) name17867 (
		_w23509_,
		_w23510_,
		_w23511_,
		_w23694_
	);
	LUT2 #(
		.INIT('h8)
	) name17868 (
		_w23507_,
		_w23508_,
		_w23695_
	);
	LUT2 #(
		.INIT('h4)
	) name17869 (
		_w23694_,
		_w23695_,
		_w23696_
	);
	LUT3 #(
		.INIT('h04)
	) name17870 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23697_
	);
	LUT3 #(
		.INIT('h01)
	) name17871 (
		_w23512_,
		_w23522_,
		_w23697_,
		_w23698_
	);
	LUT2 #(
		.INIT('h4)
	) name17872 (
		_w23696_,
		_w23698_,
		_w23699_
	);
	LUT3 #(
		.INIT('h79)
	) name17873 (
		_w23508_,
		_w23509_,
		_w23511_,
		_w23700_
	);
	LUT2 #(
		.INIT('h2)
	) name17874 (
		_w23524_,
		_w23700_,
		_w23701_
	);
	LUT3 #(
		.INIT('h20)
	) name17875 (
		_w23507_,
		_w23510_,
		_w23511_,
		_w23702_
	);
	LUT4 #(
		.INIT('hefaa)
	) name17876 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23703_
	);
	LUT2 #(
		.INIT('h1)
	) name17877 (
		_w23507_,
		_w23522_,
		_w23704_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name17878 (
		_w23523_,
		_w23702_,
		_w23703_,
		_w23704_,
		_w23705_
	);
	LUT2 #(
		.INIT('h4)
	) name17879 (
		_w23701_,
		_w23705_,
		_w23706_
	);
	LUT4 #(
		.INIT('ha955)
	) name17880 (
		\u1_L0_reg[26]/NET0131 ,
		_w23693_,
		_w23699_,
		_w23706_,
		_w23707_
	);
	LUT4 #(
		.INIT('h440c)
	) name17881 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23708_
	);
	LUT3 #(
		.INIT('h01)
	) name17882 (
		_w23509_,
		_w23510_,
		_w23511_,
		_w23709_
	);
	LUT4 #(
		.INIT('hfad8)
	) name17883 (
		_w23507_,
		_w23516_,
		_w23708_,
		_w23709_,
		_w23710_
	);
	LUT4 #(
		.INIT('h7df7)
	) name17884 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23711_
	);
	LUT3 #(
		.INIT('h45)
	) name17885 (
		_w23522_,
		_w23710_,
		_w23711_,
		_w23712_
	);
	LUT2 #(
		.INIT('h4)
	) name17886 (
		_w23507_,
		_w23508_,
		_w23713_
	);
	LUT2 #(
		.INIT('h8)
	) name17887 (
		_w23694_,
		_w23713_,
		_w23714_
	);
	LUT4 #(
		.INIT('h1090)
	) name17888 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23715_
	);
	LUT4 #(
		.INIT('haafb)
	) name17889 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23716_
	);
	LUT3 #(
		.INIT('h31)
	) name17890 (
		_w23507_,
		_w23715_,
		_w23716_,
		_w23717_
	);
	LUT3 #(
		.INIT('h8a)
	) name17891 (
		_w23522_,
		_w23714_,
		_w23717_,
		_w23718_
	);
	LUT4 #(
		.INIT('h6fdf)
	) name17892 (
		_w23508_,
		_w23509_,
		_w23510_,
		_w23511_,
		_w23719_
	);
	LUT2 #(
		.INIT('h2)
	) name17893 (
		_w23507_,
		_w23719_,
		_w23720_
	);
	LUT4 #(
		.INIT('h0777)
	) name17894 (
		_w23520_,
		_w23521_,
		_w23531_,
		_w23713_,
		_w23721_
	);
	LUT2 #(
		.INIT('h4)
	) name17895 (
		_w23720_,
		_w23721_,
		_w23722_
	);
	LUT4 #(
		.INIT('h5655)
	) name17896 (
		\u1_L0_reg[1]/NET0131 ,
		_w23718_,
		_w23712_,
		_w23722_,
		_w23723_
	);
	LUT4 #(
		.INIT('haa2a)
	) name17897 (
		_w23546_,
		_w23543_,
		_w23544_,
		_w23542_,
		_w23724_
	);
	LUT4 #(
		.INIT('h3fdd)
	) name17898 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23725_
	);
	LUT4 #(
		.INIT('h5545)
	) name17899 (
		_w23546_,
		_w23543_,
		_w23542_,
		_w23541_,
		_w23726_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name17900 (
		_w23670_,
		_w23724_,
		_w23725_,
		_w23726_,
		_w23727_
	);
	LUT4 #(
		.INIT('h4100)
	) name17901 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23728_
	);
	LUT3 #(
		.INIT('h02)
	) name17902 (
		_w23540_,
		_w23678_,
		_w23728_,
		_w23729_
	);
	LUT2 #(
		.INIT('h4)
	) name17903 (
		_w23727_,
		_w23729_,
		_w23730_
	);
	LUT4 #(
		.INIT('h002e)
	) name17904 (
		_w23546_,
		_w23543_,
		_w23542_,
		_w23541_,
		_w23731_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name17905 (
		_w23546_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23732_
	);
	LUT3 #(
		.INIT('h10)
	) name17906 (
		_w23562_,
		_w23731_,
		_w23732_,
		_w23733_
	);
	LUT2 #(
		.INIT('h1)
	) name17907 (
		_w23540_,
		_w23553_,
		_w23734_
	);
	LUT3 #(
		.INIT('h70)
	) name17908 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23735_
	);
	LUT3 #(
		.INIT('ha8)
	) name17909 (
		_w23546_,
		_w23544_,
		_w23541_,
		_w23736_
	);
	LUT3 #(
		.INIT('h15)
	) name17910 (
		_w23566_,
		_w23735_,
		_w23736_,
		_w23737_
	);
	LUT3 #(
		.INIT('h40)
	) name17911 (
		_w23733_,
		_w23734_,
		_w23737_,
		_w23738_
	);
	LUT4 #(
		.INIT('h0002)
	) name17912 (
		_w23546_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23739_
	);
	LUT3 #(
		.INIT('h07)
	) name17913 (
		_w23664_,
		_w23666_,
		_w23739_,
		_w23740_
	);
	LUT4 #(
		.INIT('ha955)
	) name17914 (
		\u1_L0_reg[21]/NET0131 ,
		_w23730_,
		_w23738_,
		_w23740_,
		_w23741_
	);
	LUT4 #(
		.INIT('h5eb0)
	) name17915 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23742_
	);
	LUT4 #(
		.INIT('h9fdf)
	) name17916 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23743_
	);
	LUT4 #(
		.INIT('he200)
	) name17917 (
		_w23648_,
		_w23630_,
		_w23742_,
		_w23743_,
		_w23744_
	);
	LUT2 #(
		.INIT('h2)
	) name17918 (
		_w23629_,
		_w23744_,
		_w23745_
	);
	LUT4 #(
		.INIT('hbff9)
	) name17919 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23746_
	);
	LUT2 #(
		.INIT('h2)
	) name17920 (
		_w23630_,
		_w23746_,
		_w23747_
	);
	LUT2 #(
		.INIT('h4)
	) name17921 (
		_w23631_,
		_w23630_,
		_w23748_
	);
	LUT4 #(
		.INIT('hfa3f)
	) name17922 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23749_
	);
	LUT3 #(
		.INIT('hb0)
	) name17923 (
		_w23631_,
		_w23632_,
		_w23630_,
		_w23750_
	);
	LUT4 #(
		.INIT('h5501)
	) name17924 (
		_w23634_,
		_w23632_,
		_w23633_,
		_w23630_,
		_w23751_
	);
	LUT4 #(
		.INIT('he0ee)
	) name17925 (
		_w23748_,
		_w23749_,
		_w23750_,
		_w23751_,
		_w23752_
	);
	LUT4 #(
		.INIT('h0020)
	) name17926 (
		_w23634_,
		_w23632_,
		_w23633_,
		_w23630_,
		_w23753_
	);
	LUT2 #(
		.INIT('h1)
	) name17927 (
		_w23650_,
		_w23753_,
		_w23754_
	);
	LUT4 #(
		.INIT('h0e00)
	) name17928 (
		_w23629_,
		_w23752_,
		_w23747_,
		_w23754_,
		_w23755_
	);
	LUT3 #(
		.INIT('h65)
	) name17929 (
		\u1_L0_reg[25]/NET0131 ,
		_w23745_,
		_w23755_,
		_w23756_
	);
	LUT4 #(
		.INIT('hc693)
	) name17930 (
		decrypt_pad,
		\u1_R0_reg[9]/NET0131 ,
		\u1_uk_K_r0_reg[26]/NET0131 ,
		\u1_uk_K_r0_reg[5]/NET0131 ,
		_w23757_
	);
	LUT4 #(
		.INIT('hc693)
	) name17931 (
		decrypt_pad,
		\u1_R0_reg[5]/NET0131 ,
		\u1_uk_K_r0_reg[13]/NET0131 ,
		\u1_uk_K_r0_reg[17]/NET0131 ,
		_w23758_
	);
	LUT4 #(
		.INIT('hc963)
	) name17932 (
		decrypt_pad,
		\u1_R0_reg[4]/NET0131 ,
		\u1_uk_K_r0_reg[13]/NET0131 ,
		\u1_uk_K_r0_reg[34]/NET0131 ,
		_w23759_
	);
	LUT3 #(
		.INIT('h8a)
	) name17933 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23760_
	);
	LUT3 #(
		.INIT('h82)
	) name17934 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23761_
	);
	LUT4 #(
		.INIT('hc963)
	) name17935 (
		decrypt_pad,
		\u1_R0_reg[7]/NET0131 ,
		\u1_uk_K_r0_reg[34]/NET0131 ,
		\u1_uk_K_r0_reg[55]/NET0131 ,
		_w23762_
	);
	LUT4 #(
		.INIT('hc963)
	) name17936 (
		decrypt_pad,
		\u1_R0_reg[6]/NET0131 ,
		\u1_uk_K_r0_reg[40]/NET0131 ,
		\u1_uk_K_r0_reg[4]/NET0131 ,
		_w23763_
	);
	LUT4 #(
		.INIT('h1000)
	) name17937 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23764_
	);
	LUT3 #(
		.INIT('h02)
	) name17938 (
		_w23762_,
		_w23764_,
		_w23761_,
		_w23765_
	);
	LUT3 #(
		.INIT('h10)
	) name17939 (
		_w23759_,
		_w23758_,
		_w23763_,
		_w23766_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name17940 (
		_w23759_,
		_w23758_,
		_w23762_,
		_w23763_,
		_w23767_
	);
	LUT4 #(
		.INIT('hbfae)
	) name17941 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23768_
	);
	LUT4 #(
		.INIT('h2000)
	) name17942 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23769_
	);
	LUT4 #(
		.INIT('h9fae)
	) name17943 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23770_
	);
	LUT2 #(
		.INIT('h8)
	) name17944 (
		_w23767_,
		_w23770_,
		_w23771_
	);
	LUT3 #(
		.INIT('h0d)
	) name17945 (
		_w23757_,
		_w23758_,
		_w23762_,
		_w23772_
	);
	LUT2 #(
		.INIT('h2)
	) name17946 (
		_w23759_,
		_w23763_,
		_w23773_
	);
	LUT4 #(
		.INIT('hc963)
	) name17947 (
		decrypt_pad,
		\u1_R0_reg[8]/NET0131 ,
		\u1_uk_K_r0_reg[25]/P0001 ,
		\u1_uk_K_r0_reg[46]/NET0131 ,
		_w23774_
	);
	LUT4 #(
		.INIT('h0400)
	) name17948 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23775_
	);
	LUT4 #(
		.INIT('h008a)
	) name17949 (
		_w23774_,
		_w23772_,
		_w23773_,
		_w23775_,
		_w23776_
	);
	LUT3 #(
		.INIT('he0)
	) name17950 (
		_w23765_,
		_w23771_,
		_w23776_,
		_w23777_
	);
	LUT4 #(
		.INIT('h0b08)
	) name17951 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23778_
	);
	LUT4 #(
		.INIT('ha4a6)
	) name17952 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23779_
	);
	LUT4 #(
		.INIT('h7772)
	) name17953 (
		_w23762_,
		_w23768_,
		_w23766_,
		_w23779_,
		_w23780_
	);
	LUT4 #(
		.INIT('h0900)
	) name17954 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23781_
	);
	LUT3 #(
		.INIT('h01)
	) name17955 (
		_w23774_,
		_w23769_,
		_w23781_,
		_w23782_
	);
	LUT2 #(
		.INIT('h4)
	) name17956 (
		_w23780_,
		_w23782_,
		_w23783_
	);
	LUT3 #(
		.INIT('ha9)
	) name17957 (
		\u1_L0_reg[28]/NET0131 ,
		_w23777_,
		_w23783_,
		_w23784_
	);
	LUT4 #(
		.INIT('h7d7c)
	) name17958 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23785_
	);
	LUT2 #(
		.INIT('h1)
	) name17959 (
		_w23480_,
		_w23785_,
		_w23786_
	);
	LUT4 #(
		.INIT('hc6ff)
	) name17960 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23787_
	);
	LUT2 #(
		.INIT('h2)
	) name17961 (
		_w23480_,
		_w23787_,
		_w23788_
	);
	LUT4 #(
		.INIT('h0012)
	) name17962 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23789_
	);
	LUT3 #(
		.INIT('h01)
	) name17963 (
		_w23495_,
		_w23496_,
		_w23789_,
		_w23790_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name17964 (
		_w23474_,
		_w23788_,
		_w23786_,
		_w23790_,
		_w23791_
	);
	LUT4 #(
		.INIT('h3df2)
	) name17965 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23792_
	);
	LUT4 #(
		.INIT('ha6bf)
	) name17966 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23793_
	);
	LUT4 #(
		.INIT('h0020)
	) name17967 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23794_
	);
	LUT4 #(
		.INIT('h00d8)
	) name17968 (
		_w23480_,
		_w23792_,
		_w23793_,
		_w23794_,
		_w23795_
	);
	LUT4 #(
		.INIT('h4000)
	) name17969 (
		_w23475_,
		_w23480_,
		_w23478_,
		_w23477_,
		_w23796_
	);
	LUT2 #(
		.INIT('h1)
	) name17970 (
		_w23483_,
		_w23796_,
		_w23797_
	);
	LUT3 #(
		.INIT('he0)
	) name17971 (
		_w23474_,
		_w23795_,
		_w23797_,
		_w23798_
	);
	LUT3 #(
		.INIT('h9a)
	) name17972 (
		\u1_L0_reg[29]/NET0131 ,
		_w23791_,
		_w23798_,
		_w23799_
	);
	LUT4 #(
		.INIT('h0800)
	) name17973 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23800_
	);
	LUT2 #(
		.INIT('h8)
	) name17974 (
		_w23762_,
		_w23800_,
		_w23801_
	);
	LUT2 #(
		.INIT('h1)
	) name17975 (
		_w23758_,
		_w23762_,
		_w23802_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name17976 (
		_w23759_,
		_w23758_,
		_w23762_,
		_w23763_,
		_w23803_
	);
	LUT3 #(
		.INIT('h8a)
	) name17977 (
		_w23757_,
		_w23758_,
		_w23763_,
		_w23804_
	);
	LUT3 #(
		.INIT('h45)
	) name17978 (
		_w23774_,
		_w23803_,
		_w23804_,
		_w23805_
	);
	LUT4 #(
		.INIT('h0034)
	) name17979 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23806_
	);
	LUT3 #(
		.INIT('h08)
	) name17980 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23807_
	);
	LUT4 #(
		.INIT('h51f3)
	) name17981 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23808_
	);
	LUT4 #(
		.INIT('h3332)
	) name17982 (
		_w23762_,
		_w23806_,
		_w23808_,
		_w23807_,
		_w23809_
	);
	LUT3 #(
		.INIT('h01)
	) name17983 (
		_w23757_,
		_w23758_,
		_w23763_,
		_w23810_
	);
	LUT4 #(
		.INIT('h0002)
	) name17984 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23811_
	);
	LUT4 #(
		.INIT('h0080)
	) name17985 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23812_
	);
	LUT4 #(
		.INIT('h80c0)
	) name17986 (
		_w23759_,
		_w23758_,
		_w23762_,
		_w23763_,
		_w23813_
	);
	LUT4 #(
		.INIT('h0002)
	) name17987 (
		_w23774_,
		_w23813_,
		_w23812_,
		_w23811_,
		_w23814_
	);
	LUT4 #(
		.INIT('h00bf)
	) name17988 (
		_w23801_,
		_w23805_,
		_w23809_,
		_w23814_,
		_w23815_
	);
	LUT4 #(
		.INIT('h0100)
	) name17989 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23816_
	);
	LUT4 #(
		.INIT('hf070)
	) name17990 (
		_w23759_,
		_w23758_,
		_w23762_,
		_w23763_,
		_w23817_
	);
	LUT2 #(
		.INIT('h4)
	) name17991 (
		_w23816_,
		_w23817_,
		_w23818_
	);
	LUT4 #(
		.INIT('he6fe)
	) name17992 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23819_
	);
	LUT4 #(
		.INIT('h4004)
	) name17993 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23820_
	);
	LUT4 #(
		.INIT('h0301)
	) name17994 (
		_w23774_,
		_w23762_,
		_w23820_,
		_w23819_,
		_w23821_
	);
	LUT2 #(
		.INIT('h1)
	) name17995 (
		_w23818_,
		_w23821_,
		_w23822_
	);
	LUT3 #(
		.INIT('h56)
	) name17996 (
		\u1_L0_reg[2]/NET0131 ,
		_w23815_,
		_w23822_,
		_w23823_
	);
	LUT4 #(
		.INIT('hfcdf)
	) name17997 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23824_
	);
	LUT2 #(
		.INIT('h1)
	) name17998 (
		_w23480_,
		_w23824_,
		_w23825_
	);
	LUT4 #(
		.INIT('he36f)
	) name17999 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23826_
	);
	LUT4 #(
		.INIT('h0301)
	) name18000 (
		_w23480_,
		_w23483_,
		_w23486_,
		_w23826_,
		_w23827_
	);
	LUT3 #(
		.INIT('h45)
	) name18001 (
		_w23474_,
		_w23825_,
		_w23827_,
		_w23828_
	);
	LUT4 #(
		.INIT('h4000)
	) name18002 (
		_w23475_,
		_w23480_,
		_w23476_,
		_w23478_,
		_w23829_
	);
	LUT4 #(
		.INIT('h5eff)
	) name18003 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23830_
	);
	LUT4 #(
		.INIT('h0d00)
	) name18004 (
		_w23485_,
		_w23489_,
		_w23829_,
		_w23830_,
		_w23831_
	);
	LUT3 #(
		.INIT('h9e)
	) name18005 (
		_w23476_,
		_w23478_,
		_w23477_,
		_w23832_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name18006 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23833_
	);
	LUT4 #(
		.INIT('h2223)
	) name18007 (
		_w23475_,
		_w23480_,
		_w23476_,
		_w23478_,
		_w23834_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name18008 (
		_w23492_,
		_w23832_,
		_w23833_,
		_w23834_,
		_w23835_
	);
	LUT3 #(
		.INIT('hd0)
	) name18009 (
		_w23474_,
		_w23831_,
		_w23835_,
		_w23836_
	);
	LUT3 #(
		.INIT('h65)
	) name18010 (
		\u1_L0_reg[4]/NET0131 ,
		_w23828_,
		_w23836_,
		_w23837_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name18011 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23838_
	);
	LUT4 #(
		.INIT('hebed)
	) name18012 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23839_
	);
	LUT4 #(
		.INIT('h0313)
	) name18013 (
		_w23774_,
		_w23762_,
		_w23838_,
		_w23839_,
		_w23840_
	);
	LUT4 #(
		.INIT('h74d6)
	) name18014 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23841_
	);
	LUT2 #(
		.INIT('h2)
	) name18015 (
		_w23762_,
		_w23841_,
		_w23842_
	);
	LUT3 #(
		.INIT('h04)
	) name18016 (
		_w23759_,
		_w23757_,
		_w23763_,
		_w23843_
	);
	LUT3 #(
		.INIT('h45)
	) name18017 (
		_w23774_,
		_w23802_,
		_w23843_,
		_w23844_
	);
	LUT3 #(
		.INIT('h40)
	) name18018 (
		_w23759_,
		_w23757_,
		_w23763_,
		_w23845_
	);
	LUT4 #(
		.INIT('heee4)
	) name18019 (
		_w23762_,
		_w23778_,
		_w23810_,
		_w23845_,
		_w23846_
	);
	LUT4 #(
		.INIT('hdf6f)
	) name18020 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w23847_
	);
	LUT4 #(
		.INIT('h8a00)
	) name18021 (
		_w23774_,
		_w23803_,
		_w23804_,
		_w23847_,
		_w23848_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name18022 (
		_w23842_,
		_w23844_,
		_w23846_,
		_w23848_,
		_w23849_
	);
	LUT3 #(
		.INIT('ha9)
	) name18023 (
		\u1_L0_reg[13]/NET0131 ,
		_w23840_,
		_w23849_,
		_w23850_
	);
	LUT4 #(
		.INIT('hf3ec)
	) name18024 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23851_
	);
	LUT3 #(
		.INIT('h7d)
	) name18025 (
		_w23576_,
		_w23573_,
		_w23574_,
		_w23852_
	);
	LUT4 #(
		.INIT('hfd7f)
	) name18026 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23853_
	);
	LUT4 #(
		.INIT('he400)
	) name18027 (
		_w23572_,
		_w23851_,
		_w23852_,
		_w23853_,
		_w23854_
	);
	LUT4 #(
		.INIT('h4555)
	) name18028 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23855_
	);
	LUT4 #(
		.INIT('haa8a)
	) name18029 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23856_
	);
	LUT3 #(
		.INIT('h02)
	) name18030 (
		_w23572_,
		_w23856_,
		_w23855_,
		_w23857_
	);
	LUT4 #(
		.INIT('h0400)
	) name18031 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23858_
	);
	LUT4 #(
		.INIT('hc9cd)
	) name18032 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23859_
	);
	LUT4 #(
		.INIT('h4041)
	) name18033 (
		_w23572_,
		_w23575_,
		_w23576_,
		_w23573_,
		_w23860_
	);
	LUT4 #(
		.INIT('h0040)
	) name18034 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23861_
	);
	LUT4 #(
		.INIT('h5fbf)
	) name18035 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23862_
	);
	LUT4 #(
		.INIT('h0d00)
	) name18036 (
		_w23572_,
		_w23859_,
		_w23860_,
		_w23862_,
		_w23863_
	);
	LUT4 #(
		.INIT('h0e04)
	) name18037 (
		_w23571_,
		_w23854_,
		_w23857_,
		_w23863_,
		_w23864_
	);
	LUT2 #(
		.INIT('h9)
	) name18038 (
		\u1_L0_reg[17]/NET0131 ,
		_w23864_,
		_w23865_
	);
	LUT4 #(
		.INIT('h1001)
	) name18039 (
		_w23480_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23866_
	);
	LUT4 #(
		.INIT('h0200)
	) name18040 (
		_w23480_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23867_
	);
	LUT3 #(
		.INIT('h15)
	) name18041 (
		_w23480_,
		_w23478_,
		_w23477_,
		_w23868_
	);
	LUT3 #(
		.INIT('h8c)
	) name18042 (
		_w23475_,
		_w23476_,
		_w23477_,
		_w23869_
	);
	LUT4 #(
		.INIT('h0045)
	) name18043 (
		_w23474_,
		_w23868_,
		_w23869_,
		_w23867_,
		_w23870_
	);
	LUT4 #(
		.INIT('h2000)
	) name18044 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23871_
	);
	LUT3 #(
		.INIT('h04)
	) name18045 (
		_w23480_,
		_w23476_,
		_w23477_,
		_w23872_
	);
	LUT4 #(
		.INIT('hef00)
	) name18046 (
		_w23475_,
		_w23478_,
		_w23477_,
		_w23474_,
		_w23873_
	);
	LUT3 #(
		.INIT('h10)
	) name18047 (
		_w23872_,
		_w23871_,
		_w23873_,
		_w23874_
	);
	LUT4 #(
		.INIT('hbbcf)
	) name18048 (
		_w23475_,
		_w23476_,
		_w23478_,
		_w23477_,
		_w23875_
	);
	LUT3 #(
		.INIT('h31)
	) name18049 (
		_w23480_,
		_w23789_,
		_w23875_,
		_w23876_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name18050 (
		_w23866_,
		_w23870_,
		_w23874_,
		_w23876_,
		_w23877_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name18051 (
		_w23475_,
		_w23477_,
		_w23486_,
		_w23500_,
		_w23878_
	);
	LUT3 #(
		.INIT('h65)
	) name18052 (
		\u1_L0_reg[19]/NET0131 ,
		_w23877_,
		_w23878_,
		_w23879_
	);
	LUT4 #(
		.INIT('hb7b4)
	) name18053 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23880_
	);
	LUT2 #(
		.INIT('h1)
	) name18054 (
		_w23546_,
		_w23880_,
		_w23881_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name18055 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23882_
	);
	LUT4 #(
		.INIT('h80aa)
	) name18056 (
		_w23546_,
		_w23543_,
		_w23544_,
		_w23542_,
		_w23883_
	);
	LUT4 #(
		.INIT('he7dd)
	) name18057 (
		_w23543_,
		_w23544_,
		_w23542_,
		_w23541_,
		_w23884_
	);
	LUT3 #(
		.INIT('hb0)
	) name18058 (
		_w23882_,
		_w23883_,
		_w23884_,
		_w23885_
	);
	LUT3 #(
		.INIT('h8a)
	) name18059 (
		_w23540_,
		_w23881_,
		_w23885_,
		_w23886_
	);
	LUT4 #(
		.INIT('haa8a)
	) name18060 (
		_w23546_,
		_w23543_,
		_w23544_,
		_w23541_,
		_w23887_
	);
	LUT4 #(
		.INIT('h4544)
	) name18061 (
		_w23540_,
		_w23565_,
		_w23563_,
		_w23887_,
		_w23888_
	);
	LUT2 #(
		.INIT('h4)
	) name18062 (
		_w23546_,
		_w23564_,
		_w23889_
	);
	LUT3 #(
		.INIT('h10)
	) name18063 (
		_w23559_,
		_w23562_,
		_w23680_,
		_w23890_
	);
	LUT4 #(
		.INIT('h0200)
	) name18064 (
		_w23546_,
		_w23543_,
		_w23544_,
		_w23541_,
		_w23891_
	);
	LUT3 #(
		.INIT('h07)
	) name18065 (
		_w23558_,
		_w23550_,
		_w23891_,
		_w23892_
	);
	LUT4 #(
		.INIT('h0100)
	) name18066 (
		_w23888_,
		_w23890_,
		_w23889_,
		_w23892_,
		_w23893_
	);
	LUT3 #(
		.INIT('h65)
	) name18067 (
		\u1_L0_reg[27]/NET0131 ,
		_w23886_,
		_w23893_,
		_w23894_
	);
	LUT4 #(
		.INIT('hdbe9)
	) name18068 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23895_
	);
	LUT4 #(
		.INIT('h4000)
	) name18069 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23896_
	);
	LUT4 #(
		.INIT('hae76)
	) name18070 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23897_
	);
	LUT4 #(
		.INIT('h3210)
	) name18071 (
		_w23447_,
		_w23896_,
		_w23895_,
		_w23897_,
		_w23898_
	);
	LUT2 #(
		.INIT('h2)
	) name18072 (
		_w23451_,
		_w23898_,
		_w23899_
	);
	LUT4 #(
		.INIT('h79bf)
	) name18073 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23900_
	);
	LUT4 #(
		.INIT('h5507)
	) name18074 (
		_w23447_,
		_w23467_,
		_w23614_,
		_w23618_,
		_w23901_
	);
	LUT4 #(
		.INIT('h008c)
	) name18075 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23447_,
		_w23902_
	);
	LUT4 #(
		.INIT('h153f)
	) name18076 (
		_w23461_,
		_w23453_,
		_w23619_,
		_w23902_,
		_w23903_
	);
	LUT4 #(
		.INIT('hea00)
	) name18077 (
		_w23451_,
		_w23900_,
		_w23901_,
		_w23903_,
		_w23904_
	);
	LUT3 #(
		.INIT('h65)
	) name18078 (
		\u1_L0_reg[32]/NET0131 ,
		_w23899_,
		_w23904_,
		_w23905_
	);
	LUT4 #(
		.INIT('hc963)
	) name18079 (
		decrypt_pad,
		\u1_R0_reg[11]/NET0131 ,
		\u1_uk_K_r0_reg[20]/NET0131 ,
		\u1_uk_K_r0_reg[41]/NET0131 ,
		_w23906_
	);
	LUT4 #(
		.INIT('hc693)
	) name18080 (
		decrypt_pad,
		\u1_R0_reg[12]/NET0131 ,
		\u1_uk_K_r0_reg[24]/NET0131 ,
		\u1_uk_K_r0_reg[3]/NET0131 ,
		_w23907_
	);
	LUT4 #(
		.INIT('hc693)
	) name18081 (
		decrypt_pad,
		\u1_R0_reg[13]/NET0131 ,
		\u1_uk_K_r0_reg[12]/NET0131 ,
		\u1_uk_K_r0_reg[48]/NET0131 ,
		_w23908_
	);
	LUT4 #(
		.INIT('hc963)
	) name18082 (
		decrypt_pad,
		\u1_R0_reg[9]/NET0131 ,
		\u1_uk_K_r0_reg[11]/NET0131 ,
		\u1_uk_K_r0_reg[32]/NET0131 ,
		_w23909_
	);
	LUT4 #(
		.INIT('hc963)
	) name18083 (
		decrypt_pad,
		\u1_R0_reg[10]/NET0131 ,
		\u1_uk_K_r0_reg[19]/NET0131 ,
		\u1_uk_K_r0_reg[40]/NET0131 ,
		_w23910_
	);
	LUT4 #(
		.INIT('hc963)
	) name18084 (
		decrypt_pad,
		\u1_R0_reg[8]/NET0131 ,
		\u1_uk_K_r0_reg[39]/NET0131 ,
		\u1_uk_K_r0_reg[3]/NET0131 ,
		_w23911_
	);
	LUT2 #(
		.INIT('h2)
	) name18085 (
		_w23908_,
		_w23911_,
		_w23912_
	);
	LUT2 #(
		.INIT('h4)
	) name18086 (
		_w23908_,
		_w23911_,
		_w23913_
	);
	LUT4 #(
		.INIT('hc733)
	) name18087 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23914_
	);
	LUT2 #(
		.INIT('h1)
	) name18088 (
		_w23910_,
		_w23909_,
		_w23915_
	);
	LUT4 #(
		.INIT('h0001)
	) name18089 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23916_
	);
	LUT4 #(
		.INIT('hff76)
	) name18090 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23917_
	);
	LUT4 #(
		.INIT('h08cc)
	) name18091 (
		_w23907_,
		_w23906_,
		_w23914_,
		_w23917_,
		_w23918_
	);
	LUT2 #(
		.INIT('h9)
	) name18092 (
		_w23910_,
		_w23909_,
		_w23919_
	);
	LUT2 #(
		.INIT('h8)
	) name18093 (
		_w23908_,
		_w23911_,
		_w23920_
	);
	LUT3 #(
		.INIT('h46)
	) name18094 (
		_w23908_,
		_w23911_,
		_w23906_,
		_w23921_
	);
	LUT2 #(
		.INIT('h2)
	) name18095 (
		_w23919_,
		_w23921_,
		_w23922_
	);
	LUT3 #(
		.INIT('h10)
	) name18096 (
		_w23910_,
		_w23911_,
		_w23906_,
		_w23923_
	);
	LUT4 #(
		.INIT('h1428)
	) name18097 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23924_
	);
	LUT3 #(
		.INIT('h45)
	) name18098 (
		_w23907_,
		_w23923_,
		_w23924_,
		_w23925_
	);
	LUT2 #(
		.INIT('h8)
	) name18099 (
		_w23907_,
		_w23910_,
		_w23926_
	);
	LUT3 #(
		.INIT('h10)
	) name18100 (
		_w23908_,
		_w23911_,
		_w23909_,
		_w23927_
	);
	LUT4 #(
		.INIT('h0acf)
	) name18101 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23928_
	);
	LUT4 #(
		.INIT('h008a)
	) name18102 (
		_w23907_,
		_w23908_,
		_w23909_,
		_w23906_,
		_w23929_
	);
	LUT4 #(
		.INIT('h7077)
	) name18103 (
		_w23926_,
		_w23927_,
		_w23928_,
		_w23929_,
		_w23930_
	);
	LUT4 #(
		.INIT('h4500)
	) name18104 (
		_w23918_,
		_w23922_,
		_w23925_,
		_w23930_,
		_w23931_
	);
	LUT2 #(
		.INIT('h9)
	) name18105 (
		\u1_L0_reg[6]/NET0131 ,
		_w23931_,
		_w23932_
	);
	LUT4 #(
		.INIT('ha3b4)
	) name18106 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23933_
	);
	LUT2 #(
		.INIT('h1)
	) name18107 (
		_w23447_,
		_w23933_,
		_w23934_
	);
	LUT4 #(
		.INIT('h6800)
	) name18108 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23935_
	);
	LUT3 #(
		.INIT('h09)
	) name18109 (
		_w23449_,
		_w23448_,
		_w23452_,
		_w23936_
	);
	LUT4 #(
		.INIT('h00a4)
	) name18110 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23937_
	);
	LUT4 #(
		.INIT('h002a)
	) name18111 (
		_w23451_,
		_w23447_,
		_w23937_,
		_w23935_,
		_w23938_
	);
	LUT4 #(
		.INIT('h4800)
	) name18112 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23452_,
		_w23939_
	);
	LUT4 #(
		.INIT('hdf00)
	) name18113 (
		_w23449_,
		_w23450_,
		_w23448_,
		_w23447_,
		_w23940_
	);
	LUT4 #(
		.INIT('h5455)
	) name18114 (
		_w23451_,
		_w23936_,
		_w23939_,
		_w23940_,
		_w23941_
	);
	LUT3 #(
		.INIT('h0b)
	) name18115 (
		_w23934_,
		_w23938_,
		_w23941_,
		_w23942_
	);
	LUT2 #(
		.INIT('h4)
	) name18116 (
		_w23447_,
		_w23935_,
		_w23943_
	);
	LUT2 #(
		.INIT('h2)
	) name18117 (
		_w23451_,
		_w23447_,
		_w23944_
	);
	LUT4 #(
		.INIT('h00dc)
	) name18118 (
		_w23447_,
		_w23458_,
		_w23937_,
		_w23944_,
		_w23945_
	);
	LUT2 #(
		.INIT('h1)
	) name18119 (
		_w23943_,
		_w23945_,
		_w23946_
	);
	LUT3 #(
		.INIT('h65)
	) name18120 (
		\u1_L0_reg[7]/NET0131 ,
		_w23942_,
		_w23946_,
		_w23947_
	);
	LUT4 #(
		.INIT('hf55d)
	) name18121 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23948_
	);
	LUT4 #(
		.INIT('h5eff)
	) name18122 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23949_
	);
	LUT4 #(
		.INIT('hbfcb)
	) name18123 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23950_
	);
	LUT4 #(
		.INIT('he400)
	) name18124 (
		_w23630_,
		_w23948_,
		_w23949_,
		_w23950_,
		_w23951_
	);
	LUT4 #(
		.INIT('h0001)
	) name18125 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23952_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name18126 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23953_
	);
	LUT3 #(
		.INIT('h04)
	) name18127 (
		_w23634_,
		_w23633_,
		_w23630_,
		_w23954_
	);
	LUT4 #(
		.INIT('h0031)
	) name18128 (
		_w23630_,
		_w23660_,
		_w23953_,
		_w23954_,
		_w23955_
	);
	LUT4 #(
		.INIT('hbf97)
	) name18129 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w23956_
	);
	LUT3 #(
		.INIT('hb1)
	) name18130 (
		_w23630_,
		_w23641_,
		_w23956_,
		_w23957_
	);
	LUT4 #(
		.INIT('he400)
	) name18131 (
		_w23629_,
		_w23951_,
		_w23955_,
		_w23957_,
		_w23958_
	);
	LUT2 #(
		.INIT('h9)
	) name18132 (
		\u1_L0_reg[8]/NET0131 ,
		_w23958_,
		_w23959_
	);
	LUT3 #(
		.INIT('h80)
	) name18133 (
		_w23908_,
		_w23911_,
		_w23909_,
		_w23960_
	);
	LUT4 #(
		.INIT('h3ef2)
	) name18134 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23961_
	);
	LUT4 #(
		.INIT('h6800)
	) name18135 (
		_w23908_,
		_w23911_,
		_w23909_,
		_w23906_,
		_w23962_
	);
	LUT4 #(
		.INIT('h0032)
	) name18136 (
		_w23906_,
		_w23916_,
		_w23961_,
		_w23962_,
		_w23963_
	);
	LUT4 #(
		.INIT('h6979)
	) name18137 (
		_w23908_,
		_w23911_,
		_w23909_,
		_w23906_,
		_w23964_
	);
	LUT3 #(
		.INIT('h20)
	) name18138 (
		_w23908_,
		_w23911_,
		_w23909_,
		_w23965_
	);
	LUT4 #(
		.INIT('h0012)
	) name18139 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23906_,
		_w23966_
	);
	LUT4 #(
		.INIT('h0702)
	) name18140 (
		_w23910_,
		_w23965_,
		_w23966_,
		_w23964_,
		_w23967_
	);
	LUT4 #(
		.INIT('h0008)
	) name18141 (
		_w23910_,
		_w23911_,
		_w23909_,
		_w23906_,
		_w23968_
	);
	LUT4 #(
		.INIT('hdffd)
	) name18142 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23969_
	);
	LUT3 #(
		.INIT('h31)
	) name18143 (
		_w23906_,
		_w23968_,
		_w23969_,
		_w23970_
	);
	LUT4 #(
		.INIT('hd800)
	) name18144 (
		_w23907_,
		_w23967_,
		_w23963_,
		_w23970_,
		_w23971_
	);
	LUT2 #(
		.INIT('h9)
	) name18145 (
		\u1_L0_reg[16]/NET0131 ,
		_w23971_,
		_w23972_
	);
	LUT4 #(
		.INIT('hfcc7)
	) name18146 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23973_
	);
	LUT2 #(
		.INIT('h1)
	) name18147 (
		_w23572_,
		_w23973_,
		_w23974_
	);
	LUT3 #(
		.INIT('ha8)
	) name18148 (
		_w23572_,
		_w23575_,
		_w23574_,
		_w23975_
	);
	LUT2 #(
		.INIT('h8)
	) name18149 (
		_w23588_,
		_w23975_,
		_w23976_
	);
	LUT3 #(
		.INIT('h07)
	) name18150 (
		_w23587_,
		_w23595_,
		_w23858_,
		_w23977_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name18151 (
		_w23571_,
		_w23974_,
		_w23976_,
		_w23977_,
		_w23978_
	);
	LUT4 #(
		.INIT('h373f)
	) name18152 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23979_
	);
	LUT2 #(
		.INIT('h1)
	) name18153 (
		_w23572_,
		_w23979_,
		_w23980_
	);
	LUT4 #(
		.INIT('h0020)
	) name18154 (
		_w23572_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23981_
	);
	LUT4 #(
		.INIT('h0800)
	) name18155 (
		_w23572_,
		_w23575_,
		_w23576_,
		_w23574_,
		_w23982_
	);
	LUT3 #(
		.INIT('h7e)
	) name18156 (
		_w23575_,
		_w23573_,
		_w23574_,
		_w23983_
	);
	LUT3 #(
		.INIT('h10)
	) name18157 (
		_w23981_,
		_w23982_,
		_w23983_,
		_w23984_
	);
	LUT3 #(
		.INIT('hd9)
	) name18158 (
		_w23576_,
		_w23573_,
		_w23574_,
		_w23985_
	);
	LUT4 #(
		.INIT('h7ebf)
	) name18159 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w23986_
	);
	LUT4 #(
		.INIT('hfda8)
	) name18160 (
		_w23572_,
		_w23575_,
		_w23985_,
		_w23986_,
		_w23987_
	);
	LUT4 #(
		.INIT('hba00)
	) name18161 (
		_w23571_,
		_w23980_,
		_w23984_,
		_w23987_,
		_w23988_
	);
	LUT3 #(
		.INIT('h9a)
	) name18162 (
		\u1_L0_reg[23]/NET0131 ,
		_w23978_,
		_w23988_,
		_w23989_
	);
	LUT4 #(
		.INIT('hf859)
	) name18163 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23990_
	);
	LUT4 #(
		.INIT('h0020)
	) name18164 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23991_
	);
	LUT4 #(
		.INIT('h5504)
	) name18165 (
		_w23907_,
		_w23906_,
		_w23990_,
		_w23991_,
		_w23992_
	);
	LUT3 #(
		.INIT('h0e)
	) name18166 (
		_w23910_,
		_w23909_,
		_w23906_,
		_w23993_
	);
	LUT3 #(
		.INIT('h10)
	) name18167 (
		_w23910_,
		_w23909_,
		_w23906_,
		_w23994_
	);
	LUT4 #(
		.INIT('h5510)
	) name18168 (
		_w23912_,
		_w23913_,
		_w23993_,
		_w23994_,
		_w23995_
	);
	LUT4 #(
		.INIT('h57f7)
	) name18169 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23996_
	);
	LUT4 #(
		.INIT('h3f15)
	) name18170 (
		_w23906_,
		_w23915_,
		_w23921_,
		_w23996_,
		_w23997_
	);
	LUT3 #(
		.INIT('h8a)
	) name18171 (
		_w23907_,
		_w23995_,
		_w23997_,
		_w23998_
	);
	LUT4 #(
		.INIT('h0041)
	) name18172 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w23999_
	);
	LUT4 #(
		.INIT('hc7b6)
	) name18173 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w24000_
	);
	LUT2 #(
		.INIT('h1)
	) name18174 (
		_w23907_,
		_w23906_,
		_w24001_
	);
	LUT2 #(
		.INIT('h4)
	) name18175 (
		_w24000_,
		_w24001_,
		_w24002_
	);
	LUT3 #(
		.INIT('hdb)
	) name18176 (
		_w23908_,
		_w23911_,
		_w23909_,
		_w24003_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name18177 (
		_w23910_,
		_w23906_,
		_w23960_,
		_w24003_,
		_w24004_
	);
	LUT2 #(
		.INIT('h4)
	) name18178 (
		_w24002_,
		_w24004_,
		_w24005_
	);
	LUT4 #(
		.INIT('h5655)
	) name18179 (
		\u1_L0_reg[24]/NET0131 ,
		_w23998_,
		_w23992_,
		_w24005_,
		_w24006_
	);
	LUT4 #(
		.INIT('h0010)
	) name18180 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w24007_
	);
	LUT4 #(
		.INIT('hf900)
	) name18181 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23906_,
		_w24008_
	);
	LUT3 #(
		.INIT('h07)
	) name18182 (
		_w23910_,
		_w23911_,
		_w23906_,
		_w24009_
	);
	LUT4 #(
		.INIT('h8acf)
	) name18183 (
		_w23927_,
		_w24007_,
		_w24008_,
		_w24009_,
		_w24010_
	);
	LUT2 #(
		.INIT('h2)
	) name18184 (
		_w23907_,
		_w24010_,
		_w24011_
	);
	LUT3 #(
		.INIT('h10)
	) name18185 (
		_w23910_,
		_w23908_,
		_w23909_,
		_w24012_
	);
	LUT4 #(
		.INIT('h80a0)
	) name18186 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w24013_
	);
	LUT3 #(
		.INIT('h02)
	) name18187 (
		_w23906_,
		_w24013_,
		_w24012_,
		_w24014_
	);
	LUT4 #(
		.INIT('h4050)
	) name18188 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w24015_
	);
	LUT4 #(
		.INIT('h00df)
	) name18189 (
		_w23908_,
		_w23911_,
		_w23909_,
		_w23906_,
		_w24016_
	);
	LUT2 #(
		.INIT('h4)
	) name18190 (
		_w24015_,
		_w24016_,
		_w24017_
	);
	LUT4 #(
		.INIT('h0008)
	) name18191 (
		_w23910_,
		_w23908_,
		_w23911_,
		_w23909_,
		_w24018_
	);
	LUT3 #(
		.INIT('h01)
	) name18192 (
		_w23907_,
		_w23999_,
		_w24018_,
		_w24019_
	);
	LUT3 #(
		.INIT('he0)
	) name18193 (
		_w24014_,
		_w24017_,
		_w24019_,
		_w24020_
	);
	LUT3 #(
		.INIT('h80)
	) name18194 (
		_w23907_,
		_w23910_,
		_w23909_,
		_w24021_
	);
	LUT4 #(
		.INIT('h0020)
	) name18195 (
		_w23910_,
		_w23908_,
		_w23909_,
		_w23906_,
		_w24022_
	);
	LUT3 #(
		.INIT('h20)
	) name18196 (
		_w23910_,
		_w23909_,
		_w23906_,
		_w24023_
	);
	LUT4 #(
		.INIT('h0213)
	) name18197 (
		_w23920_,
		_w24022_,
		_w24023_,
		_w24021_,
		_w24024_
	);
	LUT4 #(
		.INIT('h56aa)
	) name18198 (
		\u1_L0_reg[30]/NET0131 ,
		_w24011_,
		_w24020_,
		_w24024_,
		_w24025_
	);
	LUT4 #(
		.INIT('h0004)
	) name18199 (
		_w23650_,
		_w23629_,
		_w23641_,
		_w23638_,
		_w24026_
	);
	LUT4 #(
		.INIT('h080c)
	) name18200 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w24027_
	);
	LUT4 #(
		.INIT('h7522)
	) name18201 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w24028_
	);
	LUT3 #(
		.INIT('h10)
	) name18202 (
		_w23629_,
		_w24027_,
		_w24028_,
		_w24029_
	);
	LUT4 #(
		.INIT('h0800)
	) name18203 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w24030_
	);
	LUT4 #(
		.INIT('h0001)
	) name18204 (
		_w23630_,
		_w23644_,
		_w23952_,
		_w24030_,
		_w24031_
	);
	LUT3 #(
		.INIT('he0)
	) name18205 (
		_w24026_,
		_w24029_,
		_w24031_,
		_w24032_
	);
	LUT4 #(
		.INIT('hddaf)
	) name18206 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w24033_
	);
	LUT4 #(
		.INIT('h0400)
	) name18207 (
		_w23650_,
		_w23629_,
		_w23641_,
		_w24033_,
		_w24034_
	);
	LUT4 #(
		.INIT('hafdd)
	) name18208 (
		_w23631_,
		_w23634_,
		_w23632_,
		_w23633_,
		_w24035_
	);
	LUT3 #(
		.INIT('h10)
	) name18209 (
		_w23629_,
		_w24027_,
		_w24035_,
		_w24036_
	);
	LUT3 #(
		.INIT('h04)
	) name18210 (
		_w23652_,
		_w23630_,
		_w23659_,
		_w24037_
	);
	LUT3 #(
		.INIT('he0)
	) name18211 (
		_w24034_,
		_w24036_,
		_w24037_,
		_w24038_
	);
	LUT3 #(
		.INIT('ha9)
	) name18212 (
		\u1_L0_reg[3]/NET0131 ,
		_w24032_,
		_w24038_,
		_w24039_
	);
	LUT4 #(
		.INIT('hf04f)
	) name18213 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w24040_
	);
	LUT3 #(
		.INIT('hbc)
	) name18214 (
		_w23576_,
		_w23573_,
		_w23574_,
		_w24041_
	);
	LUT4 #(
		.INIT('hb7fd)
	) name18215 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w24042_
	);
	LUT4 #(
		.INIT('hd800)
	) name18216 (
		_w23572_,
		_w24040_,
		_w24041_,
		_w24042_,
		_w24043_
	);
	LUT4 #(
		.INIT('h9fff)
	) name18217 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w24044_
	);
	LUT2 #(
		.INIT('h1)
	) name18218 (
		_w23572_,
		_w24044_,
		_w24045_
	);
	LUT4 #(
		.INIT('h8228)
	) name18219 (
		_w23575_,
		_w23576_,
		_w23573_,
		_w23574_,
		_w24046_
	);
	LUT4 #(
		.INIT('h0031)
	) name18220 (
		_w23580_,
		_w23861_,
		_w24041_,
		_w24046_,
		_w24047_
	);
	LUT4 #(
		.INIT('h0e04)
	) name18221 (
		_w23571_,
		_w24043_,
		_w24045_,
		_w24047_,
		_w24048_
	);
	LUT2 #(
		.INIT('h9)
	) name18222 (
		\u1_L0_reg[9]/NET0131 ,
		_w24048_,
		_w24049_
	);
	LUT4 #(
		.INIT('h3400)
	) name18223 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23762_,
		_w24050_
	);
	LUT3 #(
		.INIT('h13)
	) name18224 (
		_w23757_,
		_w23762_,
		_w23763_,
		_w24051_
	);
	LUT4 #(
		.INIT('h0103)
	) name18225 (
		_w23760_,
		_w23816_,
		_w24050_,
		_w24051_,
		_w24052_
	);
	LUT4 #(
		.INIT('h2800)
	) name18226 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w24053_
	);
	LUT4 #(
		.INIT('h0411)
	) name18227 (
		_w23759_,
		_w23758_,
		_w23762_,
		_w23763_,
		_w24054_
	);
	LUT4 #(
		.INIT('h8000)
	) name18228 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23762_,
		_w24055_
	);
	LUT4 #(
		.INIT('h0001)
	) name18229 (
		_w23810_,
		_w24054_,
		_w24053_,
		_w24055_,
		_w24056_
	);
	LUT4 #(
		.INIT('h0040)
	) name18230 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23762_,
		_w24057_
	);
	LUT4 #(
		.INIT('h77ef)
	) name18231 (
		_w23759_,
		_w23757_,
		_w23758_,
		_w23763_,
		_w24058_
	);
	LUT3 #(
		.INIT('h31)
	) name18232 (
		_w23762_,
		_w24057_,
		_w24058_,
		_w24059_
	);
	LUT4 #(
		.INIT('he400)
	) name18233 (
		_w23774_,
		_w24056_,
		_w24052_,
		_w24059_,
		_w24060_
	);
	LUT2 #(
		.INIT('h9)
	) name18234 (
		\u1_L0_reg[18]/NET0131 ,
		_w24060_,
		_w24061_
	);
	LUT4 #(
		.INIT('hc693)
	) name18235 (
		decrypt_pad,
		\u1_desIn_r_reg[31]/NET0131 ,
		\u1_key_r_reg[13]/NET0131 ,
		\u1_key_r_reg[6]/NET0131 ,
		_w24062_
	);
	LUT4 #(
		.INIT('hc963)
	) name18236 (
		decrypt_pad,
		\u1_desIn_r_reg[57]/NET0131 ,
		\u1_key_r_reg[40]/NET0131 ,
		\u1_key_r_reg[47]/NET0131 ,
		_w24063_
	);
	LUT4 #(
		.INIT('hc693)
	) name18237 (
		decrypt_pad,
		\u1_desIn_r_reg[7]/NET0131 ,
		\u1_key_r_reg[11]/NET0131 ,
		\u1_key_r_reg[4]/NET0131 ,
		_w24064_
	);
	LUT4 #(
		.INIT('hc963)
	) name18238 (
		decrypt_pad,
		\u1_desIn_r_reg[15]/NET0131 ,
		\u1_key_r_reg[19]/NET0131 ,
		\u1_key_r_reg[26]/NET0131 ,
		_w24065_
	);
	LUT4 #(
		.INIT('hc963)
	) name18239 (
		decrypt_pad,
		\u1_desIn_r_reg[39]/NET0131 ,
		\u1_key_r_reg[34]/NET0131 ,
		\u1_key_r_reg[41]/NET0131 ,
		_w24066_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name18240 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24067_
	);
	LUT2 #(
		.INIT('h1)
	) name18241 (
		_w24066_,
		_w24063_,
		_w24068_
	);
	LUT4 #(
		.INIT('hc693)
	) name18242 (
		decrypt_pad,
		\u1_desIn_r_reg[23]/NET0131 ,
		\u1_key_r_reg[3]/NET0131 ,
		\u1_key_r_reg[53]/NET0131 ,
		_w24069_
	);
	LUT2 #(
		.INIT('h4)
	) name18243 (
		_w24065_,
		_w24069_,
		_w24070_
	);
	LUT3 #(
		.INIT('hb0)
	) name18244 (
		_w24065_,
		_w24069_,
		_w24064_,
		_w24071_
	);
	LUT3 #(
		.INIT('h01)
	) name18245 (
		_w24068_,
		_w24071_,
		_w24067_,
		_w24072_
	);
	LUT3 #(
		.INIT('h02)
	) name18246 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24073_
	);
	LUT4 #(
		.INIT('hfd31)
	) name18247 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24074_
	);
	LUT4 #(
		.INIT('h300a)
	) name18248 (
		_w24065_,
		_w24069_,
		_w24063_,
		_w24064_,
		_w24075_
	);
	LUT3 #(
		.INIT('h0d)
	) name18249 (
		_w24069_,
		_w24074_,
		_w24075_,
		_w24076_
	);
	LUT3 #(
		.INIT('h8a)
	) name18250 (
		_w24062_,
		_w24072_,
		_w24076_,
		_w24077_
	);
	LUT3 #(
		.INIT('he6)
	) name18251 (
		_w24065_,
		_w24063_,
		_w24064_,
		_w24078_
	);
	LUT3 #(
		.INIT('h51)
	) name18252 (
		_w24069_,
		_w24066_,
		_w24064_,
		_w24079_
	);
	LUT2 #(
		.INIT('h4)
	) name18253 (
		_w24078_,
		_w24079_,
		_w24080_
	);
	LUT2 #(
		.INIT('h8)
	) name18254 (
		_w24065_,
		_w24069_,
		_w24081_
	);
	LUT3 #(
		.INIT('h60)
	) name18255 (
		_w24066_,
		_w24063_,
		_w24064_,
		_w24082_
	);
	LUT4 #(
		.INIT('h7c3f)
	) name18256 (
		_w24069_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24083_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name18257 (
		_w24065_,
		_w24069_,
		_w24082_,
		_w24083_,
		_w24084_
	);
	LUT2 #(
		.INIT('h2)
	) name18258 (
		_w24069_,
		_w24064_,
		_w24085_
	);
	LUT3 #(
		.INIT('had)
	) name18259 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24086_
	);
	LUT4 #(
		.INIT('h8000)
	) name18260 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24087_
	);
	LUT4 #(
		.INIT('h0008)
	) name18261 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24088_
	);
	LUT4 #(
		.INIT('h6ef7)
	) name18262 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24089_
	);
	LUT4 #(
		.INIT('hfda8)
	) name18263 (
		_w24069_,
		_w24064_,
		_w24086_,
		_w24089_,
		_w24090_
	);
	LUT4 #(
		.INIT('hba00)
	) name18264 (
		_w24062_,
		_w24080_,
		_w24084_,
		_w24090_,
		_w24091_
	);
	LUT3 #(
		.INIT('h65)
	) name18265 (
		\u1_desIn_r_reg[48]/NET0131 ,
		_w24077_,
		_w24091_,
		_w24092_
	);
	LUT4 #(
		.INIT('hc963)
	) name18266 (
		decrypt_pad,
		\u1_desIn_r_reg[51]/NET0131 ,
		\u1_key_r_reg[2]/NET0131 ,
		\u1_key_r_reg[9]/NET0131 ,
		_w24093_
	);
	LUT4 #(
		.INIT('hc963)
	) name18267 (
		decrypt_pad,
		\u1_desIn_r_reg[59]/NET0131 ,
		\u1_key_r_reg[28]/NET0131 ,
		\u1_key_r_reg[35]/P0001 ,
		_w24094_
	);
	LUT4 #(
		.INIT('hc963)
	) name18268 (
		decrypt_pad,
		\u1_desIn_r_reg[35]/NET0131 ,
		\u1_key_r_reg[22]/NET0131 ,
		\u1_key_r_reg[29]/NET0131 ,
		_w24095_
	);
	LUT4 #(
		.INIT('hc963)
	) name18269 (
		decrypt_pad,
		\u1_desIn_r_reg[43]/NET0131 ,
		\u1_key_r_reg[44]/NET0131 ,
		\u1_key_r_reg[51]/NET0131 ,
		_w24096_
	);
	LUT4 #(
		.INIT('hc693)
	) name18270 (
		decrypt_pad,
		\u1_desIn_r_reg[27]/NET0131 ,
		\u1_key_r_reg[14]/NET0131 ,
		\u1_key_r_reg[7]/NET0131 ,
		_w24097_
	);
	LUT4 #(
		.INIT('hc963)
	) name18271 (
		decrypt_pad,
		\u1_desIn_r_reg[1]/NET0131 ,
		\u1_key_r_reg[23]/NET0131 ,
		\u1_key_r_reg[30]/NET0131 ,
		_w24098_
	);
	LUT4 #(
		.INIT('h57e7)
	) name18272 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24099_
	);
	LUT4 #(
		.INIT('h0002)
	) name18273 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24100_
	);
	LUT4 #(
		.INIT('h3efd)
	) name18274 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24101_
	);
	LUT4 #(
		.INIT('h08aa)
	) name18275 (
		_w24093_,
		_w24094_,
		_w24099_,
		_w24101_,
		_w24102_
	);
	LUT4 #(
		.INIT('h00f7)
	) name18276 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24093_,
		_w24103_
	);
	LUT4 #(
		.INIT('h00d7)
	) name18277 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24093_,
		_w24104_
	);
	LUT3 #(
		.INIT('h54)
	) name18278 (
		_w24095_,
		_w24097_,
		_w24098_,
		_w24105_
	);
	LUT4 #(
		.INIT('h4440)
	) name18279 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24106_
	);
	LUT3 #(
		.INIT('he0)
	) name18280 (
		_w24096_,
		_w24097_,
		_w24093_,
		_w24107_
	);
	LUT3 #(
		.INIT('h45)
	) name18281 (
		_w24104_,
		_w24106_,
		_w24107_,
		_w24108_
	);
	LUT4 #(
		.INIT('h4000)
	) name18282 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24109_
	);
	LUT2 #(
		.INIT('h1)
	) name18283 (
		_w24096_,
		_w24093_,
		_w24110_
	);
	LUT4 #(
		.INIT('h0004)
	) name18284 (
		_w24096_,
		_w24097_,
		_w24093_,
		_w24098_,
		_w24111_
	);
	LUT4 #(
		.INIT('h0020)
	) name18285 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24112_
	);
	LUT3 #(
		.INIT('h01)
	) name18286 (
		_w24109_,
		_w24111_,
		_w24112_,
		_w24113_
	);
	LUT3 #(
		.INIT('h0b)
	) name18287 (
		_w24108_,
		_w24113_,
		_w24094_,
		_w24114_
	);
	LUT4 #(
		.INIT('h2133)
	) name18288 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24115_
	);
	LUT4 #(
		.INIT('h7f00)
	) name18289 (
		_w24096_,
		_w24097_,
		_w24098_,
		_w24094_,
		_w24116_
	);
	LUT3 #(
		.INIT('h20)
	) name18290 (
		_w24103_,
		_w24115_,
		_w24116_,
		_w24117_
	);
	LUT3 #(
		.INIT('ha2)
	) name18291 (
		_w24095_,
		_w24097_,
		_w24098_,
		_w24118_
	);
	LUT3 #(
		.INIT('h04)
	) name18292 (
		_w24105_,
		_w24110_,
		_w24118_,
		_w24119_
	);
	LUT2 #(
		.INIT('h1)
	) name18293 (
		_w24117_,
		_w24119_,
		_w24120_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name18294 (
		\u1_desIn_r_reg[20]/NET0131 ,
		_w24114_,
		_w24102_,
		_w24120_,
		_w24121_
	);
	LUT4 #(
		.INIT('hc963)
	) name18295 (
		decrypt_pad,
		\u1_desIn_r_reg[9]/NET0131 ,
		\u1_key_r_reg[15]/NET0131 ,
		\u1_key_r_reg[22]/NET0131 ,
		_w24122_
	);
	LUT4 #(
		.INIT('hc963)
	) name18296 (
		decrypt_pad,
		\u1_desIn_r_reg[1]/NET0131 ,
		\u1_key_r_reg[30]/NET0131 ,
		\u1_key_r_reg[37]/NET0131 ,
		_w24123_
	);
	LUT4 #(
		.INIT('hc693)
	) name18297 (
		decrypt_pad,
		\u1_desIn_r_reg[59]/NET0131 ,
		\u1_key_r_reg[2]/NET0131 ,
		\u1_key_r_reg[50]/NET0131 ,
		_w24124_
	);
	LUT4 #(
		.INIT('hc963)
	) name18298 (
		decrypt_pad,
		\u1_desIn_r_reg[33]/NET0131 ,
		\u1_key_r_reg[31]/NET0131 ,
		\u1_key_r_reg[38]/NET0131 ,
		_w24125_
	);
	LUT2 #(
		.INIT('h4)
	) name18299 (
		_w24124_,
		_w24125_,
		_w24126_
	);
	LUT4 #(
		.INIT('h0200)
	) name18300 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24127_
	);
	LUT4 #(
		.INIT('h0008)
	) name18301 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24128_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name18302 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24129_
	);
	LUT4 #(
		.INIT('hc963)
	) name18303 (
		decrypt_pad,
		\u1_desIn_r_reg[25]/NET0131 ,
		\u1_key_r_reg[35]/P0001 ,
		\u1_key_r_reg[42]/P0001 ,
		_w24130_
	);
	LUT4 #(
		.INIT('h9cfc)
	) name18304 (
		_w24122_,
		_w24123_,
		_w24125_,
		_w24130_,
		_w24131_
	);
	LUT4 #(
		.INIT('hc693)
	) name18305 (
		decrypt_pad,
		\u1_desIn_r_reg[17]/NET0131 ,
		\u1_key_r_reg[0]/NET0131 ,
		\u1_key_r_reg[52]/NET0131 ,
		_w24132_
	);
	LUT4 #(
		.INIT('h3b00)
	) name18306 (
		_w24124_,
		_w24129_,
		_w24131_,
		_w24132_,
		_w24133_
	);
	LUT4 #(
		.INIT('hee72)
	) name18307 (
		_w24122_,
		_w24123_,
		_w24125_,
		_w24132_,
		_w24134_
	);
	LUT2 #(
		.INIT('h2)
	) name18308 (
		_w24124_,
		_w24134_,
		_w24135_
	);
	LUT4 #(
		.INIT('h0002)
	) name18309 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24136_
	);
	LUT2 #(
		.INIT('h6)
	) name18310 (
		_w24122_,
		_w24124_,
		_w24137_
	);
	LUT3 #(
		.INIT('h8c)
	) name18311 (
		_w24123_,
		_w24125_,
		_w24132_,
		_w24138_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name18312 (
		_w24132_,
		_w24136_,
		_w24137_,
		_w24138_,
		_w24139_
	);
	LUT3 #(
		.INIT('h45)
	) name18313 (
		_w24130_,
		_w24135_,
		_w24139_,
		_w24140_
	);
	LUT4 #(
		.INIT('h1000)
	) name18314 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24141_
	);
	LUT4 #(
		.INIT('he3ff)
	) name18315 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24142_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name18316 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24143_
	);
	LUT4 #(
		.INIT('h02aa)
	) name18317 (
		_w24130_,
		_w24132_,
		_w24142_,
		_w24143_,
		_w24144_
	);
	LUT4 #(
		.INIT('h0084)
	) name18318 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24132_,
		_w24145_
	);
	LUT4 #(
		.INIT('h0100)
	) name18319 (
		_w24122_,
		_w24123_,
		_w24125_,
		_w24132_,
		_w24146_
	);
	LUT2 #(
		.INIT('h1)
	) name18320 (
		_w24145_,
		_w24146_,
		_w24147_
	);
	LUT2 #(
		.INIT('h4)
	) name18321 (
		_w24144_,
		_w24147_,
		_w24148_
	);
	LUT4 #(
		.INIT('h5655)
	) name18322 (
		\u1_desIn_r_reg[42]/NET0131 ,
		_w24133_,
		_w24140_,
		_w24148_,
		_w24149_
	);
	LUT4 #(
		.INIT('hfe3c)
	) name18323 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24150_
	);
	LUT2 #(
		.INIT('h1)
	) name18324 (
		_w24069_,
		_w24150_,
		_w24151_
	);
	LUT4 #(
		.INIT('h35f3)
	) name18325 (
		_w24065_,
		_w24069_,
		_w24066_,
		_w24064_,
		_w24152_
	);
	LUT4 #(
		.INIT('h0501)
	) name18326 (
		_w24062_,
		_w24063_,
		_w24088_,
		_w24152_,
		_w24153_
	);
	LUT4 #(
		.INIT('h0040)
	) name18327 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24154_
	);
	LUT4 #(
		.INIT('hf0b5)
	) name18328 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24155_
	);
	LUT2 #(
		.INIT('h2)
	) name18329 (
		_w24069_,
		_w24155_,
		_w24156_
	);
	LUT4 #(
		.INIT('h1000)
	) name18330 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24157_
	);
	LUT4 #(
		.INIT('h2021)
	) name18331 (
		_w24065_,
		_w24069_,
		_w24063_,
		_w24064_,
		_w24158_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name18332 (
		_w24062_,
		_w24065_,
		_w24066_,
		_w24064_,
		_w24159_
	);
	LUT3 #(
		.INIT('h10)
	) name18333 (
		_w24158_,
		_w24157_,
		_w24159_,
		_w24160_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name18334 (
		_w24151_,
		_w24153_,
		_w24156_,
		_w24160_,
		_w24161_
	);
	LUT3 #(
		.INIT('he0)
	) name18335 (
		_w24065_,
		_w24066_,
		_w24064_,
		_w24162_
	);
	LUT4 #(
		.INIT('h004c)
	) name18336 (
		_w24065_,
		_w24069_,
		_w24066_,
		_w24063_,
		_w24163_
	);
	LUT2 #(
		.INIT('h8)
	) name18337 (
		_w24162_,
		_w24163_,
		_w24164_
	);
	LUT3 #(
		.INIT('h56)
	) name18338 (
		\u1_desIn_r_reg[2]/NET0131 ,
		_w24161_,
		_w24164_,
		_w24165_
	);
	LUT4 #(
		.INIT('h2e25)
	) name18339 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24166_
	);
	LUT2 #(
		.INIT('h2)
	) name18340 (
		_w24093_,
		_w24166_,
		_w24167_
	);
	LUT2 #(
		.INIT('h6)
	) name18341 (
		_w24095_,
		_w24098_,
		_w24168_
	);
	LUT4 #(
		.INIT('h0201)
	) name18342 (
		_w24095_,
		_w24097_,
		_w24093_,
		_w24098_,
		_w24169_
	);
	LUT4 #(
		.INIT('h8000)
	) name18343 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24170_
	);
	LUT3 #(
		.INIT('h01)
	) name18344 (
		_w24094_,
		_w24170_,
		_w24169_,
		_w24171_
	);
	LUT4 #(
		.INIT('hdadf)
	) name18345 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24172_
	);
	LUT2 #(
		.INIT('h2)
	) name18346 (
		_w24093_,
		_w24172_,
		_w24173_
	);
	LUT3 #(
		.INIT('h04)
	) name18347 (
		_w24095_,
		_w24097_,
		_w24093_,
		_w24174_
	);
	LUT4 #(
		.INIT('hfd00)
	) name18348 (
		_w24095_,
		_w24096_,
		_w24098_,
		_w24094_,
		_w24175_
	);
	LUT4 #(
		.INIT('hf6fb)
	) name18349 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24176_
	);
	LUT3 #(
		.INIT('h40)
	) name18350 (
		_w24174_,
		_w24175_,
		_w24176_,
		_w24177_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name18351 (
		_w24167_,
		_w24171_,
		_w24173_,
		_w24177_,
		_w24178_
	);
	LUT3 #(
		.INIT('h04)
	) name18352 (
		_w24096_,
		_w24097_,
		_w24093_,
		_w24179_
	);
	LUT2 #(
		.INIT('h8)
	) name18353 (
		_w24168_,
		_w24179_,
		_w24180_
	);
	LUT3 #(
		.INIT('h56)
	) name18354 (
		\u1_desIn_r_reg[18]/P0001 ,
		_w24178_,
		_w24180_,
		_w24181_
	);
	LUT4 #(
		.INIT('hc963)
	) name18355 (
		decrypt_pad,
		\u1_desIn_r_reg[37]/NET0131 ,
		\u1_key_r_reg[48]/NET0131 ,
		\u1_key_r_reg[55]/NET0131 ,
		_w24182_
	);
	LUT4 #(
		.INIT('hc693)
	) name18356 (
		decrypt_pad,
		\u1_desIn_r_reg[29]/NET0131 ,
		\u1_key_r_reg[4]/NET0131 ,
		\u1_key_r_reg[54]/NET0131 ,
		_w24183_
	);
	LUT2 #(
		.INIT('h2)
	) name18357 (
		_w24182_,
		_w24183_,
		_w24184_
	);
	LUT2 #(
		.INIT('h9)
	) name18358 (
		_w24182_,
		_w24183_,
		_w24185_
	);
	LUT4 #(
		.INIT('hc963)
	) name18359 (
		decrypt_pad,
		\u1_desIn_r_reg[53]/NET0131 ,
		\u1_key_r_reg[25]/NET0131 ,
		\u1_key_r_reg[32]/NET0131 ,
		_w24186_
	);
	LUT4 #(
		.INIT('hc963)
	) name18360 (
		decrypt_pad,
		\u1_desIn_r_reg[45]/NET0131 ,
		\u1_key_r_reg[17]/NET0131 ,
		\u1_key_r_reg[24]/NET0131 ,
		_w24187_
	);
	LUT4 #(
		.INIT('h0012)
	) name18361 (
		_w24182_,
		_w24186_,
		_w24183_,
		_w24187_,
		_w24188_
	);
	LUT4 #(
		.INIT('hc963)
	) name18362 (
		decrypt_pad,
		\u1_desIn_r_reg[3]/NET0131 ,
		\u1_key_r_reg[13]/NET0131 ,
		\u1_key_r_reg[20]/NET0131 ,
		_w24189_
	);
	LUT2 #(
		.INIT('h8)
	) name18363 (
		_w24182_,
		_w24186_,
		_w24190_
	);
	LUT4 #(
		.INIT('h0080)
	) name18364 (
		_w24182_,
		_w24186_,
		_w24183_,
		_w24189_,
		_w24191_
	);
	LUT2 #(
		.INIT('h4)
	) name18365 (
		_w24182_,
		_w24186_,
		_w24192_
	);
	LUT2 #(
		.INIT('h4)
	) name18366 (
		_w24183_,
		_w24189_,
		_w24193_
	);
	LUT4 #(
		.INIT('h0400)
	) name18367 (
		_w24182_,
		_w24186_,
		_w24183_,
		_w24189_,
		_w24194_
	);
	LUT4 #(
		.INIT('hc963)
	) name18368 (
		decrypt_pad,
		\u1_desIn_r_reg[61]/NET0131 ,
		\u1_key_r_reg[33]/NET0131 ,
		\u1_key_r_reg[40]/NET0131 ,
		_w24195_
	);
	LUT4 #(
		.INIT('h0010)
	) name18369 (
		_w24194_,
		_w24191_,
		_w24195_,
		_w24188_,
		_w24196_
	);
	LUT4 #(
		.INIT('h0001)
	) name18370 (
		_w24182_,
		_w24186_,
		_w24183_,
		_w24189_,
		_w24197_
	);
	LUT4 #(
		.INIT('h0020)
	) name18371 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24198_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name18372 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24199_
	);
	LUT3 #(
		.INIT('h70)
	) name18373 (
		_w24197_,
		_w24187_,
		_w24199_,
		_w24200_
	);
	LUT2 #(
		.INIT('h8)
	) name18374 (
		_w24196_,
		_w24200_,
		_w24201_
	);
	LUT3 #(
		.INIT('h04)
	) name18375 (
		_w24182_,
		_w24183_,
		_w24187_,
		_w24202_
	);
	LUT4 #(
		.INIT('h0040)
	) name18376 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24203_
	);
	LUT4 #(
		.INIT('h8000)
	) name18377 (
		_w24182_,
		_w24186_,
		_w24183_,
		_w24189_,
		_w24204_
	);
	LUT3 #(
		.INIT('h01)
	) name18378 (
		_w24195_,
		_w24203_,
		_w24204_,
		_w24205_
	);
	LUT4 #(
		.INIT('h0004)
	) name18379 (
		_w24182_,
		_w24186_,
		_w24183_,
		_w24189_,
		_w24206_
	);
	LUT3 #(
		.INIT('h80)
	) name18380 (
		_w24182_,
		_w24186_,
		_w24187_,
		_w24207_
	);
	LUT4 #(
		.INIT('h0800)
	) name18381 (
		_w24182_,
		_w24186_,
		_w24183_,
		_w24187_,
		_w24208_
	);
	LUT2 #(
		.INIT('h1)
	) name18382 (
		_w24206_,
		_w24208_,
		_w24209_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name18383 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24210_
	);
	LUT4 #(
		.INIT('ha3af)
	) name18384 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24211_
	);
	LUT3 #(
		.INIT('hc8)
	) name18385 (
		_w24186_,
		_w24210_,
		_w24211_,
		_w24212_
	);
	LUT3 #(
		.INIT('h80)
	) name18386 (
		_w24205_,
		_w24209_,
		_w24212_,
		_w24213_
	);
	LUT3 #(
		.INIT('hde)
	) name18387 (
		_w24183_,
		_w24189_,
		_w24187_,
		_w24214_
	);
	LUT2 #(
		.INIT('h2)
	) name18388 (
		_w24192_,
		_w24214_,
		_w24215_
	);
	LUT2 #(
		.INIT('h2)
	) name18389 (
		_w24189_,
		_w24187_,
		_w24216_
	);
	LUT3 #(
		.INIT('h04)
	) name18390 (
		_w24186_,
		_w24189_,
		_w24187_,
		_w24217_
	);
	LUT3 #(
		.INIT('h02)
	) name18391 (
		_w24183_,
		_w24189_,
		_w24187_,
		_w24218_
	);
	LUT4 #(
		.INIT('h153f)
	) name18392 (
		_w24190_,
		_w24184_,
		_w24217_,
		_w24218_,
		_w24219_
	);
	LUT2 #(
		.INIT('h4)
	) name18393 (
		_w24215_,
		_w24219_,
		_w24220_
	);
	LUT4 #(
		.INIT('ha955)
	) name18394 (
		\u1_desIn_r_reg[26]/NET0131 ,
		_w24201_,
		_w24213_,
		_w24220_,
		_w24221_
	);
	LUT4 #(
		.INIT('hcd7d)
	) name18395 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24222_
	);
	LUT4 #(
		.INIT('h5fa6)
	) name18396 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24223_
	);
	LUT4 #(
		.INIT('h0400)
	) name18397 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24224_
	);
	LUT4 #(
		.INIT('h00d8)
	) name18398 (
		_w24093_,
		_w24223_,
		_w24222_,
		_w24224_,
		_w24225_
	);
	LUT2 #(
		.INIT('h1)
	) name18399 (
		_w24094_,
		_w24225_,
		_w24226_
	);
	LUT4 #(
		.INIT('hf57d)
	) name18400 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24227_
	);
	LUT2 #(
		.INIT('h2)
	) name18401 (
		_w24093_,
		_w24227_,
		_w24228_
	);
	LUT2 #(
		.INIT('h6)
	) name18402 (
		_w24097_,
		_w24098_,
		_w24229_
	);
	LUT4 #(
		.INIT('h0c0d)
	) name18403 (
		_w24095_,
		_w24096_,
		_w24093_,
		_w24098_,
		_w24230_
	);
	LUT2 #(
		.INIT('h4)
	) name18404 (
		_w24229_,
		_w24230_,
		_w24231_
	);
	LUT4 #(
		.INIT('hfefb)
	) name18405 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24232_
	);
	LUT3 #(
		.INIT('h10)
	) name18406 (
		_w24109_,
		_w24111_,
		_w24232_,
		_w24233_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name18407 (
		_w24094_,
		_w24228_,
		_w24231_,
		_w24233_,
		_w24234_
	);
	LUT4 #(
		.INIT('h0010)
	) name18408 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24235_
	);
	LUT4 #(
		.INIT('h2000)
	) name18409 (
		_w24095_,
		_w24096_,
		_w24093_,
		_w24098_,
		_w24236_
	);
	LUT2 #(
		.INIT('h1)
	) name18410 (
		_w24235_,
		_w24236_,
		_w24237_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name18411 (
		\u1_desIn_r_reg[32]/NET0131 ,
		_w24234_,
		_w24226_,
		_w24237_,
		_w24238_
	);
	LUT4 #(
		.INIT('hc963)
	) name18412 (
		decrypt_pad,
		\u1_desIn_r_reg[63]/NET0131 ,
		\u1_key_r_reg[32]/NET0131 ,
		\u1_key_r_reg[39]/P0001 ,
		_w24239_
	);
	LUT4 #(
		.INIT('hc963)
	) name18413 (
		decrypt_pad,
		\u1_desIn_r_reg[55]/NET0131 ,
		\u1_key_r_reg[41]/NET0131 ,
		\u1_key_r_reg[48]/NET0131 ,
		_w24240_
	);
	LUT4 #(
		.INIT('hc963)
	) name18414 (
		decrypt_pad,
		\u1_desIn_r_reg[39]/NET0131 ,
		\u1_key_r_reg[24]/NET0131 ,
		\u1_key_r_reg[6]/NET0131 ,
		_w24241_
	);
	LUT4 #(
		.INIT('hc963)
	) name18415 (
		decrypt_pad,
		\u1_desIn_r_reg[31]/NET0131 ,
		\u1_key_r_reg[20]/NET0131 ,
		\u1_key_r_reg[27]/NET0131 ,
		_w24242_
	);
	LUT4 #(
		.INIT('hc963)
	) name18416 (
		decrypt_pad,
		\u1_desIn_r_reg[5]/NET0131 ,
		\u1_key_r_reg[12]/NET0131 ,
		\u1_key_r_reg[19]/NET0131 ,
		_w24243_
	);
	LUT4 #(
		.INIT('hc963)
	) name18417 (
		decrypt_pad,
		\u1_desIn_r_reg[47]/NET0131 ,
		\u1_key_r_reg[47]/NET0131 ,
		\u1_key_r_reg[54]/NET0131 ,
		_w24244_
	);
	LUT4 #(
		.INIT('h59fb)
	) name18418 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24245_
	);
	LUT2 #(
		.INIT('h1)
	) name18419 (
		_w24240_,
		_w24245_,
		_w24246_
	);
	LUT4 #(
		.INIT('h0034)
	) name18420 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24247_
	);
	LUT4 #(
		.INIT('h0800)
	) name18421 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24248_
	);
	LUT2 #(
		.INIT('h2)
	) name18422 (
		_w24243_,
		_w24244_,
		_w24249_
	);
	LUT4 #(
		.INIT('h0004)
	) name18423 (
		_w24240_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24250_
	);
	LUT4 #(
		.INIT('h4000)
	) name18424 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24251_
	);
	LUT4 #(
		.INIT('h0007)
	) name18425 (
		_w24240_,
		_w24248_,
		_w24250_,
		_w24251_,
		_w24252_
	);
	LUT4 #(
		.INIT('h5455)
	) name18426 (
		_w24239_,
		_w24246_,
		_w24247_,
		_w24252_,
		_w24253_
	);
	LUT4 #(
		.INIT('he6ee)
	) name18427 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24254_
	);
	LUT4 #(
		.INIT('h4044)
	) name18428 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24255_
	);
	LUT3 #(
		.INIT('h51)
	) name18429 (
		_w24240_,
		_w24241_,
		_w24244_,
		_w24256_
	);
	LUT4 #(
		.INIT('hf200)
	) name18430 (
		_w24239_,
		_w24254_,
		_w24255_,
		_w24256_,
		_w24257_
	);
	LUT3 #(
		.INIT('h10)
	) name18431 (
		_w24243_,
		_w24241_,
		_w24244_,
		_w24258_
	);
	LUT4 #(
		.INIT('h0100)
	) name18432 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24259_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name18433 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24260_
	);
	LUT2 #(
		.INIT('h2)
	) name18434 (
		_w24240_,
		_w24260_,
		_w24261_
	);
	LUT4 #(
		.INIT('h0082)
	) name18435 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24262_
	);
	LUT4 #(
		.INIT('h80a0)
	) name18436 (
		_w24240_,
		_w24242_,
		_w24241_,
		_w24244_,
		_w24263_
	);
	LUT3 #(
		.INIT('ha8)
	) name18437 (
		_w24239_,
		_w24262_,
		_w24263_,
		_w24264_
	);
	LUT3 #(
		.INIT('h01)
	) name18438 (
		_w24261_,
		_w24264_,
		_w24257_,
		_w24265_
	);
	LUT3 #(
		.INIT('h65)
	) name18439 (
		\u1_desIn_r_reg[14]/NET0131 ,
		_w24253_,
		_w24265_,
		_w24266_
	);
	LUT4 #(
		.INIT('h2090)
	) name18440 (
		_w24095_,
		_w24097_,
		_w24093_,
		_w24098_,
		_w24267_
	);
	LUT4 #(
		.INIT('h0804)
	) name18441 (
		_w24095_,
		_w24097_,
		_w24093_,
		_w24098_,
		_w24268_
	);
	LUT3 #(
		.INIT('h80)
	) name18442 (
		_w24095_,
		_w24098_,
		_w24094_,
		_w24269_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18443 (
		_w24096_,
		_w24268_,
		_w24269_,
		_w24267_,
		_w24270_
	);
	LUT4 #(
		.INIT('hfcdc)
	) name18444 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24271_
	);
	LUT3 #(
		.INIT('h0d)
	) name18445 (
		_w24093_,
		_w24100_,
		_w24271_,
		_w24272_
	);
	LUT4 #(
		.INIT('h4000)
	) name18446 (
		_w24096_,
		_w24097_,
		_w24093_,
		_w24098_,
		_w24273_
	);
	LUT2 #(
		.INIT('h2)
	) name18447 (
		_w24094_,
		_w24273_,
		_w24274_
	);
	LUT2 #(
		.INIT('h4)
	) name18448 (
		_w24272_,
		_w24274_,
		_w24275_
	);
	LUT3 #(
		.INIT('h41)
	) name18449 (
		_w24096_,
		_w24097_,
		_w24098_,
		_w24276_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name18450 (
		_w24095_,
		_w24097_,
		_w24093_,
		_w24098_,
		_w24277_
	);
	LUT3 #(
		.INIT('h10)
	) name18451 (
		_w24224_,
		_w24276_,
		_w24277_,
		_w24278_
	);
	LUT4 #(
		.INIT('h03a0)
	) name18452 (
		_w24095_,
		_w24096_,
		_w24097_,
		_w24098_,
		_w24279_
	);
	LUT3 #(
		.INIT('h02)
	) name18453 (
		_w24093_,
		_w24109_,
		_w24279_,
		_w24280_
	);
	LUT2 #(
		.INIT('h1)
	) name18454 (
		_w24094_,
		_w24235_,
		_w24281_
	);
	LUT3 #(
		.INIT('he0)
	) name18455 (
		_w24278_,
		_w24280_,
		_w24281_,
		_w24282_
	);
	LUT4 #(
		.INIT('h6665)
	) name18456 (
		\u1_desIn_r_reg[30]/NET0131 ,
		_w24270_,
		_w24275_,
		_w24282_,
		_w24283_
	);
	LUT3 #(
		.INIT('h09)
	) name18457 (
		_w24123_,
		_w24125_,
		_w24132_,
		_w24284_
	);
	LUT4 #(
		.INIT('h0004)
	) name18458 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24285_
	);
	LUT3 #(
		.INIT('h47)
	) name18459 (
		_w24122_,
		_w24123_,
		_w24132_,
		_w24286_
	);
	LUT4 #(
		.INIT('h0031)
	) name18460 (
		_w24126_,
		_w24285_,
		_w24286_,
		_w24284_,
		_w24287_
	);
	LUT3 #(
		.INIT('h04)
	) name18461 (
		_w24122_,
		_w24124_,
		_w24125_,
		_w24288_
	);
	LUT4 #(
		.INIT('h2010)
	) name18462 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24289_
	);
	LUT4 #(
		.INIT('h0f07)
	) name18463 (
		_w24122_,
		_w24124_,
		_w24130_,
		_w24132_,
		_w24290_
	);
	LUT3 #(
		.INIT('h10)
	) name18464 (
		_w24136_,
		_w24289_,
		_w24290_,
		_w24291_
	);
	LUT2 #(
		.INIT('h8)
	) name18465 (
		_w24287_,
		_w24291_,
		_w24292_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name18466 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24293_
	);
	LUT2 #(
		.INIT('h2)
	) name18467 (
		_w24132_,
		_w24293_,
		_w24294_
	);
	LUT3 #(
		.INIT('h04)
	) name18468 (
		_w24128_,
		_w24130_,
		_w24141_,
		_w24295_
	);
	LUT4 #(
		.INIT('h0400)
	) name18469 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24296_
	);
	LUT2 #(
		.INIT('h6)
	) name18470 (
		_w24124_,
		_w24125_,
		_w24297_
	);
	LUT4 #(
		.INIT('h2022)
	) name18471 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24132_,
		_w24298_
	);
	LUT3 #(
		.INIT('h15)
	) name18472 (
		_w24296_,
		_w24297_,
		_w24298_,
		_w24299_
	);
	LUT3 #(
		.INIT('h40)
	) name18473 (
		_w24294_,
		_w24295_,
		_w24299_,
		_w24300_
	);
	LUT3 #(
		.INIT('ha9)
	) name18474 (
		\u1_desIn_r_reg[28]/NET0131 ,
		_w24292_,
		_w24300_,
		_w24301_
	);
	LUT4 #(
		.INIT('h5515)
	) name18475 (
		_w24240_,
		_w24242_,
		_w24243_,
		_w24241_,
		_w24302_
	);
	LUT3 #(
		.INIT('h40)
	) name18476 (
		_w24242_,
		_w24243_,
		_w24244_,
		_w24303_
	);
	LUT3 #(
		.INIT('h01)
	) name18477 (
		_w24243_,
		_w24241_,
		_w24244_,
		_w24304_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18478 (
		_w24240_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24305_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name18479 (
		_w24258_,
		_w24302_,
		_w24303_,
		_w24305_,
		_w24306_
	);
	LUT4 #(
		.INIT('h0010)
	) name18480 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24307_
	);
	LUT4 #(
		.INIT('h0002)
	) name18481 (
		_w24239_,
		_w24250_,
		_w24251_,
		_w24307_,
		_w24308_
	);
	LUT2 #(
		.INIT('h4)
	) name18482 (
		_w24306_,
		_w24308_,
		_w24309_
	);
	LUT3 #(
		.INIT('h32)
	) name18483 (
		_w24240_,
		_w24242_,
		_w24241_,
		_w24310_
	);
	LUT2 #(
		.INIT('h8)
	) name18484 (
		_w24249_,
		_w24310_,
		_w24311_
	);
	LUT2 #(
		.INIT('h8)
	) name18485 (
		_w24240_,
		_w24242_,
		_w24312_
	);
	LUT3 #(
		.INIT('hb0)
	) name18486 (
		_w24243_,
		_w24241_,
		_w24244_,
		_w24313_
	);
	LUT3 #(
		.INIT('h15)
	) name18487 (
		_w24239_,
		_w24312_,
		_w24313_,
		_w24314_
	);
	LUT4 #(
		.INIT('h5455)
	) name18488 (
		_w24240_,
		_w24242_,
		_w24243_,
		_w24241_,
		_w24315_
	);
	LUT4 #(
		.INIT('h0400)
	) name18489 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24316_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name18490 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24317_
	);
	LUT2 #(
		.INIT('h8)
	) name18491 (
		_w24315_,
		_w24317_,
		_w24318_
	);
	LUT3 #(
		.INIT('h40)
	) name18492 (
		_w24311_,
		_w24314_,
		_w24318_,
		_w24319_
	);
	LUT4 #(
		.INIT('h2000)
	) name18493 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24320_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name18494 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24321_
	);
	LUT3 #(
		.INIT('h09)
	) name18495 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24322_
	);
	LUT3 #(
		.INIT('h02)
	) name18496 (
		_w24242_,
		_w24243_,
		_w24244_,
		_w24323_
	);
	LUT4 #(
		.INIT('h0020)
	) name18497 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24324_
	);
	LUT3 #(
		.INIT('h02)
	) name18498 (
		_w24240_,
		_w24324_,
		_w24322_,
		_w24325_
	);
	LUT3 #(
		.INIT('h40)
	) name18499 (
		_w24311_,
		_w24314_,
		_w24325_,
		_w24326_
	);
	LUT4 #(
		.INIT('h001f)
	) name18500 (
		_w24309_,
		_w24319_,
		_w24321_,
		_w24326_,
		_w24327_
	);
	LUT2 #(
		.INIT('h9)
	) name18501 (
		\u1_desIn_r_reg[36]/NET0131 ,
		_w24327_,
		_w24328_
	);
	LUT4 #(
		.INIT('hc963)
	) name18502 (
		decrypt_pad,
		\u1_desIn_r_reg[41]/NET0131 ,
		\u1_key_r_reg[37]/NET0131 ,
		\u1_key_r_reg[44]/NET0131 ,
		_w24329_
	);
	LUT4 #(
		.INIT('hc693)
	) name18503 (
		decrypt_pad,
		\u1_desIn_r_reg[25]/NET0131 ,
		\u1_key_r_reg[16]/NET0131 ,
		\u1_key_r_reg[9]/NET0131 ,
		_w24330_
	);
	LUT4 #(
		.INIT('hc963)
	) name18504 (
		decrypt_pad,
		\u1_desIn_r_reg[33]/NET0131 ,
		\u1_key_r_reg[36]/NET0131 ,
		\u1_key_r_reg[43]/NET0131 ,
		_w24331_
	);
	LUT4 #(
		.INIT('hc963)
	) name18505 (
		decrypt_pad,
		\u1_desIn_r_reg[7]/NET0131 ,
		\u1_key_r_reg[21]/NET0131 ,
		\u1_key_r_reg[28]/NET0131 ,
		_w24332_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name18506 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24333_
	);
	LUT4 #(
		.INIT('hc693)
	) name18507 (
		decrypt_pad,
		\u1_desIn_r_reg[49]/NET0131 ,
		\u1_key_r_reg[1]/NET0131 ,
		\u1_key_r_reg[49]/NET0131 ,
		_w24334_
	);
	LUT2 #(
		.INIT('h4)
	) name18508 (
		_w24331_,
		_w24329_,
		_w24335_
	);
	LUT4 #(
		.INIT('h2240)
	) name18509 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24336_
	);
	LUT3 #(
		.INIT('h10)
	) name18510 (
		_w24334_,
		_w24336_,
		_w24333_,
		_w24337_
	);
	LUT4 #(
		.INIT('h0010)
	) name18511 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24338_
	);
	LUT4 #(
		.INIT('h4000)
	) name18512 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24339_
	);
	LUT3 #(
		.INIT('h02)
	) name18513 (
		_w24334_,
		_w24339_,
		_w24338_,
		_w24340_
	);
	LUT2 #(
		.INIT('h1)
	) name18514 (
		_w24337_,
		_w24340_,
		_w24341_
	);
	LUT4 #(
		.INIT('hc963)
	) name18515 (
		decrypt_pad,
		\u1_desIn_r_reg[57]/NET0131 ,
		\u1_key_r_reg[0]/NET0131 ,
		\u1_key_r_reg[7]/NET0131 ,
		_w24342_
	);
	LUT4 #(
		.INIT('h6763)
	) name18516 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24343_
	);
	LUT4 #(
		.INIT('h0002)
	) name18517 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24344_
	);
	LUT4 #(
		.INIT('h5504)
	) name18518 (
		_w24342_,
		_w24334_,
		_w24343_,
		_w24344_,
		_w24345_
	);
	LUT4 #(
		.INIT('h0488)
	) name18519 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24346_
	);
	LUT4 #(
		.INIT('h0002)
	) name18520 (
		_w24334_,
		_w24330_,
		_w24331_,
		_w24332_,
		_w24347_
	);
	LUT3 #(
		.INIT('h2f)
	) name18521 (
		_w24334_,
		_w24330_,
		_w24332_,
		_w24348_
	);
	LUT4 #(
		.INIT('h1101)
	) name18522 (
		_w24347_,
		_w24346_,
		_w24335_,
		_w24348_,
		_w24349_
	);
	LUT4 #(
		.INIT('h0010)
	) name18523 (
		_w24342_,
		_w24334_,
		_w24330_,
		_w24331_,
		_w24350_
	);
	LUT4 #(
		.INIT('h0031)
	) name18524 (
		_w24342_,
		_w24345_,
		_w24349_,
		_w24350_,
		_w24351_
	);
	LUT3 #(
		.INIT('h65)
	) name18525 (
		\u1_desIn_r_reg[52]/P0001 ,
		_w24341_,
		_w24351_,
		_w24352_
	);
	LUT4 #(
		.INIT('hc963)
	) name18526 (
		decrypt_pad,
		\u1_desIn_r_reg[27]/NET0131 ,
		\u1_key_r_reg[16]/NET0131 ,
		\u1_key_r_reg[23]/NET0131 ,
		_w24353_
	);
	LUT4 #(
		.INIT('hc963)
	) name18527 (
		decrypt_pad,
		\u1_desIn_r_reg[19]/NET0131 ,
		\u1_key_r_reg[1]/NET0131 ,
		\u1_key_r_reg[8]/NET0131 ,
		_w24354_
	);
	LUT4 #(
		.INIT('hc693)
	) name18528 (
		decrypt_pad,
		\u1_desIn_r_reg[3]/NET0131 ,
		\u1_key_r_reg[31]/NET0131 ,
		\u1_key_r_reg[51]/NET0131 ,
		_w24355_
	);
	LUT4 #(
		.INIT('hc963)
	) name18529 (
		decrypt_pad,
		\u1_desIn_r_reg[61]/NET0131 ,
		\u1_key_r_reg[29]/NET0131 ,
		\u1_key_r_reg[36]/NET0131 ,
		_w24356_
	);
	LUT4 #(
		.INIT('hc963)
	) name18530 (
		decrypt_pad,
		\u1_desIn_r_reg[35]/NET0131 ,
		\u1_key_r_reg[45]/NET0131 ,
		\u1_key_r_reg[52]/NET0131 ,
		_w24357_
	);
	LUT4 #(
		.INIT('hc963)
	) name18531 (
		decrypt_pad,
		\u1_desIn_r_reg[11]/NET0131 ,
		\u1_key_r_reg[14]/NET0131 ,
		\u1_key_r_reg[21]/NET0131 ,
		_w24358_
	);
	LUT4 #(
		.INIT('hc25f)
	) name18532 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24359_
	);
	LUT2 #(
		.INIT('h2)
	) name18533 (
		_w24354_,
		_w24359_,
		_w24360_
	);
	LUT2 #(
		.INIT('h1)
	) name18534 (
		_w24358_,
		_w24354_,
		_w24361_
	);
	LUT3 #(
		.INIT('h20)
	) name18535 (
		_w24355_,
		_w24356_,
		_w24357_,
		_w24362_
	);
	LUT3 #(
		.INIT('hde)
	) name18536 (
		_w24355_,
		_w24356_,
		_w24357_,
		_w24363_
	);
	LUT2 #(
		.INIT('h2)
	) name18537 (
		_w24361_,
		_w24363_,
		_w24364_
	);
	LUT3 #(
		.INIT('hc4)
	) name18538 (
		_w24355_,
		_w24358_,
		_w24354_,
		_w24365_
	);
	LUT4 #(
		.INIT('hd000)
	) name18539 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24366_
	);
	LUT4 #(
		.INIT('h0020)
	) name18540 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24367_
	);
	LUT4 #(
		.INIT('h0040)
	) name18541 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24368_
	);
	LUT4 #(
		.INIT('hff9f)
	) name18542 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24369_
	);
	LUT3 #(
		.INIT('hb0)
	) name18543 (
		_w24365_,
		_w24366_,
		_w24369_,
		_w24370_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name18544 (
		_w24353_,
		_w24364_,
		_w24360_,
		_w24370_,
		_w24371_
	);
	LUT4 #(
		.INIT('h0010)
	) name18545 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24372_
	);
	LUT4 #(
		.INIT('hda67)
	) name18546 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24373_
	);
	LUT3 #(
		.INIT('h02)
	) name18547 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24374_
	);
	LUT4 #(
		.INIT('h3df8)
	) name18548 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24375_
	);
	LUT4 #(
		.INIT('h4000)
	) name18549 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24376_
	);
	LUT4 #(
		.INIT('hbffd)
	) name18550 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24377_
	);
	LUT4 #(
		.INIT('he400)
	) name18551 (
		_w24354_,
		_w24373_,
		_w24375_,
		_w24377_,
		_w24378_
	);
	LUT4 #(
		.INIT('hffdb)
	) name18552 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24379_
	);
	LUT4 #(
		.INIT('h0400)
	) name18553 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24380_
	);
	LUT4 #(
		.INIT('hfbf7)
	) name18554 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24381_
	);
	LUT3 #(
		.INIT('hd8)
	) name18555 (
		_w24354_,
		_w24379_,
		_w24381_,
		_w24382_
	);
	LUT3 #(
		.INIT('he0)
	) name18556 (
		_w24353_,
		_w24378_,
		_w24382_,
		_w24383_
	);
	LUT3 #(
		.INIT('h65)
	) name18557 (
		\u1_desIn_r_reg[44]/NET0131 ,
		_w24371_,
		_w24383_,
		_w24384_
	);
	LUT4 #(
		.INIT('h0400)
	) name18558 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24385_
	);
	LUT4 #(
		.INIT('haaa8)
	) name18559 (
		_w24186_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24386_
	);
	LUT3 #(
		.INIT('h40)
	) name18560 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24387_
	);
	LUT4 #(
		.INIT('h5551)
	) name18561 (
		_w24186_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24388_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name18562 (
		_w24385_,
		_w24386_,
		_w24387_,
		_w24388_,
		_w24389_
	);
	LUT4 #(
		.INIT('h7fd7)
	) name18563 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24390_
	);
	LUT3 #(
		.INIT('h45)
	) name18564 (
		_w24195_,
		_w24389_,
		_w24390_,
		_w24391_
	);
	LUT4 #(
		.INIT('hdf5d)
	) name18565 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24392_
	);
	LUT4 #(
		.INIT('h0800)
	) name18566 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24393_
	);
	LUT4 #(
		.INIT('he6ff)
	) name18567 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24394_
	);
	LUT4 #(
		.INIT('h04cc)
	) name18568 (
		_w24186_,
		_w24195_,
		_w24392_,
		_w24394_,
		_w24395_
	);
	LUT4 #(
		.INIT('h6fff)
	) name18569 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24396_
	);
	LUT4 #(
		.INIT('h6dff)
	) name18570 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24397_
	);
	LUT2 #(
		.INIT('h2)
	) name18571 (
		_w24186_,
		_w24397_,
		_w24398_
	);
	LUT2 #(
		.INIT('h4)
	) name18572 (
		_w24186_,
		_w24393_,
		_w24399_
	);
	LUT4 #(
		.INIT('hafab)
	) name18573 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24400_
	);
	LUT2 #(
		.INIT('h8)
	) name18574 (
		_w24186_,
		_w24195_,
		_w24401_
	);
	LUT4 #(
		.INIT('h7077)
	) name18575 (
		_w24197_,
		_w24187_,
		_w24400_,
		_w24401_,
		_w24402_
	);
	LUT4 #(
		.INIT('h0100)
	) name18576 (
		_w24398_,
		_w24399_,
		_w24395_,
		_w24402_,
		_w24403_
	);
	LUT3 #(
		.INIT('h65)
	) name18577 (
		\u1_desIn_r_reg[6]/NET0131 ,
		_w24391_,
		_w24403_,
		_w24404_
	);
	LUT4 #(
		.INIT('hab5b)
	) name18578 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24405_
	);
	LUT2 #(
		.INIT('h1)
	) name18579 (
		_w24334_,
		_w24405_,
		_w24406_
	);
	LUT4 #(
		.INIT('h0080)
	) name18580 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24407_
	);
	LUT4 #(
		.INIT('hbb7e)
	) name18581 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24408_
	);
	LUT3 #(
		.INIT('h2a)
	) name18582 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24409_
	);
	LUT3 #(
		.INIT('ha8)
	) name18583 (
		_w24334_,
		_w24331_,
		_w24329_,
		_w24410_
	);
	LUT3 #(
		.INIT('h10)
	) name18584 (
		_w24331_,
		_w24332_,
		_w24329_,
		_w24411_
	);
	LUT4 #(
		.INIT('h0200)
	) name18585 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24412_
	);
	LUT4 #(
		.INIT('h0700)
	) name18586 (
		_w24409_,
		_w24410_,
		_w24412_,
		_w24408_,
		_w24413_
	);
	LUT3 #(
		.INIT('h45)
	) name18587 (
		_w24342_,
		_w24406_,
		_w24413_,
		_w24414_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name18588 (
		_w24334_,
		_w24330_,
		_w24331_,
		_w24332_,
		_w24415_
	);
	LUT4 #(
		.INIT('h77cf)
	) name18589 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24416_
	);
	LUT4 #(
		.INIT('h2000)
	) name18590 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24417_
	);
	LUT4 #(
		.INIT('h5551)
	) name18591 (
		_w24334_,
		_w24330_,
		_w24332_,
		_w24329_,
		_w24418_
	);
	LUT4 #(
		.INIT('h7077)
	) name18592 (
		_w24415_,
		_w24416_,
		_w24417_,
		_w24418_,
		_w24419_
	);
	LUT4 #(
		.INIT('hf6ef)
	) name18593 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24420_
	);
	LUT4 #(
		.INIT('h0002)
	) name18594 (
		_w24334_,
		_w24330_,
		_w24331_,
		_w24329_,
		_w24421_
	);
	LUT3 #(
		.INIT('h0b)
	) name18595 (
		_w24334_,
		_w24407_,
		_w24421_,
		_w24422_
	);
	LUT4 #(
		.INIT('h7500)
	) name18596 (
		_w24342_,
		_w24419_,
		_w24420_,
		_w24422_,
		_w24423_
	);
	LUT3 #(
		.INIT('h65)
	) name18597 (
		\u1_desIn_r_reg[34]/NET0131 ,
		_w24414_,
		_w24423_,
		_w24424_
	);
	LUT4 #(
		.INIT('hfcd3)
	) name18598 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24425_
	);
	LUT4 #(
		.INIT('heffb)
	) name18599 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24426_
	);
	LUT4 #(
		.INIT('h0233)
	) name18600 (
		_w24062_,
		_w24069_,
		_w24425_,
		_w24426_,
		_w24427_
	);
	LUT4 #(
		.INIT('h02a0)
	) name18601 (
		_w24069_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24428_
	);
	LUT3 #(
		.INIT('h54)
	) name18602 (
		_w24081_,
		_w24087_,
		_w24428_,
		_w24429_
	);
	LUT3 #(
		.INIT('h8c)
	) name18603 (
		_w24065_,
		_w24069_,
		_w24063_,
		_w24430_
	);
	LUT2 #(
		.INIT('h8)
	) name18604 (
		_w24082_,
		_w24430_,
		_w24431_
	);
	LUT4 #(
		.INIT('h002a)
	) name18605 (
		_w24062_,
		_w24073_,
		_w24085_,
		_w24154_,
		_w24432_
	);
	LUT4 #(
		.INIT('h1554)
	) name18606 (
		_w24062_,
		_w24065_,
		_w24066_,
		_w24064_,
		_w24433_
	);
	LUT3 #(
		.INIT('h47)
	) name18607 (
		_w24065_,
		_w24066_,
		_w24064_,
		_w24434_
	);
	LUT3 #(
		.INIT('h07)
	) name18608 (
		_w24065_,
		_w24066_,
		_w24064_,
		_w24435_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name18609 (
		_w24069_,
		_w24063_,
		_w24434_,
		_w24435_,
		_w24436_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name18610 (
		_w24431_,
		_w24432_,
		_w24433_,
		_w24436_,
		_w24437_
	);
	LUT4 #(
		.INIT('haaa9)
	) name18611 (
		\u1_desIn_r_reg[50]/NET0131 ,
		_w24429_,
		_w24437_,
		_w24427_,
		_w24438_
	);
	LUT4 #(
		.INIT('h00bf)
	) name18612 (
		_w24355_,
		_w24356_,
		_w24357_,
		_w24354_,
		_w24439_
	);
	LUT4 #(
		.INIT('h7f00)
	) name18613 (
		_w24355_,
		_w24356_,
		_w24357_,
		_w24354_,
		_w24440_
	);
	LUT4 #(
		.INIT('hfae2)
	) name18614 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24441_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name18615 (
		_w24374_,
		_w24439_,
		_w24440_,
		_w24441_,
		_w24442_
	);
	LUT4 #(
		.INIT('h0080)
	) name18616 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24443_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name18617 (
		_w24353_,
		_w24355_,
		_w24358_,
		_w24357_,
		_w24444_
	);
	LUT2 #(
		.INIT('h4)
	) name18618 (
		_w24443_,
		_w24444_,
		_w24445_
	);
	LUT4 #(
		.INIT('hf5ee)
	) name18619 (
		_w24355_,
		_w24356_,
		_w24357_,
		_w24354_,
		_w24446_
	);
	LUT2 #(
		.INIT('h1)
	) name18620 (
		_w24358_,
		_w24446_,
		_w24447_
	);
	LUT2 #(
		.INIT('h4)
	) name18621 (
		_w24357_,
		_w24354_,
		_w24448_
	);
	LUT3 #(
		.INIT('h08)
	) name18622 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24449_
	);
	LUT4 #(
		.INIT('h0004)
	) name18623 (
		_w24355_,
		_w24356_,
		_w24357_,
		_w24354_,
		_w24450_
	);
	LUT4 #(
		.INIT('h1011)
	) name18624 (
		_w24353_,
		_w24450_,
		_w24448_,
		_w24449_,
		_w24451_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name18625 (
		_w24442_,
		_w24445_,
		_w24447_,
		_w24451_,
		_w24452_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name18626 (
		_w24355_,
		_w24358_,
		_w24357_,
		_w24354_,
		_w24453_
	);
	LUT4 #(
		.INIT('hff7b)
	) name18627 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24454_
	);
	LUT4 #(
		.INIT('hfe7b)
	) name18628 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24455_
	);
	LUT4 #(
		.INIT('hf531)
	) name18629 (
		_w24356_,
		_w24354_,
		_w24453_,
		_w24455_,
		_w24456_
	);
	LUT3 #(
		.INIT('h65)
	) name18630 (
		\u1_desIn_r_reg[0]/NET0131 ,
		_w24452_,
		_w24456_,
		_w24457_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name18631 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24458_
	);
	LUT2 #(
		.INIT('h2)
	) name18632 (
		_w24240_,
		_w24458_,
		_w24459_
	);
	LUT4 #(
		.INIT('hbfae)
	) name18633 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24460_
	);
	LUT2 #(
		.INIT('h1)
	) name18634 (
		_w24240_,
		_w24460_,
		_w24461_
	);
	LUT4 #(
		.INIT('h7737)
	) name18635 (
		_w24240_,
		_w24242_,
		_w24243_,
		_w24241_,
		_w24462_
	);
	LUT3 #(
		.INIT('h32)
	) name18636 (
		_w24244_,
		_w24316_,
		_w24462_,
		_w24463_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name18637 (
		_w24239_,
		_w24461_,
		_w24459_,
		_w24463_,
		_w24464_
	);
	LUT4 #(
		.INIT('hdaff)
	) name18638 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24465_
	);
	LUT2 #(
		.INIT('h1)
	) name18639 (
		_w24240_,
		_w24465_,
		_w24466_
	);
	LUT4 #(
		.INIT('h1145)
	) name18640 (
		_w24240_,
		_w24242_,
		_w24243_,
		_w24241_,
		_w24467_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name18641 (
		_w24240_,
		_w24323_,
		_w24460_,
		_w24467_,
		_w24468_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name18642 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24469_
	);
	LUT4 #(
		.INIT('h2322)
	) name18643 (
		_w24239_,
		_w24466_,
		_w24468_,
		_w24469_,
		_w24470_
	);
	LUT3 #(
		.INIT('h65)
	) name18644 (
		\u1_desIn_r_reg[24]/NET0131 ,
		_w24464_,
		_w24470_,
		_w24471_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name18645 (
		_w24182_,
		_w24186_,
		_w24183_,
		_w24189_,
		_w24472_
	);
	LUT3 #(
		.INIT('h31)
	) name18646 (
		_w24187_,
		_w24206_,
		_w24472_,
		_w24473_
	);
	LUT4 #(
		.INIT('h0802)
	) name18647 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24474_
	);
	LUT4 #(
		.INIT('h3fef)
	) name18648 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24475_
	);
	LUT3 #(
		.INIT('h32)
	) name18649 (
		_w24186_,
		_w24474_,
		_w24475_,
		_w24476_
	);
	LUT3 #(
		.INIT('h2a)
	) name18650 (
		_w24195_,
		_w24473_,
		_w24476_,
		_w24477_
	);
	LUT4 #(
		.INIT('heafa)
	) name18651 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24478_
	);
	LUT4 #(
		.INIT('h0086)
	) name18652 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24479_
	);
	LUT4 #(
		.INIT('h5501)
	) name18653 (
		_w24186_,
		_w24195_,
		_w24478_,
		_w24479_,
		_w24480_
	);
	LUT2 #(
		.INIT('h4)
	) name18654 (
		_w24193_,
		_w24207_,
		_w24481_
	);
	LUT3 #(
		.INIT('h01)
	) name18655 (
		_w24198_,
		_w24191_,
		_w24202_,
		_w24482_
	);
	LUT3 #(
		.INIT('h08)
	) name18656 (
		_w24186_,
		_w24189_,
		_w24187_,
		_w24483_
	);
	LUT2 #(
		.INIT('h4)
	) name18657 (
		_w24185_,
		_w24483_,
		_w24484_
	);
	LUT4 #(
		.INIT('h00ba)
	) name18658 (
		_w24195_,
		_w24481_,
		_w24482_,
		_w24484_,
		_w24485_
	);
	LUT4 #(
		.INIT('h5655)
	) name18659 (
		\u1_desIn_r_reg[8]/NET0131 ,
		_w24480_,
		_w24477_,
		_w24485_,
		_w24486_
	);
	LUT4 #(
		.INIT('h0144)
	) name18660 (
		_w24334_,
		_w24330_,
		_w24332_,
		_w24329_,
		_w24487_
	);
	LUT4 #(
		.INIT('h2fa3)
	) name18661 (
		_w24334_,
		_w24330_,
		_w24332_,
		_w24329_,
		_w24488_
	);
	LUT4 #(
		.INIT('h5054)
	) name18662 (
		_w24342_,
		_w24331_,
		_w24487_,
		_w24488_,
		_w24489_
	);
	LUT4 #(
		.INIT('hedef)
	) name18663 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24490_
	);
	LUT4 #(
		.INIT('hebde)
	) name18664 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24491_
	);
	LUT4 #(
		.INIT('h04cc)
	) name18665 (
		_w24342_,
		_w24334_,
		_w24490_,
		_w24491_,
		_w24492_
	);
	LUT4 #(
		.INIT('h0008)
	) name18666 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24493_
	);
	LUT2 #(
		.INIT('h4)
	) name18667 (
		_w24334_,
		_w24493_,
		_w24494_
	);
	LUT4 #(
		.INIT('hf351)
	) name18668 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24495_
	);
	LUT3 #(
		.INIT('h02)
	) name18669 (
		_w24334_,
		_w24493_,
		_w24495_,
		_w24496_
	);
	LUT4 #(
		.INIT('h0401)
	) name18670 (
		_w24334_,
		_w24330_,
		_w24331_,
		_w24329_,
		_w24497_
	);
	LUT2 #(
		.INIT('h1)
	) name18671 (
		_w24339_,
		_w24497_,
		_w24498_
	);
	LUT4 #(
		.INIT('h1311)
	) name18672 (
		_w24342_,
		_w24494_,
		_w24496_,
		_w24498_,
		_w24499_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name18673 (
		\u1_desIn_r_reg[38]/NET0131 ,
		_w24492_,
		_w24489_,
		_w24499_,
		_w24500_
	);
	LUT4 #(
		.INIT('hfd77)
	) name18674 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24501_
	);
	LUT4 #(
		.INIT('he4ee)
	) name18675 (
		_w24354_,
		_w24368_,
		_w24380_,
		_w24501_,
		_w24502_
	);
	LUT4 #(
		.INIT('h0001)
	) name18676 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24503_
	);
	LUT4 #(
		.INIT('haffe)
	) name18677 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24504_
	);
	LUT4 #(
		.INIT('haa8a)
	) name18678 (
		_w24353_,
		_w24358_,
		_w24356_,
		_w24354_,
		_w24505_
	);
	LUT4 #(
		.INIT('hc400)
	) name18679 (
		_w24354_,
		_w24381_,
		_w24504_,
		_w24505_,
		_w24506_
	);
	LUT4 #(
		.INIT('h0b00)
	) name18680 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24507_
	);
	LUT4 #(
		.INIT('haf23)
	) name18681 (
		_w24372_,
		_w24439_,
		_w24440_,
		_w24507_,
		_w24508_
	);
	LUT4 #(
		.INIT('h5551)
	) name18682 (
		_w24353_,
		_w24355_,
		_w24358_,
		_w24356_,
		_w24509_
	);
	LUT2 #(
		.INIT('h8)
	) name18683 (
		_w24454_,
		_w24509_,
		_w24510_
	);
	LUT4 #(
		.INIT('h4544)
	) name18684 (
		_w24502_,
		_w24506_,
		_w24508_,
		_w24510_,
		_w24511_
	);
	LUT2 #(
		.INIT('h9)
	) name18685 (
		\u1_desIn_r_reg[62]/NET0131 ,
		_w24511_,
		_w24512_
	);
	LUT4 #(
		.INIT('h0020)
	) name18686 (
		_w24186_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24513_
	);
	LUT3 #(
		.INIT('h40)
	) name18687 (
		_w24182_,
		_w24186_,
		_w24183_,
		_w24514_
	);
	LUT4 #(
		.INIT('h0045)
	) name18688 (
		_w24197_,
		_w24216_,
		_w24514_,
		_w24513_,
		_w24515_
	);
	LUT4 #(
		.INIT('hff45)
	) name18689 (
		_w24182_,
		_w24186_,
		_w24189_,
		_w24187_,
		_w24516_
	);
	LUT3 #(
		.INIT('hc4)
	) name18690 (
		_w24183_,
		_w24210_,
		_w24516_,
		_w24517_
	);
	LUT3 #(
		.INIT('h15)
	) name18691 (
		_w24195_,
		_w24515_,
		_w24517_,
		_w24518_
	);
	LUT4 #(
		.INIT('hfdbd)
	) name18692 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24519_
	);
	LUT4 #(
		.INIT('hf3db)
	) name18693 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24520_
	);
	LUT4 #(
		.INIT('hc840)
	) name18694 (
		_w24186_,
		_w24396_,
		_w24520_,
		_w24519_,
		_w24521_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name18695 (
		_w24182_,
		_w24183_,
		_w24189_,
		_w24187_,
		_w24522_
	);
	LUT2 #(
		.INIT('h1)
	) name18696 (
		_w24186_,
		_w24522_,
		_w24523_
	);
	LUT3 #(
		.INIT('h13)
	) name18697 (
		_w24190_,
		_w24208_,
		_w24218_,
		_w24524_
	);
	LUT4 #(
		.INIT('h0d00)
	) name18698 (
		_w24195_,
		_w24521_,
		_w24523_,
		_w24524_,
		_w24525_
	);
	LUT3 #(
		.INIT('h65)
	) name18699 (
		\u1_desIn_r_reg[12]/NET0131 ,
		_w24518_,
		_w24525_,
		_w24526_
	);
	LUT4 #(
		.INIT('hb7a6)
	) name18700 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24527_
	);
	LUT2 #(
		.INIT('h1)
	) name18701 (
		_w24334_,
		_w24527_,
		_w24528_
	);
	LUT4 #(
		.INIT('h5551)
	) name18702 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24529_
	);
	LUT4 #(
		.INIT('ha222)
	) name18703 (
		_w24334_,
		_w24330_,
		_w24331_,
		_w24332_,
		_w24530_
	);
	LUT4 #(
		.INIT('hbdcf)
	) name18704 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24531_
	);
	LUT3 #(
		.INIT('hb0)
	) name18705 (
		_w24529_,
		_w24530_,
		_w24531_,
		_w24532_
	);
	LUT3 #(
		.INIT('h8a)
	) name18706 (
		_w24342_,
		_w24528_,
		_w24532_,
		_w24533_
	);
	LUT4 #(
		.INIT('h5551)
	) name18707 (
		_w24342_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24534_
	);
	LUT4 #(
		.INIT('h0bcf)
	) name18708 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24535_
	);
	LUT4 #(
		.INIT('ha888)
	) name18709 (
		_w24334_,
		_w24411_,
		_w24534_,
		_w24535_,
		_w24536_
	);
	LUT4 #(
		.INIT('h5bfb)
	) name18710 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24537_
	);
	LUT4 #(
		.INIT('h1000)
	) name18711 (
		_w24330_,
		_w24331_,
		_w24332_,
		_w24329_,
		_w24538_
	);
	LUT4 #(
		.INIT('h5501)
	) name18712 (
		_w24342_,
		_w24334_,
		_w24537_,
		_w24538_,
		_w24539_
	);
	LUT2 #(
		.INIT('h6)
	) name18713 (
		_w24331_,
		_w24332_,
		_w24540_
	);
	LUT2 #(
		.INIT('h8)
	) name18714 (
		_w24487_,
		_w24540_,
		_w24541_
	);
	LUT3 #(
		.INIT('h01)
	) name18715 (
		_w24539_,
		_w24536_,
		_w24541_,
		_w24542_
	);
	LUT3 #(
		.INIT('h65)
	) name18716 (
		\u1_desIn_r_reg[16]/NET0131 ,
		_w24533_,
		_w24542_,
		_w24543_
	);
	LUT3 #(
		.INIT('h41)
	) name18717 (
		_w24122_,
		_w24124_,
		_w24125_,
		_w24544_
	);
	LUT3 #(
		.INIT('h40)
	) name18718 (
		_w24123_,
		_w24124_,
		_w24125_,
		_w24545_
	);
	LUT4 #(
		.INIT('hdee3)
	) name18719 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24546_
	);
	LUT4 #(
		.INIT('h0080)
	) name18720 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24547_
	);
	LUT4 #(
		.INIT('hbb5c)
	) name18721 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24548_
	);
	LUT4 #(
		.INIT('h3210)
	) name18722 (
		_w24132_,
		_w24547_,
		_w24546_,
		_w24548_,
		_w24549_
	);
	LUT2 #(
		.INIT('h2)
	) name18723 (
		_w24130_,
		_w24549_,
		_w24550_
	);
	LUT4 #(
		.INIT('h7db7)
	) name18724 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24551_
	);
	LUT4 #(
		.INIT('h4547)
	) name18725 (
		_w24132_,
		_w24288_,
		_w24284_,
		_w24545_,
		_w24552_
	);
	LUT4 #(
		.INIT('h00a2)
	) name18726 (
		_w24123_,
		_w24124_,
		_w24125_,
		_w24132_,
		_w24553_
	);
	LUT4 #(
		.INIT('h0777)
	) name18727 (
		_w24127_,
		_w24132_,
		_w24137_,
		_w24553_,
		_w24554_
	);
	LUT4 #(
		.INIT('hea00)
	) name18728 (
		_w24130_,
		_w24551_,
		_w24552_,
		_w24554_,
		_w24555_
	);
	LUT3 #(
		.INIT('h65)
	) name18729 (
		\u1_desIn_r_reg[56]/NET0131 ,
		_w24550_,
		_w24555_,
		_w24556_
	);
	LUT4 #(
		.INIT('hcff5)
	) name18730 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24557_
	);
	LUT4 #(
		.INIT('hdfbf)
	) name18731 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24558_
	);
	LUT4 #(
		.INIT('hb100)
	) name18732 (
		_w24354_,
		_w24362_,
		_w24557_,
		_w24558_,
		_w24559_
	);
	LUT2 #(
		.INIT('h2)
	) name18733 (
		_w24353_,
		_w24559_,
		_w24560_
	);
	LUT4 #(
		.INIT('hb85b)
	) name18734 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24561_
	);
	LUT2 #(
		.INIT('h1)
	) name18735 (
		_w24353_,
		_w24561_,
		_w24562_
	);
	LUT3 #(
		.INIT('h02)
	) name18736 (
		_w24354_,
		_w24372_,
		_w24380_,
		_w24563_
	);
	LUT4 #(
		.INIT('h23f0)
	) name18737 (
		_w24355_,
		_w24358_,
		_w24356_,
		_w24357_,
		_w24564_
	);
	LUT3 #(
		.INIT('h0d)
	) name18738 (
		_w24353_,
		_w24376_,
		_w24564_,
		_w24565_
	);
	LUT3 #(
		.INIT('h01)
	) name18739 (
		_w24354_,
		_w24367_,
		_w24503_,
		_w24566_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name18740 (
		_w24562_,
		_w24563_,
		_w24565_,
		_w24566_,
		_w24567_
	);
	LUT3 #(
		.INIT('h56)
	) name18741 (
		\u1_desIn_r_reg[22]/NET0131 ,
		_w24560_,
		_w24567_,
		_w24568_
	);
	LUT4 #(
		.INIT('hc963)
	) name18742 (
		decrypt_pad,
		\u1_desIn_r_reg[5]/NET0131 ,
		\u1_key_r_reg[18]/NET0131 ,
		\u1_key_r_reg[25]/NET0131 ,
		_w24569_
	);
	LUT4 #(
		.INIT('hc963)
	) name18743 (
		decrypt_pad,
		\u1_desIn_r_reg[13]/NET0131 ,
		\u1_key_r_reg[26]/NET0131 ,
		\u1_key_r_reg[33]/NET0131 ,
		_w24570_
	);
	LUT2 #(
		.INIT('h8)
	) name18744 (
		_w24569_,
		_w24570_,
		_w24571_
	);
	LUT4 #(
		.INIT('hc963)
	) name18745 (
		decrypt_pad,
		\u1_desIn_r_reg[37]/NET0131 ,
		\u1_key_r_reg[55]/NET0131 ,
		\u1_key_r_reg[5]/NET0131 ,
		_w24572_
	);
	LUT4 #(
		.INIT('hc963)
	) name18746 (
		decrypt_pad,
		\u1_desIn_r_reg[63]/NET0131 ,
		\u1_key_r_reg[46]/NET0131 ,
		\u1_key_r_reg[53]/NET0131 ,
		_w24573_
	);
	LUT2 #(
		.INIT('h8)
	) name18747 (
		_w24572_,
		_w24573_,
		_w24574_
	);
	LUT4 #(
		.INIT('he00e)
	) name18748 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24575_
	);
	LUT2 #(
		.INIT('h2)
	) name18749 (
		_w24572_,
		_w24573_,
		_w24576_
	);
	LUT4 #(
		.INIT('hc963)
	) name18750 (
		decrypt_pad,
		\u1_desIn_r_reg[21]/NET0131 ,
		\u1_key_r_reg[27]/NET0131 ,
		\u1_key_r_reg[34]/NET0131 ,
		_w24577_
	);
	LUT4 #(
		.INIT('hefeb)
	) name18751 (
		_w24570_,
		_w24572_,
		_w24573_,
		_w24577_,
		_w24578_
	);
	LUT2 #(
		.INIT('h1)
	) name18752 (
		_w24569_,
		_w24578_,
		_w24579_
	);
	LUT4 #(
		.INIT('h3031)
	) name18753 (
		_w24569_,
		_w24571_,
		_w24575_,
		_w24578_,
		_w24580_
	);
	LUT3 #(
		.INIT('h08)
	) name18754 (
		_w24569_,
		_w24570_,
		_w24577_,
		_w24581_
	);
	LUT2 #(
		.INIT('h4)
	) name18755 (
		_w24570_,
		_w24577_,
		_w24582_
	);
	LUT4 #(
		.INIT('h0200)
	) name18756 (
		_w24569_,
		_w24570_,
		_w24573_,
		_w24577_,
		_w24583_
	);
	LUT4 #(
		.INIT('h0800)
	) name18757 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24584_
	);
	LUT4 #(
		.INIT('h0013)
	) name18758 (
		_w24576_,
		_w24583_,
		_w24581_,
		_w24584_,
		_w24585_
	);
	LUT4 #(
		.INIT('hc963)
	) name18759 (
		decrypt_pad,
		\u1_desIn_r_reg[29]/NET0131 ,
		\u1_key_r_reg[10]/NET0131 ,
		\u1_key_r_reg[17]/NET0131 ,
		_w24586_
	);
	LUT3 #(
		.INIT('h0b)
	) name18760 (
		_w24580_,
		_w24585_,
		_w24586_,
		_w24587_
	);
	LUT4 #(
		.INIT('hf53f)
	) name18761 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24588_
	);
	LUT4 #(
		.INIT('ha52f)
	) name18762 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24589_
	);
	LUT2 #(
		.INIT('h2)
	) name18763 (
		_w24577_,
		_w24589_,
		_w24590_
	);
	LUT4 #(
		.INIT('h0008)
	) name18764 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24591_
	);
	LUT3 #(
		.INIT('hd8)
	) name18765 (
		_w24569_,
		_w24572_,
		_w24573_,
		_w24592_
	);
	LUT4 #(
		.INIT('h00d8)
	) name18766 (
		_w24569_,
		_w24572_,
		_w24573_,
		_w24577_,
		_w24593_
	);
	LUT4 #(
		.INIT('h50dd)
	) name18767 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24594_
	);
	LUT3 #(
		.INIT('h51)
	) name18768 (
		_w24591_,
		_w24593_,
		_w24594_,
		_w24595_
	);
	LUT4 #(
		.INIT('h0001)
	) name18769 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24596_
	);
	LUT2 #(
		.INIT('h4)
	) name18770 (
		_w24569_,
		_w24570_,
		_w24597_
	);
	LUT4 #(
		.INIT('hbfbe)
	) name18771 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24598_
	);
	LUT2 #(
		.INIT('h2)
	) name18772 (
		_w24577_,
		_w24598_,
		_w24599_
	);
	LUT4 #(
		.INIT('h0075)
	) name18773 (
		_w24586_,
		_w24590_,
		_w24595_,
		_w24599_,
		_w24600_
	);
	LUT3 #(
		.INIT('h65)
	) name18774 (
		\u1_desIn_r_reg[46]/NET0131 ,
		_w24587_,
		_w24600_,
		_w24601_
	);
	LUT4 #(
		.INIT('h5004)
	) name18775 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24602_
	);
	LUT2 #(
		.INIT('h2)
	) name18776 (
		_w24132_,
		_w24602_,
		_w24603_
	);
	LUT3 #(
		.INIT('h09)
	) name18777 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24604_
	);
	LUT3 #(
		.INIT('h28)
	) name18778 (
		_w24123_,
		_w24124_,
		_w24125_,
		_w24605_
	);
	LUT4 #(
		.INIT('h00f7)
	) name18779 (
		_w24122_,
		_w24124_,
		_w24125_,
		_w24132_,
		_w24606_
	);
	LUT3 #(
		.INIT('h10)
	) name18780 (
		_w24605_,
		_w24604_,
		_w24606_,
		_w24607_
	);
	LUT4 #(
		.INIT('h2880)
	) name18781 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24608_
	);
	LUT2 #(
		.INIT('h2)
	) name18782 (
		_w24130_,
		_w24608_,
		_w24609_
	);
	LUT4 #(
		.INIT('h0880)
	) name18783 (
		_w24122_,
		_w24123_,
		_w24124_,
		_w24125_,
		_w24610_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18784 (
		_w24123_,
		_w24124_,
		_w24125_,
		_w24132_,
		_w24611_
	);
	LUT4 #(
		.INIT('h5455)
	) name18785 (
		_w24130_,
		_w24544_,
		_w24610_,
		_w24611_,
		_w24612_
	);
	LUT4 #(
		.INIT('h001f)
	) name18786 (
		_w24603_,
		_w24607_,
		_w24609_,
		_w24612_,
		_w24613_
	);
	LUT2 #(
		.INIT('h4)
	) name18787 (
		_w24132_,
		_w24608_,
		_w24614_
	);
	LUT2 #(
		.INIT('h2)
	) name18788 (
		_w24130_,
		_w24132_,
		_w24615_
	);
	LUT4 #(
		.INIT('h00dc)
	) name18789 (
		_w24132_,
		_w24136_,
		_w24602_,
		_w24615_,
		_w24616_
	);
	LUT2 #(
		.INIT('h1)
	) name18790 (
		_w24614_,
		_w24616_,
		_w24617_
	);
	LUT3 #(
		.INIT('h65)
	) name18791 (
		\u1_desIn_r_reg[54]/NET0131 ,
		_w24613_,
		_w24617_,
		_w24618_
	);
	LUT4 #(
		.INIT('hdc33)
	) name18792 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24619_
	);
	LUT2 #(
		.INIT('h2)
	) name18793 (
		_w24069_,
		_w24619_,
		_w24620_
	);
	LUT4 #(
		.INIT('h0082)
	) name18794 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24621_
	);
	LUT3 #(
		.INIT('h25)
	) name18795 (
		_w24066_,
		_w24063_,
		_w24064_,
		_w24622_
	);
	LUT4 #(
		.INIT('h0411)
	) name18796 (
		_w24069_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24623_
	);
	LUT4 #(
		.INIT('h4000)
	) name18797 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24624_
	);
	LUT3 #(
		.INIT('h01)
	) name18798 (
		_w24623_,
		_w24621_,
		_w24624_,
		_w24625_
	);
	LUT3 #(
		.INIT('h45)
	) name18799 (
		_w24062_,
		_w24620_,
		_w24625_,
		_w24626_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name18800 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24627_
	);
	LUT2 #(
		.INIT('h1)
	) name18801 (
		_w24069_,
		_w24627_,
		_w24628_
	);
	LUT4 #(
		.INIT('h8228)
	) name18802 (
		_w24065_,
		_w24066_,
		_w24063_,
		_w24064_,
		_w24629_
	);
	LUT4 #(
		.INIT('h0013)
	) name18803 (
		_w24070_,
		_w24157_,
		_w24622_,
		_w24629_,
		_w24630_
	);
	LUT3 #(
		.INIT('h31)
	) name18804 (
		_w24062_,
		_w24628_,
		_w24630_,
		_w24631_
	);
	LUT3 #(
		.INIT('h65)
	) name18805 (
		\u1_desIn_r_reg[4]/NET0131 ,
		_w24626_,
		_w24631_,
		_w24632_
	);
	LUT3 #(
		.INIT('h84)
	) name18806 (
		_w24569_,
		_w24572_,
		_w24573_,
		_w24633_
	);
	LUT3 #(
		.INIT('h68)
	) name18807 (
		_w24569_,
		_w24572_,
		_w24573_,
		_w24634_
	);
	LUT4 #(
		.INIT('h0103)
	) name18808 (
		_w24569_,
		_w24572_,
		_w24573_,
		_w24577_,
		_w24635_
	);
	LUT3 #(
		.INIT('h01)
	) name18809 (
		_w24570_,
		_w24634_,
		_w24635_,
		_w24636_
	);
	LUT4 #(
		.INIT('h0012)
	) name18810 (
		_w24570_,
		_w24572_,
		_w24573_,
		_w24577_,
		_w24637_
	);
	LUT4 #(
		.INIT('h0080)
	) name18811 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24638_
	);
	LUT3 #(
		.INIT('h02)
	) name18812 (
		_w24586_,
		_w24638_,
		_w24637_,
		_w24639_
	);
	LUT4 #(
		.INIT('h9700)
	) name18813 (
		_w24569_,
		_w24572_,
		_w24573_,
		_w24577_,
		_w24640_
	);
	LUT4 #(
		.INIT('h00fe)
	) name18814 (
		_w24570_,
		_w24572_,
		_w24573_,
		_w24577_,
		_w24641_
	);
	LUT3 #(
		.INIT('h23)
	) name18815 (
		_w24633_,
		_w24640_,
		_w24641_,
		_w24642_
	);
	LUT2 #(
		.INIT('h1)
	) name18816 (
		_w24586_,
		_w24596_,
		_w24643_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name18817 (
		_w24636_,
		_w24639_,
		_w24642_,
		_w24643_,
		_w24644_
	);
	LUT2 #(
		.INIT('h8)
	) name18818 (
		_w24570_,
		_w24573_,
		_w24645_
	);
	LUT4 #(
		.INIT('h0040)
	) name18819 (
		_w24569_,
		_w24570_,
		_w24573_,
		_w24577_,
		_w24646_
	);
	LUT4 #(
		.INIT('hf7fb)
	) name18820 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24647_
	);
	LUT3 #(
		.INIT('h31)
	) name18821 (
		_w24577_,
		_w24646_,
		_w24647_,
		_w24648_
	);
	LUT3 #(
		.INIT('h65)
	) name18822 (
		\u1_desIn_r_reg[60]/NET0131 ,
		_w24644_,
		_w24648_,
		_w24649_
	);
	LUT4 #(
		.INIT('hfd75)
	) name18823 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24650_
	);
	LUT2 #(
		.INIT('h1)
	) name18824 (
		_w24240_,
		_w24650_,
		_w24651_
	);
	LUT4 #(
		.INIT('h0a20)
	) name18825 (
		_w24240_,
		_w24242_,
		_w24243_,
		_w24241_,
		_w24652_
	);
	LUT3 #(
		.INIT('h02)
	) name18826 (
		_w24239_,
		_w24259_,
		_w24652_,
		_w24653_
	);
	LUT2 #(
		.INIT('h4)
	) name18827 (
		_w24651_,
		_w24653_,
		_w24654_
	);
	LUT4 #(
		.INIT('h1003)
	) name18828 (
		_w24240_,
		_w24242_,
		_w24241_,
		_w24244_,
		_w24655_
	);
	LUT3 #(
		.INIT('h01)
	) name18829 (
		_w24239_,
		_w24320_,
		_w24304_,
		_w24656_
	);
	LUT4 #(
		.INIT('h8000)
	) name18830 (
		_w24240_,
		_w24242_,
		_w24243_,
		_w24241_,
		_w24657_
	);
	LUT2 #(
		.INIT('h1)
	) name18831 (
		_w24248_,
		_w24657_,
		_w24658_
	);
	LUT3 #(
		.INIT('h40)
	) name18832 (
		_w24655_,
		_w24656_,
		_w24658_,
		_w24659_
	);
	LUT4 #(
		.INIT('h1000)
	) name18833 (
		_w24240_,
		_w24242_,
		_w24243_,
		_w24241_,
		_w24660_
	);
	LUT4 #(
		.INIT('h77ef)
	) name18834 (
		_w24242_,
		_w24243_,
		_w24241_,
		_w24244_,
		_w24661_
	);
	LUT3 #(
		.INIT('h31)
	) name18835 (
		_w24240_,
		_w24660_,
		_w24661_,
		_w24662_
	);
	LUT4 #(
		.INIT('ha955)
	) name18836 (
		\u1_desIn_r_reg[10]/NET0131 ,
		_w24654_,
		_w24659_,
		_w24662_,
		_w24663_
	);
	LUT4 #(
		.INIT('hf900)
	) name18837 (
		_w24570_,
		_w24572_,
		_w24573_,
		_w24577_,
		_w24664_
	);
	LUT3 #(
		.INIT('h02)
	) name18838 (
		_w24569_,
		_w24572_,
		_w24573_,
		_w24665_
	);
	LUT4 #(
		.INIT('hbbf5)
	) name18839 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24666_
	);
	LUT2 #(
		.INIT('h8)
	) name18840 (
		_w24664_,
		_w24666_,
		_w24667_
	);
	LUT4 #(
		.INIT('h1001)
	) name18841 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24668_
	);
	LUT3 #(
		.INIT('h04)
	) name18842 (
		_w24577_,
		_w24588_,
		_w24668_,
		_w24669_
	);
	LUT4 #(
		.INIT('h0400)
	) name18843 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24670_
	);
	LUT2 #(
		.INIT('h1)
	) name18844 (
		_w24586_,
		_w24670_,
		_w24671_
	);
	LUT3 #(
		.INIT('he0)
	) name18845 (
		_w24667_,
		_w24669_,
		_w24671_,
		_w24672_
	);
	LUT2 #(
		.INIT('h2)
	) name18846 (
		_w24575_,
		_w24577_,
		_w24673_
	);
	LUT3 #(
		.INIT('h51)
	) name18847 (
		_w24569_,
		_w24572_,
		_w24573_,
		_w24674_
	);
	LUT2 #(
		.INIT('h8)
	) name18848 (
		_w24582_,
		_w24674_,
		_w24675_
	);
	LUT3 #(
		.INIT('h53)
	) name18849 (
		_w24569_,
		_w24572_,
		_w24573_,
		_w24676_
	);
	LUT2 #(
		.INIT('h8)
	) name18850 (
		_w24570_,
		_w24577_,
		_w24677_
	);
	LUT3 #(
		.INIT('h8a)
	) name18851 (
		_w24586_,
		_w24676_,
		_w24677_,
		_w24678_
	);
	LUT4 #(
		.INIT('h0100)
	) name18852 (
		_w24579_,
		_w24675_,
		_w24673_,
		_w24678_,
		_w24679_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name18853 (
		_w24574_,
		_w24582_,
		_w24581_,
		_w24592_,
		_w24680_
	);
	LUT4 #(
		.INIT('ha955)
	) name18854 (
		\u1_desIn_r_reg[58]/NET0131 ,
		_w24672_,
		_w24679_,
		_w24680_,
		_w24681_
	);
	LUT4 #(
		.INIT('h0100)
	) name18855 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24682_
	);
	LUT3 #(
		.INIT('h07)
	) name18856 (
		_w24570_,
		_w24573_,
		_w24577_,
		_w24683_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name18857 (
		_w24665_,
		_w24664_,
		_w24682_,
		_w24683_,
		_w24684_
	);
	LUT4 #(
		.INIT('h0040)
	) name18858 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24685_
	);
	LUT3 #(
		.INIT('h01)
	) name18859 (
		_w24586_,
		_w24668_,
		_w24685_,
		_w24686_
	);
	LUT4 #(
		.INIT('h39fd)
	) name18860 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24573_,
		_w24687_
	);
	LUT4 #(
		.INIT('hfb51)
	) name18861 (
		_w24577_,
		_w24592_,
		_w24645_,
		_w24687_,
		_w24688_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name18862 (
		_w24586_,
		_w24684_,
		_w24686_,
		_w24688_,
		_w24689_
	);
	LUT3 #(
		.INIT('h80)
	) name18863 (
		_w24572_,
		_w24573_,
		_w24577_,
		_w24690_
	);
	LUT2 #(
		.INIT('h8)
	) name18864 (
		_w24597_,
		_w24690_,
		_w24691_
	);
	LUT4 #(
		.INIT('h0008)
	) name18865 (
		_w24569_,
		_w24570_,
		_w24572_,
		_w24577_,
		_w24692_
	);
	LUT3 #(
		.INIT('h80)
	) name18866 (
		_w24569_,
		_w24570_,
		_w24586_,
		_w24693_
	);
	LUT3 #(
		.INIT('h23)
	) name18867 (
		_w24574_,
		_w24692_,
		_w24693_,
		_w24694_
	);
	LUT2 #(
		.INIT('h4)
	) name18868 (
		_w24691_,
		_w24694_,
		_w24695_
	);
	LUT3 #(
		.INIT('h9a)
	) name18869 (
		\u1_desIn_r_reg[40]/NET0131 ,
		_w24689_,
		_w24695_,
		_w24696_
	);
	LUT4 #(
		.INIT('hc963)
	) name18870 (
		decrypt_pad,
		\u0_R14_reg[29]/NET0131 ,
		\u0_uk_K_r14_reg[36]/NET0131 ,
		\u0_uk_K_r14_reg[43]/NET0131 ,
		_w24697_
	);
	LUT4 #(
		.INIT('hc963)
	) name18871 (
		decrypt_pad,
		\u0_R14_reg[30]/NET0131 ,
		\u0_uk_K_r14_reg[37]/NET0131 ,
		\u0_uk_K_r14_reg[44]/NET0131 ,
		_w24698_
	);
	LUT2 #(
		.INIT('h9)
	) name18872 (
		_w24697_,
		_w24698_,
		_w24699_
	);
	LUT4 #(
		.INIT('hc693)
	) name18873 (
		decrypt_pad,
		\u0_R14_reg[28]/NET0131 ,
		\u0_uk_K_r14_reg[16]/NET0131 ,
		\u0_uk_K_r14_reg[9]/NET0131 ,
		_w24700_
	);
	LUT4 #(
		.INIT('hc963)
	) name18874 (
		decrypt_pad,
		\u0_R14_reg[1]/NET0131 ,
		\u0_uk_K_r14_reg[21]/NET0131 ,
		\u0_uk_K_r14_reg[28]/NET0131 ,
		_w24701_
	);
	LUT4 #(
		.INIT('h0400)
	) name18875 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24702_
	);
	LUT4 #(
		.INIT('hebf6)
	) name18876 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24703_
	);
	LUT4 #(
		.INIT('h0200)
	) name18877 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24704_
	);
	LUT4 #(
		.INIT('hc693)
	) name18878 (
		decrypt_pad,
		\u0_R14_reg[31]/P0001 ,
		\u0_uk_K_r14_reg[1]/NET0131 ,
		\u0_uk_K_r14_reg[49]/NET0131 ,
		_w24705_
	);
	LUT4 #(
		.INIT('hfb00)
	) name18879 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24705_,
		_w24706_
	);
	LUT3 #(
		.INIT('h20)
	) name18880 (
		_w24703_,
		_w24704_,
		_w24706_,
		_w24707_
	);
	LUT4 #(
		.INIT('h0020)
	) name18881 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24708_
	);
	LUT2 #(
		.INIT('h8)
	) name18882 (
		_w24701_,
		_w24697_,
		_w24709_
	);
	LUT4 #(
		.INIT('h2e3f)
	) name18883 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24710_
	);
	LUT3 #(
		.INIT('h10)
	) name18884 (
		_w24705_,
		_w24708_,
		_w24710_,
		_w24711_
	);
	LUT4 #(
		.INIT('hc963)
	) name18885 (
		decrypt_pad,
		\u0_R14_reg[32]/NET0131 ,
		\u0_uk_K_r14_reg[0]/NET0131 ,
		\u0_uk_K_r14_reg[7]/NET0131 ,
		_w24712_
	);
	LUT3 #(
		.INIT('h02)
	) name18886 (
		_w24700_,
		_w24698_,
		_w24705_,
		_w24713_
	);
	LUT4 #(
		.INIT('h8000)
	) name18887 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24714_
	);
	LUT4 #(
		.INIT('h0001)
	) name18888 (
		_w24708_,
		_w24712_,
		_w24713_,
		_w24714_,
		_w24715_
	);
	LUT3 #(
		.INIT('he0)
	) name18889 (
		_w24707_,
		_w24711_,
		_w24715_,
		_w24716_
	);
	LUT3 #(
		.INIT('hde)
	) name18890 (
		_w24700_,
		_w24697_,
		_w24698_,
		_w24717_
	);
	LUT3 #(
		.INIT('h10)
	) name18891 (
		_w24705_,
		_w24708_,
		_w24717_,
		_w24718_
	);
	LUT4 #(
		.INIT('h309a)
	) name18892 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24719_
	);
	LUT3 #(
		.INIT('h08)
	) name18893 (
		_w24703_,
		_w24705_,
		_w24719_,
		_w24720_
	);
	LUT4 #(
		.INIT('h4000)
	) name18894 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24721_
	);
	LUT2 #(
		.INIT('h2)
	) name18895 (
		_w24712_,
		_w24721_,
		_w24722_
	);
	LUT3 #(
		.INIT('he0)
	) name18896 (
		_w24718_,
		_w24720_,
		_w24722_,
		_w24723_
	);
	LUT3 #(
		.INIT('h56)
	) name18897 (
		\u0_L14_reg[5]/P0001 ,
		_w24716_,
		_w24723_,
		_w24724_
	);
	LUT4 #(
		.INIT('hc693)
	) name18898 (
		decrypt_pad,
		\u0_R14_reg[4]/NET0131 ,
		\u0_uk_K_r14_reg[13]/NET0131 ,
		\u0_uk_K_r14_reg[6]/NET0131 ,
		_w24725_
	);
	LUT4 #(
		.INIT('hc693)
	) name18899 (
		decrypt_pad,
		\u0_R14_reg[3]/NET0131 ,
		\u0_uk_K_r14_reg[3]/NET0131 ,
		\u0_uk_K_r14_reg[53]/NET0131 ,
		_w24726_
	);
	LUT4 #(
		.INIT('hc963)
	) name18900 (
		decrypt_pad,
		\u0_R14_reg[32]/NET0131 ,
		\u0_uk_K_r14_reg[40]/NET0131 ,
		\u0_uk_K_r14_reg[47]/NET0131 ,
		_w24727_
	);
	LUT4 #(
		.INIT('hc693)
	) name18901 (
		decrypt_pad,
		\u0_R14_reg[1]/NET0131 ,
		\u0_uk_K_r14_reg[11]/NET0131 ,
		\u0_uk_K_r14_reg[4]/NET0131 ,
		_w24728_
	);
	LUT4 #(
		.INIT('hc963)
	) name18902 (
		decrypt_pad,
		\u0_R14_reg[5]/NET0131 ,
		\u0_uk_K_r14_reg[34]/NET0131 ,
		\u0_uk_K_r14_reg[41]/NET0131 ,
		_w24729_
	);
	LUT4 #(
		.INIT('hc963)
	) name18903 (
		decrypt_pad,
		\u0_R14_reg[2]/NET0131 ,
		\u0_uk_K_r14_reg[19]/NET0131 ,
		\u0_uk_K_r14_reg[26]/NET0131 ,
		_w24730_
	);
	LUT4 #(
		.INIT('h0800)
	) name18904 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24731_
	);
	LUT4 #(
		.INIT('hd7df)
	) name18905 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24732_
	);
	LUT2 #(
		.INIT('h2)
	) name18906 (
		_w24726_,
		_w24732_,
		_w24733_
	);
	LUT2 #(
		.INIT('h2)
	) name18907 (
		_w24726_,
		_w24728_,
		_w24734_
	);
	LUT3 #(
		.INIT('h10)
	) name18908 (
		_w24727_,
		_w24729_,
		_w24730_,
		_w24735_
	);
	LUT4 #(
		.INIT('h0040)
	) name18909 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24736_
	);
	LUT3 #(
		.INIT('h07)
	) name18910 (
		_w24734_,
		_w24735_,
		_w24736_,
		_w24737_
	);
	LUT3 #(
		.INIT('h8a)
	) name18911 (
		_w24725_,
		_w24733_,
		_w24737_,
		_w24738_
	);
	LUT4 #(
		.INIT('h23ff)
	) name18912 (
		_w24726_,
		_w24728_,
		_w24727_,
		_w24729_,
		_w24739_
	);
	LUT2 #(
		.INIT('h2)
	) name18913 (
		_w24730_,
		_w24739_,
		_w24740_
	);
	LUT3 #(
		.INIT('h02)
	) name18914 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24741_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name18915 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24742_
	);
	LUT2 #(
		.INIT('h4)
	) name18916 (
		_w24726_,
		_w24728_,
		_w24743_
	);
	LUT3 #(
		.INIT('h40)
	) name18917 (
		_w24726_,
		_w24728_,
		_w24727_,
		_w24744_
	);
	LUT3 #(
		.INIT('h01)
	) name18918 (
		_w24728_,
		_w24729_,
		_w24730_,
		_w24745_
	);
	LUT4 #(
		.INIT('h0031)
	) name18919 (
		_w24726_,
		_w24744_,
		_w24742_,
		_w24745_,
		_w24746_
	);
	LUT3 #(
		.INIT('h45)
	) name18920 (
		_w24725_,
		_w24740_,
		_w24746_,
		_w24747_
	);
	LUT3 #(
		.INIT('h80)
	) name18921 (
		_w24728_,
		_w24729_,
		_w24730_,
		_w24748_
	);
	LUT4 #(
		.INIT('h0008)
	) name18922 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24749_
	);
	LUT4 #(
		.INIT('h7fe7)
	) name18923 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24750_
	);
	LUT2 #(
		.INIT('h1)
	) name18924 (
		_w24726_,
		_w24750_,
		_w24751_
	);
	LUT4 #(
		.INIT('he9ed)
	) name18925 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24752_
	);
	LUT2 #(
		.INIT('h2)
	) name18926 (
		_w24725_,
		_w24726_,
		_w24753_
	);
	LUT2 #(
		.INIT('h4)
	) name18927 (
		_w24752_,
		_w24753_,
		_w24754_
	);
	LUT2 #(
		.INIT('h2)
	) name18928 (
		_w24726_,
		_w24730_,
		_w24755_
	);
	LUT4 #(
		.INIT('h0020)
	) name18929 (
		_w24726_,
		_w24728_,
		_w24727_,
		_w24730_,
		_w24756_
	);
	LUT3 #(
		.INIT('h07)
	) name18930 (
		_w24741_,
		_w24755_,
		_w24756_,
		_w24757_
	);
	LUT3 #(
		.INIT('h10)
	) name18931 (
		_w24751_,
		_w24754_,
		_w24757_,
		_w24758_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name18932 (
		\u0_L14_reg[23]/P0001 ,
		_w24747_,
		_w24738_,
		_w24758_,
		_w24759_
	);
	LUT4 #(
		.INIT('h0002)
	) name18933 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24760_
	);
	LUT4 #(
		.INIT('h5b4b)
	) name18934 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24761_
	);
	LUT4 #(
		.INIT('h3032)
	) name18935 (
		_w24705_,
		_w24712_,
		_w24760_,
		_w24761_,
		_w24762_
	);
	LUT4 #(
		.INIT('h10a0)
	) name18936 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24763_
	);
	LUT4 #(
		.INIT('h0800)
	) name18937 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24764_
	);
	LUT4 #(
		.INIT('h0020)
	) name18938 (
		_w24701_,
		_w24697_,
		_w24698_,
		_w24705_,
		_w24765_
	);
	LUT4 #(
		.INIT('h0100)
	) name18939 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24705_,
		_w24766_
	);
	LUT4 #(
		.INIT('h0001)
	) name18940 (
		_w24765_,
		_w24763_,
		_w24766_,
		_w24764_,
		_w24767_
	);
	LUT4 #(
		.INIT('he5be)
	) name18941 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24768_
	);
	LUT2 #(
		.INIT('h1)
	) name18942 (
		_w24705_,
		_w24768_,
		_w24769_
	);
	LUT4 #(
		.INIT('h0002)
	) name18943 (
		_w24700_,
		_w24697_,
		_w24705_,
		_w24712_,
		_w24770_
	);
	LUT3 #(
		.INIT('h40)
	) name18944 (
		_w24700_,
		_w24701_,
		_w24705_,
		_w24771_
	);
	LUT3 #(
		.INIT('h13)
	) name18945 (
		_w24699_,
		_w24770_,
		_w24771_,
		_w24772_
	);
	LUT4 #(
		.INIT('h0d00)
	) name18946 (
		_w24712_,
		_w24767_,
		_w24769_,
		_w24772_,
		_w24773_
	);
	LUT3 #(
		.INIT('h65)
	) name18947 (
		\u0_L14_reg[15]/P0001 ,
		_w24762_,
		_w24773_,
		_w24774_
	);
	LUT4 #(
		.INIT('h9f9a)
	) name18948 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24775_
	);
	LUT4 #(
		.INIT('h7f6f)
	) name18949 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24776_
	);
	LUT4 #(
		.INIT('hbdf3)
	) name18950 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24777_
	);
	LUT4 #(
		.INIT('hd800)
	) name18951 (
		_w24705_,
		_w24776_,
		_w24775_,
		_w24777_,
		_w24778_
	);
	LUT2 #(
		.INIT('h2)
	) name18952 (
		_w24712_,
		_w24778_,
		_w24779_
	);
	LUT4 #(
		.INIT('hbf00)
	) name18953 (
		_w24700_,
		_w24697_,
		_w24698_,
		_w24705_,
		_w24780_
	);
	LUT3 #(
		.INIT('h59)
	) name18954 (
		_w24701_,
		_w24697_,
		_w24698_,
		_w24781_
	);
	LUT2 #(
		.INIT('h8)
	) name18955 (
		_w24780_,
		_w24781_,
		_w24782_
	);
	LUT4 #(
		.INIT('h0010)
	) name18956 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24705_,
		_w24783_
	);
	LUT4 #(
		.INIT('h0080)
	) name18957 (
		_w24700_,
		_w24701_,
		_w24698_,
		_w24705_,
		_w24784_
	);
	LUT3 #(
		.INIT('h01)
	) name18958 (
		_w24702_,
		_w24784_,
		_w24783_,
		_w24785_
	);
	LUT4 #(
		.INIT('h1000)
	) name18959 (
		_w24701_,
		_w24697_,
		_w24698_,
		_w24705_,
		_w24786_
	);
	LUT4 #(
		.INIT('hefd7)
	) name18960 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w24787_
	);
	LUT3 #(
		.INIT('h32)
	) name18961 (
		_w24705_,
		_w24786_,
		_w24787_,
		_w24788_
	);
	LUT4 #(
		.INIT('hba00)
	) name18962 (
		_w24712_,
		_w24782_,
		_w24785_,
		_w24788_,
		_w24789_
	);
	LUT3 #(
		.INIT('h65)
	) name18963 (
		\u0_L14_reg[27]/P0001 ,
		_w24779_,
		_w24789_,
		_w24790_
	);
	LUT4 #(
		.INIT('hc963)
	) name18964 (
		decrypt_pad,
		\u0_R14_reg[20]/NET0131 ,
		\u0_uk_K_r14_reg[16]/NET0131 ,
		\u0_uk_K_r14_reg[23]/NET0131 ,
		_w24791_
	);
	LUT4 #(
		.INIT('hc963)
	) name18965 (
		decrypt_pad,
		\u0_R14_reg[19]/NET0131 ,
		\u0_uk_K_r14_reg[1]/NET0131 ,
		\u0_uk_K_r14_reg[8]/NET0131 ,
		_w24792_
	);
	LUT4 #(
		.INIT('hc693)
	) name18966 (
		decrypt_pad,
		\u0_R14_reg[17]/NET0131 ,
		\u0_uk_K_r14_reg[31]/NET0131 ,
		\u0_uk_K_r14_reg[51]/NET0131 ,
		_w24793_
	);
	LUT4 #(
		.INIT('hc963)
	) name18967 (
		decrypt_pad,
		\u0_R14_reg[21]/NET0131 ,
		\u0_uk_K_r14_reg[45]/NET0131 ,
		\u0_uk_K_r14_reg[52]/NET0131 ,
		_w24794_
	);
	LUT4 #(
		.INIT('hc963)
	) name18968 (
		decrypt_pad,
		\u0_R14_reg[16]/NET0131 ,
		\u0_uk_K_r14_reg[29]/NET0131 ,
		\u0_uk_K_r14_reg[36]/NET0131 ,
		_w24795_
	);
	LUT4 #(
		.INIT('hc963)
	) name18969 (
		decrypt_pad,
		\u0_R14_reg[18]/NET0131 ,
		\u0_uk_K_r14_reg[14]/NET0131 ,
		\u0_uk_K_r14_reg[21]/NET0131 ,
		_w24796_
	);
	LUT4 #(
		.INIT('h44e6)
	) name18970 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24797_
	);
	LUT4 #(
		.INIT('h0b00)
	) name18971 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24798_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name18972 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24799_
	);
	LUT4 #(
		.INIT('h4540)
	) name18973 (
		_w24798_,
		_w24799_,
		_w24792_,
		_w24797_,
		_w24800_
	);
	LUT2 #(
		.INIT('h1)
	) name18974 (
		_w24791_,
		_w24800_,
		_w24801_
	);
	LUT4 #(
		.INIT('h0004)
	) name18975 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24802_
	);
	LUT4 #(
		.INIT('h0200)
	) name18976 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24803_
	);
	LUT3 #(
		.INIT('h02)
	) name18977 (
		_w24792_,
		_w24802_,
		_w24803_,
		_w24804_
	);
	LUT4 #(
		.INIT('h0001)
	) name18978 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24805_
	);
	LUT4 #(
		.INIT('h0800)
	) name18979 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24806_
	);
	LUT4 #(
		.INIT('h0040)
	) name18980 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24807_
	);
	LUT4 #(
		.INIT('h0001)
	) name18981 (
		_w24792_,
		_w24807_,
		_w24806_,
		_w24805_,
		_w24808_
	);
	LUT2 #(
		.INIT('h1)
	) name18982 (
		_w24804_,
		_w24808_,
		_w24809_
	);
	LUT4 #(
		.INIT('hef67)
	) name18983 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24810_
	);
	LUT2 #(
		.INIT('h2)
	) name18984 (
		_w24792_,
		_w24810_,
		_w24811_
	);
	LUT4 #(
		.INIT('h0080)
	) name18985 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24812_
	);
	LUT4 #(
		.INIT('h0400)
	) name18986 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w24813_
	);
	LUT2 #(
		.INIT('h2)
	) name18987 (
		_w24793_,
		_w24792_,
		_w24814_
	);
	LUT4 #(
		.INIT('h0020)
	) name18988 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24792_,
		_w24815_
	);
	LUT3 #(
		.INIT('h01)
	) name18989 (
		_w24813_,
		_w24815_,
		_w24812_,
		_w24816_
	);
	LUT3 #(
		.INIT('h8a)
	) name18990 (
		_w24791_,
		_w24811_,
		_w24816_,
		_w24817_
	);
	LUT4 #(
		.INIT('h5556)
	) name18991 (
		\u0_L14_reg[3]/P0001 ,
		_w24801_,
		_w24809_,
		_w24817_,
		_w24818_
	);
	LUT3 #(
		.INIT('hb7)
	) name18992 (
		_w24727_,
		_w24729_,
		_w24730_,
		_w24819_
	);
	LUT2 #(
		.INIT('h2)
	) name18993 (
		_w24743_,
		_w24819_,
		_w24820_
	);
	LUT2 #(
		.INIT('h4)
	) name18994 (
		_w24727_,
		_w24729_,
		_w24821_
	);
	LUT3 #(
		.INIT('h41)
	) name18995 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24822_
	);
	LUT4 #(
		.INIT('h4180)
	) name18996 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24823_
	);
	LUT4 #(
		.INIT('ha5ad)
	) name18997 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24824_
	);
	LUT3 #(
		.INIT('h25)
	) name18998 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24825_
	);
	LUT4 #(
		.INIT('h4501)
	) name18999 (
		_w24725_,
		_w24726_,
		_w24825_,
		_w24824_,
		_w24826_
	);
	LUT4 #(
		.INIT('h9600)
	) name19000 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w24827_
	);
	LUT4 #(
		.INIT('h020a)
	) name19001 (
		_w24725_,
		_w24755_,
		_w24749_,
		_w24825_,
		_w24828_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name19002 (
		_w24823_,
		_w24826_,
		_w24827_,
		_w24828_,
		_w24829_
	);
	LUT3 #(
		.INIT('h56)
	) name19003 (
		\u0_L14_reg[9]/P0001 ,
		_w24820_,
		_w24829_,
		_w24830_
	);
	LUT4 #(
		.INIT('hc963)
	) name19004 (
		decrypt_pad,
		\u0_R14_reg[8]/NET0131 ,
		\u0_uk_K_r14_reg[32]/NET0131 ,
		\u0_uk_K_r14_reg[39]/P0001 ,
		_w24831_
	);
	LUT4 #(
		.INIT('hc963)
	) name19005 (
		decrypt_pad,
		\u0_R14_reg[7]/NET0131 ,
		\u0_uk_K_r14_reg[41]/NET0131 ,
		\u0_uk_K_r14_reg[48]/NET0131 ,
		_w24832_
	);
	LUT4 #(
		.INIT('hc963)
	) name19006 (
		decrypt_pad,
		\u0_R14_reg[5]/NET0131 ,
		\u0_uk_K_r14_reg[24]/NET0131 ,
		\u0_uk_K_r14_reg[6]/NET0131 ,
		_w24833_
	);
	LUT4 #(
		.INIT('hc963)
	) name19007 (
		decrypt_pad,
		\u0_R14_reg[4]/NET0131 ,
		\u0_uk_K_r14_reg[20]/NET0131 ,
		\u0_uk_K_r14_reg[27]/NET0131 ,
		_w24834_
	);
	LUT4 #(
		.INIT('hc963)
	) name19008 (
		decrypt_pad,
		\u0_R14_reg[9]/NET0131 ,
		\u0_uk_K_r14_reg[12]/NET0131 ,
		\u0_uk_K_r14_reg[19]/NET0131 ,
		_w24835_
	);
	LUT4 #(
		.INIT('hc963)
	) name19009 (
		decrypt_pad,
		\u0_R14_reg[6]/NET0131 ,
		\u0_uk_K_r14_reg[47]/NET0131 ,
		\u0_uk_K_r14_reg[54]/NET0131 ,
		_w24836_
	);
	LUT4 #(
		.INIT('hfd75)
	) name19010 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w24837_
	);
	LUT3 #(
		.INIT('hcb)
	) name19011 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24838_
	);
	LUT3 #(
		.INIT('h10)
	) name19012 (
		_w24834_,
		_w24833_,
		_w24836_,
		_w24839_
	);
	LUT4 #(
		.INIT('h0100)
	) name19013 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w24840_
	);
	LUT4 #(
		.INIT('h00d8)
	) name19014 (
		_w24832_,
		_w24838_,
		_w24837_,
		_w24840_,
		_w24841_
	);
	LUT4 #(
		.INIT('h0411)
	) name19015 (
		_w24834_,
		_w24833_,
		_w24832_,
		_w24836_,
		_w24842_
	);
	LUT4 #(
		.INIT('h8000)
	) name19016 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24832_,
		_w24843_
	);
	LUT4 #(
		.INIT('h0800)
	) name19017 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w24844_
	);
	LUT4 #(
		.INIT('h2000)
	) name19018 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w24845_
	);
	LUT4 #(
		.INIT('hd7fc)
	) name19019 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w24846_
	);
	LUT3 #(
		.INIT('h10)
	) name19020 (
		_w24842_,
		_w24843_,
		_w24846_,
		_w24847_
	);
	LUT4 #(
		.INIT('h0040)
	) name19021 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24832_,
		_w24848_
	);
	LUT4 #(
		.INIT('h0010)
	) name19022 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w24849_
	);
	LUT4 #(
		.INIT('h77ef)
	) name19023 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w24850_
	);
	LUT3 #(
		.INIT('h31)
	) name19024 (
		_w24832_,
		_w24848_,
		_w24850_,
		_w24851_
	);
	LUT4 #(
		.INIT('he400)
	) name19025 (
		_w24831_,
		_w24847_,
		_w24841_,
		_w24851_,
		_w24852_
	);
	LUT2 #(
		.INIT('h9)
	) name19026 (
		\u0_L14_reg[18]/P0001 ,
		_w24852_,
		_w24853_
	);
	LUT4 #(
		.INIT('hc963)
	) name19027 (
		decrypt_pad,
		\u0_R14_reg[12]/NET0131 ,
		\u0_uk_K_r14_reg[10]/P0001 ,
		\u0_uk_K_r14_reg[17]/NET0131 ,
		_w24854_
	);
	LUT4 #(
		.INIT('hc963)
	) name19028 (
		decrypt_pad,
		\u0_R14_reg[9]/NET0131 ,
		\u0_uk_K_r14_reg[18]/NET0131 ,
		\u0_uk_K_r14_reg[25]/NET0131 ,
		_w24855_
	);
	LUT4 #(
		.INIT('hc963)
	) name19029 (
		decrypt_pad,
		\u0_R14_reg[10]/NET0131 ,
		\u0_uk_K_r14_reg[26]/NET0131 ,
		\u0_uk_K_r14_reg[33]/NET0131 ,
		_w24856_
	);
	LUT4 #(
		.INIT('hc963)
	) name19030 (
		decrypt_pad,
		\u0_R14_reg[13]/NET0131 ,
		\u0_uk_K_r14_reg[55]/NET0131 ,
		\u0_uk_K_r14_reg[5]/NET0131 ,
		_w24857_
	);
	LUT4 #(
		.INIT('hc963)
	) name19031 (
		decrypt_pad,
		\u0_R14_reg[8]/NET0131 ,
		\u0_uk_K_r14_reg[46]/NET0131 ,
		\u0_uk_K_r14_reg[53]/NET0131 ,
		_w24858_
	);
	LUT4 #(
		.INIT('h0100)
	) name19032 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24859_
	);
	LUT4 #(
		.INIT('hc963)
	) name19033 (
		decrypt_pad,
		\u0_R14_reg[11]/P0001 ,
		\u0_uk_K_r14_reg[27]/NET0131 ,
		\u0_uk_K_r14_reg[34]/NET0131 ,
		_w24860_
	);
	LUT2 #(
		.INIT('h2)
	) name19034 (
		_w24857_,
		_w24858_,
		_w24861_
	);
	LUT3 #(
		.INIT('h02)
	) name19035 (
		_w24857_,
		_w24856_,
		_w24858_,
		_w24862_
	);
	LUT4 #(
		.INIT('hcc84)
	) name19036 (
		_w24857_,
		_w24860_,
		_w24856_,
		_w24858_,
		_w24863_
	);
	LUT3 #(
		.INIT('h04)
	) name19037 (
		_w24857_,
		_w24855_,
		_w24858_,
		_w24864_
	);
	LUT3 #(
		.INIT('h15)
	) name19038 (
		_w24860_,
		_w24856_,
		_w24858_,
		_w24865_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name19039 (
		_w24859_,
		_w24863_,
		_w24864_,
		_w24865_,
		_w24866_
	);
	LUT2 #(
		.INIT('h2)
	) name19040 (
		_w24854_,
		_w24866_,
		_w24867_
	);
	LUT4 #(
		.INIT('h4bfb)
	) name19041 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24868_
	);
	LUT2 #(
		.INIT('h2)
	) name19042 (
		_w24860_,
		_w24868_,
		_w24869_
	);
	LUT3 #(
		.INIT('h0b)
	) name19043 (
		_w24857_,
		_w24855_,
		_w24860_,
		_w24870_
	);
	LUT3 #(
		.INIT('h3a)
	) name19044 (
		_w24855_,
		_w24856_,
		_w24858_,
		_w24871_
	);
	LUT2 #(
		.INIT('h8)
	) name19045 (
		_w24870_,
		_w24871_,
		_w24872_
	);
	LUT2 #(
		.INIT('h8)
	) name19046 (
		_w24857_,
		_w24858_,
		_w24873_
	);
	LUT4 #(
		.INIT('h0201)
	) name19047 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24874_
	);
	LUT4 #(
		.INIT('h0020)
	) name19048 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24875_
	);
	LUT3 #(
		.INIT('h01)
	) name19049 (
		_w24854_,
		_w24875_,
		_w24874_,
		_w24876_
	);
	LUT3 #(
		.INIT('h10)
	) name19050 (
		_w24869_,
		_w24872_,
		_w24876_,
		_w24877_
	);
	LUT2 #(
		.INIT('h8)
	) name19051 (
		_w24857_,
		_w24860_,
		_w24878_
	);
	LUT3 #(
		.INIT('h40)
	) name19052 (
		_w24855_,
		_w24856_,
		_w24858_,
		_w24879_
	);
	LUT2 #(
		.INIT('h8)
	) name19053 (
		_w24878_,
		_w24879_,
		_w24880_
	);
	LUT4 #(
		.INIT('h0400)
	) name19054 (
		_w24857_,
		_w24855_,
		_w24860_,
		_w24856_,
		_w24881_
	);
	LUT2 #(
		.INIT('h8)
	) name19055 (
		_w24856_,
		_w24854_,
		_w24882_
	);
	LUT3 #(
		.INIT('h4c)
	) name19056 (
		_w24857_,
		_w24855_,
		_w24858_,
		_w24883_
	);
	LUT3 #(
		.INIT('h15)
	) name19057 (
		_w24881_,
		_w24882_,
		_w24883_,
		_w24884_
	);
	LUT2 #(
		.INIT('h4)
	) name19058 (
		_w24880_,
		_w24884_,
		_w24885_
	);
	LUT4 #(
		.INIT('h56aa)
	) name19059 (
		\u0_L14_reg[30]/P0001 ,
		_w24867_,
		_w24877_,
		_w24885_,
		_w24886_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name19060 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24887_
	);
	LUT3 #(
		.INIT('hc8)
	) name19061 (
		_w24855_,
		_w24860_,
		_w24856_,
		_w24888_
	);
	LUT4 #(
		.INIT('h0302)
	) name19062 (
		_w24860_,
		_w24861_,
		_w24888_,
		_w24887_,
		_w24889_
	);
	LUT2 #(
		.INIT('h1)
	) name19063 (
		_w24855_,
		_w24860_,
		_w24890_
	);
	LUT3 #(
		.INIT('h15)
	) name19064 (
		_w24859_,
		_w24862_,
		_w24890_,
		_w24891_
	);
	LUT2 #(
		.INIT('h4)
	) name19065 (
		_w24855_,
		_w24858_,
		_w24892_
	);
	LUT4 #(
		.INIT('hc080)
	) name19066 (
		_w24857_,
		_w24860_,
		_w24856_,
		_w24858_,
		_w24893_
	);
	LUT2 #(
		.INIT('h4)
	) name19067 (
		_w24892_,
		_w24893_,
		_w24894_
	);
	LUT4 #(
		.INIT('haaa2)
	) name19068 (
		_w24854_,
		_w24891_,
		_w24894_,
		_w24889_,
		_w24895_
	);
	LUT4 #(
		.INIT('hcfa1)
	) name19069 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24896_
	);
	LUT4 #(
		.INIT('h1000)
	) name19070 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24897_
	);
	LUT4 #(
		.INIT('h3302)
	) name19071 (
		_w24860_,
		_w24854_,
		_w24896_,
		_w24897_,
		_w24898_
	);
	LUT4 #(
		.INIT('hb95e)
	) name19072 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24899_
	);
	LUT2 #(
		.INIT('h1)
	) name19073 (
		_w24860_,
		_w24854_,
		_w24900_
	);
	LUT2 #(
		.INIT('h4)
	) name19074 (
		_w24899_,
		_w24900_,
		_w24901_
	);
	LUT4 #(
		.INIT('h0008)
	) name19075 (
		_w24855_,
		_w24860_,
		_w24856_,
		_w24858_,
		_w24902_
	);
	LUT2 #(
		.INIT('h8)
	) name19076 (
		_w24857_,
		_w24902_,
		_w24903_
	);
	LUT3 #(
		.INIT('h20)
	) name19077 (
		_w24855_,
		_w24860_,
		_w24856_,
		_w24904_
	);
	LUT4 #(
		.INIT('h0777)
	) name19078 (
		_w24860_,
		_w24859_,
		_w24873_,
		_w24904_,
		_w24905_
	);
	LUT4 #(
		.INIT('h0100)
	) name19079 (
		_w24898_,
		_w24903_,
		_w24901_,
		_w24905_,
		_w24906_
	);
	LUT3 #(
		.INIT('h65)
	) name19080 (
		\u0_L14_reg[24]/P0001 ,
		_w24895_,
		_w24906_,
		_w24907_
	);
	LUT4 #(
		.INIT('h669d)
	) name19081 (
		_w24857_,
		_w24855_,
		_w24860_,
		_w24858_,
		_w24908_
	);
	LUT4 #(
		.INIT('h0080)
	) name19082 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24909_
	);
	LUT4 #(
		.INIT('h0110)
	) name19083 (
		_w24857_,
		_w24860_,
		_w24856_,
		_w24858_,
		_w24910_
	);
	LUT4 #(
		.INIT('h0032)
	) name19084 (
		_w24856_,
		_w24909_,
		_w24908_,
		_w24910_,
		_w24911_
	);
	LUT4 #(
		.INIT('h77d8)
	) name19085 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24912_
	);
	LUT4 #(
		.INIT('h0001)
	) name19086 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24913_
	);
	LUT4 #(
		.INIT('h9f7f)
	) name19087 (
		_w24857_,
		_w24855_,
		_w24860_,
		_w24858_,
		_w24914_
	);
	LUT4 #(
		.INIT('h0e00)
	) name19088 (
		_w24860_,
		_w24912_,
		_w24913_,
		_w24914_,
		_w24915_
	);
	LUT4 #(
		.INIT('h4000)
	) name19089 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24916_
	);
	LUT4 #(
		.INIT('hbfef)
	) name19090 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w24917_
	);
	LUT4 #(
		.INIT('h1000)
	) name19091 (
		_w24855_,
		_w24860_,
		_w24856_,
		_w24858_,
		_w24918_
	);
	LUT3 #(
		.INIT('h0d)
	) name19092 (
		_w24860_,
		_w24917_,
		_w24918_,
		_w24919_
	);
	LUT4 #(
		.INIT('he400)
	) name19093 (
		_w24854_,
		_w24915_,
		_w24911_,
		_w24919_,
		_w24920_
	);
	LUT2 #(
		.INIT('h9)
	) name19094 (
		\u0_L14_reg[16]/P0001 ,
		_w24920_,
		_w24921_
	);
	LUT4 #(
		.INIT('hc963)
	) name19095 (
		decrypt_pad,
		\u0_R13_reg[27]/P0001 ,
		\u0_uk_K_r13_reg[45]/NET0131 ,
		\u0_uk_K_r13_reg[7]/NET0131 ,
		_w24922_
	);
	LUT4 #(
		.INIT('hc693)
	) name19096 (
		decrypt_pad,
		\u0_R13_reg[29]/NET0131 ,
		\u0_uk_K_r13_reg[45]/NET0131 ,
		\u0_uk_K_r13_reg[51]/NET0131 ,
		_w24923_
	);
	LUT4 #(
		.INIT('hc963)
	) name19097 (
		decrypt_pad,
		\u0_R13_reg[25]/NET0131 ,
		\u0_uk_K_r13_reg[23]/NET0131 ,
		\u0_uk_K_r13_reg[44]/NET0131 ,
		_w24924_
	);
	LUT4 #(
		.INIT('hc693)
	) name19098 (
		decrypt_pad,
		\u0_R13_reg[26]/NET0131 ,
		\u0_uk_K_r13_reg[29]/NET0131 ,
		\u0_uk_K_r13_reg[8]/NET0131 ,
		_w24925_
	);
	LUT4 #(
		.INIT('hc963)
	) name19099 (
		decrypt_pad,
		\u0_R13_reg[24]/NET0131 ,
		\u0_uk_K_r13_reg[43]/NET0131 ,
		\u0_uk_K_r13_reg[9]/NET0131 ,
		_w24926_
	);
	LUT2 #(
		.INIT('h9)
	) name19100 (
		_w24924_,
		_w24926_,
		_w24927_
	);
	LUT4 #(
		.INIT('h0020)
	) name19101 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w24928_
	);
	LUT4 #(
		.INIT('hee9e)
	) name19102 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w24929_
	);
	LUT2 #(
		.INIT('h2)
	) name19103 (
		_w24922_,
		_w24929_,
		_w24930_
	);
	LUT4 #(
		.INIT('hc7ff)
	) name19104 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w24931_
	);
	LUT2 #(
		.INIT('h4)
	) name19105 (
		_w24931_,
		_w24922_,
		_w24932_
	);
	LUT4 #(
		.INIT('h002a)
	) name19106 (
		_w24923_,
		_w24925_,
		_w24926_,
		_w24922_,
		_w24933_
	);
	LUT4 #(
		.INIT('h0021)
	) name19107 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w24934_
	);
	LUT4 #(
		.INIT('hc963)
	) name19108 (
		decrypt_pad,
		\u0_R13_reg[28]/NET0131 ,
		\u0_uk_K_r13_reg[28]/NET0131 ,
		\u0_uk_K_r13_reg[49]/NET0131 ,
		_w24935_
	);
	LUT4 #(
		.INIT('h4044)
	) name19109 (
		_w24934_,
		_w24935_,
		_w24927_,
		_w24933_,
		_w24936_
	);
	LUT2 #(
		.INIT('h4)
	) name19110 (
		_w24932_,
		_w24936_,
		_w24937_
	);
	LUT4 #(
		.INIT('h0010)
	) name19111 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w24938_
	);
	LUT4 #(
		.INIT('h1bef)
	) name19112 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w24939_
	);
	LUT2 #(
		.INIT('h1)
	) name19113 (
		_w24922_,
		_w24939_,
		_w24940_
	);
	LUT3 #(
		.INIT('h08)
	) name19114 (
		_w24923_,
		_w24926_,
		_w24922_,
		_w24941_
	);
	LUT4 #(
		.INIT('hcf45)
	) name19115 (
		_w24923_,
		_w24924_,
		_w24926_,
		_w24922_,
		_w24942_
	);
	LUT3 #(
		.INIT('h01)
	) name19116 (
		_w24925_,
		_w24942_,
		_w24941_,
		_w24943_
	);
	LUT4 #(
		.INIT('h8008)
	) name19117 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w24944_
	);
	LUT2 #(
		.INIT('h1)
	) name19118 (
		_w24935_,
		_w24944_,
		_w24945_
	);
	LUT3 #(
		.INIT('h10)
	) name19119 (
		_w24943_,
		_w24940_,
		_w24945_,
		_w24946_
	);
	LUT4 #(
		.INIT('h0082)
	) name19120 (
		_w24924_,
		_w24925_,
		_w24926_,
		_w24922_,
		_w24947_
	);
	LUT4 #(
		.INIT('h000e)
	) name19121 (
		_w24937_,
		_w24946_,
		_w24930_,
		_w24947_,
		_w24948_
	);
	LUT2 #(
		.INIT('h9)
	) name19122 (
		\u0_L13_reg[22]/NET0131 ,
		_w24948_,
		_w24949_
	);
	LUT4 #(
		.INIT('hc693)
	) name19123 (
		decrypt_pad,
		\u0_R13_reg[4]/NET0131 ,
		\u0_uk_K_r13_reg[20]/NET0131 ,
		\u0_uk_K_r13_reg[24]/NET0131 ,
		_w24950_
	);
	LUT4 #(
		.INIT('hc963)
	) name19124 (
		decrypt_pad,
		\u0_R13_reg[5]/NET0131 ,
		\u0_uk_K_r13_reg[27]/NET0131 ,
		\u0_uk_K_r13_reg[48]/NET0131 ,
		_w24951_
	);
	LUT4 #(
		.INIT('hc963)
	) name19125 (
		decrypt_pad,
		\u0_R13_reg[32]/NET0131 ,
		\u0_uk_K_r13_reg[33]/NET0131 ,
		\u0_uk_K_r13_reg[54]/NET0131 ,
		_w24952_
	);
	LUT2 #(
		.INIT('h1)
	) name19126 (
		_w24951_,
		_w24952_,
		_w24953_
	);
	LUT4 #(
		.INIT('hc693)
	) name19127 (
		decrypt_pad,
		\u0_R13_reg[1]/NET0131 ,
		\u0_uk_K_r13_reg[18]/NET0131 ,
		\u0_uk_K_r13_reg[54]/NET0131 ,
		_w24954_
	);
	LUT4 #(
		.INIT('hc693)
	) name19128 (
		decrypt_pad,
		\u0_R13_reg[3]/NET0131 ,
		\u0_uk_K_r13_reg[10]/NET0131 ,
		\u0_uk_K_r13_reg[46]/NET0131 ,
		_w24955_
	);
	LUT4 #(
		.INIT('hc963)
	) name19129 (
		decrypt_pad,
		\u0_R13_reg[2]/NET0131 ,
		\u0_uk_K_r13_reg[12]/NET0131 ,
		\u0_uk_K_r13_reg[33]/NET0131 ,
		_w24956_
	);
	LUT2 #(
		.INIT('h2)
	) name19130 (
		_w24955_,
		_w24956_,
		_w24957_
	);
	LUT4 #(
		.INIT('h020f)
	) name19131 (
		_w24955_,
		_w24956_,
		_w24952_,
		_w24954_,
		_w24958_
	);
	LUT3 #(
		.INIT('h01)
	) name19132 (
		_w24956_,
		_w24951_,
		_w24954_,
		_w24959_
	);
	LUT3 #(
		.INIT('h54)
	) name19133 (
		_w24953_,
		_w24958_,
		_w24959_,
		_w24960_
	);
	LUT3 #(
		.INIT('h02)
	) name19134 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24961_
	);
	LUT4 #(
		.INIT('hfd31)
	) name19135 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w24962_
	);
	LUT2 #(
		.INIT('h4)
	) name19136 (
		_w24955_,
		_w24952_,
		_w24963_
	);
	LUT4 #(
		.INIT('h500c)
	) name19137 (
		_w24955_,
		_w24956_,
		_w24952_,
		_w24954_,
		_w24964_
	);
	LUT3 #(
		.INIT('h0d)
	) name19138 (
		_w24955_,
		_w24962_,
		_w24964_,
		_w24965_
	);
	LUT3 #(
		.INIT('h8a)
	) name19139 (
		_w24950_,
		_w24960_,
		_w24965_,
		_w24966_
	);
	LUT4 #(
		.INIT('hfade)
	) name19140 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w24967_
	);
	LUT2 #(
		.INIT('h1)
	) name19141 (
		_w24955_,
		_w24967_,
		_w24968_
	);
	LUT3 #(
		.INIT('h60)
	) name19142 (
		_w24951_,
		_w24952_,
		_w24954_,
		_w24969_
	);
	LUT4 #(
		.INIT('h7c3f)
	) name19143 (
		_w24955_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w24970_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name19144 (
		_w24955_,
		_w24956_,
		_w24969_,
		_w24970_,
		_w24971_
	);
	LUT2 #(
		.INIT('h2)
	) name19145 (
		_w24955_,
		_w24954_,
		_w24972_
	);
	LUT3 #(
		.INIT('had)
	) name19146 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24973_
	);
	LUT4 #(
		.INIT('h6ef7)
	) name19147 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w24974_
	);
	LUT4 #(
		.INIT('hfda8)
	) name19148 (
		_w24955_,
		_w24954_,
		_w24973_,
		_w24974_,
		_w24975_
	);
	LUT4 #(
		.INIT('hba00)
	) name19149 (
		_w24950_,
		_w24968_,
		_w24971_,
		_w24975_,
		_w24976_
	);
	LUT3 #(
		.INIT('h65)
	) name19150 (
		\u0_L13_reg[31]/NET0131 ,
		_w24966_,
		_w24976_,
		_w24977_
	);
	LUT4 #(
		.INIT('hc693)
	) name19151 (
		decrypt_pad,
		\u0_R13_reg[32]/NET0131 ,
		\u0_uk_K_r13_reg[14]/NET0131 ,
		\u0_uk_K_r13_reg[52]/P0001 ,
		_w24978_
	);
	LUT4 #(
		.INIT('hc963)
	) name19152 (
		decrypt_pad,
		\u0_R13_reg[31]/NET0131 ,
		\u0_uk_K_r13_reg[42]/NET0131 ,
		\u0_uk_K_r13_reg[8]/NET0131 ,
		_w24979_
	);
	LUT4 #(
		.INIT('hc963)
	) name19153 (
		decrypt_pad,
		\u0_R13_reg[29]/NET0131 ,
		\u0_uk_K_r13_reg[29]/NET0131 ,
		\u0_uk_K_r13_reg[50]/NET0131 ,
		_w24980_
	);
	LUT4 #(
		.INIT('hc963)
	) name19154 (
		decrypt_pad,
		\u0_R13_reg[1]/NET0131 ,
		\u0_uk_K_r13_reg[14]/NET0131 ,
		\u0_uk_K_r13_reg[35]/NET0131 ,
		_w24981_
	);
	LUT4 #(
		.INIT('hc963)
	) name19155 (
		decrypt_pad,
		\u0_R13_reg[30]/NET0131 ,
		\u0_uk_K_r13_reg[30]/NET0131 ,
		\u0_uk_K_r13_reg[51]/NET0131 ,
		_w24982_
	);
	LUT4 #(
		.INIT('hc693)
	) name19156 (
		decrypt_pad,
		\u0_R13_reg[28]/NET0131 ,
		\u0_uk_K_r13_reg[23]/NET0131 ,
		\u0_uk_K_r13_reg[2]/NET0131 ,
		_w24983_
	);
	LUT4 #(
		.INIT('h0040)
	) name19157 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w24984_
	);
	LUT2 #(
		.INIT('h2)
	) name19158 (
		_w24980_,
		_w24981_,
		_w24985_
	);
	LUT4 #(
		.INIT('h44b4)
	) name19159 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w24986_
	);
	LUT4 #(
		.INIT('h00f7)
	) name19160 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24979_,
		_w24987_
	);
	LUT4 #(
		.INIT('h00f6)
	) name19161 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24979_,
		_w24988_
	);
	LUT3 #(
		.INIT('h20)
	) name19162 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24989_
	);
	LUT4 #(
		.INIT('h2000)
	) name19163 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w24990_
	);
	LUT4 #(
		.INIT('h00f2)
	) name19164 (
		_w24979_,
		_w24986_,
		_w24988_,
		_w24990_,
		_w24991_
	);
	LUT2 #(
		.INIT('h2)
	) name19165 (
		_w24978_,
		_w24991_,
		_w24992_
	);
	LUT4 #(
		.INIT('h0008)
	) name19166 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w24993_
	);
	LUT4 #(
		.INIT('hfcf7)
	) name19167 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w24994_
	);
	LUT2 #(
		.INIT('h4)
	) name19168 (
		_w24994_,
		_w24979_,
		_w24995_
	);
	LUT4 #(
		.INIT('h8000)
	) name19169 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w24996_
	);
	LUT3 #(
		.INIT('h04)
	) name19170 (
		_w24982_,
		_w24983_,
		_w24979_,
		_w24997_
	);
	LUT2 #(
		.INIT('h1)
	) name19171 (
		_w24996_,
		_w24997_,
		_w24998_
	);
	LUT3 #(
		.INIT('h0d)
	) name19172 (
		_w24982_,
		_w24983_,
		_w24981_,
		_w24999_
	);
	LUT3 #(
		.INIT('h0b)
	) name19173 (
		_w24980_,
		_w24981_,
		_w24979_,
		_w25000_
	);
	LUT3 #(
		.INIT('h45)
	) name19174 (
		_w24984_,
		_w24999_,
		_w25000_,
		_w25001_
	);
	LUT4 #(
		.INIT('h4555)
	) name19175 (
		_w24978_,
		_w24995_,
		_w24998_,
		_w25001_,
		_w25002_
	);
	LUT4 #(
		.INIT('h0001)
	) name19176 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25003_
	);
	LUT4 #(
		.INIT('hffde)
	) name19177 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25004_
	);
	LUT4 #(
		.INIT('h0200)
	) name19178 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25005_
	);
	LUT4 #(
		.INIT('hf9de)
	) name19179 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25006_
	);
	LUT4 #(
		.INIT('h3f15)
	) name19180 (
		_w24979_,
		_w24997_,
		_w24985_,
		_w25006_,
		_w25007_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name19181 (
		\u0_L13_reg[5]/NET0131 ,
		_w25002_,
		_w24992_,
		_w25007_,
		_w25008_
	);
	LUT4 #(
		.INIT('hc693)
	) name19182 (
		decrypt_pad,
		\u0_R13_reg[17]/NET0131 ,
		\u0_uk_K_r13_reg[27]/NET0131 ,
		\u0_uk_K_r13_reg[6]/NET0131 ,
		_w25009_
	);
	LUT4 #(
		.INIT('hc963)
	) name19183 (
		decrypt_pad,
		\u0_R13_reg[13]/NET0131 ,
		\u0_uk_K_r13_reg[41]/NET0131 ,
		\u0_uk_K_r13_reg[5]/NET0131 ,
		_w25010_
	);
	LUT4 #(
		.INIT('hc693)
	) name19184 (
		decrypt_pad,
		\u0_R13_reg[12]/NET0131 ,
		\u0_uk_K_r13_reg[11]/NET0131 ,
		\u0_uk_K_r13_reg[47]/NET0131 ,
		_w25011_
	);
	LUT4 #(
		.INIT('hc963)
	) name19185 (
		decrypt_pad,
		\u0_R13_reg[14]/NET0131 ,
		\u0_uk_K_r13_reg[10]/NET0131 ,
		\u0_uk_K_r13_reg[6]/NET0131 ,
		_w25012_
	);
	LUT4 #(
		.INIT('h0008)
	) name19186 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25013_
	);
	LUT4 #(
		.INIT('hc963)
	) name19187 (
		decrypt_pad,
		\u0_R13_reg[15]/NET0131 ,
		\u0_uk_K_r13_reg[18]/NET0131 ,
		\u0_uk_K_r13_reg[39]/NET0131 ,
		_w25014_
	);
	LUT3 #(
		.INIT('h80)
	) name19188 (
		_w25010_,
		_w25012_,
		_w25014_,
		_w25015_
	);
	LUT4 #(
		.INIT('h4000)
	) name19189 (
		_w25011_,
		_w25010_,
		_w25012_,
		_w25014_,
		_w25016_
	);
	LUT4 #(
		.INIT('hc963)
	) name19190 (
		decrypt_pad,
		\u0_R13_reg[16]/NET0131 ,
		\u0_uk_K_r13_reg[26]/NET0131 ,
		\u0_uk_K_r13_reg[47]/NET0131 ,
		_w25017_
	);
	LUT3 #(
		.INIT('h01)
	) name19191 (
		_w25016_,
		_w25013_,
		_w25017_,
		_w25018_
	);
	LUT2 #(
		.INIT('h4)
	) name19192 (
		_w25011_,
		_w25009_,
		_w25019_
	);
	LUT4 #(
		.INIT('h8100)
	) name19193 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25014_,
		_w25020_
	);
	LUT4 #(
		.INIT('heffe)
	) name19194 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25021_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name19195 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25022_
	);
	LUT4 #(
		.INIT('h00a8)
	) name19196 (
		_w25021_,
		_w25022_,
		_w25014_,
		_w25020_,
		_w25023_
	);
	LUT2 #(
		.INIT('h8)
	) name19197 (
		_w25018_,
		_w25023_,
		_w25024_
	);
	LUT4 #(
		.INIT('hfe00)
	) name19198 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25025_
	);
	LUT4 #(
		.INIT('h00f6)
	) name19199 (
		_w25011_,
		_w25010_,
		_w25012_,
		_w25014_,
		_w25026_
	);
	LUT2 #(
		.INIT('h4)
	) name19200 (
		_w25025_,
		_w25026_,
		_w25027_
	);
	LUT4 #(
		.INIT('h2000)
	) name19201 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25014_,
		_w25028_
	);
	LUT4 #(
		.INIT('h0040)
	) name19202 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25029_
	);
	LUT2 #(
		.INIT('h1)
	) name19203 (
		_w25028_,
		_w25029_,
		_w25030_
	);
	LUT4 #(
		.INIT('h0400)
	) name19204 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25014_,
		_w25031_
	);
	LUT4 #(
		.INIT('h8000)
	) name19205 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25032_
	);
	LUT3 #(
		.INIT('h02)
	) name19206 (
		_w25017_,
		_w25032_,
		_w25031_,
		_w25033_
	);
	LUT3 #(
		.INIT('h20)
	) name19207 (
		_w25030_,
		_w25027_,
		_w25033_,
		_w25034_
	);
	LUT2 #(
		.INIT('h4)
	) name19208 (
		_w25014_,
		_w25029_,
		_w25035_
	);
	LUT2 #(
		.INIT('h4)
	) name19209 (
		_w25010_,
		_w25014_,
		_w25036_
	);
	LUT3 #(
		.INIT('hde)
	) name19210 (
		_w25011_,
		_w25009_,
		_w25012_,
		_w25037_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name19211 (
		_w25012_,
		_w25028_,
		_w25036_,
		_w25037_,
		_w25038_
	);
	LUT2 #(
		.INIT('h4)
	) name19212 (
		_w25035_,
		_w25038_,
		_w25039_
	);
	LUT4 #(
		.INIT('ha955)
	) name19213 (
		\u0_L13_reg[20]/NET0131 ,
		_w25024_,
		_w25034_,
		_w25039_,
		_w25040_
	);
	LUT4 #(
		.INIT('hc963)
	) name19214 (
		decrypt_pad,
		\u0_R13_reg[24]/NET0131 ,
		\u0_uk_K_r13_reg[21]/NET0131 ,
		\u0_uk_K_r13_reg[42]/NET0131 ,
		_w25041_
	);
	LUT4 #(
		.INIT('hc693)
	) name19215 (
		decrypt_pad,
		\u0_R13_reg[22]/P0001 ,
		\u0_uk_K_r13_reg[31]/NET0131 ,
		\u0_uk_K_r13_reg[37]/NET0131 ,
		_w25042_
	);
	LUT4 #(
		.INIT('hc963)
	) name19216 (
		decrypt_pad,
		\u0_R13_reg[21]/NET0131 ,
		\u0_uk_K_r13_reg[15]/NET0131 ,
		\u0_uk_K_r13_reg[36]/NET0131 ,
		_w25043_
	);
	LUT4 #(
		.INIT('hc963)
	) name19217 (
		decrypt_pad,
		\u0_R13_reg[20]/NET0131 ,
		\u0_uk_K_r13_reg[0]/NET0131 ,
		\u0_uk_K_r13_reg[21]/NET0131 ,
		_w25044_
	);
	LUT4 #(
		.INIT('hc963)
	) name19218 (
		decrypt_pad,
		\u0_R13_reg[25]/NET0131 ,
		\u0_uk_K_r13_reg[16]/NET0131 ,
		\u0_uk_K_r13_reg[37]/NET0131 ,
		_w25045_
	);
	LUT4 #(
		.INIT('hca00)
	) name19219 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25046_
	);
	LUT4 #(
		.INIT('hc693)
	) name19220 (
		decrypt_pad,
		\u0_R13_reg[23]/NET0131 ,
		\u0_uk_K_r13_reg[16]/NET0131 ,
		\u0_uk_K_r13_reg[50]/NET0131 ,
		_w25047_
	);
	LUT4 #(
		.INIT('h00f7)
	) name19221 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25048_
	);
	LUT3 #(
		.INIT('h01)
	) name19222 (
		_w25047_,
		_w25048_,
		_w25046_,
		_w25049_
	);
	LUT4 #(
		.INIT('h0010)
	) name19223 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25050_
	);
	LUT4 #(
		.INIT('h756f)
	) name19224 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25051_
	);
	LUT2 #(
		.INIT('h1)
	) name19225 (
		_w25047_,
		_w25042_,
		_w25052_
	);
	LUT4 #(
		.INIT('h0008)
	) name19226 (
		_w25045_,
		_w25044_,
		_w25047_,
		_w25042_,
		_w25053_
	);
	LUT2 #(
		.INIT('h4)
	) name19227 (
		_w25043_,
		_w25053_,
		_w25054_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name19228 (
		_w25043_,
		_w25047_,
		_w25051_,
		_w25053_,
		_w25055_
	);
	LUT3 #(
		.INIT('h8a)
	) name19229 (
		_w25041_,
		_w25049_,
		_w25055_,
		_w25056_
	);
	LUT3 #(
		.INIT('hd0)
	) name19230 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25057_
	);
	LUT2 #(
		.INIT('h2)
	) name19231 (
		_w25047_,
		_w25042_,
		_w25058_
	);
	LUT4 #(
		.INIT('h0020)
	) name19232 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25059_
	);
	LUT3 #(
		.INIT('h54)
	) name19233 (
		_w25057_,
		_w25058_,
		_w25059_,
		_w25060_
	);
	LUT4 #(
		.INIT('h0208)
	) name19234 (
		_w25043_,
		_w25044_,
		_w25047_,
		_w25042_,
		_w25061_
	);
	LUT3 #(
		.INIT('hc4)
	) name19235 (
		_w25044_,
		_w25047_,
		_w25042_,
		_w25062_
	);
	LUT3 #(
		.INIT('h54)
	) name19236 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25063_
	);
	LUT4 #(
		.INIT('h4000)
	) name19237 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25064_
	);
	LUT4 #(
		.INIT('h0004)
	) name19238 (
		_w25045_,
		_w25044_,
		_w25047_,
		_w25042_,
		_w25065_
	);
	LUT4 #(
		.INIT('h0007)
	) name19239 (
		_w25062_,
		_w25063_,
		_w25064_,
		_w25065_,
		_w25066_
	);
	LUT4 #(
		.INIT('h00ef)
	) name19240 (
		_w25060_,
		_w25061_,
		_w25066_,
		_w25041_,
		_w25067_
	);
	LUT4 #(
		.INIT('hfb00)
	) name19241 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25047_,
		_w25068_
	);
	LUT3 #(
		.INIT('h0e)
	) name19242 (
		_w25058_,
		_w25059_,
		_w25068_,
		_w25069_
	);
	LUT3 #(
		.INIT('h01)
	) name19243 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25070_
	);
	LUT4 #(
		.INIT('h3f1d)
	) name19244 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25071_
	);
	LUT4 #(
		.INIT('h3f15)
	) name19245 (
		_w25062_,
		_w25052_,
		_w25070_,
		_w25071_,
		_w25072_
	);
	LUT2 #(
		.INIT('h4)
	) name19246 (
		_w25069_,
		_w25072_,
		_w25073_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name19247 (
		\u0_L13_reg[11]/NET0131 ,
		_w25067_,
		_w25056_,
		_w25073_,
		_w25074_
	);
	LUT4 #(
		.INIT('h0040)
	) name19248 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25075_
	);
	LUT4 #(
		.INIT('hf0b5)
	) name19249 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25076_
	);
	LUT4 #(
		.INIT('h4041)
	) name19250 (
		_w24955_,
		_w24956_,
		_w24952_,
		_w24954_,
		_w25077_
	);
	LUT4 #(
		.INIT('h1000)
	) name19251 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25078_
	);
	LUT4 #(
		.INIT('h67ff)
	) name19252 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25079_
	);
	LUT4 #(
		.INIT('h0d00)
	) name19253 (
		_w24955_,
		_w25076_,
		_w25077_,
		_w25079_,
		_w25080_
	);
	LUT4 #(
		.INIT('hfe3c)
	) name19254 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25081_
	);
	LUT3 #(
		.INIT('h7b)
	) name19255 (
		_w24951_,
		_w24952_,
		_w24954_,
		_w25082_
	);
	LUT4 #(
		.INIT('hdff7)
	) name19256 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25083_
	);
	LUT4 #(
		.INIT('he400)
	) name19257 (
		_w24955_,
		_w25081_,
		_w25082_,
		_w25083_,
		_w25084_
	);
	LUT3 #(
		.INIT('hf9)
	) name19258 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w25085_
	);
	LUT2 #(
		.INIT('h8)
	) name19259 (
		_w24955_,
		_w24954_,
		_w25086_
	);
	LUT2 #(
		.INIT('h4)
	) name19260 (
		_w25085_,
		_w25086_,
		_w25087_
	);
	LUT4 #(
		.INIT('h00e4)
	) name19261 (
		_w24950_,
		_w25084_,
		_w25080_,
		_w25087_,
		_w25088_
	);
	LUT2 #(
		.INIT('h9)
	) name19262 (
		\u0_L13_reg[17]/NET0131 ,
		_w25088_,
		_w25089_
	);
	LUT4 #(
		.INIT('hddbd)
	) name19263 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25090_
	);
	LUT4 #(
		.INIT('hefe7)
	) name19264 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25091_
	);
	LUT4 #(
		.INIT('h8400)
	) name19265 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25092_
	);
	LUT4 #(
		.INIT('h0d08)
	) name19266 (
		_w25014_,
		_w25091_,
		_w25092_,
		_w25090_,
		_w25093_
	);
	LUT2 #(
		.INIT('h2)
	) name19267 (
		_w25017_,
		_w25093_,
		_w25094_
	);
	LUT3 #(
		.INIT('ha2)
	) name19268 (
		_w25011_,
		_w25009_,
		_w25012_,
		_w25095_
	);
	LUT3 #(
		.INIT('h2a)
	) name19269 (
		_w25021_,
		_w25036_,
		_w25095_,
		_w25096_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name19270 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25014_,
		_w25097_
	);
	LUT4 #(
		.INIT('h00ab)
	) name19271 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25014_,
		_w25098_
	);
	LUT4 #(
		.INIT('he0ee)
	) name19272 (
		_w25012_,
		_w25097_,
		_w25095_,
		_w25098_,
		_w25099_
	);
	LUT3 #(
		.INIT('h15)
	) name19273 (
		_w25017_,
		_w25096_,
		_w25099_,
		_w25100_
	);
	LUT4 #(
		.INIT('h7bfe)
	) name19274 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25101_
	);
	LUT2 #(
		.INIT('h1)
	) name19275 (
		_w25014_,
		_w25101_,
		_w25102_
	);
	LUT3 #(
		.INIT('h23)
	) name19276 (
		_w25012_,
		_w25016_,
		_w25028_,
		_w25103_
	);
	LUT2 #(
		.INIT('h4)
	) name19277 (
		_w25102_,
		_w25103_,
		_w25104_
	);
	LUT4 #(
		.INIT('h5655)
	) name19278 (
		\u0_L13_reg[10]/NET0131 ,
		_w25100_,
		_w25094_,
		_w25104_,
		_w25105_
	);
	LUT4 #(
		.INIT('h3c2f)
	) name19279 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25106_
	);
	LUT4 #(
		.INIT('h0004)
	) name19280 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25107_
	);
	LUT4 #(
		.INIT('h0501)
	) name19281 (
		_w24978_,
		_w24979_,
		_w25107_,
		_w25106_,
		_w25108_
	);
	LUT4 #(
		.INIT('h0020)
	) name19282 (
		_w24982_,
		_w24980_,
		_w24981_,
		_w24979_,
		_w25109_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name19283 (
		_w24978_,
		_w24982_,
		_w24983_,
		_w24980_,
		_w25110_
	);
	LUT4 #(
		.INIT('h0100)
	) name19284 (
		_w24983_,
		_w24980_,
		_w24981_,
		_w24979_,
		_w25111_
	);
	LUT4 #(
		.INIT('hf7df)
	) name19285 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25112_
	);
	LUT4 #(
		.INIT('h1000)
	) name19286 (
		_w25111_,
		_w25109_,
		_w25110_,
		_w25112_,
		_w25113_
	);
	LUT2 #(
		.INIT('h1)
	) name19287 (
		_w25108_,
		_w25113_,
		_w25114_
	);
	LUT4 #(
		.INIT('h1000)
	) name19288 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25115_
	);
	LUT3 #(
		.INIT('h08)
	) name19289 (
		_w24987_,
		_w25004_,
		_w25115_,
		_w25116_
	);
	LUT4 #(
		.INIT('h0100)
	) name19290 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25117_
	);
	LUT3 #(
		.INIT('h02)
	) name19291 (
		_w24979_,
		_w24990_,
		_w25117_,
		_w25118_
	);
	LUT4 #(
		.INIT('h0004)
	) name19292 (
		_w24978_,
		_w24983_,
		_w24980_,
		_w24979_,
		_w25119_
	);
	LUT3 #(
		.INIT('h0e)
	) name19293 (
		_w25116_,
		_w25118_,
		_w25119_,
		_w25120_
	);
	LUT3 #(
		.INIT('h65)
	) name19294 (
		\u0_L13_reg[15]/P0001 ,
		_w25114_,
		_w25120_,
		_w25121_
	);
	LUT4 #(
		.INIT('h4a7f)
	) name19295 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25122_
	);
	LUT4 #(
		.INIT('hf7bb)
	) name19296 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25123_
	);
	LUT4 #(
		.INIT('hfe7d)
	) name19297 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25124_
	);
	LUT4 #(
		.INIT('he400)
	) name19298 (
		_w24979_,
		_w25123_,
		_w25122_,
		_w25124_,
		_w25125_
	);
	LUT2 #(
		.INIT('h2)
	) name19299 (
		_w24978_,
		_w25125_,
		_w25126_
	);
	LUT4 #(
		.INIT('h0004)
	) name19300 (
		_w24983_,
		_w24980_,
		_w24981_,
		_w24979_,
		_w25127_
	);
	LUT3 #(
		.INIT('h01)
	) name19301 (
		_w24993_,
		_w24989_,
		_w25127_,
		_w25128_
	);
	LUT4 #(
		.INIT('h0040)
	) name19302 (
		_w24982_,
		_w24983_,
		_w24981_,
		_w24979_,
		_w25129_
	);
	LUT2 #(
		.INIT('h1)
	) name19303 (
		_w25003_,
		_w25129_,
		_w25130_
	);
	LUT4 #(
		.INIT('hf737)
	) name19304 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25131_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name19305 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24979_,
		_w25132_
	);
	LUT4 #(
		.INIT('hf351)
	) name19306 (
		_w24981_,
		_w24979_,
		_w25131_,
		_w25132_,
		_w25133_
	);
	LUT4 #(
		.INIT('h1555)
	) name19307 (
		_w24978_,
		_w25128_,
		_w25130_,
		_w25133_,
		_w25134_
	);
	LUT4 #(
		.INIT('h0100)
	) name19308 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24979_,
		_w25135_
	);
	LUT3 #(
		.INIT('h07)
	) name19309 (
		_w24980_,
		_w25129_,
		_w25135_,
		_w25136_
	);
	LUT4 #(
		.INIT('h5655)
	) name19310 (
		\u0_L13_reg[21]/NET0131 ,
		_w25134_,
		_w25126_,
		_w25136_,
		_w25137_
	);
	LUT4 #(
		.INIT('hfe0e)
	) name19311 (
		_w24923_,
		_w24924_,
		_w24926_,
		_w24922_,
		_w25138_
	);
	LUT2 #(
		.INIT('h2)
	) name19312 (
		_w24925_,
		_w25138_,
		_w25139_
	);
	LUT4 #(
		.INIT('h2184)
	) name19313 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25140_
	);
	LUT3 #(
		.INIT('h09)
	) name19314 (
		_w24923_,
		_w24924_,
		_w24922_,
		_w25141_
	);
	LUT4 #(
		.INIT('h0200)
	) name19315 (
		_w24923_,
		_w24924_,
		_w24926_,
		_w24922_,
		_w25142_
	);
	LUT4 #(
		.INIT('h0001)
	) name19316 (
		_w24935_,
		_w25142_,
		_w25141_,
		_w25140_,
		_w25143_
	);
	LUT4 #(
		.INIT('hcd00)
	) name19317 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24922_,
		_w25144_
	);
	LUT3 #(
		.INIT('h31)
	) name19318 (
		_w24927_,
		_w25140_,
		_w25144_,
		_w25145_
	);
	LUT3 #(
		.INIT('h8c)
	) name19319 (
		_w24922_,
		_w24935_,
		_w24928_,
		_w25146_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name19320 (
		_w25139_,
		_w25143_,
		_w25145_,
		_w25146_,
		_w25147_
	);
	LUT2 #(
		.INIT('h6)
	) name19321 (
		\u0_L13_reg[12]/NET0131 ,
		_w25147_,
		_w25148_
	);
	LUT4 #(
		.INIT('hc693)
	) name19322 (
		decrypt_pad,
		\u0_R13_reg[20]/NET0131 ,
		\u0_uk_K_r13_reg[30]/NET0131 ,
		\u0_uk_K_r13_reg[9]/NET0131 ,
		_w25149_
	);
	LUT4 #(
		.INIT('hc693)
	) name19323 (
		decrypt_pad,
		\u0_R13_reg[19]/NET0131 ,
		\u0_uk_K_r13_reg[15]/NET0131 ,
		\u0_uk_K_r13_reg[49]/NET0131 ,
		_w25150_
	);
	LUT4 #(
		.INIT('hc693)
	) name19324 (
		decrypt_pad,
		\u0_R13_reg[21]/NET0131 ,
		\u0_uk_K_r13_reg[0]/NET0131 ,
		\u0_uk_K_r13_reg[38]/NET0131 ,
		_w25151_
	);
	LUT4 #(
		.INIT('hc963)
	) name19325 (
		decrypt_pad,
		\u0_R13_reg[16]/NET0131 ,
		\u0_uk_K_r13_reg[22]/NET0131 ,
		\u0_uk_K_r13_reg[43]/NET0131 ,
		_w25152_
	);
	LUT4 #(
		.INIT('hc693)
	) name19326 (
		decrypt_pad,
		\u0_R13_reg[18]/NET0131 ,
		\u0_uk_K_r13_reg[28]/NET0131 ,
		\u0_uk_K_r13_reg[7]/NET0131 ,
		_w25153_
	);
	LUT4 #(
		.INIT('hc693)
	) name19327 (
		decrypt_pad,
		\u0_R13_reg[17]/NET0131 ,
		\u0_uk_K_r13_reg[38]/NET0131 ,
		\u0_uk_K_r13_reg[44]/NET0131 ,
		_w25154_
	);
	LUT3 #(
		.INIT('h80)
	) name19328 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25155_
	);
	LUT4 #(
		.INIT('h6c6a)
	) name19329 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25156_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name19330 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25157_
	);
	LUT4 #(
		.INIT('h08a0)
	) name19331 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25158_
	);
	LUT4 #(
		.INIT('h0e02)
	) name19332 (
		_w25157_,
		_w25150_,
		_w25158_,
		_w25156_,
		_w25159_
	);
	LUT2 #(
		.INIT('h2)
	) name19333 (
		_w25149_,
		_w25159_,
		_w25160_
	);
	LUT4 #(
		.INIT('hf6ef)
	) name19334 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25161_
	);
	LUT2 #(
		.INIT('h2)
	) name19335 (
		_w25150_,
		_w25161_,
		_w25162_
	);
	LUT2 #(
		.INIT('h4)
	) name19336 (
		_w25151_,
		_w25150_,
		_w25163_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name19337 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25164_
	);
	LUT3 #(
		.INIT('hd0)
	) name19338 (
		_w25154_,
		_w25151_,
		_w25150_,
		_w25165_
	);
	LUT4 #(
		.INIT('h0f01)
	) name19339 (
		_w25154_,
		_w25152_,
		_w25153_,
		_w25150_,
		_w25166_
	);
	LUT4 #(
		.INIT('he0ee)
	) name19340 (
		_w25163_,
		_w25164_,
		_w25165_,
		_w25166_,
		_w25167_
	);
	LUT4 #(
		.INIT('h0040)
	) name19341 (
		_w25154_,
		_w25152_,
		_w25153_,
		_w25150_,
		_w25168_
	);
	LUT4 #(
		.INIT('h0080)
	) name19342 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25169_
	);
	LUT2 #(
		.INIT('h1)
	) name19343 (
		_w25168_,
		_w25169_,
		_w25170_
	);
	LUT4 #(
		.INIT('h0e00)
	) name19344 (
		_w25149_,
		_w25167_,
		_w25162_,
		_w25170_,
		_w25171_
	);
	LUT3 #(
		.INIT('h65)
	) name19345 (
		\u0_L13_reg[25]/NET0131 ,
		_w25160_,
		_w25171_,
		_w25172_
	);
	LUT3 #(
		.INIT('h10)
	) name19346 (
		_w25011_,
		_w25010_,
		_w25012_,
		_w25173_
	);
	LUT4 #(
		.INIT('hf8fc)
	) name19347 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25174_
	);
	LUT4 #(
		.INIT('h0092)
	) name19348 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25175_
	);
	LUT4 #(
		.INIT('h0504)
	) name19349 (
		_w25014_,
		_w25017_,
		_w25175_,
		_w25174_,
		_w25176_
	);
	LUT3 #(
		.INIT('h02)
	) name19350 (
		_w25014_,
		_w25013_,
		_w25029_,
		_w25177_
	);
	LUT2 #(
		.INIT('h1)
	) name19351 (
		_w25176_,
		_w25177_,
		_w25178_
	);
	LUT4 #(
		.INIT('h2010)
	) name19352 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25179_
	);
	LUT4 #(
		.INIT('h0100)
	) name19353 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25014_,
		_w25180_
	);
	LUT3 #(
		.INIT('h02)
	) name19354 (
		_w25017_,
		_w25179_,
		_w25180_,
		_w25181_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name19355 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25014_,
		_w25182_
	);
	LUT4 #(
		.INIT('h7773)
	) name19356 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25183_
	);
	LUT3 #(
		.INIT('h0d)
	) name19357 (
		_w25011_,
		_w25012_,
		_w25014_,
		_w25184_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name19358 (
		_w25012_,
		_w25182_,
		_w25183_,
		_w25184_,
		_w25185_
	);
	LUT4 #(
		.INIT('h00fd)
	) name19359 (
		_w25011_,
		_w25010_,
		_w25012_,
		_w25017_,
		_w25186_
	);
	LUT3 #(
		.INIT('hb0)
	) name19360 (
		_w25019_,
		_w25015_,
		_w25186_,
		_w25187_
	);
	LUT4 #(
		.INIT('h153f)
	) name19361 (
		_w25030_,
		_w25181_,
		_w25185_,
		_w25187_,
		_w25188_
	);
	LUT3 #(
		.INIT('h56)
	) name19362 (
		\u0_L13_reg[26]/NET0131 ,
		_w25178_,
		_w25188_,
		_w25189_
	);
	LUT4 #(
		.INIT('hc963)
	) name19363 (
		decrypt_pad,
		\u0_R13_reg[8]/NET0131 ,
		\u0_uk_K_r13_reg[25]/P0001 ,
		\u0_uk_K_r13_reg[46]/NET0131 ,
		_w25190_
	);
	LUT4 #(
		.INIT('hc963)
	) name19364 (
		decrypt_pad,
		\u0_R13_reg[7]/NET0131 ,
		\u0_uk_K_r13_reg[34]/NET0131 ,
		\u0_uk_K_r13_reg[55]/NET0131 ,
		_w25191_
	);
	LUT4 #(
		.INIT('hc963)
	) name19365 (
		decrypt_pad,
		\u0_R13_reg[6]/NET0131 ,
		\u0_uk_K_r13_reg[40]/NET0131 ,
		\u0_uk_K_r13_reg[4]/NET0131 ,
		_w25192_
	);
	LUT4 #(
		.INIT('hc693)
	) name19366 (
		decrypt_pad,
		\u0_R13_reg[5]/NET0131 ,
		\u0_uk_K_r13_reg[13]/NET0131 ,
		\u0_uk_K_r13_reg[17]/NET0131 ,
		_w25193_
	);
	LUT4 #(
		.INIT('hc963)
	) name19367 (
		decrypt_pad,
		\u0_R13_reg[4]/NET0131 ,
		\u0_uk_K_r13_reg[13]/NET0131 ,
		\u0_uk_K_r13_reg[34]/NET0131 ,
		_w25194_
	);
	LUT4 #(
		.INIT('hc693)
	) name19368 (
		decrypt_pad,
		\u0_R13_reg[9]/NET0131 ,
		\u0_uk_K_r13_reg[26]/NET0131 ,
		\u0_uk_K_r13_reg[5]/NET0131 ,
		_w25195_
	);
	LUT4 #(
		.INIT('h797d)
	) name19369 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25196_
	);
	LUT2 #(
		.INIT('h2)
	) name19370 (
		_w25191_,
		_w25196_,
		_w25197_
	);
	LUT4 #(
		.INIT('h00df)
	) name19371 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25191_,
		_w25198_
	);
	LUT2 #(
		.INIT('h2)
	) name19372 (
		_w25194_,
		_w25192_,
		_w25199_
	);
	LUT2 #(
		.INIT('h4)
	) name19373 (
		_w25198_,
		_w25199_,
		_w25200_
	);
	LUT4 #(
		.INIT('hbfba)
	) name19374 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25201_
	);
	LUT4 #(
		.INIT('h1000)
	) name19375 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25202_
	);
	LUT3 #(
		.INIT('h0e)
	) name19376 (
		_w25191_,
		_w25201_,
		_w25202_,
		_w25203_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name19377 (
		_w25190_,
		_w25200_,
		_w25197_,
		_w25203_,
		_w25204_
	);
	LUT4 #(
		.INIT('h6765)
	) name19378 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25205_
	);
	LUT4 #(
		.INIT('h2900)
	) name19379 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25206_
	);
	LUT4 #(
		.INIT('h5404)
	) name19380 (
		_w25206_,
		_w25205_,
		_w25191_,
		_w25201_,
		_w25207_
	);
	LUT4 #(
		.INIT('h0800)
	) name19381 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25208_
	);
	LUT4 #(
		.INIT('he6ff)
	) name19382 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25209_
	);
	LUT2 #(
		.INIT('h1)
	) name19383 (
		_w25191_,
		_w25209_,
		_w25210_
	);
	LUT3 #(
		.INIT('h0e)
	) name19384 (
		_w25190_,
		_w25207_,
		_w25210_,
		_w25211_
	);
	LUT3 #(
		.INIT('h65)
	) name19385 (
		\u0_L13_reg[28]/NET0131 ,
		_w25204_,
		_w25211_,
		_w25212_
	);
	LUT4 #(
		.INIT('h3cfe)
	) name19386 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25213_
	);
	LUT2 #(
		.INIT('h1)
	) name19387 (
		_w25047_,
		_w25213_,
		_w25214_
	);
	LUT4 #(
		.INIT('hd7f5)
	) name19388 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25215_
	);
	LUT2 #(
		.INIT('h2)
	) name19389 (
		_w25047_,
		_w25215_,
		_w25216_
	);
	LUT4 #(
		.INIT('h0104)
	) name19390 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25217_
	);
	LUT3 #(
		.INIT('h01)
	) name19391 (
		_w25064_,
		_w25065_,
		_w25217_,
		_w25218_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name19392 (
		_w25041_,
		_w25216_,
		_w25214_,
		_w25218_,
		_w25219_
	);
	LUT4 #(
		.INIT('h6d6e)
	) name19393 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25220_
	);
	LUT4 #(
		.INIT('hdf35)
	) name19394 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25221_
	);
	LUT4 #(
		.INIT('h0400)
	) name19395 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25222_
	);
	LUT4 #(
		.INIT('h00d8)
	) name19396 (
		_w25047_,
		_w25220_,
		_w25221_,
		_w25222_,
		_w25223_
	);
	LUT4 #(
		.INIT('h0080)
	) name19397 (
		_w25043_,
		_w25045_,
		_w25047_,
		_w25042_,
		_w25224_
	);
	LUT2 #(
		.INIT('h1)
	) name19398 (
		_w25050_,
		_w25224_,
		_w25225_
	);
	LUT3 #(
		.INIT('he0)
	) name19399 (
		_w25041_,
		_w25223_,
		_w25225_,
		_w25226_
	);
	LUT3 #(
		.INIT('h9a)
	) name19400 (
		\u0_L13_reg[29]/NET0131 ,
		_w25219_,
		_w25226_,
		_w25227_
	);
	LUT4 #(
		.INIT('h65ef)
	) name19401 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25228_
	);
	LUT2 #(
		.INIT('h1)
	) name19402 (
		_w25191_,
		_w25228_,
		_w25229_
	);
	LUT4 #(
		.INIT('h001c)
	) name19403 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25230_
	);
	LUT4 #(
		.INIT('h2000)
	) name19404 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25231_
	);
	LUT2 #(
		.INIT('h2)
	) name19405 (
		_w25195_,
		_w25192_,
		_w25232_
	);
	LUT4 #(
		.INIT('h0004)
	) name19406 (
		_w25193_,
		_w25195_,
		_w25192_,
		_w25191_,
		_w25233_
	);
	LUT4 #(
		.INIT('h4000)
	) name19407 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25234_
	);
	LUT4 #(
		.INIT('h0007)
	) name19408 (
		_w25191_,
		_w25231_,
		_w25233_,
		_w25234_,
		_w25235_
	);
	LUT4 #(
		.INIT('h5455)
	) name19409 (
		_w25190_,
		_w25229_,
		_w25230_,
		_w25235_,
		_w25236_
	);
	LUT4 #(
		.INIT('hda7c)
	) name19410 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25237_
	);
	LUT4 #(
		.INIT('h4010)
	) name19411 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25238_
	);
	LUT4 #(
		.INIT('h0031)
	) name19412 (
		_w25190_,
		_w25191_,
		_w25237_,
		_w25238_,
		_w25239_
	);
	LUT4 #(
		.INIT('h7731)
	) name19413 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25240_
	);
	LUT4 #(
		.INIT('h0100)
	) name19414 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25241_
	);
	LUT4 #(
		.INIT('hf700)
	) name19415 (
		_w25194_,
		_w25193_,
		_w25192_,
		_w25191_,
		_w25242_
	);
	LUT4 #(
		.INIT('h3100)
	) name19416 (
		_w25190_,
		_w25241_,
		_w25240_,
		_w25242_,
		_w25243_
	);
	LUT2 #(
		.INIT('h1)
	) name19417 (
		_w25239_,
		_w25243_,
		_w25244_
	);
	LUT3 #(
		.INIT('h56)
	) name19418 (
		\u0_L13_reg[2]/NET0131 ,
		_w25236_,
		_w25244_,
		_w25245_
	);
	LUT4 #(
		.INIT('h0004)
	) name19419 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25246_
	);
	LUT4 #(
		.INIT('he56b)
	) name19420 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25247_
	);
	LUT4 #(
		.INIT('h4002)
	) name19421 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25248_
	);
	LUT4 #(
		.INIT('h3fdd)
	) name19422 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25249_
	);
	LUT4 #(
		.INIT('h3edc)
	) name19423 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25250_
	);
	LUT4 #(
		.INIT('h3120)
	) name19424 (
		_w25150_,
		_w25248_,
		_w25250_,
		_w25247_,
		_w25251_
	);
	LUT2 #(
		.INIT('h1)
	) name19425 (
		_w25149_,
		_w25251_,
		_w25252_
	);
	LUT3 #(
		.INIT('h20)
	) name19426 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25253_
	);
	LUT4 #(
		.INIT('hb796)
	) name19427 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25150_,
		_w25254_
	);
	LUT2 #(
		.INIT('h1)
	) name19428 (
		_w25153_,
		_w25254_,
		_w25255_
	);
	LUT4 #(
		.INIT('hf800)
	) name19429 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25150_,
		_w25256_
	);
	LUT2 #(
		.INIT('h8)
	) name19430 (
		_w25249_,
		_w25256_,
		_w25257_
	);
	LUT2 #(
		.INIT('h2)
	) name19431 (
		_w25153_,
		_w25150_,
		_w25258_
	);
	LUT4 #(
		.INIT('h0400)
	) name19432 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25259_
	);
	LUT3 #(
		.INIT('h07)
	) name19433 (
		_w25155_,
		_w25258_,
		_w25259_,
		_w25260_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name19434 (
		_w25149_,
		_w25257_,
		_w25255_,
		_w25260_,
		_w25261_
	);
	LUT4 #(
		.INIT('h0108)
	) name19435 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25262_
	);
	LUT4 #(
		.INIT('h1000)
	) name19436 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25263_
	);
	LUT4 #(
		.INIT('hedff)
	) name19437 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25264_
	);
	LUT3 #(
		.INIT('h8d)
	) name19438 (
		_w25150_,
		_w25262_,
		_w25264_,
		_w25265_
	);
	LUT4 #(
		.INIT('h5556)
	) name19439 (
		\u0_L13_reg[14]/NET0131 ,
		_w25261_,
		_w25252_,
		_w25265_,
		_w25266_
	);
	LUT4 #(
		.INIT('hffd0)
	) name19440 (
		_w25043_,
		_w25045_,
		_w25047_,
		_w25042_,
		_w25267_
	);
	LUT2 #(
		.INIT('h1)
	) name19441 (
		_w25044_,
		_w25267_,
		_w25268_
	);
	LUT4 #(
		.INIT('h8802)
	) name19442 (
		_w25043_,
		_w25045_,
		_w25047_,
		_w25042_,
		_w25269_
	);
	LUT4 #(
		.INIT('h0080)
	) name19443 (
		_w25045_,
		_w25044_,
		_w25047_,
		_w25042_,
		_w25270_
	);
	LUT3 #(
		.INIT('h02)
	) name19444 (
		_w25041_,
		_w25270_,
		_w25269_,
		_w25271_
	);
	LUT4 #(
		.INIT('hdf00)
	) name19445 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25047_,
		_w25272_
	);
	LUT4 #(
		.INIT('hbff3)
	) name19446 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25273_
	);
	LUT4 #(
		.INIT('h00fd)
	) name19447 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25047_,
		_w25274_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name19448 (
		_w25222_,
		_w25272_,
		_w25273_,
		_w25274_,
		_w25275_
	);
	LUT3 #(
		.INIT('h01)
	) name19449 (
		_w25041_,
		_w25050_,
		_w25053_,
		_w25276_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name19450 (
		_w25268_,
		_w25271_,
		_w25275_,
		_w25276_,
		_w25277_
	);
	LUT4 #(
		.INIT('h006f)
	) name19451 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25047_,
		_w25278_
	);
	LUT4 #(
		.INIT('hd600)
	) name19452 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25047_,
		_w25279_
	);
	LUT4 #(
		.INIT('h0001)
	) name19453 (
		_w25045_,
		_w25044_,
		_w25047_,
		_w25042_,
		_w25280_
	);
	LUT4 #(
		.INIT('h00fd)
	) name19454 (
		_w25042_,
		_w25279_,
		_w25278_,
		_w25280_,
		_w25281_
	);
	LUT3 #(
		.INIT('h65)
	) name19455 (
		\u0_L13_reg[4]/NET0131 ,
		_w25277_,
		_w25281_,
		_w25282_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name19456 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25283_
	);
	LUT4 #(
		.INIT('h2100)
	) name19457 (
		_w25011_,
		_w25009_,
		_w25012_,
		_w25014_,
		_w25284_
	);
	LUT2 #(
		.INIT('h4)
	) name19458 (
		_w25283_,
		_w25284_,
		_w25285_
	);
	LUT3 #(
		.INIT('hd8)
	) name19459 (
		_w25009_,
		_w25010_,
		_w25012_,
		_w25286_
	);
	LUT2 #(
		.INIT('h2)
	) name19460 (
		_w25011_,
		_w25014_,
		_w25287_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name19461 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25288_
	);
	LUT3 #(
		.INIT('hb0)
	) name19462 (
		_w25286_,
		_w25287_,
		_w25288_,
		_w25289_
	);
	LUT3 #(
		.INIT('h45)
	) name19463 (
		_w25017_,
		_w25285_,
		_w25289_,
		_w25290_
	);
	LUT4 #(
		.INIT('h2000)
	) name19464 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25291_
	);
	LUT3 #(
		.INIT('h31)
	) name19465 (
		_w25011_,
		_w25009_,
		_w25012_,
		_w25292_
	);
	LUT4 #(
		.INIT('h0031)
	) name19466 (
		_w25036_,
		_w25173_,
		_w25292_,
		_w25291_,
		_w25293_
	);
	LUT4 #(
		.INIT('h6bff)
	) name19467 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25294_
	);
	LUT2 #(
		.INIT('h2)
	) name19468 (
		_w25014_,
		_w25294_,
		_w25295_
	);
	LUT4 #(
		.INIT('h2100)
	) name19469 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25296_
	);
	LUT4 #(
		.INIT('hbf2f)
	) name19470 (
		_w25011_,
		_w25009_,
		_w25010_,
		_w25012_,
		_w25297_
	);
	LUT4 #(
		.INIT('h5054)
	) name19471 (
		_w25014_,
		_w25017_,
		_w25296_,
		_w25297_,
		_w25298_
	);
	LUT4 #(
		.INIT('h0301)
	) name19472 (
		_w25017_,
		_w25295_,
		_w25298_,
		_w25293_,
		_w25299_
	);
	LUT3 #(
		.INIT('h65)
	) name19473 (
		\u0_L13_reg[1]/NET0131 ,
		_w25290_,
		_w25299_,
		_w25300_
	);
	LUT4 #(
		.INIT('hf77f)
	) name19474 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25301_
	);
	LUT3 #(
		.INIT('h01)
	) name19475 (
		_w25193_,
		_w25195_,
		_w25192_,
		_w25302_
	);
	LUT4 #(
		.INIT('hebf9)
	) name19476 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25303_
	);
	LUT4 #(
		.INIT('h0313)
	) name19477 (
		_w25190_,
		_w25191_,
		_w25301_,
		_w25303_,
		_w25304_
	);
	LUT4 #(
		.INIT('hded6)
	) name19478 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25305_
	);
	LUT2 #(
		.INIT('h2)
	) name19479 (
		_w25191_,
		_w25305_,
		_w25306_
	);
	LUT2 #(
		.INIT('h8)
	) name19480 (
		_w25192_,
		_w25191_,
		_w25307_
	);
	LUT3 #(
		.INIT('ha2)
	) name19481 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25308_
	);
	LUT2 #(
		.INIT('h8)
	) name19482 (
		_w25307_,
		_w25308_,
		_w25309_
	);
	LUT3 #(
		.INIT('h54)
	) name19483 (
		_w25194_,
		_w25193_,
		_w25191_,
		_w25310_
	);
	LUT3 #(
		.INIT('h15)
	) name19484 (
		_w25190_,
		_w25232_,
		_w25310_,
		_w25311_
	);
	LUT3 #(
		.INIT('h10)
	) name19485 (
		_w25306_,
		_w25309_,
		_w25311_,
		_w25312_
	);
	LUT3 #(
		.INIT('h10)
	) name19486 (
		_w25193_,
		_w25195_,
		_w25192_,
		_w25313_
	);
	LUT4 #(
		.INIT('hbf00)
	) name19487 (
		_w25194_,
		_w25195_,
		_w25192_,
		_w25191_,
		_w25314_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name19488 (
		_w25198_,
		_w25302_,
		_w25313_,
		_w25314_,
		_w25315_
	);
	LUT4 #(
		.INIT('h0004)
	) name19489 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25316_
	);
	LUT4 #(
		.INIT('h0002)
	) name19490 (
		_w25190_,
		_w25233_,
		_w25234_,
		_w25316_,
		_w25317_
	);
	LUT3 #(
		.INIT('h20)
	) name19491 (
		_w25301_,
		_w25315_,
		_w25317_,
		_w25318_
	);
	LUT4 #(
		.INIT('h999a)
	) name19492 (
		\u0_L13_reg[13]/NET0131 ,
		_w25304_,
		_w25312_,
		_w25318_,
		_w25319_
	);
	LUT3 #(
		.INIT('h0d)
	) name19493 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25320_
	);
	LUT4 #(
		.INIT('hf070)
	) name19494 (
		_w25043_,
		_w25044_,
		_w25047_,
		_w25042_,
		_w25321_
	);
	LUT2 #(
		.INIT('h4)
	) name19495 (
		_w25320_,
		_w25321_,
		_w25322_
	);
	LUT4 #(
		.INIT('h0009)
	) name19496 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25047_,
		_w25323_
	);
	LUT4 #(
		.INIT('h8000)
	) name19497 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25324_
	);
	LUT3 #(
		.INIT('h01)
	) name19498 (
		_w25041_,
		_w25323_,
		_w25324_,
		_w25325_
	);
	LUT4 #(
		.INIT('hfb5b)
	) name19499 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25326_
	);
	LUT2 #(
		.INIT('h2)
	) name19500 (
		_w25047_,
		_w25326_,
		_w25327_
	);
	LUT4 #(
		.INIT('hfd00)
	) name19501 (
		_w25043_,
		_w25045_,
		_w25042_,
		_w25041_,
		_w25328_
	);
	LUT4 #(
		.INIT('h0800)
	) name19502 (
		_w25043_,
		_w25045_,
		_w25044_,
		_w25042_,
		_w25329_
	);
	LUT3 #(
		.INIT('h04)
	) name19503 (
		_w25043_,
		_w25044_,
		_w25047_,
		_w25330_
	);
	LUT4 #(
		.INIT('h0100)
	) name19504 (
		_w25217_,
		_w25329_,
		_w25330_,
		_w25328_,
		_w25331_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name19505 (
		_w25322_,
		_w25325_,
		_w25327_,
		_w25331_,
		_w25332_
	);
	LUT2 #(
		.INIT('h1)
	) name19506 (
		_w25069_,
		_w25054_,
		_w25333_
	);
	LUT3 #(
		.INIT('h65)
	) name19507 (
		\u0_L13_reg[19]/NET0131 ,
		_w25332_,
		_w25333_,
		_w25334_
	);
	LUT4 #(
		.INIT('hfcd3)
	) name19508 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25335_
	);
	LUT2 #(
		.INIT('h1)
	) name19509 (
		_w24955_,
		_w25335_,
		_w25336_
	);
	LUT3 #(
		.INIT('h8a)
	) name19510 (
		_w24955_,
		_w24956_,
		_w24952_,
		_w25337_
	);
	LUT2 #(
		.INIT('h8)
	) name19511 (
		_w24969_,
		_w25337_,
		_w25338_
	);
	LUT3 #(
		.INIT('h07)
	) name19512 (
		_w24961_,
		_w24972_,
		_w25075_,
		_w25339_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name19513 (
		_w24950_,
		_w25336_,
		_w25338_,
		_w25339_,
		_w25340_
	);
	LUT4 #(
		.INIT('h0080)
	) name19514 (
		_w24955_,
		_w24956_,
		_w24951_,
		_w24952_,
		_w25341_
	);
	LUT3 #(
		.INIT('h7e)
	) name19515 (
		_w24956_,
		_w24951_,
		_w24954_,
		_w25342_
	);
	LUT2 #(
		.INIT('h4)
	) name19516 (
		_w25341_,
		_w25342_,
		_w25343_
	);
	LUT4 #(
		.INIT('h0200)
	) name19517 (
		_w24955_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25344_
	);
	LUT3 #(
		.INIT('h07)
	) name19518 (
		_w24956_,
		_w24951_,
		_w24954_,
		_w25345_
	);
	LUT3 #(
		.INIT('h31)
	) name19519 (
		_w24963_,
		_w25344_,
		_w25345_,
		_w25346_
	);
	LUT3 #(
		.INIT('he3)
	) name19520 (
		_w24951_,
		_w24952_,
		_w24954_,
		_w25347_
	);
	LUT4 #(
		.INIT('h6ffb)
	) name19521 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25348_
	);
	LUT4 #(
		.INIT('hfda8)
	) name19522 (
		_w24955_,
		_w24956_,
		_w25347_,
		_w25348_,
		_w25349_
	);
	LUT4 #(
		.INIT('hea00)
	) name19523 (
		_w24950_,
		_w25343_,
		_w25346_,
		_w25349_,
		_w25350_
	);
	LUT3 #(
		.INIT('h9a)
	) name19524 (
		\u0_L13_reg[23]/NET0131 ,
		_w25340_,
		_w25350_,
		_w25351_
	);
	LUT4 #(
		.INIT('h3fef)
	) name19525 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25352_
	);
	LUT4 #(
		.INIT('hce3e)
	) name19526 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25353_
	);
	LUT4 #(
		.INIT('hdaf7)
	) name19527 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25354_
	);
	LUT4 #(
		.INIT('he400)
	) name19528 (
		_w24979_,
		_w25353_,
		_w25352_,
		_w25354_,
		_w25355_
	);
	LUT2 #(
		.INIT('h2)
	) name19529 (
		_w24978_,
		_w25355_,
		_w25356_
	);
	LUT4 #(
		.INIT('hdf00)
	) name19530 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24979_,
		_w25357_
	);
	LUT3 #(
		.INIT('h4b)
	) name19531 (
		_w24982_,
		_w24980_,
		_w24981_,
		_w25358_
	);
	LUT2 #(
		.INIT('h8)
	) name19532 (
		_w25357_,
		_w25358_,
		_w25359_
	);
	LUT4 #(
		.INIT('h0080)
	) name19533 (
		_w24982_,
		_w24983_,
		_w24981_,
		_w24979_,
		_w25360_
	);
	LUT3 #(
		.INIT('h01)
	) name19534 (
		_w25005_,
		_w25127_,
		_w25360_,
		_w25361_
	);
	LUT3 #(
		.INIT('h45)
	) name19535 (
		_w24978_,
		_w25359_,
		_w25361_,
		_w25362_
	);
	LUT4 #(
		.INIT('hfbdf)
	) name19536 (
		_w24982_,
		_w24983_,
		_w24980_,
		_w24981_,
		_w25363_
	);
	LUT2 #(
		.INIT('h1)
	) name19537 (
		_w24979_,
		_w25363_,
		_w25364_
	);
	LUT4 #(
		.INIT('h0200)
	) name19538 (
		_w24982_,
		_w24980_,
		_w24981_,
		_w24979_,
		_w25365_
	);
	LUT3 #(
		.INIT('h07)
	) name19539 (
		_w24997_,
		_w24985_,
		_w25365_,
		_w25366_
	);
	LUT2 #(
		.INIT('h4)
	) name19540 (
		_w25364_,
		_w25366_,
		_w25367_
	);
	LUT4 #(
		.INIT('h5655)
	) name19541 (
		\u0_L13_reg[27]/NET0131 ,
		_w25362_,
		_w25356_,
		_w25367_,
		_w25368_
	);
	LUT3 #(
		.INIT('h40)
	) name19542 (
		_w24923_,
		_w24925_,
		_w24926_,
		_w25369_
	);
	LUT4 #(
		.INIT('ha7e6)
	) name19543 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25370_
	);
	LUT2 #(
		.INIT('h2)
	) name19544 (
		_w24922_,
		_w25370_,
		_w25371_
	);
	LUT4 #(
		.INIT('h8a11)
	) name19545 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25372_
	);
	LUT4 #(
		.INIT('h54a8)
	) name19546 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25373_
	);
	LUT3 #(
		.INIT('h01)
	) name19547 (
		_w24922_,
		_w25373_,
		_w25372_,
		_w25374_
	);
	LUT4 #(
		.INIT('h4000)
	) name19548 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25375_
	);
	LUT2 #(
		.INIT('h2)
	) name19549 (
		_w24935_,
		_w25375_,
		_w25376_
	);
	LUT3 #(
		.INIT('h10)
	) name19550 (
		_w25374_,
		_w25371_,
		_w25376_,
		_w25377_
	);
	LUT3 #(
		.INIT('h10)
	) name19551 (
		_w24923_,
		_w24925_,
		_w24926_,
		_w25378_
	);
	LUT4 #(
		.INIT('hd8ff)
	) name19552 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25379_
	);
	LUT4 #(
		.INIT('h8040)
	) name19553 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25380_
	);
	LUT4 #(
		.INIT('h0301)
	) name19554 (
		_w24922_,
		_w24935_,
		_w25380_,
		_w25379_,
		_w25381_
	);
	LUT4 #(
		.INIT('h0420)
	) name19555 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25382_
	);
	LUT3 #(
		.INIT('h0d)
	) name19556 (
		_w25141_,
		_w25378_,
		_w25382_,
		_w25383_
	);
	LUT2 #(
		.INIT('h8)
	) name19557 (
		_w25381_,
		_w25383_,
		_w25384_
	);
	LUT3 #(
		.INIT('h08)
	) name19558 (
		_w24924_,
		_w24925_,
		_w24926_,
		_w25385_
	);
	LUT4 #(
		.INIT('hf73f)
	) name19559 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25386_
	);
	LUT3 #(
		.INIT('h72)
	) name19560 (
		_w24922_,
		_w24928_,
		_w25386_,
		_w25387_
	);
	LUT4 #(
		.INIT('ha955)
	) name19561 (
		\u0_L13_reg[32]/NET0131 ,
		_w25377_,
		_w25384_,
		_w25387_,
		_w25388_
	);
	LUT4 #(
		.INIT('hc963)
	) name19562 (
		decrypt_pad,
		\u0_R13_reg[8]/NET0131 ,
		\u0_uk_K_r13_reg[39]/NET0131 ,
		\u0_uk_K_r13_reg[3]/NET0131 ,
		_w25389_
	);
	LUT4 #(
		.INIT('hc963)
	) name19563 (
		decrypt_pad,
		\u0_R13_reg[9]/NET0131 ,
		\u0_uk_K_r13_reg[11]/NET0131 ,
		\u0_uk_K_r13_reg[32]/NET0131 ,
		_w25390_
	);
	LUT4 #(
		.INIT('hc963)
	) name19564 (
		decrypt_pad,
		\u0_R13_reg[10]/NET0131 ,
		\u0_uk_K_r13_reg[19]/NET0131 ,
		\u0_uk_K_r13_reg[40]/NET0131 ,
		_w25391_
	);
	LUT3 #(
		.INIT('h51)
	) name19565 (
		_w25389_,
		_w25390_,
		_w25391_,
		_w25392_
	);
	LUT4 #(
		.INIT('hc963)
	) name19566 (
		decrypt_pad,
		\u0_R13_reg[11]/NET0131 ,
		\u0_uk_K_r13_reg[20]/NET0131 ,
		\u0_uk_K_r13_reg[41]/NET0131 ,
		_w25393_
	);
	LUT4 #(
		.INIT('hc693)
	) name19567 (
		decrypt_pad,
		\u0_R13_reg[13]/NET0131 ,
		\u0_uk_K_r13_reg[12]/NET0131 ,
		\u0_uk_K_r13_reg[48]/NET0131 ,
		_w25394_
	);
	LUT3 #(
		.INIT('h09)
	) name19568 (
		_w25394_,
		_w25390_,
		_w25393_,
		_w25395_
	);
	LUT4 #(
		.INIT('h1000)
	) name19569 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25396_
	);
	LUT4 #(
		.INIT('hc693)
	) name19570 (
		decrypt_pad,
		\u0_R13_reg[12]/NET0131 ,
		\u0_uk_K_r13_reg[24]/NET0131 ,
		\u0_uk_K_r13_reg[3]/NET0131 ,
		_w25397_
	);
	LUT4 #(
		.INIT('h4500)
	) name19571 (
		_w25396_,
		_w25392_,
		_w25395_,
		_w25397_,
		_w25398_
	);
	LUT2 #(
		.INIT('h6)
	) name19572 (
		_w25394_,
		_w25389_,
		_w25399_
	);
	LUT2 #(
		.INIT('h8)
	) name19573 (
		_w25394_,
		_w25393_,
		_w25400_
	);
	LUT4 #(
		.INIT('h0103)
	) name19574 (
		_w25394_,
		_w25390_,
		_w25391_,
		_w25393_,
		_w25401_
	);
	LUT2 #(
		.INIT('h8)
	) name19575 (
		_w25399_,
		_w25401_,
		_w25402_
	);
	LUT4 #(
		.INIT('h4000)
	) name19576 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25403_
	);
	LUT4 #(
		.INIT('h0400)
	) name19577 (
		_w25389_,
		_w25390_,
		_w25391_,
		_w25393_,
		_w25404_
	);
	LUT3 #(
		.INIT('h01)
	) name19578 (
		_w25397_,
		_w25404_,
		_w25403_,
		_w25405_
	);
	LUT4 #(
		.INIT('h9990)
	) name19579 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25406_
	);
	LUT4 #(
		.INIT('h0990)
	) name19580 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25407_
	);
	LUT2 #(
		.INIT('h2)
	) name19581 (
		_w25394_,
		_w25389_,
		_w25408_
	);
	LUT4 #(
		.INIT('h2000)
	) name19582 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25409_
	);
	LUT3 #(
		.INIT('h23)
	) name19583 (
		_w25393_,
		_w25407_,
		_w25409_,
		_w25410_
	);
	LUT4 #(
		.INIT('h4555)
	) name19584 (
		_w25398_,
		_w25402_,
		_w25405_,
		_w25410_,
		_w25411_
	);
	LUT4 #(
		.INIT('h95b5)
	) name19585 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25412_
	);
	LUT4 #(
		.INIT('h0001)
	) name19586 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25413_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name19587 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25414_
	);
	LUT4 #(
		.INIT('h08aa)
	) name19588 (
		_w25393_,
		_w25397_,
		_w25412_,
		_w25414_,
		_w25415_
	);
	LUT3 #(
		.INIT('h56)
	) name19589 (
		\u0_L13_reg[6]/NET0131 ,
		_w25411_,
		_w25415_,
		_w25416_
	);
	LUT2 #(
		.INIT('h2)
	) name19590 (
		_w24922_,
		_w24935_,
		_w25417_
	);
	LUT4 #(
		.INIT('h4080)
	) name19591 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25418_
	);
	LUT4 #(
		.INIT('h957a)
	) name19592 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25419_
	);
	LUT2 #(
		.INIT('h2)
	) name19593 (
		_w25417_,
		_w25419_,
		_w25420_
	);
	LUT4 #(
		.INIT('h2a04)
	) name19594 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25421_
	);
	LUT2 #(
		.INIT('h4)
	) name19595 (
		_w24922_,
		_w24935_,
		_w25422_
	);
	LUT2 #(
		.INIT('h9)
	) name19596 (
		_w24922_,
		_w24935_,
		_w25423_
	);
	LUT3 #(
		.INIT('h10)
	) name19597 (
		_w25418_,
		_w25421_,
		_w25423_,
		_w25424_
	);
	LUT4 #(
		.INIT('h8b74)
	) name19598 (
		_w24923_,
		_w24924_,
		_w24925_,
		_w24926_,
		_w25425_
	);
	LUT4 #(
		.INIT('h1000)
	) name19599 (
		_w25369_,
		_w25385_,
		_w25422_,
		_w25425_,
		_w25426_
	);
	LUT4 #(
		.INIT('h00ab)
	) name19600 (
		_w24938_,
		_w25420_,
		_w25424_,
		_w25426_,
		_w25427_
	);
	LUT2 #(
		.INIT('h6)
	) name19601 (
		\u0_L13_reg[7]/NET0131 ,
		_w25427_,
		_w25428_
	);
	LUT3 #(
		.INIT('h04)
	) name19602 (
		_w25152_,
		_w25151_,
		_w25153_,
		_w25429_
	);
	LUT4 #(
		.INIT('h9f8f)
	) name19603 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25430_
	);
	LUT4 #(
		.INIT('h7f7b)
	) name19604 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25431_
	);
	LUT4 #(
		.INIT('hf6dd)
	) name19605 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25432_
	);
	LUT4 #(
		.INIT('hd800)
	) name19606 (
		_w25150_,
		_w25431_,
		_w25430_,
		_w25432_,
		_w25433_
	);
	LUT2 #(
		.INIT('h1)
	) name19607 (
		_w25149_,
		_w25433_,
		_w25434_
	);
	LUT3 #(
		.INIT('hbe)
	) name19608 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25435_
	);
	LUT4 #(
		.INIT('hbf00)
	) name19609 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25436_
	);
	LUT3 #(
		.INIT('h02)
	) name19610 (
		_w25150_,
		_w25436_,
		_w25435_,
		_w25437_
	);
	LUT3 #(
		.INIT('h02)
	) name19611 (
		_w25152_,
		_w25153_,
		_w25150_,
		_w25438_
	);
	LUT2 #(
		.INIT('h2)
	) name19612 (
		_w25264_,
		_w25438_,
		_w25439_
	);
	LUT4 #(
		.INIT('hf5df)
	) name19613 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25440_
	);
	LUT4 #(
		.INIT('he4ee)
	) name19614 (
		_w25150_,
		_w25259_,
		_w25263_,
		_w25440_,
		_w25441_
	);
	LUT4 #(
		.INIT('h0075)
	) name19615 (
		_w25149_,
		_w25437_,
		_w25439_,
		_w25441_,
		_w25442_
	);
	LUT3 #(
		.INIT('h65)
	) name19616 (
		\u0_L13_reg[8]/NET0131 ,
		_w25434_,
		_w25442_,
		_w25443_
	);
	LUT3 #(
		.INIT('hed)
	) name19617 (
		_w25394_,
		_w25389_,
		_w25391_,
		_w25444_
	);
	LUT3 #(
		.INIT('h20)
	) name19618 (
		_w25389_,
		_w25390_,
		_w25391_,
		_w25445_
	);
	LUT3 #(
		.INIT('h10)
	) name19619 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25446_
	);
	LUT4 #(
		.INIT('he2cd)
	) name19620 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25447_
	);
	LUT2 #(
		.INIT('h1)
	) name19621 (
		_w25397_,
		_w25447_,
		_w25448_
	);
	LUT4 #(
		.INIT('h0020)
	) name19622 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25449_
	);
	LUT4 #(
		.INIT('h0004)
	) name19623 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25450_
	);
	LUT3 #(
		.INIT('h02)
	) name19624 (
		_w25393_,
		_w25449_,
		_w25450_,
		_w25451_
	);
	LUT4 #(
		.INIT('h0026)
	) name19625 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25452_
	);
	LUT3 #(
		.INIT('h01)
	) name19626 (
		_w25397_,
		_w25406_,
		_w25452_,
		_w25453_
	);
	LUT4 #(
		.INIT('h8000)
	) name19627 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25454_
	);
	LUT2 #(
		.INIT('h1)
	) name19628 (
		_w25393_,
		_w25454_,
		_w25455_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name19629 (
		_w25448_,
		_w25451_,
		_w25453_,
		_w25455_,
		_w25456_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name19630 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25457_
	);
	LUT3 #(
		.INIT('he0)
	) name19631 (
		_w25390_,
		_w25391_,
		_w25393_,
		_w25458_
	);
	LUT4 #(
		.INIT('h0302)
	) name19632 (
		_w25393_,
		_w25408_,
		_w25458_,
		_w25457_,
		_w25459_
	);
	LUT4 #(
		.INIT('h1dff)
	) name19633 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25460_
	);
	LUT4 #(
		.INIT('h3f15)
	) name19634 (
		_w25393_,
		_w25399_,
		_w25401_,
		_w25460_,
		_w25461_
	);
	LUT3 #(
		.INIT('h8a)
	) name19635 (
		_w25397_,
		_w25459_,
		_w25461_,
		_w25462_
	);
	LUT3 #(
		.INIT('h56)
	) name19636 (
		\u0_L13_reg[24]/NET0131 ,
		_w25456_,
		_w25462_,
		_w25463_
	);
	LUT4 #(
		.INIT('h6979)
	) name19637 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25393_,
		_w25464_
	);
	LUT2 #(
		.INIT('h1)
	) name19638 (
		_w25391_,
		_w25464_,
		_w25465_
	);
	LUT4 #(
		.INIT('h0014)
	) name19639 (
		_w25394_,
		_w25389_,
		_w25391_,
		_w25393_,
		_w25466_
	);
	LUT3 #(
		.INIT('h02)
	) name19640 (
		_w25397_,
		_w25409_,
		_w25466_,
		_w25467_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name19641 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25468_
	);
	LUT2 #(
		.INIT('h1)
	) name19642 (
		_w25393_,
		_w25468_,
		_w25469_
	);
	LUT4 #(
		.INIT('h6800)
	) name19643 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25393_,
		_w25470_
	);
	LUT3 #(
		.INIT('h01)
	) name19644 (
		_w25397_,
		_w25413_,
		_w25470_,
		_w25471_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name19645 (
		_w25465_,
		_w25467_,
		_w25469_,
		_w25471_,
		_w25472_
	);
	LUT4 #(
		.INIT('h0020)
	) name19646 (
		_w25389_,
		_w25390_,
		_w25391_,
		_w25393_,
		_w25473_
	);
	LUT4 #(
		.INIT('hbeff)
	) name19647 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25474_
	);
	LUT3 #(
		.INIT('h31)
	) name19648 (
		_w25393_,
		_w25473_,
		_w25474_,
		_w25475_
	);
	LUT3 #(
		.INIT('h65)
	) name19649 (
		\u0_L13_reg[16]/NET0131 ,
		_w25472_,
		_w25475_,
		_w25476_
	);
	LUT4 #(
		.INIT('h0209)
	) name19650 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25477_
	);
	LUT4 #(
		.INIT('h73af)
	) name19651 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25478_
	);
	LUT3 #(
		.INIT('h07)
	) name19652 (
		_w25389_,
		_w25391_,
		_w25393_,
		_w25479_
	);
	LUT3 #(
		.INIT('hac)
	) name19653 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25480_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name19654 (
		_w25393_,
		_w25478_,
		_w25479_,
		_w25480_,
		_w25481_
	);
	LUT3 #(
		.INIT('h45)
	) name19655 (
		_w25397_,
		_w25477_,
		_w25481_,
		_w25482_
	);
	LUT3 #(
		.INIT('h08)
	) name19656 (
		_w25393_,
		_w25444_,
		_w25450_,
		_w25483_
	);
	LUT3 #(
		.INIT('h8a)
	) name19657 (
		_w25397_,
		_w25446_,
		_w25479_,
		_w25484_
	);
	LUT3 #(
		.INIT('h0e)
	) name19658 (
		_w25394_,
		_w25393_,
		_w25397_,
		_w25485_
	);
	LUT4 #(
		.INIT('h7000)
	) name19659 (
		_w25394_,
		_w25389_,
		_w25390_,
		_w25391_,
		_w25486_
	);
	LUT4 #(
		.INIT('h7077)
	) name19660 (
		_w25400_,
		_w25445_,
		_w25485_,
		_w25486_,
		_w25487_
	);
	LUT3 #(
		.INIT('hb0)
	) name19661 (
		_w25483_,
		_w25484_,
		_w25487_,
		_w25488_
	);
	LUT3 #(
		.INIT('h9a)
	) name19662 (
		\u0_L13_reg[30]/NET0131 ,
		_w25482_,
		_w25488_,
		_w25489_
	);
	LUT4 #(
		.INIT('hdc33)
	) name19663 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25490_
	);
	LUT3 #(
		.INIT('h25)
	) name19664 (
		_w24951_,
		_w24952_,
		_w24954_,
		_w25491_
	);
	LUT4 #(
		.INIT('hbf7d)
	) name19665 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25492_
	);
	LUT4 #(
		.INIT('h8d00)
	) name19666 (
		_w24955_,
		_w25490_,
		_w25491_,
		_w25492_,
		_w25493_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name19667 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25494_
	);
	LUT2 #(
		.INIT('h1)
	) name19668 (
		_w24955_,
		_w25494_,
		_w25495_
	);
	LUT4 #(
		.INIT('h8228)
	) name19669 (
		_w24956_,
		_w24951_,
		_w24952_,
		_w24954_,
		_w25496_
	);
	LUT4 #(
		.INIT('h0013)
	) name19670 (
		_w24957_,
		_w25078_,
		_w25491_,
		_w25496_,
		_w25497_
	);
	LUT4 #(
		.INIT('h0e04)
	) name19671 (
		_w24950_,
		_w25493_,
		_w25495_,
		_w25497_,
		_w25498_
	);
	LUT2 #(
		.INIT('h9)
	) name19672 (
		\u0_L13_reg[9]/NET0131 ,
		_w25498_,
		_w25499_
	);
	LUT4 #(
		.INIT('hfd3d)
	) name19673 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25500_
	);
	LUT4 #(
		.INIT('hfb7f)
	) name19674 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25501_
	);
	LUT4 #(
		.INIT('hb100)
	) name19675 (
		_w25150_,
		_w25253_,
		_w25500_,
		_w25501_,
		_w25502_
	);
	LUT2 #(
		.INIT('h2)
	) name19676 (
		_w25149_,
		_w25502_,
		_w25503_
	);
	LUT4 #(
		.INIT('h4009)
	) name19677 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25504_
	);
	LUT4 #(
		.INIT('hfda8)
	) name19678 (
		_w25150_,
		_w25246_,
		_w25263_,
		_w25504_,
		_w25505_
	);
	LUT4 #(
		.INIT('hf7c7)
	) name19679 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25506_
	);
	LUT2 #(
		.INIT('h2)
	) name19680 (
		_w25150_,
		_w25506_,
		_w25507_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name19681 (
		_w25154_,
		_w25152_,
		_w25151_,
		_w25153_,
		_w25508_
	);
	LUT3 #(
		.INIT('hb0)
	) name19682 (
		_w25154_,
		_w25153_,
		_w25150_,
		_w25509_
	);
	LUT3 #(
		.INIT('h01)
	) name19683 (
		_w25429_,
		_w25509_,
		_w25508_,
		_w25510_
	);
	LUT4 #(
		.INIT('h2223)
	) name19684 (
		_w25149_,
		_w25505_,
		_w25507_,
		_w25510_,
		_w25511_
	);
	LUT3 #(
		.INIT('h65)
	) name19685 (
		\u0_L13_reg[3]/NET0131 ,
		_w25503_,
		_w25511_,
		_w25512_
	);
	LUT4 #(
		.INIT('h1c00)
	) name19686 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25191_,
		_w25513_
	);
	LUT3 #(
		.INIT('h07)
	) name19687 (
		_w25195_,
		_w25192_,
		_w25191_,
		_w25514_
	);
	LUT4 #(
		.INIT('h0222)
	) name19688 (
		_w25190_,
		_w25241_,
		_w25308_,
		_w25514_,
		_w25515_
	);
	LUT4 #(
		.INIT('h5554)
	) name19689 (
		_w25190_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25516_
	);
	LUT2 #(
		.INIT('h4)
	) name19690 (
		_w25208_,
		_w25516_,
		_w25517_
	);
	LUT4 #(
		.INIT('h0141)
	) name19691 (
		_w25194_,
		_w25193_,
		_w25192_,
		_w25191_,
		_w25518_
	);
	LUT4 #(
		.INIT('h8000)
	) name19692 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25191_,
		_w25519_
	);
	LUT3 #(
		.INIT('h01)
	) name19693 (
		_w25231_,
		_w25519_,
		_w25518_,
		_w25520_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name19694 (
		_w25513_,
		_w25515_,
		_w25517_,
		_w25520_,
		_w25521_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name19695 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25192_,
		_w25522_
	);
	LUT4 #(
		.INIT('h0040)
	) name19696 (
		_w25194_,
		_w25193_,
		_w25195_,
		_w25191_,
		_w25523_
	);
	LUT3 #(
		.INIT('h0d)
	) name19697 (
		_w25191_,
		_w25522_,
		_w25523_,
		_w25524_
	);
	LUT3 #(
		.INIT('h65)
	) name19698 (
		\u0_L13_reg[18]/NET0131 ,
		_w25521_,
		_w25524_,
		_w25525_
	);
	LUT4 #(
		.INIT('hc693)
	) name19699 (
		decrypt_pad,
		\u0_R12_reg[3]/NET0131 ,
		\u0_uk_K_r12_reg[24]/NET0131 ,
		\u0_uk_K_r12_reg[32]/NET0131 ,
		_w25526_
	);
	LUT4 #(
		.INIT('hc693)
	) name19700 (
		decrypt_pad,
		\u0_R12_reg[32]/NET0131 ,
		\u0_uk_K_r12_reg[11]/NET0131 ,
		\u0_uk_K_r12_reg[19]/NET0131 ,
		_w25527_
	);
	LUT4 #(
		.INIT('hc963)
	) name19701 (
		decrypt_pad,
		\u0_R12_reg[5]/NET0131 ,
		\u0_uk_K_r12_reg[13]/NET0131 ,
		\u0_uk_K_r12_reg[5]/NET0131 ,
		_w25528_
	);
	LUT4 #(
		.INIT('hc693)
	) name19702 (
		decrypt_pad,
		\u0_R12_reg[2]/NET0131 ,
		\u0_uk_K_r12_reg[47]/NET0131 ,
		\u0_uk_K_r12_reg[55]/NET0131 ,
		_w25529_
	);
	LUT4 #(
		.INIT('hc693)
	) name19703 (
		decrypt_pad,
		\u0_R12_reg[1]/NET0131 ,
		\u0_uk_K_r12_reg[32]/NET0131 ,
		\u0_uk_K_r12_reg[40]/NET0131 ,
		_w25530_
	);
	LUT4 #(
		.INIT('hd7df)
	) name19704 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25531_
	);
	LUT2 #(
		.INIT('h2)
	) name19705 (
		_w25526_,
		_w25531_,
		_w25532_
	);
	LUT3 #(
		.INIT('h40)
	) name19706 (
		_w25527_,
		_w25529_,
		_w25526_,
		_w25533_
	);
	LUT4 #(
		.INIT('h4000)
	) name19707 (
		_w25527_,
		_w25529_,
		_w25526_,
		_w25528_,
		_w25534_
	);
	LUT4 #(
		.INIT('hbfee)
	) name19708 (
		_w25527_,
		_w25529_,
		_w25526_,
		_w25528_,
		_w25535_
	);
	LUT2 #(
		.INIT('h4)
	) name19709 (
		_w25535_,
		_w25530_,
		_w25536_
	);
	LUT2 #(
		.INIT('h9)
	) name19710 (
		_w25527_,
		_w25529_,
		_w25537_
	);
	LUT4 #(
		.INIT('h1103)
	) name19711 (
		_w25529_,
		_w25526_,
		_w25528_,
		_w25530_,
		_w25538_
	);
	LUT4 #(
		.INIT('h0020)
	) name19712 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25539_
	);
	LUT3 #(
		.INIT('h07)
	) name19713 (
		_w25537_,
		_w25538_,
		_w25539_,
		_w25540_
	);
	LUT4 #(
		.INIT('hc963)
	) name19714 (
		decrypt_pad,
		\u0_R12_reg[4]/NET0131 ,
		\u0_uk_K_r12_reg[10]/P0001 ,
		\u0_uk_K_r12_reg[34]/NET0131 ,
		_w25541_
	);
	LUT4 #(
		.INIT('h00ef)
	) name19715 (
		_w25536_,
		_w25532_,
		_w25540_,
		_w25541_,
		_w25542_
	);
	LUT2 #(
		.INIT('h1)
	) name19716 (
		_w25528_,
		_w25530_,
		_w25543_
	);
	LUT4 #(
		.INIT('hccfa)
	) name19717 (
		_w25529_,
		_w25526_,
		_w25528_,
		_w25530_,
		_w25544_
	);
	LUT2 #(
		.INIT('h2)
	) name19718 (
		_w25527_,
		_w25544_,
		_w25545_
	);
	LUT4 #(
		.INIT('hfb0b)
	) name19719 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25546_
	);
	LUT2 #(
		.INIT('h4)
	) name19720 (
		_w25529_,
		_w25526_,
		_w25547_
	);
	LUT3 #(
		.INIT('hb0)
	) name19721 (
		_w25529_,
		_w25526_,
		_w25530_,
		_w25548_
	);
	LUT3 #(
		.INIT('h54)
	) name19722 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25549_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name19723 (
		_w25526_,
		_w25546_,
		_w25548_,
		_w25549_,
		_w25550_
	);
	LUT3 #(
		.INIT('h8a)
	) name19724 (
		_w25541_,
		_w25545_,
		_w25550_,
		_w25551_
	);
	LUT4 #(
		.INIT('h7cbf)
	) name19725 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25552_
	);
	LUT2 #(
		.INIT('h1)
	) name19726 (
		_w25526_,
		_w25552_,
		_w25553_
	);
	LUT4 #(
		.INIT('h0020)
	) name19727 (
		_w25527_,
		_w25529_,
		_w25526_,
		_w25530_,
		_w25554_
	);
	LUT3 #(
		.INIT('h07)
	) name19728 (
		_w25533_,
		_w25543_,
		_w25554_,
		_w25555_
	);
	LUT2 #(
		.INIT('h4)
	) name19729 (
		_w25553_,
		_w25555_,
		_w25556_
	);
	LUT4 #(
		.INIT('h5655)
	) name19730 (
		\u0_L12_reg[31]/NET0131 ,
		_w25542_,
		_w25551_,
		_w25556_,
		_w25557_
	);
	LUT4 #(
		.INIT('hc693)
	) name19731 (
		decrypt_pad,
		\u0_R12_reg[24]/NET0131 ,
		\u0_uk_K_r12_reg[1]/NET0131 ,
		\u0_uk_K_r12_reg[7]/P0001 ,
		_w25558_
	);
	LUT4 #(
		.INIT('hc693)
	) name19732 (
		decrypt_pad,
		\u0_R12_reg[23]/NET0131 ,
		\u0_uk_K_r12_reg[30]/NET0131 ,
		\u0_uk_K_r12_reg[36]/NET0131 ,
		_w25559_
	);
	LUT4 #(
		.INIT('hc963)
	) name19733 (
		decrypt_pad,
		\u0_R12_reg[21]/NET0131 ,
		\u0_uk_K_r12_reg[1]/NET0131 ,
		\u0_uk_K_r12_reg[50]/NET0131 ,
		_w25560_
	);
	LUT4 #(
		.INIT('hc963)
	) name19734 (
		decrypt_pad,
		\u0_R12_reg[22]/NET0131 ,
		\u0_uk_K_r12_reg[23]/NET0131 ,
		\u0_uk_K_r12_reg[45]/NET0131 ,
		_w25561_
	);
	LUT4 #(
		.INIT('hc693)
	) name19735 (
		decrypt_pad,
		\u0_R12_reg[20]/NET0131 ,
		\u0_uk_K_r12_reg[35]/NET0131 ,
		\u0_uk_K_r12_reg[45]/NET0131 ,
		_w25562_
	);
	LUT4 #(
		.INIT('hc963)
	) name19736 (
		decrypt_pad,
		\u0_R12_reg[25]/NET0131 ,
		\u0_uk_K_r12_reg[2]/NET0131 ,
		\u0_uk_K_r12_reg[51]/NET0131 ,
		_w25563_
	);
	LUT4 #(
		.INIT('h1000)
	) name19737 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25564_
	);
	LUT4 #(
		.INIT('he93b)
	) name19738 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25565_
	);
	LUT3 #(
		.INIT('h54)
	) name19739 (
		_w25560_,
		_w25561_,
		_w25563_,
		_w25566_
	);
	LUT4 #(
		.INIT('h888a)
	) name19740 (
		_w25559_,
		_w25560_,
		_w25561_,
		_w25563_,
		_w25567_
	);
	LUT4 #(
		.INIT('hfc5c)
	) name19741 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25568_
	);
	LUT4 #(
		.INIT('he4ee)
	) name19742 (
		_w25559_,
		_w25565_,
		_w25566_,
		_w25568_,
		_w25569_
	);
	LUT2 #(
		.INIT('h2)
	) name19743 (
		_w25558_,
		_w25569_,
		_w25570_
	);
	LUT4 #(
		.INIT('hc9db)
	) name19744 (
		_w25559_,
		_w25560_,
		_w25562_,
		_w25563_,
		_w25571_
	);
	LUT3 #(
		.INIT('hc4)
	) name19745 (
		_w25560_,
		_w25562_,
		_w25563_,
		_w25572_
	);
	LUT4 #(
		.INIT('ha020)
	) name19746 (
		_w25559_,
		_w25560_,
		_w25562_,
		_w25563_,
		_w25573_
	);
	LUT4 #(
		.INIT('h1505)
	) name19747 (
		_w25559_,
		_w25560_,
		_w25562_,
		_w25563_,
		_w25574_
	);
	LUT4 #(
		.INIT('hddd8)
	) name19748 (
		_w25561_,
		_w25571_,
		_w25574_,
		_w25573_,
		_w25575_
	);
	LUT4 #(
		.INIT('h0200)
	) name19749 (
		_w25559_,
		_w25560_,
		_w25562_,
		_w25563_,
		_w25576_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name19750 (
		_w25559_,
		_w25560_,
		_w25562_,
		_w25563_,
		_w25577_
	);
	LUT2 #(
		.INIT('h1)
	) name19751 (
		_w25561_,
		_w25577_,
		_w25578_
	);
	LUT2 #(
		.INIT('h1)
	) name19752 (
		_w25562_,
		_w25563_,
		_w25579_
	);
	LUT2 #(
		.INIT('h1)
	) name19753 (
		_w25559_,
		_w25561_,
		_w25580_
	);
	LUT3 #(
		.INIT('h01)
	) name19754 (
		_w25559_,
		_w25560_,
		_w25561_,
		_w25581_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name19755 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25582_
	);
	LUT4 #(
		.INIT('h3f15)
	) name19756 (
		_w25559_,
		_w25579_,
		_w25581_,
		_w25582_,
		_w25583_
	);
	LUT4 #(
		.INIT('h0e00)
	) name19757 (
		_w25558_,
		_w25575_,
		_w25578_,
		_w25583_,
		_w25584_
	);
	LUT3 #(
		.INIT('h9a)
	) name19758 (
		\u0_L12_reg[11]/NET0131 ,
		_w25570_,
		_w25584_,
		_w25585_
	);
	LUT4 #(
		.INIT('hc693)
	) name19759 (
		decrypt_pad,
		\u0_R12_reg[27]/NET0131 ,
		\u0_uk_K_r12_reg[21]/NET0131 ,
		\u0_uk_K_r12_reg[31]/NET0131 ,
		_w25586_
	);
	LUT4 #(
		.INIT('hc693)
	) name19760 (
		decrypt_pad,
		\u0_R12_reg[25]/NET0131 ,
		\u0_uk_K_r12_reg[31]/NET0131 ,
		\u0_uk_K_r12_reg[9]/NET0131 ,
		_w25587_
	);
	LUT4 #(
		.INIT('hc693)
	) name19761 (
		decrypt_pad,
		\u0_R12_reg[24]/NET0131 ,
		\u0_uk_K_r12_reg[23]/NET0131 ,
		\u0_uk_K_r12_reg[29]/NET0131 ,
		_w25588_
	);
	LUT4 #(
		.INIT('hc693)
	) name19762 (
		decrypt_pad,
		\u0_R12_reg[29]/NET0131 ,
		\u0_uk_K_r12_reg[0]/NET0131 ,
		\u0_uk_K_r12_reg[37]/NET0131 ,
		_w25589_
	);
	LUT4 #(
		.INIT('hc693)
	) name19763 (
		decrypt_pad,
		\u0_R12_reg[26]/NET0131 ,
		\u0_uk_K_r12_reg[43]/NET0131 ,
		\u0_uk_K_r12_reg[49]/NET0131 ,
		_w25590_
	);
	LUT4 #(
		.INIT('h0004)
	) name19764 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25591_
	);
	LUT4 #(
		.INIT('h757b)
	) name19765 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25592_
	);
	LUT2 #(
		.INIT('h1)
	) name19766 (
		_w25586_,
		_w25592_,
		_w25593_
	);
	LUT4 #(
		.INIT('hb5b9)
	) name19767 (
		_w25588_,
		_w25589_,
		_w25587_,
		_w25586_,
		_w25594_
	);
	LUT4 #(
		.INIT('h8000)
	) name19768 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25595_
	);
	LUT4 #(
		.INIT('hc963)
	) name19769 (
		decrypt_pad,
		\u0_R12_reg[28]/NET0131 ,
		\u0_uk_K_r12_reg[14]/NET0131 ,
		\u0_uk_K_r12_reg[8]/NET0131 ,
		_w25596_
	);
	LUT4 #(
		.INIT('h0032)
	) name19770 (
		_w25590_,
		_w25595_,
		_w25594_,
		_w25596_,
		_w25597_
	);
	LUT4 #(
		.INIT('h2088)
	) name19771 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25598_
	);
	LUT3 #(
		.INIT('h08)
	) name19772 (
		_w25588_,
		_w25589_,
		_w25587_,
		_w25599_
	);
	LUT4 #(
		.INIT('h0020)
	) name19773 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25600_
	);
	LUT3 #(
		.INIT('h40)
	) name19774 (
		_w25588_,
		_w25589_,
		_w25587_,
		_w25601_
	);
	LUT4 #(
		.INIT('hddd8)
	) name19775 (
		_w25586_,
		_w25598_,
		_w25600_,
		_w25601_,
		_w25602_
	);
	LUT4 #(
		.INIT('h0001)
	) name19776 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25603_
	);
	LUT4 #(
		.INIT('h0040)
	) name19777 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25604_
	);
	LUT3 #(
		.INIT('h02)
	) name19778 (
		_w25596_,
		_w25603_,
		_w25604_,
		_w25605_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name19779 (
		_w25593_,
		_w25597_,
		_w25602_,
		_w25605_,
		_w25606_
	);
	LUT4 #(
		.INIT('h007f)
	) name19780 (
		_w25588_,
		_w25590_,
		_w25587_,
		_w25586_,
		_w25607_
	);
	LUT4 #(
		.INIT('h006f)
	) name19781 (
		_w25588_,
		_w25590_,
		_w25587_,
		_w25586_,
		_w25608_
	);
	LUT4 #(
		.INIT('h0400)
	) name19782 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25609_
	);
	LUT4 #(
		.INIT('hfbbf)
	) name19783 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25610_
	);
	LUT4 #(
		.INIT('h000b)
	) name19784 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25611_
	);
	LUT4 #(
		.INIT('h3313)
	) name19785 (
		_w25586_,
		_w25608_,
		_w25610_,
		_w25611_,
		_w25612_
	);
	LUT3 #(
		.INIT('h56)
	) name19786 (
		\u0_L12_reg[22]/NET0131 ,
		_w25606_,
		_w25612_,
		_w25613_
	);
	LUT4 #(
		.INIT('hfe5a)
	) name19787 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25614_
	);
	LUT2 #(
		.INIT('h9)
	) name19788 (
		_w25528_,
		_w25530_,
		_w25615_
	);
	LUT3 #(
		.INIT('h82)
	) name19789 (
		_w25527_,
		_w25528_,
		_w25530_,
		_w25616_
	);
	LUT4 #(
		.INIT('hf7bf)
	) name19790 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25617_
	);
	LUT4 #(
		.INIT('h4e00)
	) name19791 (
		_w25526_,
		_w25614_,
		_w25616_,
		_w25617_,
		_w25618_
	);
	LUT4 #(
		.INIT('haa9b)
	) name19792 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25619_
	);
	LUT4 #(
		.INIT('h0809)
	) name19793 (
		_w25527_,
		_w25529_,
		_w25526_,
		_w25530_,
		_w25620_
	);
	LUT4 #(
		.INIT('h0200)
	) name19794 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25621_
	);
	LUT4 #(
		.INIT('h3dff)
	) name19795 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25622_
	);
	LUT4 #(
		.INIT('h0d00)
	) name19796 (
		_w25526_,
		_w25619_,
		_w25620_,
		_w25622_,
		_w25623_
	);
	LUT3 #(
		.INIT('h10)
	) name19797 (
		_w25527_,
		_w25528_,
		_w25530_,
		_w25624_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name19798 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25625_
	);
	LUT4 #(
		.INIT('h2333)
	) name19799 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25626_
	);
	LUT3 #(
		.INIT('h02)
	) name19800 (
		_w25526_,
		_w25626_,
		_w25625_,
		_w25627_
	);
	LUT4 #(
		.INIT('h0d08)
	) name19801 (
		_w25541_,
		_w25623_,
		_w25627_,
		_w25618_,
		_w25628_
	);
	LUT2 #(
		.INIT('h9)
	) name19802 (
		\u0_L12_reg[17]/NET0131 ,
		_w25628_,
		_w25629_
	);
	LUT4 #(
		.INIT('hc693)
	) name19803 (
		decrypt_pad,
		\u0_R12_reg[13]/NET0131 ,
		\u0_uk_K_r12_reg[19]/NET0131 ,
		\u0_uk_K_r12_reg[27]/NET0131 ,
		_w25630_
	);
	LUT4 #(
		.INIT('hc963)
	) name19804 (
		decrypt_pad,
		\u0_R12_reg[17]/NET0131 ,
		\u0_uk_K_r12_reg[17]/NET0131 ,
		\u0_uk_K_r12_reg[41]/NET0131 ,
		_w25631_
	);
	LUT4 #(
		.INIT('hc693)
	) name19805 (
		decrypt_pad,
		\u0_R12_reg[14]/NET0131 ,
		\u0_uk_K_r12_reg[20]/NET0131 ,
		\u0_uk_K_r12_reg[53]/NET0131 ,
		_w25632_
	);
	LUT4 #(
		.INIT('hc693)
	) name19806 (
		decrypt_pad,
		\u0_R12_reg[12]/NET0131 ,
		\u0_uk_K_r12_reg[25]/NET0131 ,
		\u0_uk_K_r12_reg[33]/NET0131 ,
		_w25633_
	);
	LUT4 #(
		.INIT('h8000)
	) name19807 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25634_
	);
	LUT4 #(
		.INIT('hc963)
	) name19808 (
		decrypt_pad,
		\u0_R12_reg[16]/NET0131 ,
		\u0_uk_K_r12_reg[12]/NET0131 ,
		\u0_uk_K_r12_reg[4]/NET0131 ,
		_w25635_
	);
	LUT4 #(
		.INIT('hc963)
	) name19809 (
		decrypt_pad,
		\u0_R12_reg[15]/NET0131 ,
		\u0_uk_K_r12_reg[4]/NET0131 ,
		\u0_uk_K_r12_reg[53]/NET0131 ,
		_w25636_
	);
	LUT2 #(
		.INIT('h2)
	) name19810 (
		_w25630_,
		_w25633_,
		_w25637_
	);
	LUT4 #(
		.INIT('h0104)
	) name19811 (
		_w25632_,
		_w25630_,
		_w25636_,
		_w25633_,
		_w25638_
	);
	LUT2 #(
		.INIT('h4)
	) name19812 (
		_w25633_,
		_w25631_,
		_w25639_
	);
	LUT4 #(
		.INIT('h0400)
	) name19813 (
		_w25630_,
		_w25636_,
		_w25633_,
		_w25631_,
		_w25640_
	);
	LUT4 #(
		.INIT('h0100)
	) name19814 (
		_w25634_,
		_w25638_,
		_w25640_,
		_w25635_,
		_w25641_
	);
	LUT4 #(
		.INIT('h0080)
	) name19815 (
		_w25630_,
		_w25636_,
		_w25633_,
		_w25631_,
		_w25642_
	);
	LUT3 #(
		.INIT('h20)
	) name19816 (
		_w25630_,
		_w25633_,
		_w25631_,
		_w25643_
	);
	LUT4 #(
		.INIT('h0400)
	) name19817 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25644_
	);
	LUT2 #(
		.INIT('h1)
	) name19818 (
		_w25642_,
		_w25644_,
		_w25645_
	);
	LUT3 #(
		.INIT('h01)
	) name19819 (
		_w25630_,
		_w25633_,
		_w25631_,
		_w25646_
	);
	LUT4 #(
		.INIT('h0001)
	) name19820 (
		_w25630_,
		_w25636_,
		_w25633_,
		_w25631_,
		_w25647_
	);
	LUT4 #(
		.INIT('h0123)
	) name19821 (
		_w25632_,
		_w25642_,
		_w25643_,
		_w25647_,
		_w25648_
	);
	LUT2 #(
		.INIT('h8)
	) name19822 (
		_w25641_,
		_w25648_,
		_w25649_
	);
	LUT3 #(
		.INIT('h80)
	) name19823 (
		_w25632_,
		_w25630_,
		_w25636_,
		_w25650_
	);
	LUT4 #(
		.INIT('h0080)
	) name19824 (
		_w25632_,
		_w25630_,
		_w25636_,
		_w25633_,
		_w25651_
	);
	LUT4 #(
		.INIT('h0004)
	) name19825 (
		_w25630_,
		_w25636_,
		_w25633_,
		_w25631_,
		_w25652_
	);
	LUT3 #(
		.INIT('h01)
	) name19826 (
		_w25635_,
		_w25652_,
		_w25651_,
		_w25653_
	);
	LUT4 #(
		.INIT('hcc5f)
	) name19827 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25654_
	);
	LUT2 #(
		.INIT('h1)
	) name19828 (
		_w25636_,
		_w25654_,
		_w25655_
	);
	LUT4 #(
		.INIT('h2eff)
	) name19829 (
		_w25632_,
		_w25630_,
		_w25636_,
		_w25633_,
		_w25656_
	);
	LUT4 #(
		.INIT('hfff6)
	) name19830 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25657_
	);
	LUT3 #(
		.INIT('hd0)
	) name19831 (
		_w25631_,
		_w25656_,
		_w25657_,
		_w25658_
	);
	LUT3 #(
		.INIT('h40)
	) name19832 (
		_w25655_,
		_w25653_,
		_w25658_,
		_w25659_
	);
	LUT4 #(
		.INIT('h0020)
	) name19833 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25660_
	);
	LUT4 #(
		.INIT('hffde)
	) name19834 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25661_
	);
	LUT2 #(
		.INIT('h2)
	) name19835 (
		_w25636_,
		_w25661_,
		_w25662_
	);
	LUT3 #(
		.INIT('h10)
	) name19836 (
		_w25632_,
		_w25636_,
		_w25631_,
		_w25663_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name19837 (
		_w25632_,
		_w25642_,
		_w25637_,
		_w25663_,
		_w25664_
	);
	LUT2 #(
		.INIT('h4)
	) name19838 (
		_w25662_,
		_w25664_,
		_w25665_
	);
	LUT4 #(
		.INIT('ha955)
	) name19839 (
		\u0_L12_reg[20]/NET0131 ,
		_w25649_,
		_w25659_,
		_w25665_,
		_w25666_
	);
	LUT4 #(
		.INIT('h5fa6)
	) name19840 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25667_
	);
	LUT4 #(
		.INIT('h0400)
	) name19841 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25668_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name19842 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25669_
	);
	LUT4 #(
		.INIT('hcd7d)
	) name19843 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25670_
	);
	LUT4 #(
		.INIT('h3120)
	) name19844 (
		_w25559_,
		_w25668_,
		_w25667_,
		_w25670_,
		_w25671_
	);
	LUT2 #(
		.INIT('h1)
	) name19845 (
		_w25558_,
		_w25671_,
		_w25672_
	);
	LUT4 #(
		.INIT('hf57d)
	) name19846 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25673_
	);
	LUT2 #(
		.INIT('h2)
	) name19847 (
		_w25559_,
		_w25673_,
		_w25674_
	);
	LUT3 #(
		.INIT('h28)
	) name19848 (
		_w25561_,
		_w25562_,
		_w25563_,
		_w25675_
	);
	LUT3 #(
		.INIT('h04)
	) name19849 (
		_w25567_,
		_w25669_,
		_w25675_,
		_w25676_
	);
	LUT4 #(
		.INIT('h0800)
	) name19850 (
		_w25559_,
		_w25560_,
		_w25561_,
		_w25563_,
		_w25677_
	);
	LUT4 #(
		.INIT('h0010)
	) name19851 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25678_
	);
	LUT2 #(
		.INIT('h1)
	) name19852 (
		_w25677_,
		_w25678_,
		_w25679_
	);
	LUT4 #(
		.INIT('h5700)
	) name19853 (
		_w25558_,
		_w25674_,
		_w25676_,
		_w25679_,
		_w25680_
	);
	LUT3 #(
		.INIT('h9a)
	) name19854 (
		\u0_L12_reg[29]/NET0131 ,
		_w25672_,
		_w25680_,
		_w25681_
	);
	LUT4 #(
		.INIT('hc693)
	) name19855 (
		decrypt_pad,
		\u0_R12_reg[32]/NET0131 ,
		\u0_uk_K_r12_reg[28]/NET0131 ,
		\u0_uk_K_r12_reg[38]/NET0131 ,
		_w25682_
	);
	LUT4 #(
		.INIT('hc693)
	) name19856 (
		decrypt_pad,
		\u0_R12_reg[31]/P0001 ,
		\u0_uk_K_r12_reg[22]/NET0131 ,
		\u0_uk_K_r12_reg[28]/NET0131 ,
		_w25683_
	);
	LUT4 #(
		.INIT('hc963)
	) name19857 (
		decrypt_pad,
		\u0_R12_reg[29]/NET0131 ,
		\u0_uk_K_r12_reg[15]/NET0131 ,
		\u0_uk_K_r12_reg[9]/NET0131 ,
		_w25684_
	);
	LUT4 #(
		.INIT('hc963)
	) name19858 (
		decrypt_pad,
		\u0_R12_reg[1]/NET0131 ,
		\u0_uk_K_r12_reg[0]/NET0131 ,
		\u0_uk_K_r12_reg[49]/NET0131 ,
		_w25685_
	);
	LUT4 #(
		.INIT('hc963)
	) name19859 (
		decrypt_pad,
		\u0_R12_reg[30]/NET0131 ,
		\u0_uk_K_r12_reg[16]/NET0131 ,
		\u0_uk_K_r12_reg[38]/NET0131 ,
		_w25686_
	);
	LUT4 #(
		.INIT('hc693)
	) name19860 (
		decrypt_pad,
		\u0_R12_reg[28]/NET0131 ,
		\u0_uk_K_r12_reg[37]/NET0131 ,
		\u0_uk_K_r12_reg[43]/NET0131 ,
		_w25687_
	);
	LUT4 #(
		.INIT('h0040)
	) name19861 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25688_
	);
	LUT2 #(
		.INIT('h2)
	) name19862 (
		_w25684_,
		_w25685_,
		_w25689_
	);
	LUT4 #(
		.INIT('h44b4)
	) name19863 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25690_
	);
	LUT4 #(
		.INIT('h00f7)
	) name19864 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25683_,
		_w25691_
	);
	LUT4 #(
		.INIT('h00f6)
	) name19865 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25683_,
		_w25692_
	);
	LUT3 #(
		.INIT('h20)
	) name19866 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25693_
	);
	LUT4 #(
		.INIT('h2000)
	) name19867 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25694_
	);
	LUT4 #(
		.INIT('h00f2)
	) name19868 (
		_w25683_,
		_w25690_,
		_w25692_,
		_w25694_,
		_w25695_
	);
	LUT2 #(
		.INIT('h2)
	) name19869 (
		_w25682_,
		_w25695_,
		_w25696_
	);
	LUT4 #(
		.INIT('h0008)
	) name19870 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25697_
	);
	LUT4 #(
		.INIT('hfcf7)
	) name19871 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25698_
	);
	LUT2 #(
		.INIT('h4)
	) name19872 (
		_w25698_,
		_w25683_,
		_w25699_
	);
	LUT4 #(
		.INIT('h8000)
	) name19873 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25700_
	);
	LUT3 #(
		.INIT('h04)
	) name19874 (
		_w25686_,
		_w25687_,
		_w25683_,
		_w25701_
	);
	LUT2 #(
		.INIT('h1)
	) name19875 (
		_w25700_,
		_w25701_,
		_w25702_
	);
	LUT3 #(
		.INIT('h0d)
	) name19876 (
		_w25686_,
		_w25687_,
		_w25685_,
		_w25703_
	);
	LUT3 #(
		.INIT('h0b)
	) name19877 (
		_w25684_,
		_w25685_,
		_w25683_,
		_w25704_
	);
	LUT3 #(
		.INIT('h45)
	) name19878 (
		_w25688_,
		_w25703_,
		_w25704_,
		_w25705_
	);
	LUT4 #(
		.INIT('h4555)
	) name19879 (
		_w25682_,
		_w25699_,
		_w25702_,
		_w25705_,
		_w25706_
	);
	LUT4 #(
		.INIT('h0001)
	) name19880 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25707_
	);
	LUT4 #(
		.INIT('hffde)
	) name19881 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25708_
	);
	LUT4 #(
		.INIT('h0200)
	) name19882 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25709_
	);
	LUT4 #(
		.INIT('hf9de)
	) name19883 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25710_
	);
	LUT4 #(
		.INIT('h3f15)
	) name19884 (
		_w25683_,
		_w25701_,
		_w25689_,
		_w25710_,
		_w25711_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name19885 (
		\u0_L12_reg[5]/NET0131 ,
		_w25706_,
		_w25696_,
		_w25711_,
		_w25712_
	);
	LUT4 #(
		.INIT('hc963)
	) name19886 (
		decrypt_pad,
		\u0_R12_reg[8]/NET0131 ,
		\u0_uk_K_r12_reg[11]/NET0131 ,
		\u0_uk_K_r12_reg[3]/NET0131 ,
		_w25713_
	);
	LUT4 #(
		.INIT('hc693)
	) name19887 (
		decrypt_pad,
		\u0_R12_reg[7]/NET0131 ,
		\u0_uk_K_r12_reg[12]/NET0131 ,
		\u0_uk_K_r12_reg[20]/NET0131 ,
		_w25714_
	);
	LUT4 #(
		.INIT('hc693)
	) name19888 (
		decrypt_pad,
		\u0_R12_reg[5]/NET0131 ,
		\u0_uk_K_r12_reg[27]/NET0131 ,
		\u0_uk_K_r12_reg[3]/NET0131 ,
		_w25715_
	);
	LUT4 #(
		.INIT('hc963)
	) name19889 (
		decrypt_pad,
		\u0_R12_reg[4]/NET0131 ,
		\u0_uk_K_r12_reg[24]/NET0131 ,
		\u0_uk_K_r12_reg[48]/NET0131 ,
		_w25716_
	);
	LUT4 #(
		.INIT('hc693)
	) name19890 (
		decrypt_pad,
		\u0_R12_reg[9]/NET0131 ,
		\u0_uk_K_r12_reg[40]/NET0131 ,
		\u0_uk_K_r12_reg[48]/NET0131 ,
		_w25717_
	);
	LUT4 #(
		.INIT('hc693)
	) name19891 (
		decrypt_pad,
		\u0_R12_reg[6]/NET0131 ,
		\u0_uk_K_r12_reg[18]/NET0131 ,
		\u0_uk_K_r12_reg[26]/NET0131 ,
		_w25718_
	);
	LUT4 #(
		.INIT('h59fb)
	) name19892 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25719_
	);
	LUT2 #(
		.INIT('h1)
	) name19893 (
		_w25714_,
		_w25719_,
		_w25720_
	);
	LUT4 #(
		.INIT('h0034)
	) name19894 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25721_
	);
	LUT4 #(
		.INIT('h0800)
	) name19895 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25722_
	);
	LUT2 #(
		.INIT('h2)
	) name19896 (
		_w25717_,
		_w25718_,
		_w25723_
	);
	LUT4 #(
		.INIT('h0004)
	) name19897 (
		_w25714_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25724_
	);
	LUT4 #(
		.INIT('h4000)
	) name19898 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25725_
	);
	LUT4 #(
		.INIT('h0007)
	) name19899 (
		_w25714_,
		_w25722_,
		_w25724_,
		_w25725_,
		_w25726_
	);
	LUT4 #(
		.INIT('h5455)
	) name19900 (
		_w25713_,
		_w25720_,
		_w25721_,
		_w25726_,
		_w25727_
	);
	LUT4 #(
		.INIT('he6ee)
	) name19901 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25728_
	);
	LUT4 #(
		.INIT('h4044)
	) name19902 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25729_
	);
	LUT3 #(
		.INIT('h51)
	) name19903 (
		_w25714_,
		_w25715_,
		_w25718_,
		_w25730_
	);
	LUT4 #(
		.INIT('hf200)
	) name19904 (
		_w25713_,
		_w25728_,
		_w25729_,
		_w25730_,
		_w25731_
	);
	LUT3 #(
		.INIT('h10)
	) name19905 (
		_w25717_,
		_w25715_,
		_w25718_,
		_w25732_
	);
	LUT4 #(
		.INIT('h0100)
	) name19906 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25733_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name19907 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25734_
	);
	LUT2 #(
		.INIT('h2)
	) name19908 (
		_w25714_,
		_w25734_,
		_w25735_
	);
	LUT4 #(
		.INIT('h0082)
	) name19909 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25736_
	);
	LUT4 #(
		.INIT('h80a0)
	) name19910 (
		_w25714_,
		_w25716_,
		_w25715_,
		_w25718_,
		_w25737_
	);
	LUT3 #(
		.INIT('ha8)
	) name19911 (
		_w25713_,
		_w25736_,
		_w25737_,
		_w25738_
	);
	LUT3 #(
		.INIT('h01)
	) name19912 (
		_w25735_,
		_w25738_,
		_w25731_,
		_w25739_
	);
	LUT3 #(
		.INIT('h65)
	) name19913 (
		\u0_L12_reg[2]/NET0131 ,
		_w25727_,
		_w25739_,
		_w25740_
	);
	LUT4 #(
		.INIT('hbc5f)
	) name19914 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25741_
	);
	LUT4 #(
		.INIT('h0884)
	) name19915 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25742_
	);
	LUT4 #(
		.INIT('hcc04)
	) name19916 (
		_w25558_,
		_w25559_,
		_w25741_,
		_w25742_,
		_w25743_
	);
	LUT4 #(
		.INIT('hcbf5)
	) name19917 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25744_
	);
	LUT4 #(
		.INIT('h5051)
	) name19918 (
		_w25558_,
		_w25559_,
		_w25678_,
		_w25744_,
		_w25745_
	);
	LUT4 #(
		.INIT('h2000)
	) name19919 (
		_w25559_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25746_
	);
	LUT4 #(
		.INIT('h77fd)
	) name19920 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25747_
	);
	LUT4 #(
		.INIT('h0b00)
	) name19921 (
		_w25572_,
		_w25580_,
		_w25746_,
		_w25747_,
		_w25748_
	);
	LUT4 #(
		.INIT('h5f8c)
	) name19922 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25749_
	);
	LUT3 #(
		.INIT('h45)
	) name19923 (
		_w25559_,
		_w25561_,
		_w25562_,
		_w25750_
	);
	LUT2 #(
		.INIT('h4)
	) name19924 (
		_w25749_,
		_w25750_,
		_w25751_
	);
	LUT4 #(
		.INIT('h0031)
	) name19925 (
		_w25558_,
		_w25745_,
		_w25748_,
		_w25751_,
		_w25752_
	);
	LUT3 #(
		.INIT('h65)
	) name19926 (
		\u0_L12_reg[4]/NET0131 ,
		_w25743_,
		_w25752_,
		_w25753_
	);
	LUT3 #(
		.INIT('h02)
	) name19927 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25754_
	);
	LUT4 #(
		.INIT('h0082)
	) name19928 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25755_
	);
	LUT3 #(
		.INIT('hb0)
	) name19929 (
		_w25588_,
		_w25590_,
		_w25586_,
		_w25756_
	);
	LUT2 #(
		.INIT('h6)
	) name19930 (
		_w25589_,
		_w25587_,
		_w25757_
	);
	LUT4 #(
		.INIT('h0770)
	) name19931 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25758_
	);
	LUT2 #(
		.INIT('h1)
	) name19932 (
		_w25756_,
		_w25758_,
		_w25759_
	);
	LUT4 #(
		.INIT('h0100)
	) name19933 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25760_
	);
	LUT4 #(
		.INIT('h0400)
	) name19934 (
		_w25588_,
		_w25589_,
		_w25587_,
		_w25586_,
		_w25761_
	);
	LUT3 #(
		.INIT('h01)
	) name19935 (
		_w25596_,
		_w25760_,
		_w25761_,
		_w25762_
	);
	LUT3 #(
		.INIT('h10)
	) name19936 (
		_w25759_,
		_w25755_,
		_w25762_,
		_w25763_
	);
	LUT4 #(
		.INIT('h55fe)
	) name19937 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25764_
	);
	LUT2 #(
		.INIT('h2)
	) name19938 (
		_w25586_,
		_w25764_,
		_w25765_
	);
	LUT4 #(
		.INIT('h1020)
	) name19939 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w25766_
	);
	LUT2 #(
		.INIT('h9)
	) name19940 (
		_w25588_,
		_w25589_,
		_w25767_
	);
	LUT4 #(
		.INIT('h080c)
	) name19941 (
		_w25588_,
		_w25590_,
		_w25587_,
		_w25586_,
		_w25768_
	);
	LUT4 #(
		.INIT('h2022)
	) name19942 (
		_w25596_,
		_w25609_,
		_w25767_,
		_w25768_,
		_w25769_
	);
	LUT3 #(
		.INIT('h10)
	) name19943 (
		_w25766_,
		_w25765_,
		_w25769_,
		_w25770_
	);
	LUT3 #(
		.INIT('ha9)
	) name19944 (
		\u0_L12_reg[12]/NET0131 ,
		_w25763_,
		_w25770_,
		_w25771_
	);
	LUT4 #(
		.INIT('hfb4f)
	) name19945 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25772_
	);
	LUT4 #(
		.INIT('h7dff)
	) name19946 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25773_
	);
	LUT4 #(
		.INIT('h1000)
	) name19947 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25774_
	);
	LUT4 #(
		.INIT('heff3)
	) name19948 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25775_
	);
	LUT4 #(
		.INIT('hc480)
	) name19949 (
		_w25636_,
		_w25773_,
		_w25775_,
		_w25772_,
		_w25776_
	);
	LUT2 #(
		.INIT('h2)
	) name19950 (
		_w25635_,
		_w25776_,
		_w25777_
	);
	LUT4 #(
		.INIT('h0400)
	) name19951 (
		_w25632_,
		_w25636_,
		_w25633_,
		_w25631_,
		_w25778_
	);
	LUT3 #(
		.INIT('hdc)
	) name19952 (
		_w25632_,
		_w25630_,
		_w25631_,
		_w25779_
	);
	LUT2 #(
		.INIT('h8)
	) name19953 (
		_w25636_,
		_w25633_,
		_w25780_
	);
	LUT4 #(
		.INIT('h0045)
	) name19954 (
		_w25647_,
		_w25779_,
		_w25780_,
		_w25778_,
		_w25781_
	);
	LUT4 #(
		.INIT('hbabb)
	) name19955 (
		_w25632_,
		_w25630_,
		_w25636_,
		_w25631_,
		_w25782_
	);
	LUT3 #(
		.INIT('hc4)
	) name19956 (
		_w25633_,
		_w25657_,
		_w25782_,
		_w25783_
	);
	LUT3 #(
		.INIT('h15)
	) name19957 (
		_w25635_,
		_w25781_,
		_w25783_,
		_w25784_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name19958 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25785_
	);
	LUT2 #(
		.INIT('h1)
	) name19959 (
		_w25636_,
		_w25785_,
		_w25786_
	);
	LUT3 #(
		.INIT('h0b)
	) name19960 (
		_w25632_,
		_w25642_,
		_w25651_,
		_w25787_
	);
	LUT2 #(
		.INIT('h4)
	) name19961 (
		_w25786_,
		_w25787_,
		_w25788_
	);
	LUT4 #(
		.INIT('h5655)
	) name19962 (
		\u0_L12_reg[10]/NET0131 ,
		_w25777_,
		_w25784_,
		_w25788_,
		_w25789_
	);
	LUT4 #(
		.INIT('h5515)
	) name19963 (
		_w25714_,
		_w25716_,
		_w25717_,
		_w25715_,
		_w25790_
	);
	LUT3 #(
		.INIT('h40)
	) name19964 (
		_w25716_,
		_w25717_,
		_w25718_,
		_w25791_
	);
	LUT3 #(
		.INIT('h01)
	) name19965 (
		_w25717_,
		_w25715_,
		_w25718_,
		_w25792_
	);
	LUT4 #(
		.INIT('haaa8)
	) name19966 (
		_w25714_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25793_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name19967 (
		_w25732_,
		_w25790_,
		_w25791_,
		_w25793_,
		_w25794_
	);
	LUT4 #(
		.INIT('h0010)
	) name19968 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25795_
	);
	LUT4 #(
		.INIT('h0002)
	) name19969 (
		_w25713_,
		_w25724_,
		_w25725_,
		_w25795_,
		_w25796_
	);
	LUT2 #(
		.INIT('h4)
	) name19970 (
		_w25794_,
		_w25796_,
		_w25797_
	);
	LUT3 #(
		.INIT('h32)
	) name19971 (
		_w25714_,
		_w25716_,
		_w25715_,
		_w25798_
	);
	LUT2 #(
		.INIT('h8)
	) name19972 (
		_w25723_,
		_w25798_,
		_w25799_
	);
	LUT2 #(
		.INIT('h8)
	) name19973 (
		_w25714_,
		_w25716_,
		_w25800_
	);
	LUT3 #(
		.INIT('hb0)
	) name19974 (
		_w25717_,
		_w25715_,
		_w25718_,
		_w25801_
	);
	LUT3 #(
		.INIT('h15)
	) name19975 (
		_w25713_,
		_w25800_,
		_w25801_,
		_w25802_
	);
	LUT4 #(
		.INIT('h5455)
	) name19976 (
		_w25714_,
		_w25716_,
		_w25717_,
		_w25715_,
		_w25803_
	);
	LUT4 #(
		.INIT('h0400)
	) name19977 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25804_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name19978 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25805_
	);
	LUT2 #(
		.INIT('h8)
	) name19979 (
		_w25803_,
		_w25805_,
		_w25806_
	);
	LUT3 #(
		.INIT('h40)
	) name19980 (
		_w25799_,
		_w25802_,
		_w25806_,
		_w25807_
	);
	LUT4 #(
		.INIT('h2000)
	) name19981 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25808_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name19982 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25809_
	);
	LUT3 #(
		.INIT('h09)
	) name19983 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25810_
	);
	LUT3 #(
		.INIT('h02)
	) name19984 (
		_w25716_,
		_w25717_,
		_w25718_,
		_w25811_
	);
	LUT4 #(
		.INIT('h0020)
	) name19985 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25812_
	);
	LUT3 #(
		.INIT('h02)
	) name19986 (
		_w25714_,
		_w25812_,
		_w25810_,
		_w25813_
	);
	LUT3 #(
		.INIT('h40)
	) name19987 (
		_w25799_,
		_w25802_,
		_w25813_,
		_w25814_
	);
	LUT4 #(
		.INIT('h001f)
	) name19988 (
		_w25797_,
		_w25807_,
		_w25809_,
		_w25814_,
		_w25815_
	);
	LUT2 #(
		.INIT('h9)
	) name19989 (
		\u0_L12_reg[13]/NET0131 ,
		_w25815_,
		_w25816_
	);
	LUT4 #(
		.INIT('hc693)
	) name19990 (
		decrypt_pad,
		\u0_R12_reg[20]/NET0131 ,
		\u0_uk_K_r12_reg[44]/P0001 ,
		\u0_uk_K_r12_reg[50]/NET0131 ,
		_w25817_
	);
	LUT4 #(
		.INIT('hc693)
	) name19991 (
		decrypt_pad,
		\u0_R12_reg[18]/NET0131 ,
		\u0_uk_K_r12_reg[42]/NET0131 ,
		\u0_uk_K_r12_reg[52]/NET0131 ,
		_w25818_
	);
	LUT4 #(
		.INIT('hc963)
	) name19992 (
		decrypt_pad,
		\u0_R12_reg[17]/NET0131 ,
		\u0_uk_K_r12_reg[30]/NET0131 ,
		\u0_uk_K_r12_reg[52]/NET0131 ,
		_w25819_
	);
	LUT4 #(
		.INIT('hc693)
	) name19993 (
		decrypt_pad,
		\u0_R12_reg[16]/NET0131 ,
		\u0_uk_K_r12_reg[2]/NET0131 ,
		\u0_uk_K_r12_reg[8]/NET0131 ,
		_w25820_
	);
	LUT4 #(
		.INIT('hc693)
	) name19994 (
		decrypt_pad,
		\u0_R12_reg[21]/NET0131 ,
		\u0_uk_K_r12_reg[14]/NET0131 ,
		\u0_uk_K_r12_reg[51]/NET0131 ,
		_w25821_
	);
	LUT4 #(
		.INIT('h0180)
	) name19995 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25822_
	);
	LUT3 #(
		.INIT('h80)
	) name19996 (
		_w25820_,
		_w25821_,
		_w25819_,
		_w25823_
	);
	LUT4 #(
		.INIT('h0800)
	) name19997 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25824_
	);
	LUT4 #(
		.INIT('hc693)
	) name19998 (
		decrypt_pad,
		\u0_R12_reg[19]/NET0131 ,
		\u0_uk_K_r12_reg[29]/NET0131 ,
		\u0_uk_K_r12_reg[35]/NET0131 ,
		_w25825_
	);
	LUT4 #(
		.INIT('h0002)
	) name19999 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25826_
	);
	LUT4 #(
		.INIT('hcfbb)
	) name20000 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25827_
	);
	LUT4 #(
		.INIT('h0100)
	) name20001 (
		_w25825_,
		_w25824_,
		_w25826_,
		_w25827_,
		_w25828_
	);
	LUT4 #(
		.INIT('haaa8)
	) name20002 (
		_w25825_,
		_w25820_,
		_w25821_,
		_w25819_,
		_w25829_
	);
	LUT4 #(
		.INIT('h7a7f)
	) name20003 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25830_
	);
	LUT2 #(
		.INIT('h8)
	) name20004 (
		_w25829_,
		_w25830_,
		_w25831_
	);
	LUT4 #(
		.INIT('h4445)
	) name20005 (
		_w25817_,
		_w25822_,
		_w25828_,
		_w25831_,
		_w25832_
	);
	LUT4 #(
		.INIT('h95b3)
	) name20006 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25833_
	);
	LUT2 #(
		.INIT('h2)
	) name20007 (
		_w25825_,
		_w25833_,
		_w25834_
	);
	LUT2 #(
		.INIT('h1)
	) name20008 (
		_w25825_,
		_w25818_,
		_w25835_
	);
	LUT3 #(
		.INIT('hbe)
	) name20009 (
		_w25820_,
		_w25821_,
		_w25819_,
		_w25836_
	);
	LUT2 #(
		.INIT('h2)
	) name20010 (
		_w25835_,
		_w25836_,
		_w25837_
	);
	LUT3 #(
		.INIT('hb0)
	) name20011 (
		_w25825_,
		_w25818_,
		_w25819_,
		_w25838_
	);
	LUT4 #(
		.INIT('h8808)
	) name20012 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25839_
	);
	LUT4 #(
		.INIT('h0020)
	) name20013 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25840_
	);
	LUT4 #(
		.INIT('h0200)
	) name20014 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25841_
	);
	LUT4 #(
		.INIT('hfddf)
	) name20015 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25842_
	);
	LUT3 #(
		.INIT('hb0)
	) name20016 (
		_w25838_,
		_w25839_,
		_w25842_,
		_w25843_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name20017 (
		_w25817_,
		_w25834_,
		_w25837_,
		_w25843_,
		_w25844_
	);
	LUT4 #(
		.INIT('h1040)
	) name20018 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25845_
	);
	LUT4 #(
		.INIT('h0010)
	) name20019 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25846_
	);
	LUT4 #(
		.INIT('hfad8)
	) name20020 (
		_w25825_,
		_w25841_,
		_w25845_,
		_w25846_,
		_w25847_
	);
	LUT4 #(
		.INIT('h5556)
	) name20021 (
		\u0_L12_reg[14]/NET0131 ,
		_w25844_,
		_w25832_,
		_w25847_,
		_w25848_
	);
	LUT4 #(
		.INIT('h3c2f)
	) name20022 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25849_
	);
	LUT4 #(
		.INIT('h0004)
	) name20023 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25850_
	);
	LUT4 #(
		.INIT('h0501)
	) name20024 (
		_w25682_,
		_w25683_,
		_w25850_,
		_w25849_,
		_w25851_
	);
	LUT4 #(
		.INIT('h0020)
	) name20025 (
		_w25686_,
		_w25684_,
		_w25685_,
		_w25683_,
		_w25852_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name20026 (
		_w25682_,
		_w25686_,
		_w25687_,
		_w25684_,
		_w25853_
	);
	LUT4 #(
		.INIT('h0100)
	) name20027 (
		_w25687_,
		_w25684_,
		_w25685_,
		_w25683_,
		_w25854_
	);
	LUT4 #(
		.INIT('hf7df)
	) name20028 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25855_
	);
	LUT4 #(
		.INIT('h1000)
	) name20029 (
		_w25854_,
		_w25852_,
		_w25853_,
		_w25855_,
		_w25856_
	);
	LUT2 #(
		.INIT('h1)
	) name20030 (
		_w25851_,
		_w25856_,
		_w25857_
	);
	LUT4 #(
		.INIT('h1000)
	) name20031 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25858_
	);
	LUT3 #(
		.INIT('h08)
	) name20032 (
		_w25691_,
		_w25708_,
		_w25858_,
		_w25859_
	);
	LUT4 #(
		.INIT('h0100)
	) name20033 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25860_
	);
	LUT3 #(
		.INIT('h02)
	) name20034 (
		_w25683_,
		_w25694_,
		_w25860_,
		_w25861_
	);
	LUT4 #(
		.INIT('h0004)
	) name20035 (
		_w25682_,
		_w25687_,
		_w25684_,
		_w25683_,
		_w25862_
	);
	LUT3 #(
		.INIT('h0e)
	) name20036 (
		_w25859_,
		_w25861_,
		_w25862_,
		_w25863_
	);
	LUT3 #(
		.INIT('h65)
	) name20037 (
		\u0_L12_reg[15]/P0001 ,
		_w25857_,
		_w25863_,
		_w25864_
	);
	LUT4 #(
		.INIT('h3050)
	) name20038 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25865_
	);
	LUT3 #(
		.INIT('h01)
	) name20039 (
		_w25632_,
		_w25633_,
		_w25631_,
		_w25866_
	);
	LUT4 #(
		.INIT('hfad8)
	) name20040 (
		_w25636_,
		_w25660_,
		_w25865_,
		_w25866_,
		_w25867_
	);
	LUT4 #(
		.INIT('h7bbf)
	) name20041 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25868_
	);
	LUT3 #(
		.INIT('h45)
	) name20042 (
		_w25635_,
		_w25867_,
		_w25868_,
		_w25869_
	);
	LUT4 #(
		.INIT('hb3fb)
	) name20043 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25870_
	);
	LUT4 #(
		.INIT('h0080)
	) name20044 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25871_
	);
	LUT4 #(
		.INIT('hfd7d)
	) name20045 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25872_
	);
	LUT4 #(
		.INIT('h04cc)
	) name20046 (
		_w25636_,
		_w25635_,
		_w25870_,
		_w25872_,
		_w25873_
	);
	LUT4 #(
		.INIT('h7df7)
	) name20047 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25874_
	);
	LUT2 #(
		.INIT('h2)
	) name20048 (
		_w25636_,
		_w25874_,
		_w25875_
	);
	LUT4 #(
		.INIT('hccef)
	) name20049 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25876_
	);
	LUT2 #(
		.INIT('h8)
	) name20050 (
		_w25636_,
		_w25635_,
		_w25877_
	);
	LUT2 #(
		.INIT('h4)
	) name20051 (
		_w25876_,
		_w25877_,
		_w25878_
	);
	LUT4 #(
		.INIT('hccdf)
	) name20052 (
		_w25632_,
		_w25636_,
		_w25646_,
		_w25871_,
		_w25879_
	);
	LUT4 #(
		.INIT('h0100)
	) name20053 (
		_w25875_,
		_w25878_,
		_w25873_,
		_w25879_,
		_w25880_
	);
	LUT3 #(
		.INIT('h65)
	) name20054 (
		\u0_L12_reg[1]/NET0131 ,
		_w25869_,
		_w25880_,
		_w25881_
	);
	LUT4 #(
		.INIT('h4a7f)
	) name20055 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25882_
	);
	LUT4 #(
		.INIT('hf7bb)
	) name20056 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25883_
	);
	LUT4 #(
		.INIT('hfe7d)
	) name20057 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25884_
	);
	LUT4 #(
		.INIT('he400)
	) name20058 (
		_w25683_,
		_w25883_,
		_w25882_,
		_w25884_,
		_w25885_
	);
	LUT2 #(
		.INIT('h2)
	) name20059 (
		_w25682_,
		_w25885_,
		_w25886_
	);
	LUT4 #(
		.INIT('h0004)
	) name20060 (
		_w25687_,
		_w25684_,
		_w25685_,
		_w25683_,
		_w25887_
	);
	LUT3 #(
		.INIT('h01)
	) name20061 (
		_w25697_,
		_w25693_,
		_w25887_,
		_w25888_
	);
	LUT4 #(
		.INIT('h0040)
	) name20062 (
		_w25686_,
		_w25687_,
		_w25685_,
		_w25683_,
		_w25889_
	);
	LUT2 #(
		.INIT('h1)
	) name20063 (
		_w25707_,
		_w25889_,
		_w25890_
	);
	LUT4 #(
		.INIT('hf737)
	) name20064 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25891_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name20065 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25683_,
		_w25892_
	);
	LUT4 #(
		.INIT('hf351)
	) name20066 (
		_w25685_,
		_w25683_,
		_w25891_,
		_w25892_,
		_w25893_
	);
	LUT4 #(
		.INIT('h1555)
	) name20067 (
		_w25682_,
		_w25888_,
		_w25890_,
		_w25893_,
		_w25894_
	);
	LUT4 #(
		.INIT('h0100)
	) name20068 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25683_,
		_w25895_
	);
	LUT3 #(
		.INIT('h07)
	) name20069 (
		_w25684_,
		_w25889_,
		_w25895_,
		_w25896_
	);
	LUT4 #(
		.INIT('h5655)
	) name20070 (
		\u0_L12_reg[21]/NET0131 ,
		_w25894_,
		_w25886_,
		_w25896_,
		_w25897_
	);
	LUT4 #(
		.INIT('h67a8)
	) name20071 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25898_
	);
	LUT4 #(
		.INIT('hfa77)
	) name20072 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25899_
	);
	LUT4 #(
		.INIT('hd3ff)
	) name20073 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25900_
	);
	LUT4 #(
		.INIT('hd800)
	) name20074 (
		_w25825_,
		_w25898_,
		_w25899_,
		_w25900_,
		_w25901_
	);
	LUT2 #(
		.INIT('h2)
	) name20075 (
		_w25817_,
		_w25901_,
		_w25902_
	);
	LUT4 #(
		.INIT('hdfef)
	) name20076 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25903_
	);
	LUT4 #(
		.INIT('hdfeb)
	) name20077 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25904_
	);
	LUT2 #(
		.INIT('h2)
	) name20078 (
		_w25825_,
		_w25904_,
		_w25905_
	);
	LUT3 #(
		.INIT('hb0)
	) name20079 (
		_w25820_,
		_w25818_,
		_w25819_,
		_w25906_
	);
	LUT4 #(
		.INIT('hf504)
	) name20080 (
		_w25825_,
		_w25820_,
		_w25821_,
		_w25819_,
		_w25907_
	);
	LUT3 #(
		.INIT('h8a)
	) name20081 (
		_w25825_,
		_w25821_,
		_w25819_,
		_w25908_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name20082 (
		_w25825_,
		_w25820_,
		_w25818_,
		_w25819_,
		_w25909_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name20083 (
		_w25906_,
		_w25907_,
		_w25908_,
		_w25909_,
		_w25910_
	);
	LUT4 #(
		.INIT('h0040)
	) name20084 (
		_w25825_,
		_w25820_,
		_w25818_,
		_w25819_,
		_w25911_
	);
	LUT2 #(
		.INIT('h1)
	) name20085 (
		_w25824_,
		_w25911_,
		_w25912_
	);
	LUT4 #(
		.INIT('h0e00)
	) name20086 (
		_w25817_,
		_w25910_,
		_w25905_,
		_w25912_,
		_w25913_
	);
	LUT3 #(
		.INIT('h65)
	) name20087 (
		\u0_L12_reg[25]/NET0131 ,
		_w25902_,
		_w25913_,
		_w25914_
	);
	LUT4 #(
		.INIT('h0004)
	) name20088 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25915_
	);
	LUT4 #(
		.INIT('h0002)
	) name20089 (
		_w25635_,
		_w25652_,
		_w25871_,
		_w25915_,
		_w25916_
	);
	LUT4 #(
		.INIT('h5eff)
	) name20090 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25917_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name20091 (
		_w25630_,
		_w25636_,
		_w25633_,
		_w25631_,
		_w25918_
	);
	LUT4 #(
		.INIT('hfc54)
	) name20092 (
		_w25632_,
		_w25636_,
		_w25917_,
		_w25918_,
		_w25919_
	);
	LUT4 #(
		.INIT('h00ef)
	) name20093 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25635_,
		_w25920_
	);
	LUT3 #(
		.INIT('hb0)
	) name20094 (
		_w25639_,
		_w25650_,
		_w25920_,
		_w25921_
	);
	LUT4 #(
		.INIT('h153f)
	) name20095 (
		_w25645_,
		_w25916_,
		_w25919_,
		_w25921_,
		_w25922_
	);
	LUT4 #(
		.INIT('h4014)
	) name20096 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25923_
	);
	LUT4 #(
		.INIT('hfdcc)
	) name20097 (
		_w25632_,
		_w25630_,
		_w25633_,
		_w25631_,
		_w25924_
	);
	LUT4 #(
		.INIT('h0054)
	) name20098 (
		_w25636_,
		_w25635_,
		_w25924_,
		_w25923_,
		_w25925_
	);
	LUT3 #(
		.INIT('h02)
	) name20099 (
		_w25636_,
		_w25644_,
		_w25774_,
		_w25926_
	);
	LUT2 #(
		.INIT('h1)
	) name20100 (
		_w25925_,
		_w25926_,
		_w25927_
	);
	LUT3 #(
		.INIT('h56)
	) name20101 (
		\u0_L12_reg[26]/NET0131 ,
		_w25922_,
		_w25927_,
		_w25928_
	);
	LUT3 #(
		.INIT('hf4)
	) name20102 (
		_w25820_,
		_w25818_,
		_w25819_,
		_w25929_
	);
	LUT3 #(
		.INIT('h82)
	) name20103 (
		_w25825_,
		_w25820_,
		_w25821_,
		_w25930_
	);
	LUT4 #(
		.INIT('haa8a)
	) name20104 (
		_w25817_,
		_w25825_,
		_w25820_,
		_w25818_,
		_w25931_
	);
	LUT4 #(
		.INIT('h4500)
	) name20105 (
		_w25845_,
		_w25929_,
		_w25930_,
		_w25931_,
		_w25932_
	);
	LUT3 #(
		.INIT('h02)
	) name20106 (
		_w25825_,
		_w25823_,
		_w25826_,
		_w25933_
	);
	LUT4 #(
		.INIT('h4404)
	) name20107 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25934_
	);
	LUT4 #(
		.INIT('h5515)
	) name20108 (
		_w25825_,
		_w25820_,
		_w25821_,
		_w25819_,
		_w25935_
	);
	LUT2 #(
		.INIT('h4)
	) name20109 (
		_w25934_,
		_w25935_,
		_w25936_
	);
	LUT4 #(
		.INIT('h5455)
	) name20110 (
		_w25817_,
		_w25820_,
		_w25818_,
		_w25819_,
		_w25937_
	);
	LUT2 #(
		.INIT('h8)
	) name20111 (
		_w25903_,
		_w25937_,
		_w25938_
	);
	LUT4 #(
		.INIT('h0155)
	) name20112 (
		_w25932_,
		_w25933_,
		_w25936_,
		_w25938_,
		_w25939_
	);
	LUT4 #(
		.INIT('h0040)
	) name20113 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25940_
	);
	LUT4 #(
		.INIT('hcbbf)
	) name20114 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w25941_
	);
	LUT3 #(
		.INIT('hb1)
	) name20115 (
		_w25825_,
		_w25840_,
		_w25941_,
		_w25942_
	);
	LUT3 #(
		.INIT('h65)
	) name20116 (
		\u0_L12_reg[8]/NET0131 ,
		_w25939_,
		_w25942_,
		_w25943_
	);
	LUT4 #(
		.INIT('hfaa7)
	) name20117 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25944_
	);
	LUT4 #(
		.INIT('h7def)
	) name20118 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25945_
	);
	LUT4 #(
		.INIT('h0455)
	) name20119 (
		_w25526_,
		_w25541_,
		_w25944_,
		_w25945_,
		_w25946_
	);
	LUT4 #(
		.INIT('ha7ff)
	) name20120 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w25947_
	);
	LUT2 #(
		.INIT('h2)
	) name20121 (
		_w25526_,
		_w25947_,
		_w25948_
	);
	LUT4 #(
		.INIT('h1030)
	) name20122 (
		_w25533_,
		_w25539_,
		_w25541_,
		_w25543_,
		_w25949_
	);
	LUT4 #(
		.INIT('h007e)
	) name20123 (
		_w25529_,
		_w25528_,
		_w25530_,
		_w25541_,
		_w25950_
	);
	LUT4 #(
		.INIT('h0400)
	) name20124 (
		_w25527_,
		_w25526_,
		_w25528_,
		_w25530_,
		_w25951_
	);
	LUT3 #(
		.INIT('h54)
	) name20125 (
		_w25526_,
		_w25528_,
		_w25530_,
		_w25952_
	);
	LUT3 #(
		.INIT('ha8)
	) name20126 (
		_w25527_,
		_w25529_,
		_w25530_,
		_w25953_
	);
	LUT4 #(
		.INIT('h0015)
	) name20127 (
		_w25534_,
		_w25952_,
		_w25953_,
		_w25951_,
		_w25954_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name20128 (
		_w25948_,
		_w25949_,
		_w25950_,
		_w25954_,
		_w25955_
	);
	LUT3 #(
		.INIT('h13)
	) name20129 (
		_w25547_,
		_w25554_,
		_w25624_,
		_w25956_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name20130 (
		\u0_L12_reg[23]/NET0131 ,
		_w25955_,
		_w25946_,
		_w25956_,
		_w25957_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name20131 (
		_w25559_,
		_w25560_,
		_w25561_,
		_w25562_,
		_w25958_
	);
	LUT4 #(
		.INIT('h1900)
	) name20132 (
		_w25559_,
		_w25560_,
		_w25561_,
		_w25562_,
		_w25959_
	);
	LUT3 #(
		.INIT('h31)
	) name20133 (
		_w25560_,
		_w25562_,
		_w25563_,
		_w25960_
	);
	LUT3 #(
		.INIT('h21)
	) name20134 (
		_w25560_,
		_w25562_,
		_w25563_,
		_w25961_
	);
	LUT4 #(
		.INIT('h3211)
	) name20135 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25962_
	);
	LUT4 #(
		.INIT('h00fd)
	) name20136 (
		_w25561_,
		_w25576_,
		_w25961_,
		_w25962_,
		_w25963_
	);
	LUT3 #(
		.INIT('ha8)
	) name20137 (
		_w25558_,
		_w25959_,
		_w25963_,
		_w25964_
	);
	LUT4 #(
		.INIT('h8000)
	) name20138 (
		_w25560_,
		_w25561_,
		_w25562_,
		_w25563_,
		_w25965_
	);
	LUT4 #(
		.INIT('h5504)
	) name20139 (
		_w25558_,
		_w25958_,
		_w25960_,
		_w25965_,
		_w25966_
	);
	LUT4 #(
		.INIT('h0401)
	) name20140 (
		_w25558_,
		_w25560_,
		_w25562_,
		_w25563_,
		_w25967_
	);
	LUT3 #(
		.INIT('h54)
	) name20141 (
		_w25559_,
		_w25564_,
		_w25967_,
		_w25968_
	);
	LUT3 #(
		.INIT('h01)
	) name20142 (
		_w25578_,
		_w25968_,
		_w25966_,
		_w25969_
	);
	LUT3 #(
		.INIT('h65)
	) name20143 (
		\u0_L12_reg[19]/P0001 ,
		_w25964_,
		_w25969_,
		_w25970_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name20144 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25971_
	);
	LUT2 #(
		.INIT('h2)
	) name20145 (
		_w25714_,
		_w25971_,
		_w25972_
	);
	LUT4 #(
		.INIT('hbfae)
	) name20146 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25973_
	);
	LUT2 #(
		.INIT('h1)
	) name20147 (
		_w25714_,
		_w25973_,
		_w25974_
	);
	LUT4 #(
		.INIT('h7737)
	) name20148 (
		_w25714_,
		_w25716_,
		_w25717_,
		_w25715_,
		_w25975_
	);
	LUT3 #(
		.INIT('h32)
	) name20149 (
		_w25718_,
		_w25804_,
		_w25975_,
		_w25976_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name20150 (
		_w25713_,
		_w25974_,
		_w25972_,
		_w25976_,
		_w25977_
	);
	LUT4 #(
		.INIT('hdaff)
	) name20151 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25978_
	);
	LUT2 #(
		.INIT('h1)
	) name20152 (
		_w25714_,
		_w25978_,
		_w25979_
	);
	LUT4 #(
		.INIT('h1145)
	) name20153 (
		_w25714_,
		_w25716_,
		_w25717_,
		_w25715_,
		_w25980_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name20154 (
		_w25714_,
		_w25811_,
		_w25973_,
		_w25980_,
		_w25981_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name20155 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w25982_
	);
	LUT4 #(
		.INIT('h2322)
	) name20156 (
		_w25713_,
		_w25979_,
		_w25981_,
		_w25982_,
		_w25983_
	);
	LUT3 #(
		.INIT('h65)
	) name20157 (
		\u0_L12_reg[28]/NET0131 ,
		_w25977_,
		_w25983_,
		_w25984_
	);
	LUT4 #(
		.INIT('h3fef)
	) name20158 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25985_
	);
	LUT4 #(
		.INIT('hce3e)
	) name20159 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25986_
	);
	LUT4 #(
		.INIT('hdaf7)
	) name20160 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25987_
	);
	LUT4 #(
		.INIT('he400)
	) name20161 (
		_w25683_,
		_w25986_,
		_w25985_,
		_w25987_,
		_w25988_
	);
	LUT2 #(
		.INIT('h2)
	) name20162 (
		_w25682_,
		_w25988_,
		_w25989_
	);
	LUT4 #(
		.INIT('hdf00)
	) name20163 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25683_,
		_w25990_
	);
	LUT3 #(
		.INIT('h4b)
	) name20164 (
		_w25686_,
		_w25684_,
		_w25685_,
		_w25991_
	);
	LUT2 #(
		.INIT('h8)
	) name20165 (
		_w25990_,
		_w25991_,
		_w25992_
	);
	LUT4 #(
		.INIT('h0080)
	) name20166 (
		_w25686_,
		_w25687_,
		_w25685_,
		_w25683_,
		_w25993_
	);
	LUT3 #(
		.INIT('h01)
	) name20167 (
		_w25709_,
		_w25887_,
		_w25993_,
		_w25994_
	);
	LUT3 #(
		.INIT('h45)
	) name20168 (
		_w25682_,
		_w25992_,
		_w25994_,
		_w25995_
	);
	LUT4 #(
		.INIT('hfbdf)
	) name20169 (
		_w25686_,
		_w25687_,
		_w25684_,
		_w25685_,
		_w25996_
	);
	LUT2 #(
		.INIT('h1)
	) name20170 (
		_w25683_,
		_w25996_,
		_w25997_
	);
	LUT4 #(
		.INIT('h0200)
	) name20171 (
		_w25686_,
		_w25684_,
		_w25685_,
		_w25683_,
		_w25998_
	);
	LUT3 #(
		.INIT('h07)
	) name20172 (
		_w25701_,
		_w25689_,
		_w25998_,
		_w25999_
	);
	LUT2 #(
		.INIT('h4)
	) name20173 (
		_w25997_,
		_w25999_,
		_w26000_
	);
	LUT4 #(
		.INIT('h5655)
	) name20174 (
		\u0_L12_reg[27]/NET0131 ,
		_w25995_,
		_w25989_,
		_w26000_,
		_w26001_
	);
	LUT4 #(
		.INIT('ha025)
	) name20175 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w26002_
	);
	LUT4 #(
		.INIT('h5a48)
	) name20176 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w26003_
	);
	LUT4 #(
		.INIT('h9bff)
	) name20177 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w26004_
	);
	LUT4 #(
		.INIT('hfd00)
	) name20178 (
		_w25596_,
		_w26003_,
		_w26002_,
		_w26004_,
		_w26005_
	);
	LUT2 #(
		.INIT('h1)
	) name20179 (
		_w25586_,
		_w26005_,
		_w26006_
	);
	LUT4 #(
		.INIT('hf700)
	) name20180 (
		_w25588_,
		_w25589_,
		_w25587_,
		_w25586_,
		_w26007_
	);
	LUT4 #(
		.INIT('haa8d)
	) name20181 (
		_w25586_,
		_w25599_,
		_w25757_,
		_w25754_,
		_w26008_
	);
	LUT4 #(
		.INIT('h79bf)
	) name20182 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w26009_
	);
	LUT3 #(
		.INIT('h45)
	) name20183 (
		_w25596_,
		_w26008_,
		_w26009_,
		_w26010_
	);
	LUT2 #(
		.INIT('h8)
	) name20184 (
		_w25586_,
		_w25604_,
		_w26011_
	);
	LUT4 #(
		.INIT('hc7f2)
	) name20185 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w26012_
	);
	LUT3 #(
		.INIT('hd0)
	) name20186 (
		_w25589_,
		_w25586_,
		_w25596_,
		_w26013_
	);
	LUT3 #(
		.INIT('h10)
	) name20187 (
		_w25607_,
		_w26012_,
		_w26013_,
		_w26014_
	);
	LUT2 #(
		.INIT('h1)
	) name20188 (
		_w26011_,
		_w26014_,
		_w26015_
	);
	LUT4 #(
		.INIT('h5655)
	) name20189 (
		\u0_L12_reg[32]/NET0131 ,
		_w26010_,
		_w26006_,
		_w26015_,
		_w26016_
	);
	LUT4 #(
		.INIT('hb3ff)
	) name20190 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w26017_
	);
	LUT3 #(
		.INIT('h20)
	) name20191 (
		_w25817_,
		_w25840_,
		_w26017_,
		_w26018_
	);
	LUT4 #(
		.INIT('h00d0)
	) name20192 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w26019_
	);
	LUT4 #(
		.INIT('h2e26)
	) name20193 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w26020_
	);
	LUT3 #(
		.INIT('h10)
	) name20194 (
		_w25817_,
		_w26019_,
		_w26020_,
		_w26021_
	);
	LUT4 #(
		.INIT('h0081)
	) name20195 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w26022_
	);
	LUT3 #(
		.INIT('h01)
	) name20196 (
		_w25825_,
		_w25841_,
		_w26022_,
		_w26023_
	);
	LUT3 #(
		.INIT('he0)
	) name20197 (
		_w26018_,
		_w26021_,
		_w26023_,
		_w26024_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name20198 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w26025_
	);
	LUT3 #(
		.INIT('h10)
	) name20199 (
		_w25817_,
		_w26019_,
		_w26025_,
		_w26026_
	);
	LUT4 #(
		.INIT('he6f7)
	) name20200 (
		_w25820_,
		_w25821_,
		_w25818_,
		_w25819_,
		_w26027_
	);
	LUT3 #(
		.INIT('h20)
	) name20201 (
		_w25817_,
		_w25840_,
		_w26027_,
		_w26028_
	);
	LUT3 #(
		.INIT('h02)
	) name20202 (
		_w25825_,
		_w25826_,
		_w25940_,
		_w26029_
	);
	LUT3 #(
		.INIT('he0)
	) name20203 (
		_w26026_,
		_w26028_,
		_w26029_,
		_w26030_
	);
	LUT3 #(
		.INIT('ha9)
	) name20204 (
		\u0_L12_reg[3]/NET0131 ,
		_w26024_,
		_w26030_,
		_w26031_
	);
	LUT4 #(
		.INIT('hc693)
	) name20205 (
		decrypt_pad,
		\u0_R12_reg[12]/NET0131 ,
		\u0_uk_K_r12_reg[13]/NET0131 ,
		\u0_uk_K_r12_reg[46]/NET0131 ,
		_w26032_
	);
	LUT4 #(
		.INIT('hc693)
	) name20206 (
		decrypt_pad,
		\u0_R12_reg[9]/NET0131 ,
		\u0_uk_K_r12_reg[46]/NET0131 ,
		\u0_uk_K_r12_reg[54]/NET0131 ,
		_w26033_
	);
	LUT4 #(
		.INIT('hc693)
	) name20207 (
		decrypt_pad,
		\u0_R12_reg[10]/NET0131 ,
		\u0_uk_K_r12_reg[54]/NET0131 ,
		\u0_uk_K_r12_reg[5]/NET0131 ,
		_w26034_
	);
	LUT2 #(
		.INIT('h8)
	) name20208 (
		_w26033_,
		_w26034_,
		_w26035_
	);
	LUT4 #(
		.INIT('hc693)
	) name20209 (
		decrypt_pad,
		\u0_R12_reg[8]/NET0131 ,
		\u0_uk_K_r12_reg[17]/NET0131 ,
		\u0_uk_K_r12_reg[25]/NET0131 ,
		_w26036_
	);
	LUT4 #(
		.INIT('hc693)
	) name20210 (
		decrypt_pad,
		\u0_R12_reg[11]/NET0131 ,
		\u0_uk_K_r12_reg[55]/NET0131 ,
		\u0_uk_K_r12_reg[6]/NET0131 ,
		_w26037_
	);
	LUT4 #(
		.INIT('hc693)
	) name20211 (
		decrypt_pad,
		\u0_R12_reg[13]/NET0131 ,
		\u0_uk_K_r12_reg[26]/NET0131 ,
		\u0_uk_K_r12_reg[34]/NET0131 ,
		_w26038_
	);
	LUT3 #(
		.INIT('h1a)
	) name20212 (
		_w26036_,
		_w26037_,
		_w26038_,
		_w26039_
	);
	LUT4 #(
		.INIT('h0200)
	) name20213 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26037_,
		_w26040_
	);
	LUT3 #(
		.INIT('h07)
	) name20214 (
		_w26035_,
		_w26039_,
		_w26040_,
		_w26041_
	);
	LUT2 #(
		.INIT('h1)
	) name20215 (
		_w26033_,
		_w26034_,
		_w26042_
	);
	LUT4 #(
		.INIT('he00e)
	) name20216 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26043_
	);
	LUT4 #(
		.INIT('h6006)
	) name20217 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26044_
	);
	LUT3 #(
		.INIT('h07)
	) name20218 (
		_w26039_,
		_w26042_,
		_w26044_,
		_w26045_
	);
	LUT3 #(
		.INIT('h15)
	) name20219 (
		_w26032_,
		_w26041_,
		_w26045_,
		_w26046_
	);
	LUT4 #(
		.INIT('ha25f)
	) name20220 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26047_
	);
	LUT2 #(
		.INIT('h8)
	) name20221 (
		_w26032_,
		_w26037_,
		_w26048_
	);
	LUT2 #(
		.INIT('h4)
	) name20222 (
		_w26047_,
		_w26048_,
		_w26049_
	);
	LUT2 #(
		.INIT('h1)
	) name20223 (
		_w26036_,
		_w26038_,
		_w26050_
	);
	LUT4 #(
		.INIT('h0001)
	) name20224 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26051_
	);
	LUT4 #(
		.INIT('hbbfe)
	) name20225 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26052_
	);
	LUT2 #(
		.INIT('h2)
	) name20226 (
		_w26037_,
		_w26052_,
		_w26053_
	);
	LUT3 #(
		.INIT('h80)
	) name20227 (
		_w26032_,
		_w26033_,
		_w26034_,
		_w26054_
	);
	LUT2 #(
		.INIT('h8)
	) name20228 (
		_w26050_,
		_w26054_,
		_w26055_
	);
	LUT3 #(
		.INIT('h31)
	) name20229 (
		_w26033_,
		_w26037_,
		_w26038_,
		_w26056_
	);
	LUT3 #(
		.INIT('h0d)
	) name20230 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26057_
	);
	LUT3 #(
		.INIT('h8a)
	) name20231 (
		_w26032_,
		_w26033_,
		_w26038_,
		_w26058_
	);
	LUT3 #(
		.INIT('h40)
	) name20232 (
		_w26057_,
		_w26056_,
		_w26058_,
		_w26059_
	);
	LUT4 #(
		.INIT('h0001)
	) name20233 (
		_w26055_,
		_w26053_,
		_w26059_,
		_w26049_,
		_w26060_
	);
	LUT3 #(
		.INIT('h65)
	) name20234 (
		\u0_L12_reg[6]/NET0131 ,
		_w26046_,
		_w26060_,
		_w26061_
	);
	LUT4 #(
		.INIT('h8448)
	) name20235 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w26062_
	);
	LUT4 #(
		.INIT('h1030)
	) name20236 (
		_w25527_,
		_w25529_,
		_w25526_,
		_w25528_,
		_w26063_
	);
	LUT4 #(
		.INIT('h0222)
	) name20237 (
		_w25541_,
		_w25621_,
		_w25615_,
		_w26063_,
		_w26064_
	);
	LUT4 #(
		.INIT('h2330)
	) name20238 (
		_w25527_,
		_w25526_,
		_w25528_,
		_w25530_,
		_w26065_
	);
	LUT4 #(
		.INIT('hc40c)
	) name20239 (
		_w25529_,
		_w25526_,
		_w25528_,
		_w25530_,
		_w26066_
	);
	LUT3 #(
		.INIT('h23)
	) name20240 (
		_w25624_,
		_w26065_,
		_w26066_,
		_w26067_
	);
	LUT4 #(
		.INIT('h0084)
	) name20241 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w26068_
	);
	LUT4 #(
		.INIT('h2000)
	) name20242 (
		_w25527_,
		_w25529_,
		_w25528_,
		_w25530_,
		_w26069_
	);
	LUT3 #(
		.INIT('h01)
	) name20243 (
		_w25541_,
		_w26068_,
		_w26069_,
		_w26070_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name20244 (
		_w26062_,
		_w26064_,
		_w26067_,
		_w26070_,
		_w26071_
	);
	LUT3 #(
		.INIT('h40)
	) name20245 (
		_w25526_,
		_w25528_,
		_w25530_,
		_w26072_
	);
	LUT2 #(
		.INIT('h4)
	) name20246 (
		_w25537_,
		_w26072_,
		_w26073_
	);
	LUT3 #(
		.INIT('h56)
	) name20247 (
		\u0_L12_reg[9]/NET0131 ,
		_w26071_,
		_w26073_,
		_w26074_
	);
	LUT4 #(
		.INIT('ha1e6)
	) name20248 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w26075_
	);
	LUT2 #(
		.INIT('h1)
	) name20249 (
		_w25586_,
		_w26075_,
		_w26076_
	);
	LUT3 #(
		.INIT('h21)
	) name20250 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w26077_
	);
	LUT4 #(
		.INIT('h2120)
	) name20251 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w26078_
	);
	LUT4 #(
		.INIT('h4880)
	) name20252 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w26079_
	);
	LUT4 #(
		.INIT('h040c)
	) name20253 (
		_w25586_,
		_w25596_,
		_w26079_,
		_w26078_,
		_w26080_
	);
	LUT4 #(
		.INIT('h4800)
	) name20254 (
		_w25588_,
		_w25590_,
		_w25589_,
		_w25587_,
		_w26081_
	);
	LUT4 #(
		.INIT('h5551)
	) name20255 (
		_w25596_,
		_w26007_,
		_w26077_,
		_w26081_,
		_w26082_
	);
	LUT3 #(
		.INIT('h0b)
	) name20256 (
		_w26076_,
		_w26080_,
		_w26082_,
		_w26083_
	);
	LUT2 #(
		.INIT('h4)
	) name20257 (
		_w25586_,
		_w26079_,
		_w26084_
	);
	LUT2 #(
		.INIT('h4)
	) name20258 (
		_w25586_,
		_w25596_,
		_w26085_
	);
	LUT4 #(
		.INIT('h00dc)
	) name20259 (
		_w25586_,
		_w25591_,
		_w26078_,
		_w26085_,
		_w26086_
	);
	LUT2 #(
		.INIT('h1)
	) name20260 (
		_w26084_,
		_w26086_,
		_w26087_
	);
	LUT3 #(
		.INIT('h65)
	) name20261 (
		\u0_L12_reg[7]/NET0131 ,
		_w26083_,
		_w26087_,
		_w26088_
	);
	LUT2 #(
		.INIT('h8)
	) name20262 (
		_w26036_,
		_w26038_,
		_w26089_
	);
	LUT3 #(
		.INIT('h80)
	) name20263 (
		_w26033_,
		_w26036_,
		_w26038_,
		_w26090_
	);
	LUT4 #(
		.INIT('h669b)
	) name20264 (
		_w26033_,
		_w26036_,
		_w26037_,
		_w26038_,
		_w26091_
	);
	LUT2 #(
		.INIT('h1)
	) name20265 (
		_w26034_,
		_w26091_,
		_w26092_
	);
	LUT4 #(
		.INIT('h0006)
	) name20266 (
		_w26034_,
		_w26036_,
		_w26037_,
		_w26038_,
		_w26093_
	);
	LUT4 #(
		.INIT('h0800)
	) name20267 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26094_
	);
	LUT3 #(
		.INIT('h02)
	) name20268 (
		_w26032_,
		_w26094_,
		_w26093_,
		_w26095_
	);
	LUT4 #(
		.INIT('h5afc)
	) name20269 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26096_
	);
	LUT2 #(
		.INIT('h1)
	) name20270 (
		_w26037_,
		_w26096_,
		_w26097_
	);
	LUT4 #(
		.INIT('h6080)
	) name20271 (
		_w26033_,
		_w26036_,
		_w26037_,
		_w26038_,
		_w26098_
	);
	LUT3 #(
		.INIT('h01)
	) name20272 (
		_w26032_,
		_w26051_,
		_w26098_,
		_w26099_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name20273 (
		_w26092_,
		_w26095_,
		_w26097_,
		_w26099_,
		_w26100_
	);
	LUT4 #(
		.INIT('h0040)
	) name20274 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26037_,
		_w26101_
	);
	LUT4 #(
		.INIT('hff7b)
	) name20275 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26102_
	);
	LUT3 #(
		.INIT('h31)
	) name20276 (
		_w26037_,
		_w26101_,
		_w26102_,
		_w26103_
	);
	LUT3 #(
		.INIT('h65)
	) name20277 (
		\u0_L12_reg[16]/NET0131 ,
		_w26100_,
		_w26103_,
		_w26104_
	);
	LUT4 #(
		.INIT('h0040)
	) name20278 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26105_
	);
	LUT4 #(
		.INIT('hbcb1)
	) name20279 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26106_
	);
	LUT4 #(
		.INIT('h5054)
	) name20280 (
		_w26032_,
		_w26037_,
		_w26105_,
		_w26106_,
		_w26107_
	);
	LUT3 #(
		.INIT('h8c)
	) name20281 (
		_w26036_,
		_w26037_,
		_w26038_,
		_w26108_
	);
	LUT3 #(
		.INIT('h37)
	) name20282 (
		_w26039_,
		_w26042_,
		_w26108_,
		_w26109_
	);
	LUT4 #(
		.INIT('h737f)
	) name20283 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26110_
	);
	LUT3 #(
		.INIT('hb1)
	) name20284 (
		_w26037_,
		_w26043_,
		_w26110_,
		_w26111_
	);
	LUT3 #(
		.INIT('h2a)
	) name20285 (
		_w26032_,
		_w26109_,
		_w26111_,
		_w26112_
	);
	LUT4 #(
		.INIT('h1001)
	) name20286 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26113_
	);
	LUT4 #(
		.INIT('he35e)
	) name20287 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26114_
	);
	LUT2 #(
		.INIT('h1)
	) name20288 (
		_w26032_,
		_w26037_,
		_w26115_
	);
	LUT2 #(
		.INIT('h4)
	) name20289 (
		_w26114_,
		_w26115_,
		_w26116_
	);
	LUT4 #(
		.INIT('h0010)
	) name20290 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26117_
	);
	LUT4 #(
		.INIT('hfdef)
	) name20291 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26118_
	);
	LUT4 #(
		.INIT('hdf13)
	) name20292 (
		_w26034_,
		_w26037_,
		_w26090_,
		_w26118_,
		_w26119_
	);
	LUT2 #(
		.INIT('h4)
	) name20293 (
		_w26116_,
		_w26119_,
		_w26120_
	);
	LUT4 #(
		.INIT('h5655)
	) name20294 (
		\u0_L12_reg[24]/NET0131 ,
		_w26112_,
		_w26107_,
		_w26120_,
		_w26121_
	);
	LUT4 #(
		.INIT('h3f35)
	) name20295 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26122_
	);
	LUT3 #(
		.INIT('h31)
	) name20296 (
		_w26032_,
		_w26037_,
		_w26122_,
		_w26123_
	);
	LUT4 #(
		.INIT('he0d0)
	) name20297 (
		_w26034_,
		_w26036_,
		_w26037_,
		_w26038_,
		_w26124_
	);
	LUT4 #(
		.INIT('h4000)
	) name20298 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26125_
	);
	LUT4 #(
		.INIT('h0075)
	) name20299 (
		_w26032_,
		_w26117_,
		_w26124_,
		_w26125_,
		_w26126_
	);
	LUT2 #(
		.INIT('h1)
	) name20300 (
		_w26123_,
		_w26126_,
		_w26127_
	);
	LUT4 #(
		.INIT('h3f9d)
	) name20301 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26128_
	);
	LUT2 #(
		.INIT('h2)
	) name20302 (
		_w26037_,
		_w26128_,
		_w26129_
	);
	LUT4 #(
		.INIT('h0400)
	) name20303 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26038_,
		_w26130_
	);
	LUT3 #(
		.INIT('h3a)
	) name20304 (
		_w26033_,
		_w26034_,
		_w26036_,
		_w26131_
	);
	LUT4 #(
		.INIT('h0013)
	) name20305 (
		_w26056_,
		_w26113_,
		_w26131_,
		_w26130_,
		_w26132_
	);
	LUT4 #(
		.INIT('h0008)
	) name20306 (
		_w26033_,
		_w26034_,
		_w26037_,
		_w26038_,
		_w26133_
	);
	LUT3 #(
		.INIT('h0d)
	) name20307 (
		_w26054_,
		_w26089_,
		_w26133_,
		_w26134_
	);
	LUT4 #(
		.INIT('hba00)
	) name20308 (
		_w26032_,
		_w26129_,
		_w26132_,
		_w26134_,
		_w26135_
	);
	LUT3 #(
		.INIT('h9a)
	) name20309 (
		\u0_L12_reg[30]/NET0131 ,
		_w26127_,
		_w26135_,
		_w26136_
	);
	LUT4 #(
		.INIT('hfd75)
	) name20310 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w26137_
	);
	LUT2 #(
		.INIT('h1)
	) name20311 (
		_w25714_,
		_w26137_,
		_w26138_
	);
	LUT4 #(
		.INIT('h0a20)
	) name20312 (
		_w25714_,
		_w25716_,
		_w25717_,
		_w25715_,
		_w26139_
	);
	LUT3 #(
		.INIT('h02)
	) name20313 (
		_w25713_,
		_w25733_,
		_w26139_,
		_w26140_
	);
	LUT2 #(
		.INIT('h4)
	) name20314 (
		_w26138_,
		_w26140_,
		_w26141_
	);
	LUT4 #(
		.INIT('h1003)
	) name20315 (
		_w25714_,
		_w25716_,
		_w25715_,
		_w25718_,
		_w26142_
	);
	LUT3 #(
		.INIT('h01)
	) name20316 (
		_w25713_,
		_w25808_,
		_w25792_,
		_w26143_
	);
	LUT4 #(
		.INIT('h8000)
	) name20317 (
		_w25714_,
		_w25716_,
		_w25717_,
		_w25715_,
		_w26144_
	);
	LUT2 #(
		.INIT('h1)
	) name20318 (
		_w25722_,
		_w26144_,
		_w26145_
	);
	LUT3 #(
		.INIT('h40)
	) name20319 (
		_w26142_,
		_w26143_,
		_w26145_,
		_w26146_
	);
	LUT4 #(
		.INIT('h1000)
	) name20320 (
		_w25714_,
		_w25716_,
		_w25717_,
		_w25715_,
		_w26147_
	);
	LUT4 #(
		.INIT('h77ef)
	) name20321 (
		_w25716_,
		_w25717_,
		_w25715_,
		_w25718_,
		_w26148_
	);
	LUT3 #(
		.INIT('h31)
	) name20322 (
		_w25714_,
		_w26147_,
		_w26148_,
		_w26149_
	);
	LUT4 #(
		.INIT('ha955)
	) name20323 (
		\u0_L12_reg[18]/NET0131 ,
		_w26141_,
		_w26146_,
		_w26149_,
		_w26150_
	);
	LUT4 #(
		.INIT('hc963)
	) name20324 (
		decrypt_pad,
		\u0_R11_reg[28]/NET0131 ,
		\u0_uk_K_r11_reg[0]/NET0131 ,
		\u0_uk_K_r11_reg[22]/NET0131 ,
		_w26151_
	);
	LUT4 #(
		.INIT('hc693)
	) name20325 (
		decrypt_pad,
		\u0_R11_reg[26]/NET0131 ,
		\u0_uk_K_r11_reg[2]/NET0131 ,
		\u0_uk_K_r11_reg[35]/NET0131 ,
		_w26152_
	);
	LUT4 #(
		.INIT('hc693)
	) name20326 (
		decrypt_pad,
		\u0_R11_reg[29]/NET0131 ,
		\u0_uk_K_r11_reg[14]/NET0131 ,
		\u0_uk_K_r11_reg[23]/NET0131 ,
		_w26153_
	);
	LUT4 #(
		.INIT('hc693)
	) name20327 (
		decrypt_pad,
		\u0_R11_reg[27]/NET0131 ,
		\u0_uk_K_r11_reg[35]/NET0131 ,
		\u0_uk_K_r11_reg[44]/NET0131 ,
		_w26154_
	);
	LUT4 #(
		.INIT('hc693)
	) name20328 (
		decrypt_pad,
		\u0_R11_reg[25]/NET0131 ,
		\u0_uk_K_r11_reg[45]/NET0131 ,
		\u0_uk_K_r11_reg[50]/NET0131 ,
		_w26155_
	);
	LUT4 #(
		.INIT('h0072)
	) name20329 (
		_w26152_,
		_w26155_,
		_w26153_,
		_w26154_,
		_w26156_
	);
	LUT4 #(
		.INIT('hc963)
	) name20330 (
		decrypt_pad,
		\u0_R11_reg[24]/NET0131 ,
		\u0_uk_K_r11_reg[15]/NET0131 ,
		\u0_uk_K_r11_reg[37]/NET0131 ,
		_w26157_
	);
	LUT4 #(
		.INIT('h04cc)
	) name20331 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26154_,
		_w26158_
	);
	LUT2 #(
		.INIT('h4)
	) name20332 (
		_w26156_,
		_w26158_,
		_w26159_
	);
	LUT4 #(
		.INIT('h0002)
	) name20333 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26160_
	);
	LUT2 #(
		.INIT('h6)
	) name20334 (
		_w26152_,
		_w26157_,
		_w26161_
	);
	LUT3 #(
		.INIT('h8c)
	) name20335 (
		_w26155_,
		_w26153_,
		_w26154_,
		_w26162_
	);
	LUT4 #(
		.INIT('h8caf)
	) name20336 (
		_w26154_,
		_w26161_,
		_w26160_,
		_w26162_,
		_w26163_
	);
	LUT3 #(
		.INIT('h45)
	) name20337 (
		_w26151_,
		_w26159_,
		_w26163_,
		_w26164_
	);
	LUT4 #(
		.INIT('h0400)
	) name20338 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26165_
	);
	LUT4 #(
		.INIT('hcbff)
	) name20339 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26166_
	);
	LUT2 #(
		.INIT('h1)
	) name20340 (
		_w26154_,
		_w26166_,
		_w26167_
	);
	LUT2 #(
		.INIT('h6)
	) name20341 (
		_w26152_,
		_w26155_,
		_w26168_
	);
	LUT4 #(
		.INIT('hc800)
	) name20342 (
		_w26152_,
		_w26157_,
		_w26153_,
		_w26154_,
		_w26169_
	);
	LUT2 #(
		.INIT('h4)
	) name20343 (
		_w26157_,
		_w26153_,
		_w26170_
	);
	LUT4 #(
		.INIT('h0200)
	) name20344 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26171_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name20345 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26172_
	);
	LUT3 #(
		.INIT('h70)
	) name20346 (
		_w26168_,
		_w26169_,
		_w26172_,
		_w26173_
	);
	LUT4 #(
		.INIT('h0020)
	) name20347 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26174_
	);
	LUT4 #(
		.INIT('hfddf)
	) name20348 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26175_
	);
	LUT4 #(
		.INIT('hfdd3)
	) name20349 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26176_
	);
	LUT4 #(
		.INIT('h0090)
	) name20350 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26154_,
		_w26177_
	);
	LUT4 #(
		.INIT('h0100)
	) name20351 (
		_w26152_,
		_w26155_,
		_w26153_,
		_w26154_,
		_w26178_
	);
	LUT4 #(
		.INIT('h0031)
	) name20352 (
		_w26154_,
		_w26177_,
		_w26176_,
		_w26178_,
		_w26179_
	);
	LUT4 #(
		.INIT('h7500)
	) name20353 (
		_w26151_,
		_w26167_,
		_w26173_,
		_w26179_,
		_w26180_
	);
	LUT3 #(
		.INIT('h65)
	) name20354 (
		\u0_L11_reg[22]/NET0131 ,
		_w26164_,
		_w26180_,
		_w26181_
	);
	LUT4 #(
		.INIT('hc693)
	) name20355 (
		decrypt_pad,
		\u0_R11_reg[3]/NET0131 ,
		\u0_uk_K_r11_reg[13]/NET0131 ,
		\u0_uk_K_r11_reg[18]/NET0131 ,
		_w26182_
	);
	LUT4 #(
		.INIT('hc693)
	) name20356 (
		decrypt_pad,
		\u0_R11_reg[5]/NET0131 ,
		\u0_uk_K_r11_reg[19]/NET0131 ,
		\u0_uk_K_r11_reg[24]/NET0131 ,
		_w26183_
	);
	LUT4 #(
		.INIT('hc963)
	) name20357 (
		decrypt_pad,
		\u0_R11_reg[1]/NET0131 ,
		\u0_uk_K_r11_reg[26]/NET0131 ,
		\u0_uk_K_r11_reg[46]/NET0131 ,
		_w26184_
	);
	LUT4 #(
		.INIT('hc963)
	) name20358 (
		decrypt_pad,
		\u0_R11_reg[2]/NET0131 ,
		\u0_uk_K_r11_reg[41]/NET0131 ,
		\u0_uk_K_r11_reg[4]/NET0131 ,
		_w26185_
	);
	LUT4 #(
		.INIT('hc693)
	) name20359 (
		decrypt_pad,
		\u0_R11_reg[32]/NET0131 ,
		\u0_uk_K_r11_reg[25]/NET0131 ,
		\u0_uk_K_r11_reg[5]/NET0131 ,
		_w26186_
	);
	LUT4 #(
		.INIT('hf3d1)
	) name20360 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26187_
	);
	LUT2 #(
		.INIT('h2)
	) name20361 (
		_w26182_,
		_w26187_,
		_w26188_
	);
	LUT4 #(
		.INIT('h500c)
	) name20362 (
		_w26182_,
		_w26185_,
		_w26184_,
		_w26186_,
		_w26189_
	);
	LUT2 #(
		.INIT('h2)
	) name20363 (
		_w26183_,
		_w26186_,
		_w26190_
	);
	LUT2 #(
		.INIT('h2)
	) name20364 (
		_w26182_,
		_w26185_,
		_w26191_
	);
	LUT3 #(
		.INIT('hd0)
	) name20365 (
		_w26182_,
		_w26185_,
		_w26184_,
		_w26192_
	);
	LUT4 #(
		.INIT('hc693)
	) name20366 (
		decrypt_pad,
		\u0_R11_reg[4]/NET0131 ,
		\u0_uk_K_r11_reg[48]/NET0131 ,
		\u0_uk_K_r11_reg[53]/P0001 ,
		_w26193_
	);
	LUT4 #(
		.INIT('h0100)
	) name20367 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26194_
	);
	LUT4 #(
		.INIT('h2202)
	) name20368 (
		_w26193_,
		_w26194_,
		_w26190_,
		_w26192_,
		_w26195_
	);
	LUT3 #(
		.INIT('h10)
	) name20369 (
		_w26188_,
		_w26189_,
		_w26195_,
		_w26196_
	);
	LUT4 #(
		.INIT('h73cf)
	) name20370 (
		_w26182_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26197_
	);
	LUT2 #(
		.INIT('h1)
	) name20371 (
		_w26185_,
		_w26197_,
		_w26198_
	);
	LUT2 #(
		.INIT('h9)
	) name20372 (
		_w26183_,
		_w26186_,
		_w26199_
	);
	LUT3 #(
		.INIT('h80)
	) name20373 (
		_w26182_,
		_w26185_,
		_w26184_,
		_w26200_
	);
	LUT3 #(
		.INIT('h45)
	) name20374 (
		_w26193_,
		_w26199_,
		_w26200_,
		_w26201_
	);
	LUT2 #(
		.INIT('h4)
	) name20375 (
		_w26198_,
		_w26201_,
		_w26202_
	);
	LUT4 #(
		.INIT('hfdae)
	) name20376 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26203_
	);
	LUT4 #(
		.INIT('h6fe7)
	) name20377 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26204_
	);
	LUT4 #(
		.INIT('h0155)
	) name20378 (
		_w26182_,
		_w26203_,
		_w26193_,
		_w26204_,
		_w26205_
	);
	LUT2 #(
		.INIT('h1)
	) name20379 (
		_w26183_,
		_w26184_,
		_w26206_
	);
	LUT3 #(
		.INIT('h08)
	) name20380 (
		_w26182_,
		_w26185_,
		_w26186_,
		_w26207_
	);
	LUT4 #(
		.INIT('h0200)
	) name20381 (
		_w26182_,
		_w26185_,
		_w26184_,
		_w26186_,
		_w26208_
	);
	LUT3 #(
		.INIT('h07)
	) name20382 (
		_w26206_,
		_w26207_,
		_w26208_,
		_w26209_
	);
	LUT2 #(
		.INIT('h4)
	) name20383 (
		_w26205_,
		_w26209_,
		_w26210_
	);
	LUT4 #(
		.INIT('ha955)
	) name20384 (
		\u0_L11_reg[31]/NET0131 ,
		_w26196_,
		_w26202_,
		_w26210_,
		_w26211_
	);
	LUT4 #(
		.INIT('hc693)
	) name20385 (
		decrypt_pad,
		\u0_R11_reg[24]/NET0131 ,
		\u0_uk_K_r11_reg[15]/NET0131 ,
		\u0_uk_K_r11_reg[52]/NET0131 ,
		_w26212_
	);
	LUT4 #(
		.INIT('hc693)
	) name20386 (
		decrypt_pad,
		\u0_R11_reg[22]/NET0131 ,
		\u0_uk_K_r11_reg[0]/NET0131 ,
		\u0_uk_K_r11_reg[9]/NET0131 ,
		_w26213_
	);
	LUT4 #(
		.INIT('hc963)
	) name20387 (
		decrypt_pad,
		\u0_R11_reg[21]/NET0131 ,
		\u0_uk_K_r11_reg[42]/NET0131 ,
		\u0_uk_K_r11_reg[9]/NET0131 ,
		_w26214_
	);
	LUT4 #(
		.INIT('hc963)
	) name20388 (
		decrypt_pad,
		\u0_R11_reg[20]/NET0131 ,
		\u0_uk_K_r11_reg[31]/NET0131 ,
		\u0_uk_K_r11_reg[49]/NET0131 ,
		_w26215_
	);
	LUT4 #(
		.INIT('hc693)
	) name20389 (
		decrypt_pad,
		\u0_R11_reg[25]/NET0131 ,
		\u0_uk_K_r11_reg[38]/NET0131 ,
		\u0_uk_K_r11_reg[43]/NET0131 ,
		_w26216_
	);
	LUT4 #(
		.INIT('ha808)
	) name20390 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26217_
	);
	LUT4 #(
		.INIT('hc963)
	) name20391 (
		decrypt_pad,
		\u0_R11_reg[23]/NET0131 ,
		\u0_uk_K_r11_reg[22]/NET0131 ,
		\u0_uk_K_r11_reg[44]/NET0131 ,
		_w26218_
	);
	LUT4 #(
		.INIT('h5155)
	) name20392 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26219_
	);
	LUT3 #(
		.INIT('h01)
	) name20393 (
		_w26218_,
		_w26219_,
		_w26217_,
		_w26220_
	);
	LUT2 #(
		.INIT('h1)
	) name20394 (
		_w26213_,
		_w26218_,
		_w26221_
	);
	LUT4 #(
		.INIT('h0400)
	) name20395 (
		_w26213_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26222_
	);
	LUT2 #(
		.INIT('h4)
	) name20396 (
		_w26214_,
		_w26222_,
		_w26223_
	);
	LUT4 #(
		.INIT('hc0d0)
	) name20397 (
		_w26213_,
		_w26214_,
		_w26218_,
		_w26216_,
		_w26224_
	);
	LUT4 #(
		.INIT('hfa3a)
	) name20398 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26225_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name20399 (
		_w26214_,
		_w26222_,
		_w26224_,
		_w26225_,
		_w26226_
	);
	LUT3 #(
		.INIT('h8a)
	) name20400 (
		_w26212_,
		_w26220_,
		_w26226_,
		_w26227_
	);
	LUT3 #(
		.INIT('hc4)
	) name20401 (
		_w26214_,
		_w26215_,
		_w26216_,
		_w26228_
	);
	LUT4 #(
		.INIT('h30b0)
	) name20402 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26229_
	);
	LUT4 #(
		.INIT('h080c)
	) name20403 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26230_
	);
	LUT3 #(
		.INIT('h01)
	) name20404 (
		_w26213_,
		_w26230_,
		_w26229_,
		_w26231_
	);
	LUT4 #(
		.INIT('h5440)
	) name20405 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26232_
	);
	LUT4 #(
		.INIT('haaa2)
	) name20406 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26218_,
		_w26233_
	);
	LUT3 #(
		.INIT('h0b)
	) name20407 (
		_w26232_,
		_w26233_,
		_w26212_,
		_w26234_
	);
	LUT3 #(
		.INIT('h10)
	) name20408 (
		_w26214_,
		_w26215_,
		_w26216_,
		_w26235_
	);
	LUT4 #(
		.INIT('he0f0)
	) name20409 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26236_
	);
	LUT4 #(
		.INIT('h0f07)
	) name20410 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26237_
	);
	LUT3 #(
		.INIT('h01)
	) name20411 (
		_w26213_,
		_w26237_,
		_w26236_,
		_w26238_
	);
	LUT3 #(
		.INIT('h01)
	) name20412 (
		_w26214_,
		_w26215_,
		_w26216_,
		_w26239_
	);
	LUT4 #(
		.INIT('h5f53)
	) name20413 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26240_
	);
	LUT3 #(
		.INIT('hc4)
	) name20414 (
		_w26213_,
		_w26218_,
		_w26216_,
		_w26241_
	);
	LUT4 #(
		.INIT('h7077)
	) name20415 (
		_w26221_,
		_w26239_,
		_w26240_,
		_w26241_,
		_w26242_
	);
	LUT4 #(
		.INIT('h0b00)
	) name20416 (
		_w26231_,
		_w26234_,
		_w26238_,
		_w26242_,
		_w26243_
	);
	LUT3 #(
		.INIT('h9a)
	) name20417 (
		\u0_L11_reg[11]/P0001 ,
		_w26227_,
		_w26243_,
		_w26244_
	);
	LUT4 #(
		.INIT('hc693)
	) name20418 (
		decrypt_pad,
		\u0_R11_reg[32]/NET0131 ,
		\u0_uk_K_r11_reg[42]/NET0131 ,
		\u0_uk_K_r11_reg[51]/NET0131 ,
		_w26245_
	);
	LUT4 #(
		.INIT('hc963)
	) name20419 (
		decrypt_pad,
		\u0_R11_reg[31]/P0001 ,
		\u0_uk_K_r11_reg[14]/NET0131 ,
		\u0_uk_K_r11_reg[36]/NET0131 ,
		_w26246_
	);
	LUT4 #(
		.INIT('hc963)
	) name20420 (
		decrypt_pad,
		\u0_R11_reg[30]/NET0131 ,
		\u0_uk_K_r11_reg[2]/NET0131 ,
		\u0_uk_K_r11_reg[52]/NET0131 ,
		_w26247_
	);
	LUT4 #(
		.INIT('hc963)
	) name20421 (
		decrypt_pad,
		\u0_R11_reg[29]/NET0131 ,
		\u0_uk_K_r11_reg[1]/NET0131 ,
		\u0_uk_K_r11_reg[23]/NET0131 ,
		_w26248_
	);
	LUT4 #(
		.INIT('hc963)
	) name20422 (
		decrypt_pad,
		\u0_R11_reg[28]/NET0131 ,
		\u0_uk_K_r11_reg[29]/NET0131 ,
		\u0_uk_K_r11_reg[51]/NET0131 ,
		_w26249_
	);
	LUT4 #(
		.INIT('hc963)
	) name20423 (
		decrypt_pad,
		\u0_R11_reg[1]/NET0131 ,
		\u0_uk_K_r11_reg[45]/NET0131 ,
		\u0_uk_K_r11_reg[8]/NET0131 ,
		_w26250_
	);
	LUT4 #(
		.INIT('ha6f3)
	) name20424 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26251_
	);
	LUT3 #(
		.INIT('h01)
	) name20425 (
		_w26247_,
		_w26248_,
		_w26249_,
		_w26252_
	);
	LUT4 #(
		.INIT('h0080)
	) name20426 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26253_
	);
	LUT4 #(
		.INIT('h0b01)
	) name20427 (
		_w26246_,
		_w26252_,
		_w26253_,
		_w26251_,
		_w26254_
	);
	LUT2 #(
		.INIT('h2)
	) name20428 (
		_w26245_,
		_w26254_,
		_w26255_
	);
	LUT2 #(
		.INIT('h1)
	) name20429 (
		_w26247_,
		_w26246_,
		_w26256_
	);
	LUT4 #(
		.INIT('h7b2a)
	) name20430 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26246_,
		_w26257_
	);
	LUT2 #(
		.INIT('h2)
	) name20431 (
		_w26249_,
		_w26257_,
		_w26258_
	);
	LUT4 #(
		.INIT('h0200)
	) name20432 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26259_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name20433 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26260_
	);
	LUT3 #(
		.INIT('h0b)
	) name20434 (
		_w26250_,
		_w26249_,
		_w26246_,
		_w26261_
	);
	LUT3 #(
		.INIT('hca)
	) name20435 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26262_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name20436 (
		_w26260_,
		_w26246_,
		_w26261_,
		_w26262_,
		_w26263_
	);
	LUT3 #(
		.INIT('h0b)
	) name20437 (
		_w26258_,
		_w26263_,
		_w26245_,
		_w26264_
	);
	LUT4 #(
		.INIT('h0008)
	) name20438 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26265_
	);
	LUT4 #(
		.INIT('heff7)
	) name20439 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26266_
	);
	LUT4 #(
		.INIT('h0020)
	) name20440 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26267_
	);
	LUT4 #(
		.INIT('h0001)
	) name20441 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26268_
	);
	LUT4 #(
		.INIT('hefd6)
	) name20442 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26269_
	);
	LUT2 #(
		.INIT('h2)
	) name20443 (
		_w26246_,
		_w26269_,
		_w26270_
	);
	LUT3 #(
		.INIT('h40)
	) name20444 (
		_w26248_,
		_w26249_,
		_w26245_,
		_w26271_
	);
	LUT3 #(
		.INIT('h20)
	) name20445 (
		_w26248_,
		_w26250_,
		_w26249_,
		_w26272_
	);
	LUT4 #(
		.INIT('hcedf)
	) name20446 (
		_w26247_,
		_w26246_,
		_w26271_,
		_w26272_,
		_w26273_
	);
	LUT2 #(
		.INIT('h4)
	) name20447 (
		_w26270_,
		_w26273_,
		_w26274_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name20448 (
		\u0_L11_reg[5]/NET0131 ,
		_w26264_,
		_w26255_,
		_w26274_,
		_w26275_
	);
	LUT4 #(
		.INIT('hc693)
	) name20449 (
		decrypt_pad,
		\u0_R11_reg[15]/NET0131 ,
		\u0_uk_K_r11_reg[10]/NET0131 ,
		\u0_uk_K_r11_reg[47]/NET0131 ,
		_w26276_
	);
	LUT4 #(
		.INIT('hc963)
	) name20450 (
		decrypt_pad,
		\u0_R11_reg[13]/NET0131 ,
		\u0_uk_K_r11_reg[13]/NET0131 ,
		\u0_uk_K_r11_reg[33]/NET0131 ,
		_w26277_
	);
	LUT4 #(
		.INIT('hc963)
	) name20451 (
		decrypt_pad,
		\u0_R11_reg[17]/NET0131 ,
		\u0_uk_K_r11_reg[3]/NET0131 ,
		\u0_uk_K_r11_reg[55]/NET0131 ,
		_w26278_
	);
	LUT4 #(
		.INIT('hc693)
	) name20452 (
		decrypt_pad,
		\u0_R11_reg[14]/NET0131 ,
		\u0_uk_K_r11_reg[34]/NET0131 ,
		\u0_uk_K_r11_reg[39]/NET0131 ,
		_w26279_
	);
	LUT4 #(
		.INIT('hc963)
	) name20453 (
		decrypt_pad,
		\u0_R11_reg[12]/NET0131 ,
		\u0_uk_K_r11_reg[19]/NET0131 ,
		\u0_uk_K_r11_reg[39]/NET0131 ,
		_w26280_
	);
	LUT3 #(
		.INIT('h20)
	) name20454 (
		_w26279_,
		_w26278_,
		_w26280_,
		_w26281_
	);
	LUT4 #(
		.INIT('ha3af)
	) name20455 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26282_
	);
	LUT2 #(
		.INIT('h1)
	) name20456 (
		_w26276_,
		_w26282_,
		_w26283_
	);
	LUT4 #(
		.INIT('h0100)
	) name20457 (
		_w26277_,
		_w26278_,
		_w26280_,
		_w26276_,
		_w26284_
	);
	LUT4 #(
		.INIT('hc693)
	) name20458 (
		decrypt_pad,
		\u0_R11_reg[16]/NET0131 ,
		\u0_uk_K_r11_reg[18]/NET0131 ,
		\u0_uk_K_r11_reg[55]/NET0131 ,
		_w26285_
	);
	LUT2 #(
		.INIT('h4)
	) name20459 (
		_w26279_,
		_w26280_,
		_w26286_
	);
	LUT4 #(
		.INIT('h1000)
	) name20460 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26287_
	);
	LUT3 #(
		.INIT('h01)
	) name20461 (
		_w26285_,
		_w26287_,
		_w26284_,
		_w26288_
	);
	LUT2 #(
		.INIT('h8)
	) name20462 (
		_w26277_,
		_w26276_,
		_w26289_
	);
	LUT3 #(
		.INIT('h35)
	) name20463 (
		_w26279_,
		_w26278_,
		_w26280_,
		_w26290_
	);
	LUT4 #(
		.INIT('hfff6)
	) name20464 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26291_
	);
	LUT3 #(
		.INIT('hd0)
	) name20465 (
		_w26289_,
		_w26290_,
		_w26291_,
		_w26292_
	);
	LUT3 #(
		.INIT('h40)
	) name20466 (
		_w26283_,
		_w26288_,
		_w26292_,
		_w26293_
	);
	LUT3 #(
		.INIT('h01)
	) name20467 (
		_w26277_,
		_w26280_,
		_w26276_,
		_w26294_
	);
	LUT4 #(
		.INIT('h0001)
	) name20468 (
		_w26277_,
		_w26278_,
		_w26280_,
		_w26276_,
		_w26295_
	);
	LUT2 #(
		.INIT('h8)
	) name20469 (
		_w26279_,
		_w26295_,
		_w26296_
	);
	LUT2 #(
		.INIT('h8)
	) name20470 (
		_w26277_,
		_w26280_,
		_w26297_
	);
	LUT3 #(
		.INIT('h47)
	) name20471 (
		_w26279_,
		_w26278_,
		_w26276_,
		_w26298_
	);
	LUT3 #(
		.INIT('ha2)
	) name20472 (
		_w26285_,
		_w26297_,
		_w26298_,
		_w26299_
	);
	LUT2 #(
		.INIT('h2)
	) name20473 (
		_w26278_,
		_w26280_,
		_w26300_
	);
	LUT2 #(
		.INIT('h4)
	) name20474 (
		_w26277_,
		_w26276_,
		_w26301_
	);
	LUT3 #(
		.INIT('h8d)
	) name20475 (
		_w26277_,
		_w26279_,
		_w26276_,
		_w26302_
	);
	LUT2 #(
		.INIT('h6)
	) name20476 (
		_w26277_,
		_w26280_,
		_w26303_
	);
	LUT4 #(
		.INIT('h0012)
	) name20477 (
		_w26277_,
		_w26279_,
		_w26280_,
		_w26276_,
		_w26304_
	);
	LUT3 #(
		.INIT('h0d)
	) name20478 (
		_w26300_,
		_w26302_,
		_w26304_,
		_w26305_
	);
	LUT3 #(
		.INIT('h40)
	) name20479 (
		_w26296_,
		_w26299_,
		_w26305_,
		_w26306_
	);
	LUT4 #(
		.INIT('h0220)
	) name20480 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26307_
	);
	LUT2 #(
		.INIT('h9)
	) name20481 (
		_w26278_,
		_w26276_,
		_w26308_
	);
	LUT2 #(
		.INIT('h9)
	) name20482 (
		_w26279_,
		_w26280_,
		_w26309_
	);
	LUT4 #(
		.INIT('h2100)
	) name20483 (
		_w26279_,
		_w26278_,
		_w26280_,
		_w26276_,
		_w26310_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name20484 (
		_w26277_,
		_w26307_,
		_w26308_,
		_w26310_,
		_w26311_
	);
	LUT4 #(
		.INIT('ha955)
	) name20485 (
		\u0_L11_reg[20]/NET0131 ,
		_w26293_,
		_w26306_,
		_w26311_,
		_w26312_
	);
	LUT2 #(
		.INIT('h2)
	) name20486 (
		_w26277_,
		_w26276_,
		_w26313_
	);
	LUT3 #(
		.INIT('h4d)
	) name20487 (
		_w26279_,
		_w26278_,
		_w26280_,
		_w26314_
	);
	LUT2 #(
		.INIT('h8)
	) name20488 (
		_w26313_,
		_w26314_,
		_w26315_
	);
	LUT4 #(
		.INIT('h0844)
	) name20489 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26316_
	);
	LUT3 #(
		.INIT('h23)
	) name20490 (
		_w26279_,
		_w26278_,
		_w26280_,
		_w26317_
	);
	LUT3 #(
		.INIT('h31)
	) name20491 (
		_w26301_,
		_w26316_,
		_w26317_,
		_w26318_
	);
	LUT3 #(
		.INIT('h8a)
	) name20492 (
		_w26285_,
		_w26315_,
		_w26318_,
		_w26319_
	);
	LUT3 #(
		.INIT('ha8)
	) name20493 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26320_
	);
	LUT2 #(
		.INIT('h2)
	) name20494 (
		_w26310_,
		_w26320_,
		_w26321_
	);
	LUT3 #(
		.INIT('hac)
	) name20495 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26322_
	);
	LUT2 #(
		.INIT('h2)
	) name20496 (
		_w26280_,
		_w26276_,
		_w26323_
	);
	LUT4 #(
		.INIT('h7ddf)
	) name20497 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26324_
	);
	LUT3 #(
		.INIT('hb0)
	) name20498 (
		_w26322_,
		_w26323_,
		_w26324_,
		_w26325_
	);
	LUT3 #(
		.INIT('h45)
	) name20499 (
		_w26285_,
		_w26321_,
		_w26325_,
		_w26326_
	);
	LUT4 #(
		.INIT('h8040)
	) name20500 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26327_
	);
	LUT4 #(
		.INIT('h7fb7)
	) name20501 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26328_
	);
	LUT2 #(
		.INIT('h2)
	) name20502 (
		_w26276_,
		_w26328_,
		_w26329_
	);
	LUT4 #(
		.INIT('h135f)
	) name20503 (
		_w26279_,
		_w26281_,
		_w26295_,
		_w26313_,
		_w26330_
	);
	LUT2 #(
		.INIT('h4)
	) name20504 (
		_w26329_,
		_w26330_,
		_w26331_
	);
	LUT4 #(
		.INIT('h5655)
	) name20505 (
		\u0_L11_reg[1]/NET0131 ,
		_w26326_,
		_w26319_,
		_w26331_,
		_w26332_
	);
	LUT4 #(
		.INIT('h0020)
	) name20506 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26333_
	);
	LUT4 #(
		.INIT('hf2df)
	) name20507 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26334_
	);
	LUT2 #(
		.INIT('h1)
	) name20508 (
		_w26276_,
		_w26334_,
		_w26335_
	);
	LUT4 #(
		.INIT('h4300)
	) name20509 (
		_w26279_,
		_w26278_,
		_w26280_,
		_w26276_,
		_w26336_
	);
	LUT3 #(
		.INIT('h13)
	) name20510 (
		_w26303_,
		_w26327_,
		_w26336_,
		_w26337_
	);
	LUT3 #(
		.INIT('h8a)
	) name20511 (
		_w26285_,
		_w26335_,
		_w26337_,
		_w26338_
	);
	LUT2 #(
		.INIT('h4)
	) name20512 (
		_w26279_,
		_w26278_,
		_w26339_
	);
	LUT4 #(
		.INIT('h0400)
	) name20513 (
		_w26279_,
		_w26278_,
		_w26280_,
		_w26276_,
		_w26340_
	);
	LUT2 #(
		.INIT('h2)
	) name20514 (
		_w26291_,
		_w26340_,
		_w26341_
	);
	LUT3 #(
		.INIT('h51)
	) name20515 (
		_w26277_,
		_w26278_,
		_w26276_,
		_w26342_
	);
	LUT2 #(
		.INIT('h2)
	) name20516 (
		_w26286_,
		_w26342_,
		_w26343_
	);
	LUT3 #(
		.INIT('h40)
	) name20517 (
		_w26277_,
		_w26280_,
		_w26276_,
		_w26344_
	);
	LUT3 #(
		.INIT('h45)
	) name20518 (
		_w26295_,
		_w26339_,
		_w26344_,
		_w26345_
	);
	LUT4 #(
		.INIT('h4555)
	) name20519 (
		_w26285_,
		_w26343_,
		_w26341_,
		_w26345_,
		_w26346_
	);
	LUT4 #(
		.INIT('h7fbe)
	) name20520 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w26347_
	);
	LUT4 #(
		.INIT('h8a00)
	) name20521 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26276_,
		_w26348_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name20522 (
		_w26276_,
		_w26309_,
		_w26347_,
		_w26348_,
		_w26349_
	);
	LUT4 #(
		.INIT('h5655)
	) name20523 (
		\u0_L11_reg[10]/NET0131 ,
		_w26346_,
		_w26338_,
		_w26349_,
		_w26350_
	);
	LUT4 #(
		.INIT('hc693)
	) name20524 (
		decrypt_pad,
		\u0_R11_reg[8]/NET0131 ,
		\u0_uk_K_r11_reg[17]/NET0131 ,
		\u0_uk_K_r11_reg[54]/NET0131 ,
		_w26351_
	);
	LUT4 #(
		.INIT('hc693)
	) name20525 (
		decrypt_pad,
		\u0_R11_reg[7]/NET0131 ,
		\u0_uk_K_r11_reg[26]/NET0131 ,
		\u0_uk_K_r11_reg[6]/NET0131 ,
		_w26352_
	);
	LUT4 #(
		.INIT('hc963)
	) name20526 (
		decrypt_pad,
		\u0_R11_reg[6]/NET0131 ,
		\u0_uk_K_r11_reg[12]/NET0131 ,
		\u0_uk_K_r11_reg[32]/NET0131 ,
		_w26353_
	);
	LUT4 #(
		.INIT('hc963)
	) name20527 (
		decrypt_pad,
		\u0_R11_reg[4]/NET0131 ,
		\u0_uk_K_r11_reg[10]/NET0131 ,
		\u0_uk_K_r11_reg[5]/NET0131 ,
		_w26354_
	);
	LUT4 #(
		.INIT('hc693)
	) name20528 (
		decrypt_pad,
		\u0_R11_reg[5]/NET0131 ,
		\u0_uk_K_r11_reg[41]/NET0131 ,
		\u0_uk_K_r11_reg[46]/NET0131 ,
		_w26355_
	);
	LUT4 #(
		.INIT('hc963)
	) name20529 (
		decrypt_pad,
		\u0_R11_reg[9]/NET0131 ,
		\u0_uk_K_r11_reg[34]/NET0131 ,
		\u0_uk_K_r11_reg[54]/NET0131 ,
		_w26356_
	);
	LUT4 #(
		.INIT('h3fc7)
	) name20530 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26357_
	);
	LUT2 #(
		.INIT('h2)
	) name20531 (
		_w26352_,
		_w26357_,
		_w26358_
	);
	LUT3 #(
		.INIT('h20)
	) name20532 (
		_w26355_,
		_w26354_,
		_w26356_,
		_w26359_
	);
	LUT4 #(
		.INIT('hf3fa)
	) name20533 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26360_
	);
	LUT2 #(
		.INIT('h1)
	) name20534 (
		_w26352_,
		_w26360_,
		_w26361_
	);
	LUT2 #(
		.INIT('h8)
	) name20535 (
		_w26354_,
		_w26352_,
		_w26362_
	);
	LUT4 #(
		.INIT('h33bf)
	) name20536 (
		_w26355_,
		_w26354_,
		_w26356_,
		_w26352_,
		_w26363_
	);
	LUT4 #(
		.INIT('h0200)
	) name20537 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26364_
	);
	LUT3 #(
		.INIT('h0e)
	) name20538 (
		_w26353_,
		_w26363_,
		_w26364_,
		_w26365_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name20539 (
		_w26351_,
		_w26361_,
		_w26358_,
		_w26365_,
		_w26366_
	);
	LUT4 #(
		.INIT('hfd7d)
	) name20540 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26367_
	);
	LUT2 #(
		.INIT('h1)
	) name20541 (
		_w26367_,
		_w26352_,
		_w26368_
	);
	LUT2 #(
		.INIT('h2)
	) name20542 (
		_w26352_,
		_w26360_,
		_w26369_
	);
	LUT3 #(
		.INIT('hd0)
	) name20543 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26370_
	);
	LUT4 #(
		.INIT('h0c2f)
	) name20544 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26371_
	);
	LUT4 #(
		.INIT('h00bf)
	) name20545 (
		_w26355_,
		_w26354_,
		_w26356_,
		_w26352_,
		_w26372_
	);
	LUT4 #(
		.INIT('hdf7d)
	) name20546 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26373_
	);
	LUT3 #(
		.INIT('hb0)
	) name20547 (
		_w26371_,
		_w26372_,
		_w26373_,
		_w26374_
	);
	LUT4 #(
		.INIT('h4544)
	) name20548 (
		_w26368_,
		_w26351_,
		_w26369_,
		_w26374_,
		_w26375_
	);
	LUT3 #(
		.INIT('h65)
	) name20549 (
		\u0_L11_reg[28]/NET0131 ,
		_w26366_,
		_w26375_,
		_w26376_
	);
	LUT4 #(
		.INIT('hff10)
	) name20550 (
		_w26247_,
		_w26250_,
		_w26249_,
		_w26246_,
		_w26377_
	);
	LUT4 #(
		.INIT('h2000)
	) name20551 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26378_
	);
	LUT4 #(
		.INIT('h7f00)
	) name20552 (
		_w26247_,
		_w26248_,
		_w26249_,
		_w26246_,
		_w26379_
	);
	LUT4 #(
		.INIT('hef2f)
	) name20553 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26380_
	);
	LUT4 #(
		.INIT('h0eee)
	) name20554 (
		_w26377_,
		_w26378_,
		_w26379_,
		_w26380_,
		_w26381_
	);
	LUT4 #(
		.INIT('h0802)
	) name20555 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26382_
	);
	LUT4 #(
		.INIT('h0010)
	) name20556 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26383_
	);
	LUT3 #(
		.INIT('h02)
	) name20557 (
		_w26245_,
		_w26383_,
		_w26382_,
		_w26384_
	);
	LUT2 #(
		.INIT('h4)
	) name20558 (
		_w26381_,
		_w26384_,
		_w26385_
	);
	LUT4 #(
		.INIT('h0040)
	) name20559 (
		_w26247_,
		_w26250_,
		_w26249_,
		_w26246_,
		_w26386_
	);
	LUT3 #(
		.INIT('h08)
	) name20560 (
		_w26247_,
		_w26248_,
		_w26249_,
		_w26387_
	);
	LUT4 #(
		.INIT('h0001)
	) name20561 (
		_w26259_,
		_w26245_,
		_w26386_,
		_w26387_,
		_w26388_
	);
	LUT4 #(
		.INIT('h0002)
	) name20562 (
		_w26248_,
		_w26250_,
		_w26249_,
		_w26246_,
		_w26389_
	);
	LUT2 #(
		.INIT('h1)
	) name20563 (
		_w26268_,
		_w26389_,
		_w26390_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name20564 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26391_
	);
	LUT3 #(
		.INIT('h40)
	) name20565 (
		_w26247_,
		_w26248_,
		_w26249_,
		_w26392_
	);
	LUT4 #(
		.INIT('hbfb5)
	) name20566 (
		_w26247_,
		_w26248_,
		_w26249_,
		_w26246_,
		_w26393_
	);
	LUT4 #(
		.INIT('hf351)
	) name20567 (
		_w26250_,
		_w26246_,
		_w26391_,
		_w26393_,
		_w26394_
	);
	LUT3 #(
		.INIT('h80)
	) name20568 (
		_w26388_,
		_w26390_,
		_w26394_,
		_w26395_
	);
	LUT4 #(
		.INIT('h0100)
	) name20569 (
		_w26247_,
		_w26248_,
		_w26249_,
		_w26246_,
		_w26396_
	);
	LUT3 #(
		.INIT('h13)
	) name20570 (
		_w26248_,
		_w26396_,
		_w26386_,
		_w26397_
	);
	LUT4 #(
		.INIT('ha955)
	) name20571 (
		\u0_L11_reg[21]/NET0131 ,
		_w26385_,
		_w26395_,
		_w26397_,
		_w26398_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name20572 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26399_
	);
	LUT2 #(
		.INIT('h2)
	) name20573 (
		_w26154_,
		_w26399_,
		_w26400_
	);
	LUT3 #(
		.INIT('h02)
	) name20574 (
		_w26151_,
		_w26165_,
		_w26174_,
		_w26401_
	);
	LUT4 #(
		.INIT('h1008)
	) name20575 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26402_
	);
	LUT3 #(
		.INIT('h0d)
	) name20576 (
		_w26171_,
		_w26154_,
		_w26402_,
		_w26403_
	);
	LUT3 #(
		.INIT('h40)
	) name20577 (
		_w26400_,
		_w26401_,
		_w26403_,
		_w26404_
	);
	LUT4 #(
		.INIT('h0014)
	) name20578 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26405_
	);
	LUT4 #(
		.INIT('h0800)
	) name20579 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26406_
	);
	LUT3 #(
		.INIT('h47)
	) name20580 (
		_w26152_,
		_w26155_,
		_w26154_,
		_w26407_
	);
	LUT4 #(
		.INIT('h0031)
	) name20581 (
		_w26170_,
		_w26406_,
		_w26407_,
		_w26405_,
		_w26408_
	);
	LUT4 #(
		.INIT('h0770)
	) name20582 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26409_
	);
	LUT4 #(
		.INIT('h0504)
	) name20583 (
		_w26151_,
		_w26154_,
		_w26160_,
		_w26409_,
		_w26410_
	);
	LUT2 #(
		.INIT('h8)
	) name20584 (
		_w26408_,
		_w26410_,
		_w26411_
	);
	LUT3 #(
		.INIT('ha9)
	) name20585 (
		\u0_L11_reg[12]/NET0131 ,
		_w26404_,
		_w26411_,
		_w26412_
	);
	LUT4 #(
		.INIT('hf3ec)
	) name20586 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26413_
	);
	LUT3 #(
		.INIT('h6f)
	) name20587 (
		_w26183_,
		_w26184_,
		_w26186_,
		_w26414_
	);
	LUT4 #(
		.INIT('hdff7)
	) name20588 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26415_
	);
	LUT4 #(
		.INIT('he400)
	) name20589 (
		_w26182_,
		_w26413_,
		_w26414_,
		_w26415_,
		_w26416_
	);
	LUT4 #(
		.INIT('hff9f)
	) name20590 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26417_
	);
	LUT2 #(
		.INIT('h2)
	) name20591 (
		_w26182_,
		_w26417_,
		_w26418_
	);
	LUT4 #(
		.INIT('h0400)
	) name20592 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26419_
	);
	LUT4 #(
		.INIT('hfb05)
	) name20593 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26420_
	);
	LUT4 #(
		.INIT('h4401)
	) name20594 (
		_w26182_,
		_w26185_,
		_w26184_,
		_w26186_,
		_w26421_
	);
	LUT4 #(
		.INIT('h1000)
	) name20595 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26422_
	);
	LUT4 #(
		.INIT('h6f7f)
	) name20596 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26423_
	);
	LUT4 #(
		.INIT('h0d00)
	) name20597 (
		_w26182_,
		_w26420_,
		_w26421_,
		_w26423_,
		_w26424_
	);
	LUT4 #(
		.INIT('h3120)
	) name20598 (
		_w26193_,
		_w26418_,
		_w26424_,
		_w26416_,
		_w26425_
	);
	LUT2 #(
		.INIT('h9)
	) name20599 (
		\u0_L11_reg[17]/NET0131 ,
		_w26425_,
		_w26426_
	);
	LUT4 #(
		.INIT('hc693)
	) name20600 (
		decrypt_pad,
		\u0_R11_reg[20]/NET0131 ,
		\u0_uk_K_r11_reg[31]/NET0131 ,
		\u0_uk_K_r11_reg[36]/NET0131 ,
		_w26427_
	);
	LUT4 #(
		.INIT('hc963)
	) name20601 (
		decrypt_pad,
		\u0_R11_reg[19]/NET0131 ,
		\u0_uk_K_r11_reg[21]/NET0131 ,
		\u0_uk_K_r11_reg[43]/NET0131 ,
		_w26428_
	);
	LUT4 #(
		.INIT('hc693)
	) name20602 (
		decrypt_pad,
		\u0_R11_reg[21]/NET0131 ,
		\u0_uk_K_r11_reg[28]/NET0131 ,
		\u0_uk_K_r11_reg[37]/NET0131 ,
		_w26429_
	);
	LUT4 #(
		.INIT('hc693)
	) name20603 (
		decrypt_pad,
		\u0_R11_reg[16]/NET0131 ,
		\u0_uk_K_r11_reg[16]/NET0131 ,
		\u0_uk_K_r11_reg[49]/NET0131 ,
		_w26430_
	);
	LUT4 #(
		.INIT('hc693)
	) name20604 (
		decrypt_pad,
		\u0_R11_reg[18]/NET0131 ,
		\u0_uk_K_r11_reg[1]/NET0131 ,
		\u0_uk_K_r11_reg[38]/NET0131 ,
		_w26431_
	);
	LUT4 #(
		.INIT('hc963)
	) name20605 (
		decrypt_pad,
		\u0_R11_reg[17]/NET0131 ,
		\u0_uk_K_r11_reg[16]/NET0131 ,
		\u0_uk_K_r11_reg[7]/NET0131 ,
		_w26432_
	);
	LUT3 #(
		.INIT('h80)
	) name20606 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26433_
	);
	LUT4 #(
		.INIT('h6c6a)
	) name20607 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26434_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name20608 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26435_
	);
	LUT4 #(
		.INIT('h08a0)
	) name20609 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26436_
	);
	LUT4 #(
		.INIT('h0e02)
	) name20610 (
		_w26435_,
		_w26428_,
		_w26436_,
		_w26434_,
		_w26437_
	);
	LUT2 #(
		.INIT('h2)
	) name20611 (
		_w26427_,
		_w26437_,
		_w26438_
	);
	LUT4 #(
		.INIT('hf6ef)
	) name20612 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26439_
	);
	LUT2 #(
		.INIT('h2)
	) name20613 (
		_w26428_,
		_w26439_,
		_w26440_
	);
	LUT2 #(
		.INIT('h4)
	) name20614 (
		_w26429_,
		_w26428_,
		_w26441_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name20615 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26442_
	);
	LUT3 #(
		.INIT('hd0)
	) name20616 (
		_w26432_,
		_w26429_,
		_w26428_,
		_w26443_
	);
	LUT4 #(
		.INIT('h0f01)
	) name20617 (
		_w26432_,
		_w26430_,
		_w26431_,
		_w26428_,
		_w26444_
	);
	LUT4 #(
		.INIT('he0ee)
	) name20618 (
		_w26441_,
		_w26442_,
		_w26443_,
		_w26444_,
		_w26445_
	);
	LUT4 #(
		.INIT('h0040)
	) name20619 (
		_w26432_,
		_w26430_,
		_w26431_,
		_w26428_,
		_w26446_
	);
	LUT4 #(
		.INIT('h0080)
	) name20620 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26447_
	);
	LUT2 #(
		.INIT('h1)
	) name20621 (
		_w26446_,
		_w26447_,
		_w26448_
	);
	LUT4 #(
		.INIT('h0e00)
	) name20622 (
		_w26427_,
		_w26445_,
		_w26440_,
		_w26448_,
		_w26449_
	);
	LUT3 #(
		.INIT('h65)
	) name20623 (
		\u0_L11_reg[25]/NET0131 ,
		_w26438_,
		_w26449_,
		_w26450_
	);
	LUT4 #(
		.INIT('h3fc6)
	) name20624 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26451_
	);
	LUT4 #(
		.INIT('h5404)
	) name20625 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26452_
	);
	LUT4 #(
		.INIT('hab7b)
	) name20626 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26453_
	);
	LUT4 #(
		.INIT('h0200)
	) name20627 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26454_
	);
	LUT4 #(
		.INIT('h00e4)
	) name20628 (
		_w26218_,
		_w26453_,
		_w26451_,
		_w26454_,
		_w26455_
	);
	LUT2 #(
		.INIT('h1)
	) name20629 (
		_w26212_,
		_w26455_,
		_w26456_
	);
	LUT4 #(
		.INIT('hf37b)
	) name20630 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26457_
	);
	LUT2 #(
		.INIT('h2)
	) name20631 (
		_w26218_,
		_w26457_,
		_w26458_
	);
	LUT3 #(
		.INIT('h28)
	) name20632 (
		_w26213_,
		_w26215_,
		_w26216_,
		_w26459_
	);
	LUT3 #(
		.INIT('h01)
	) name20633 (
		_w26224_,
		_w26452_,
		_w26459_,
		_w26460_
	);
	LUT4 #(
		.INIT('h0010)
	) name20634 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26461_
	);
	LUT4 #(
		.INIT('h4000)
	) name20635 (
		_w26213_,
		_w26214_,
		_w26218_,
		_w26216_,
		_w26462_
	);
	LUT2 #(
		.INIT('h1)
	) name20636 (
		_w26461_,
		_w26462_,
		_w26463_
	);
	LUT4 #(
		.INIT('h5700)
	) name20637 (
		_w26212_,
		_w26458_,
		_w26460_,
		_w26463_,
		_w26464_
	);
	LUT3 #(
		.INIT('h9a)
	) name20638 (
		\u0_L11_reg[29]/NET0131 ,
		_w26456_,
		_w26464_,
		_w26465_
	);
	LUT4 #(
		.INIT('h4010)
	) name20639 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26466_
	);
	LUT2 #(
		.INIT('h4)
	) name20640 (
		_w26353_,
		_w26355_,
		_w26467_
	);
	LUT4 #(
		.INIT('hc400)
	) name20641 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26352_,
		_w26468_
	);
	LUT3 #(
		.INIT('h02)
	) name20642 (
		_w26351_,
		_w26468_,
		_w26466_,
		_w26469_
	);
	LUT2 #(
		.INIT('h4)
	) name20643 (
		_w26353_,
		_w26356_,
		_w26470_
	);
	LUT4 #(
		.INIT('h0010)
	) name20644 (
		_w26353_,
		_w26355_,
		_w26356_,
		_w26352_,
		_w26471_
	);
	LUT4 #(
		.INIT('h0800)
	) name20645 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26472_
	);
	LUT2 #(
		.INIT('h1)
	) name20646 (
		_w26471_,
		_w26472_,
		_w26473_
	);
	LUT2 #(
		.INIT('h8)
	) name20647 (
		_w26356_,
		_w26352_,
		_w26474_
	);
	LUT3 #(
		.INIT('h20)
	) name20648 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26475_
	);
	LUT3 #(
		.INIT('h15)
	) name20649 (
		_w26351_,
		_w26474_,
		_w26475_,
		_w26476_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name20650 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26477_
	);
	LUT4 #(
		.INIT('h0144)
	) name20651 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26478_
	);
	LUT3 #(
		.INIT('h0d)
	) name20652 (
		_w26372_,
		_w26477_,
		_w26478_,
		_w26479_
	);
	LUT4 #(
		.INIT('h1555)
	) name20653 (
		_w26469_,
		_w26473_,
		_w26476_,
		_w26479_,
		_w26480_
	);
	LUT4 #(
		.INIT('h0d00)
	) name20654 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26481_
	);
	LUT3 #(
		.INIT('h90)
	) name20655 (
		_w26354_,
		_w26356_,
		_w26351_,
		_w26482_
	);
	LUT4 #(
		.INIT('h3130)
	) name20656 (
		_w26370_,
		_w26467_,
		_w26481_,
		_w26482_,
		_w26483_
	);
	LUT4 #(
		.INIT('h0002)
	) name20657 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26484_
	);
	LUT4 #(
		.INIT('hbf00)
	) name20658 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26352_,
		_w26485_
	);
	LUT2 #(
		.INIT('h4)
	) name20659 (
		_w26484_,
		_w26485_,
		_w26486_
	);
	LUT3 #(
		.INIT('h0e)
	) name20660 (
		_w26352_,
		_w26483_,
		_w26486_,
		_w26487_
	);
	LUT3 #(
		.INIT('h56)
	) name20661 (
		\u0_L11_reg[2]/NET0131 ,
		_w26480_,
		_w26487_,
		_w26488_
	);
	LUT4 #(
		.INIT('h0004)
	) name20662 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26489_
	);
	LUT4 #(
		.INIT('he56b)
	) name20663 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26490_
	);
	LUT4 #(
		.INIT('h4002)
	) name20664 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26491_
	);
	LUT4 #(
		.INIT('h3fdd)
	) name20665 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26492_
	);
	LUT4 #(
		.INIT('h3edc)
	) name20666 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26493_
	);
	LUT4 #(
		.INIT('h3120)
	) name20667 (
		_w26428_,
		_w26491_,
		_w26493_,
		_w26490_,
		_w26494_
	);
	LUT2 #(
		.INIT('h1)
	) name20668 (
		_w26427_,
		_w26494_,
		_w26495_
	);
	LUT3 #(
		.INIT('h20)
	) name20669 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26496_
	);
	LUT4 #(
		.INIT('hb796)
	) name20670 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26428_,
		_w26497_
	);
	LUT2 #(
		.INIT('h1)
	) name20671 (
		_w26431_,
		_w26497_,
		_w26498_
	);
	LUT4 #(
		.INIT('hf800)
	) name20672 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26428_,
		_w26499_
	);
	LUT2 #(
		.INIT('h8)
	) name20673 (
		_w26492_,
		_w26499_,
		_w26500_
	);
	LUT2 #(
		.INIT('h2)
	) name20674 (
		_w26431_,
		_w26428_,
		_w26501_
	);
	LUT4 #(
		.INIT('h0400)
	) name20675 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26502_
	);
	LUT3 #(
		.INIT('h07)
	) name20676 (
		_w26433_,
		_w26501_,
		_w26502_,
		_w26503_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name20677 (
		_w26427_,
		_w26500_,
		_w26498_,
		_w26503_,
		_w26504_
	);
	LUT4 #(
		.INIT('h0108)
	) name20678 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26505_
	);
	LUT4 #(
		.INIT('h1000)
	) name20679 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26506_
	);
	LUT4 #(
		.INIT('hedff)
	) name20680 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26507_
	);
	LUT3 #(
		.INIT('h8d)
	) name20681 (
		_w26428_,
		_w26505_,
		_w26507_,
		_w26508_
	);
	LUT4 #(
		.INIT('h5556)
	) name20682 (
		\u0_L11_reg[14]/NET0131 ,
		_w26504_,
		_w26495_,
		_w26508_,
		_w26509_
	);
	LUT4 #(
		.INIT('h2500)
	) name20683 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26510_
	);
	LUT4 #(
		.INIT('hf070)
	) name20684 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26511_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name20685 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26512_
	);
	LUT4 #(
		.INIT('h8acf)
	) name20686 (
		_w26454_,
		_w26510_,
		_w26511_,
		_w26512_,
		_w26513_
	);
	LUT2 #(
		.INIT('h1)
	) name20687 (
		_w26222_,
		_w26461_,
		_w26514_
	);
	LUT3 #(
		.INIT('h45)
	) name20688 (
		_w26212_,
		_w26513_,
		_w26514_,
		_w26515_
	);
	LUT4 #(
		.INIT('h8804)
	) name20689 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26516_
	);
	LUT4 #(
		.INIT('h4000)
	) name20690 (
		_w26213_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26517_
	);
	LUT4 #(
		.INIT('h000b)
	) name20691 (
		_w26228_,
		_w26221_,
		_w26516_,
		_w26517_,
		_w26518_
	);
	LUT4 #(
		.INIT('h2a8a)
	) name20692 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26519_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name20693 (
		_w26213_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26520_
	);
	LUT3 #(
		.INIT('h21)
	) name20694 (
		_w26214_,
		_w26215_,
		_w26216_,
		_w26521_
	);
	LUT3 #(
		.INIT('hd6)
	) name20695 (
		_w26214_,
		_w26215_,
		_w26216_,
		_w26522_
	);
	LUT2 #(
		.INIT('h8)
	) name20696 (
		_w26213_,
		_w26218_,
		_w26523_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name20697 (
		_w26519_,
		_w26520_,
		_w26522_,
		_w26523_,
		_w26524_
	);
	LUT3 #(
		.INIT('hd0)
	) name20698 (
		_w26212_,
		_w26518_,
		_w26524_,
		_w26525_
	);
	LUT3 #(
		.INIT('h65)
	) name20699 (
		\u0_L11_reg[4]/NET0131 ,
		_w26515_,
		_w26525_,
		_w26526_
	);
	LUT4 #(
		.INIT('h33fb)
	) name20700 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26527_
	);
	LUT4 #(
		.INIT('h33cb)
	) name20701 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26528_
	);
	LUT4 #(
		.INIT('h0100)
	) name20702 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26529_
	);
	LUT4 #(
		.INIT('h3302)
	) name20703 (
		_w26246_,
		_w26245_,
		_w26528_,
		_w26529_,
		_w26530_
	);
	LUT4 #(
		.INIT('h0020)
	) name20704 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26246_,
		_w26531_
	);
	LUT3 #(
		.INIT('h01)
	) name20705 (
		_w26265_,
		_w26392_,
		_w26531_,
		_w26532_
	);
	LUT4 #(
		.INIT('h0100)
	) name20706 (
		_w26248_,
		_w26250_,
		_w26249_,
		_w26246_,
		_w26533_
	);
	LUT2 #(
		.INIT('h1)
	) name20707 (
		_w26378_,
		_w26533_,
		_w26534_
	);
	LUT4 #(
		.INIT('hddb6)
	) name20708 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26535_
	);
	LUT4 #(
		.INIT('hff6f)
	) name20709 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26536_
	);
	LUT4 #(
		.INIT('h0004)
	) name20710 (
		_w26248_,
		_w26249_,
		_w26246_,
		_w26245_,
		_w26537_
	);
	LUT4 #(
		.INIT('h00e4)
	) name20711 (
		_w26246_,
		_w26535_,
		_w26536_,
		_w26537_,
		_w26538_
	);
	LUT4 #(
		.INIT('hd500)
	) name20712 (
		_w26245_,
		_w26532_,
		_w26534_,
		_w26538_,
		_w26539_
	);
	LUT3 #(
		.INIT('h65)
	) name20713 (
		\u0_L11_reg[15]/P0001 ,
		_w26530_,
		_w26539_,
		_w26540_
	);
	LUT4 #(
		.INIT('hf32e)
	) name20714 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26541_
	);
	LUT2 #(
		.INIT('h1)
	) name20715 (
		_w26246_,
		_w26541_,
		_w26542_
	);
	LUT3 #(
		.INIT('hb0)
	) name20716 (
		_w26250_,
		_w26249_,
		_w26246_,
		_w26543_
	);
	LUT4 #(
		.INIT('hed6f)
	) name20717 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26544_
	);
	LUT3 #(
		.INIT('hb0)
	) name20718 (
		_w26527_,
		_w26543_,
		_w26544_,
		_w26545_
	);
	LUT3 #(
		.INIT('h8a)
	) name20719 (
		_w26245_,
		_w26542_,
		_w26545_,
		_w26546_
	);
	LUT4 #(
		.INIT('hfb00)
	) name20720 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26246_,
		_w26547_
	);
	LUT4 #(
		.INIT('h4f47)
	) name20721 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26249_,
		_w26548_
	);
	LUT4 #(
		.INIT('h5444)
	) name20722 (
		_w26245_,
		_w26267_,
		_w26547_,
		_w26548_,
		_w26549_
	);
	LUT2 #(
		.INIT('h1)
	) name20723 (
		_w26246_,
		_w26266_,
		_w26550_
	);
	LUT4 #(
		.INIT('h0080)
	) name20724 (
		_w26247_,
		_w26250_,
		_w26249_,
		_w26246_,
		_w26551_
	);
	LUT3 #(
		.INIT('h54)
	) name20725 (
		_w26245_,
		_w26389_,
		_w26551_,
		_w26552_
	);
	LUT4 #(
		.INIT('h0200)
	) name20726 (
		_w26247_,
		_w26248_,
		_w26250_,
		_w26246_,
		_w26553_
	);
	LUT3 #(
		.INIT('h07)
	) name20727 (
		_w26256_,
		_w26272_,
		_w26553_,
		_w26554_
	);
	LUT4 #(
		.INIT('h0100)
	) name20728 (
		_w26549_,
		_w26552_,
		_w26550_,
		_w26554_,
		_w26555_
	);
	LUT3 #(
		.INIT('h65)
	) name20729 (
		\u0_L11_reg[27]/NET0131 ,
		_w26546_,
		_w26555_,
		_w26556_
	);
	LUT3 #(
		.INIT('h04)
	) name20730 (
		_w26430_,
		_w26429_,
		_w26431_,
		_w26557_
	);
	LUT4 #(
		.INIT('h9f8f)
	) name20731 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26558_
	);
	LUT4 #(
		.INIT('h7f7b)
	) name20732 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26559_
	);
	LUT4 #(
		.INIT('hf6dd)
	) name20733 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26560_
	);
	LUT4 #(
		.INIT('hd800)
	) name20734 (
		_w26428_,
		_w26559_,
		_w26558_,
		_w26560_,
		_w26561_
	);
	LUT2 #(
		.INIT('h1)
	) name20735 (
		_w26427_,
		_w26561_,
		_w26562_
	);
	LUT3 #(
		.INIT('hbe)
	) name20736 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26563_
	);
	LUT4 #(
		.INIT('hbf00)
	) name20737 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26564_
	);
	LUT3 #(
		.INIT('h02)
	) name20738 (
		_w26428_,
		_w26564_,
		_w26563_,
		_w26565_
	);
	LUT3 #(
		.INIT('h02)
	) name20739 (
		_w26430_,
		_w26431_,
		_w26428_,
		_w26566_
	);
	LUT2 #(
		.INIT('h2)
	) name20740 (
		_w26507_,
		_w26566_,
		_w26567_
	);
	LUT4 #(
		.INIT('hf5df)
	) name20741 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26568_
	);
	LUT4 #(
		.INIT('he4ee)
	) name20742 (
		_w26428_,
		_w26502_,
		_w26506_,
		_w26568_,
		_w26569_
	);
	LUT4 #(
		.INIT('h0075)
	) name20743 (
		_w26427_,
		_w26565_,
		_w26567_,
		_w26569_,
		_w26570_
	);
	LUT3 #(
		.INIT('h65)
	) name20744 (
		\u0_L11_reg[8]/NET0131 ,
		_w26562_,
		_w26570_,
		_w26571_
	);
	LUT4 #(
		.INIT('h7f55)
	) name20745 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26216_,
		_w26572_
	);
	LUT2 #(
		.INIT('h1)
	) name20746 (
		_w26213_,
		_w26572_,
		_w26573_
	);
	LUT4 #(
		.INIT('h0802)
	) name20747 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26574_
	);
	LUT2 #(
		.INIT('h2)
	) name20748 (
		_w26213_,
		_w26218_,
		_w26575_
	);
	LUT3 #(
		.INIT('h04)
	) name20749 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26576_
	);
	LUT4 #(
		.INIT('h0031)
	) name20750 (
		_w26235_,
		_w26574_,
		_w26575_,
		_w26576_,
		_w26577_
	);
	LUT3 #(
		.INIT('h8a)
	) name20751 (
		_w26212_,
		_w26573_,
		_w26577_,
		_w26578_
	);
	LUT4 #(
		.INIT('h8000)
	) name20752 (
		_w26213_,
		_w26214_,
		_w26215_,
		_w26216_,
		_w26579_
	);
	LUT3 #(
		.INIT('h01)
	) name20753 (
		_w26218_,
		_w26521_,
		_w26579_,
		_w26580_
	);
	LUT3 #(
		.INIT('hb0)
	) name20754 (
		_w26214_,
		_w26215_,
		_w26218_,
		_w26581_
	);
	LUT3 #(
		.INIT('h15)
	) name20755 (
		_w26212_,
		_w26240_,
		_w26581_,
		_w26582_
	);
	LUT4 #(
		.INIT('h1011)
	) name20756 (
		_w26238_,
		_w26223_,
		_w26580_,
		_w26582_,
		_w26583_
	);
	LUT3 #(
		.INIT('h65)
	) name20757 (
		\u0_L11_reg[19]/NET0131 ,
		_w26578_,
		_w26583_,
		_w26584_
	);
	LUT4 #(
		.INIT('hfdc3)
	) name20758 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26585_
	);
	LUT2 #(
		.INIT('h1)
	) name20759 (
		_w26182_,
		_w26585_,
		_w26586_
	);
	LUT4 #(
		.INIT('hdf3f)
	) name20760 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26587_
	);
	LUT2 #(
		.INIT('h2)
	) name20761 (
		_w26182_,
		_w26587_,
		_w26588_
	);
	LUT3 #(
		.INIT('h07)
	) name20762 (
		_w26206_,
		_w26207_,
		_w26419_,
		_w26589_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name20763 (
		_w26193_,
		_w26586_,
		_w26588_,
		_w26589_,
		_w26590_
	);
	LUT4 #(
		.INIT('h6ffb)
	) name20764 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26591_
	);
	LUT2 #(
		.INIT('h1)
	) name20765 (
		_w26182_,
		_w26591_,
		_w26592_
	);
	LUT4 #(
		.INIT('h07ff)
	) name20766 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26593_
	);
	LUT2 #(
		.INIT('h1)
	) name20767 (
		_w26182_,
		_w26593_,
		_w26594_
	);
	LUT3 #(
		.INIT('h08)
	) name20768 (
		_w26182_,
		_w26184_,
		_w26186_,
		_w26595_
	);
	LUT3 #(
		.INIT('h32)
	) name20769 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26596_
	);
	LUT3 #(
		.INIT('h4c)
	) name20770 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26597_
	);
	LUT4 #(
		.INIT('h8acf)
	) name20771 (
		_w26207_,
		_w26595_,
		_w26596_,
		_w26597_,
		_w26598_
	);
	LUT3 #(
		.INIT('hcb)
	) name20772 (
		_w26183_,
		_w26184_,
		_w26186_,
		_w26599_
	);
	LUT2 #(
		.INIT('h2)
	) name20773 (
		_w26191_,
		_w26599_,
		_w26600_
	);
	LUT4 #(
		.INIT('h00ab)
	) name20774 (
		_w26193_,
		_w26594_,
		_w26598_,
		_w26600_,
		_w26601_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name20775 (
		\u0_L11_reg[23]/NET0131 ,
		_w26590_,
		_w26592_,
		_w26601_,
		_w26602_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name20776 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26603_
	);
	LUT3 #(
		.INIT('h01)
	) name20777 (
		_w26353_,
		_w26355_,
		_w26356_,
		_w26604_
	);
	LUT4 #(
		.INIT('hfde3)
	) name20778 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26605_
	);
	LUT4 #(
		.INIT('h0515)
	) name20779 (
		_w26352_,
		_w26351_,
		_w26603_,
		_w26605_,
		_w26606_
	);
	LUT3 #(
		.INIT('h02)
	) name20780 (
		_w26353_,
		_w26355_,
		_w26356_,
		_w26607_
	);
	LUT4 #(
		.INIT('hdf00)
	) name20781 (
		_w26353_,
		_w26354_,
		_w26356_,
		_w26352_,
		_w26608_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name20782 (
		_w26372_,
		_w26604_,
		_w26607_,
		_w26608_,
		_w26609_
	);
	LUT4 #(
		.INIT('h0004)
	) name20783 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26610_
	);
	LUT4 #(
		.INIT('h0002)
	) name20784 (
		_w26351_,
		_w26471_,
		_w26472_,
		_w26610_,
		_w26611_
	);
	LUT3 #(
		.INIT('h20)
	) name20785 (
		_w26603_,
		_w26609_,
		_w26611_,
		_w26612_
	);
	LUT4 #(
		.INIT('h0fb0)
	) name20786 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26613_
	);
	LUT4 #(
		.INIT('h7d00)
	) name20787 (
		_w26355_,
		_w26354_,
		_w26356_,
		_w26352_,
		_w26614_
	);
	LUT2 #(
		.INIT('h4)
	) name20788 (
		_w26613_,
		_w26614_,
		_w26615_
	);
	LUT3 #(
		.INIT('h32)
	) name20789 (
		_w26355_,
		_w26354_,
		_w26352_,
		_w26616_
	);
	LUT2 #(
		.INIT('h8)
	) name20790 (
		_w26470_,
		_w26616_,
		_w26617_
	);
	LUT3 #(
		.INIT('ha2)
	) name20791 (
		_w26353_,
		_w26355_,
		_w26356_,
		_w26618_
	);
	LUT3 #(
		.INIT('h15)
	) name20792 (
		_w26351_,
		_w26362_,
		_w26618_,
		_w26619_
	);
	LUT3 #(
		.INIT('h10)
	) name20793 (
		_w26615_,
		_w26617_,
		_w26619_,
		_w26620_
	);
	LUT4 #(
		.INIT('h999a)
	) name20794 (
		\u0_L11_reg[13]/NET0131 ,
		_w26606_,
		_w26612_,
		_w26620_,
		_w26621_
	);
	LUT4 #(
		.INIT('hc693)
	) name20795 (
		decrypt_pad,
		\u0_R11_reg[11]/P0001 ,
		\u0_uk_K_r11_reg[12]/NET0131 ,
		\u0_uk_K_r11_reg[17]/NET0131 ,
		_w26622_
	);
	LUT4 #(
		.INIT('hc693)
	) name20796 (
		decrypt_pad,
		\u0_R11_reg[12]/NET0131 ,
		\u0_uk_K_r11_reg[27]/P0001 ,
		\u0_uk_K_r11_reg[32]/NET0131 ,
		_w26623_
	);
	LUT4 #(
		.INIT('hc963)
	) name20797 (
		decrypt_pad,
		\u0_R11_reg[13]/NET0131 ,
		\u0_uk_K_r11_reg[20]/NET0131 ,
		\u0_uk_K_r11_reg[40]/NET0131 ,
		_w26624_
	);
	LUT4 #(
		.INIT('hc693)
	) name20798 (
		decrypt_pad,
		\u0_R11_reg[9]/NET0131 ,
		\u0_uk_K_r11_reg[3]/NET0131 ,
		\u0_uk_K_r11_reg[40]/NET0131 ,
		_w26625_
	);
	LUT4 #(
		.INIT('hc693)
	) name20799 (
		decrypt_pad,
		\u0_R11_reg[10]/NET0131 ,
		\u0_uk_K_r11_reg[11]/NET0131 ,
		\u0_uk_K_r11_reg[48]/NET0131 ,
		_w26626_
	);
	LUT4 #(
		.INIT('hc963)
	) name20800 (
		decrypt_pad,
		\u0_R11_reg[8]/NET0131 ,
		\u0_uk_K_r11_reg[11]/NET0131 ,
		\u0_uk_K_r11_reg[6]/NET0131 ,
		_w26627_
	);
	LUT4 #(
		.INIT('hc733)
	) name20801 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26628_
	);
	LUT2 #(
		.INIT('h1)
	) name20802 (
		_w26626_,
		_w26625_,
		_w26629_
	);
	LUT4 #(
		.INIT('h0001)
	) name20803 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26630_
	);
	LUT4 #(
		.INIT('hff76)
	) name20804 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26631_
	);
	LUT4 #(
		.INIT('h08cc)
	) name20805 (
		_w26623_,
		_w26622_,
		_w26628_,
		_w26631_,
		_w26632_
	);
	LUT2 #(
		.INIT('h9)
	) name20806 (
		_w26626_,
		_w26625_,
		_w26633_
	);
	LUT2 #(
		.INIT('h8)
	) name20807 (
		_w26624_,
		_w26627_,
		_w26634_
	);
	LUT2 #(
		.INIT('h6)
	) name20808 (
		_w26624_,
		_w26627_,
		_w26635_
	);
	LUT3 #(
		.INIT('h46)
	) name20809 (
		_w26624_,
		_w26627_,
		_w26622_,
		_w26636_
	);
	LUT2 #(
		.INIT('h2)
	) name20810 (
		_w26633_,
		_w26636_,
		_w26637_
	);
	LUT3 #(
		.INIT('h40)
	) name20811 (
		_w26627_,
		_w26625_,
		_w26622_,
		_w26638_
	);
	LUT4 #(
		.INIT('h1428)
	) name20812 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26639_
	);
	LUT3 #(
		.INIT('h45)
	) name20813 (
		_w26623_,
		_w26638_,
		_w26639_,
		_w26640_
	);
	LUT2 #(
		.INIT('h8)
	) name20814 (
		_w26623_,
		_w26626_,
		_w26641_
	);
	LUT3 #(
		.INIT('h10)
	) name20815 (
		_w26624_,
		_w26627_,
		_w26625_,
		_w26642_
	);
	LUT4 #(
		.INIT('h0acf)
	) name20816 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26643_
	);
	LUT4 #(
		.INIT('h008a)
	) name20817 (
		_w26623_,
		_w26624_,
		_w26625_,
		_w26622_,
		_w26644_
	);
	LUT4 #(
		.INIT('h7077)
	) name20818 (
		_w26641_,
		_w26642_,
		_w26643_,
		_w26644_,
		_w26645_
	);
	LUT4 #(
		.INIT('h4500)
	) name20819 (
		_w26632_,
		_w26637_,
		_w26640_,
		_w26645_,
		_w26646_
	);
	LUT2 #(
		.INIT('h9)
	) name20820 (
		\u0_L11_reg[6]/NET0131 ,
		_w26646_,
		_w26647_
	);
	LUT4 #(
		.INIT('hf700)
	) name20821 (
		_w26152_,
		_w26157_,
		_w26153_,
		_w26154_,
		_w26648_
	);
	LUT3 #(
		.INIT('h40)
	) name20822 (
		_w26152_,
		_w26155_,
		_w26153_,
		_w26649_
	);
	LUT4 #(
		.INIT('haffc)
	) name20823 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26650_
	);
	LUT2 #(
		.INIT('h8)
	) name20824 (
		_w26648_,
		_w26650_,
		_w26651_
	);
	LUT4 #(
		.INIT('h0104)
	) name20825 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26652_
	);
	LUT4 #(
		.INIT('h00fb)
	) name20826 (
		_w26157_,
		_w26155_,
		_w26153_,
		_w26154_,
		_w26653_
	);
	LUT3 #(
		.INIT('h10)
	) name20827 (
		_w26406_,
		_w26652_,
		_w26653_,
		_w26654_
	);
	LUT4 #(
		.INIT('h0080)
	) name20828 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26655_
	);
	LUT4 #(
		.INIT('haa02)
	) name20829 (
		_w26151_,
		_w26651_,
		_w26654_,
		_w26655_,
		_w26656_
	);
	LUT4 #(
		.INIT('h0ff4)
	) name20830 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26657_
	);
	LUT2 #(
		.INIT('h1)
	) name20831 (
		_w26154_,
		_w26657_,
		_w26658_
	);
	LUT2 #(
		.INIT('h1)
	) name20832 (
		_w26155_,
		_w26154_,
		_w26659_
	);
	LUT3 #(
		.INIT('hc4)
	) name20833 (
		_w26152_,
		_w26157_,
		_w26153_,
		_w26660_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name20834 (
		_w26175_,
		_w26649_,
		_w26659_,
		_w26660_,
		_w26661_
	);
	LUT4 #(
		.INIT('h00c8)
	) name20835 (
		_w26152_,
		_w26155_,
		_w26153_,
		_w26154_,
		_w26662_
	);
	LUT4 #(
		.INIT('h0777)
	) name20836 (
		_w26171_,
		_w26154_,
		_w26161_,
		_w26662_,
		_w26663_
	);
	LUT4 #(
		.INIT('hba00)
	) name20837 (
		_w26151_,
		_w26658_,
		_w26661_,
		_w26663_,
		_w26664_
	);
	LUT3 #(
		.INIT('h65)
	) name20838 (
		\u0_L11_reg[32]/NET0131 ,
		_w26656_,
		_w26664_,
		_w26665_
	);
	LUT3 #(
		.INIT('h21)
	) name20839 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26666_
	);
	LUT4 #(
		.INIT('h30c8)
	) name20840 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26667_
	);
	LUT2 #(
		.INIT('h2)
	) name20841 (
		_w26151_,
		_w26154_,
		_w26668_
	);
	LUT3 #(
		.INIT('h10)
	) name20842 (
		_w26667_,
		_w26666_,
		_w26668_,
		_w26669_
	);
	LUT4 #(
		.INIT('h4410)
	) name20843 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26670_
	);
	LUT4 #(
		.INIT('h2080)
	) name20844 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26671_
	);
	LUT2 #(
		.INIT('h9)
	) name20845 (
		_w26151_,
		_w26154_,
		_w26672_
	);
	LUT4 #(
		.INIT('h0100)
	) name20846 (
		_w26160_,
		_w26670_,
		_w26671_,
		_w26672_,
		_w26673_
	);
	LUT4 #(
		.INIT('h936e)
	) name20847 (
		_w26152_,
		_w26157_,
		_w26155_,
		_w26153_,
		_w26674_
	);
	LUT4 #(
		.INIT('h0004)
	) name20848 (
		_w26151_,
		_w26154_,
		_w26160_,
		_w26674_,
		_w26675_
	);
	LUT4 #(
		.INIT('h00ab)
	) name20849 (
		_w26406_,
		_w26669_,
		_w26673_,
		_w26675_,
		_w26676_
	);
	LUT2 #(
		.INIT('h6)
	) name20850 (
		\u0_L11_reg[7]/NET0131 ,
		_w26676_,
		_w26677_
	);
	LUT3 #(
		.INIT('h29)
	) name20851 (
		_w26624_,
		_w26627_,
		_w26622_,
		_w26678_
	);
	LUT3 #(
		.INIT('h0e)
	) name20852 (
		_w26626_,
		_w26625_,
		_w26622_,
		_w26679_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name20853 (
		_w26629_,
		_w26635_,
		_w26678_,
		_w26679_,
		_w26680_
	);
	LUT2 #(
		.INIT('h2)
	) name20854 (
		_w26623_,
		_w26680_,
		_w26681_
	);
	LUT4 #(
		.INIT('hf859)
	) name20855 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26682_
	);
	LUT4 #(
		.INIT('h0020)
	) name20856 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26683_
	);
	LUT4 #(
		.INIT('h5504)
	) name20857 (
		_w26623_,
		_w26622_,
		_w26682_,
		_w26683_,
		_w26684_
	);
	LUT4 #(
		.INIT('h0410)
	) name20858 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26685_
	);
	LUT4 #(
		.INIT('h57f7)
	) name20859 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26686_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name20860 (
		_w26623_,
		_w26622_,
		_w26685_,
		_w26686_,
		_w26687_
	);
	LUT3 #(
		.INIT('h80)
	) name20861 (
		_w26624_,
		_w26627_,
		_w26625_,
		_w26688_
	);
	LUT2 #(
		.INIT('h2)
	) name20862 (
		_w26626_,
		_w26622_,
		_w26689_
	);
	LUT4 #(
		.INIT('h0041)
	) name20863 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26690_
	);
	LUT4 #(
		.INIT('hc7b6)
	) name20864 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26691_
	);
	LUT2 #(
		.INIT('h1)
	) name20865 (
		_w26623_,
		_w26622_,
		_w26692_
	);
	LUT4 #(
		.INIT('h7077)
	) name20866 (
		_w26688_,
		_w26689_,
		_w26691_,
		_w26692_,
		_w26693_
	);
	LUT3 #(
		.INIT('h10)
	) name20867 (
		_w26684_,
		_w26687_,
		_w26693_,
		_w26694_
	);
	LUT3 #(
		.INIT('h65)
	) name20868 (
		\u0_L11_reg[24]/NET0131 ,
		_w26681_,
		_w26694_,
		_w26695_
	);
	LUT4 #(
		.INIT('hf9e9)
	) name20869 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26696_
	);
	LUT4 #(
		.INIT('h5c5f)
	) name20870 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26697_
	);
	LUT4 #(
		.INIT('ha820)
	) name20871 (
		_w26623_,
		_w26622_,
		_w26697_,
		_w26696_,
		_w26698_
	);
	LUT4 #(
		.INIT('h80a0)
	) name20872 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26699_
	);
	LUT4 #(
		.INIT('hef00)
	) name20873 (
		_w26626_,
		_w26624_,
		_w26625_,
		_w26622_,
		_w26700_
	);
	LUT4 #(
		.INIT('h4050)
	) name20874 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26701_
	);
	LUT4 #(
		.INIT('h00df)
	) name20875 (
		_w26624_,
		_w26627_,
		_w26625_,
		_w26622_,
		_w26702_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name20876 (
		_w26699_,
		_w26700_,
		_w26701_,
		_w26702_,
		_w26703_
	);
	LUT4 #(
		.INIT('h0008)
	) name20877 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26704_
	);
	LUT3 #(
		.INIT('h01)
	) name20878 (
		_w26623_,
		_w26690_,
		_w26704_,
		_w26705_
	);
	LUT3 #(
		.INIT('h20)
	) name20879 (
		_w26626_,
		_w26625_,
		_w26622_,
		_w26706_
	);
	LUT4 #(
		.INIT('h0020)
	) name20880 (
		_w26626_,
		_w26624_,
		_w26625_,
		_w26622_,
		_w26707_
	);
	LUT3 #(
		.INIT('h80)
	) name20881 (
		_w26623_,
		_w26626_,
		_w26625_,
		_w26708_
	);
	LUT4 #(
		.INIT('h0123)
	) name20882 (
		_w26634_,
		_w26707_,
		_w26708_,
		_w26706_,
		_w26709_
	);
	LUT4 #(
		.INIT('hba00)
	) name20883 (
		_w26698_,
		_w26703_,
		_w26705_,
		_w26709_,
		_w26710_
	);
	LUT2 #(
		.INIT('h6)
	) name20884 (
		\u0_L11_reg[30]/NET0131 ,
		_w26710_,
		_w26711_
	);
	LUT4 #(
		.INIT('hfd3d)
	) name20885 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26712_
	);
	LUT4 #(
		.INIT('hfb7f)
	) name20886 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26713_
	);
	LUT4 #(
		.INIT('hb100)
	) name20887 (
		_w26428_,
		_w26496_,
		_w26712_,
		_w26713_,
		_w26714_
	);
	LUT2 #(
		.INIT('h2)
	) name20888 (
		_w26427_,
		_w26714_,
		_w26715_
	);
	LUT4 #(
		.INIT('h4009)
	) name20889 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26716_
	);
	LUT4 #(
		.INIT('hfda8)
	) name20890 (
		_w26428_,
		_w26489_,
		_w26506_,
		_w26716_,
		_w26717_
	);
	LUT4 #(
		.INIT('hf7c7)
	) name20891 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26718_
	);
	LUT2 #(
		.INIT('h2)
	) name20892 (
		_w26428_,
		_w26718_,
		_w26719_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name20893 (
		_w26432_,
		_w26430_,
		_w26429_,
		_w26431_,
		_w26720_
	);
	LUT3 #(
		.INIT('hb0)
	) name20894 (
		_w26432_,
		_w26431_,
		_w26428_,
		_w26721_
	);
	LUT3 #(
		.INIT('h01)
	) name20895 (
		_w26557_,
		_w26721_,
		_w26720_,
		_w26722_
	);
	LUT4 #(
		.INIT('h2223)
	) name20896 (
		_w26427_,
		_w26717_,
		_w26719_,
		_w26722_,
		_w26723_
	);
	LUT3 #(
		.INIT('h65)
	) name20897 (
		\u0_L11_reg[3]/NET0131 ,
		_w26715_,
		_w26723_,
		_w26724_
	);
	LUT4 #(
		.INIT('h8228)
	) name20898 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26725_
	);
	LUT3 #(
		.INIT('he6)
	) name20899 (
		_w26183_,
		_w26184_,
		_w26186_,
		_w26726_
	);
	LUT4 #(
		.INIT('h0031)
	) name20900 (
		_w26191_,
		_w26422_,
		_w26726_,
		_w26725_,
		_w26727_
	);
	LUT2 #(
		.INIT('h2)
	) name20901 (
		_w26193_,
		_w26727_,
		_w26728_
	);
	LUT4 #(
		.INIT('h4000)
	) name20902 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26729_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name20903 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26730_
	);
	LUT2 #(
		.INIT('h1)
	) name20904 (
		_w26182_,
		_w26730_,
		_w26731_
	);
	LUT4 #(
		.INIT('hd3c3)
	) name20905 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26732_
	);
	LUT2 #(
		.INIT('h2)
	) name20906 (
		_w26182_,
		_w26732_,
		_w26733_
	);
	LUT4 #(
		.INIT('h0802)
	) name20907 (
		_w26185_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26734_
	);
	LUT4 #(
		.INIT('h0141)
	) name20908 (
		_w26182_,
		_w26183_,
		_w26184_,
		_w26186_,
		_w26735_
	);
	LUT3 #(
		.INIT('h01)
	) name20909 (
		_w26729_,
		_w26735_,
		_w26734_,
		_w26736_
	);
	LUT4 #(
		.INIT('h2322)
	) name20910 (
		_w26193_,
		_w26731_,
		_w26733_,
		_w26736_,
		_w26737_
	);
	LUT3 #(
		.INIT('h65)
	) name20911 (
		\u0_L11_reg[9]/NET0131 ,
		_w26728_,
		_w26737_,
		_w26738_
	);
	LUT3 #(
		.INIT('h68)
	) name20912 (
		_w26624_,
		_w26627_,
		_w26625_,
		_w26739_
	);
	LUT4 #(
		.INIT('h6800)
	) name20913 (
		_w26624_,
		_w26627_,
		_w26625_,
		_w26622_,
		_w26740_
	);
	LUT4 #(
		.INIT('h3ef2)
	) name20914 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26741_
	);
	LUT4 #(
		.INIT('h0032)
	) name20915 (
		_w26622_,
		_w26630_,
		_w26741_,
		_w26740_,
		_w26742_
	);
	LUT2 #(
		.INIT('h1)
	) name20916 (
		_w26623_,
		_w26742_,
		_w26743_
	);
	LUT4 #(
		.INIT('h0111)
	) name20917 (
		_w26624_,
		_w26627_,
		_w26625_,
		_w26622_,
		_w26744_
	);
	LUT3 #(
		.INIT('h01)
	) name20918 (
		_w26626_,
		_w26739_,
		_w26744_,
		_w26745_
	);
	LUT4 #(
		.INIT('h0012)
	) name20919 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26622_,
		_w26746_
	);
	LUT4 #(
		.INIT('h0800)
	) name20920 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26747_
	);
	LUT2 #(
		.INIT('h1)
	) name20921 (
		_w26746_,
		_w26747_,
		_w26748_
	);
	LUT4 #(
		.INIT('h0008)
	) name20922 (
		_w26626_,
		_w26627_,
		_w26625_,
		_w26622_,
		_w26749_
	);
	LUT4 #(
		.INIT('hdffd)
	) name20923 (
		_w26626_,
		_w26624_,
		_w26627_,
		_w26625_,
		_w26750_
	);
	LUT3 #(
		.INIT('h31)
	) name20924 (
		_w26622_,
		_w26749_,
		_w26750_,
		_w26751_
	);
	LUT4 #(
		.INIT('h7500)
	) name20925 (
		_w26623_,
		_w26745_,
		_w26748_,
		_w26751_,
		_w26752_
	);
	LUT3 #(
		.INIT('h65)
	) name20926 (
		\u0_L11_reg[16]/NET0131 ,
		_w26743_,
		_w26752_,
		_w26753_
	);
	LUT4 #(
		.INIT('h1a00)
	) name20927 (
		_w26355_,
		_w26354_,
		_w26356_,
		_w26351_,
		_w26754_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name20928 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26755_
	);
	LUT3 #(
		.INIT('h8a)
	) name20929 (
		_w26352_,
		_w26754_,
		_w26755_,
		_w26756_
	);
	LUT4 #(
		.INIT('h0109)
	) name20930 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26352_,
		_w26757_
	);
	LUT4 #(
		.INIT('h2080)
	) name20931 (
		_w26353_,
		_w26355_,
		_w26354_,
		_w26356_,
		_w26758_
	);
	LUT4 #(
		.INIT('h8000)
	) name20932 (
		_w26355_,
		_w26354_,
		_w26356_,
		_w26352_,
		_w26759_
	);
	LUT4 #(
		.INIT('h0001)
	) name20933 (
		_w26604_,
		_w26759_,
		_w26758_,
		_w26757_,
		_w26760_
	);
	LUT3 #(
		.INIT('hac)
	) name20934 (
		_w26353_,
		_w26355_,
		_w26356_,
		_w26761_
	);
	LUT2 #(
		.INIT('h8)
	) name20935 (
		_w26354_,
		_w26351_,
		_w26762_
	);
	LUT4 #(
		.INIT('h4544)
	) name20936 (
		_w26352_,
		_w26359_,
		_w26761_,
		_w26762_,
		_w26763_
	);
	LUT4 #(
		.INIT('h0072)
	) name20937 (
		_w26351_,
		_w26484_,
		_w26760_,
		_w26763_,
		_w26764_
	);
	LUT3 #(
		.INIT('h65)
	) name20938 (
		\u0_L11_reg[18]/NET0131 ,
		_w26756_,
		_w26764_,
		_w26765_
	);
	LUT4 #(
		.INIT('hc963)
	) name20939 (
		decrypt_pad,
		\u0_R10_reg[4]/NET0131 ,
		\u0_uk_K_r10_reg[39]/NET0131 ,
		\u0_uk_K_r10_reg[5]/NET0131 ,
		_w26766_
	);
	LUT4 #(
		.INIT('hc693)
	) name20940 (
		decrypt_pad,
		\u0_R10_reg[32]/NET0131 ,
		\u0_uk_K_r10_reg[39]/NET0131 ,
		\u0_uk_K_r10_reg[48]/NET0131 ,
		_w26767_
	);
	LUT4 #(
		.INIT('hc963)
	) name20941 (
		decrypt_pad,
		\u0_R10_reg[5]/NET0131 ,
		\u0_uk_K_r10_reg[10]/NET0131 ,
		\u0_uk_K_r10_reg[33]/NET0131 ,
		_w26768_
	);
	LUT2 #(
		.INIT('h1)
	) name20942 (
		_w26767_,
		_w26768_,
		_w26769_
	);
	LUT4 #(
		.INIT('hc693)
	) name20943 (
		decrypt_pad,
		\u0_R10_reg[3]/NET0131 ,
		\u0_uk_K_r10_reg[27]/NET0131 ,
		\u0_uk_K_r10_reg[4]/NET0131 ,
		_w26770_
	);
	LUT4 #(
		.INIT('hc693)
	) name20944 (
		decrypt_pad,
		\u0_R10_reg[2]/NET0131 ,
		\u0_uk_K_r10_reg[18]/NET0131 ,
		\u0_uk_K_r10_reg[27]/NET0131 ,
		_w26771_
	);
	LUT3 #(
		.INIT('h02)
	) name20945 (
		_w26770_,
		_w26771_,
		_w26767_,
		_w26772_
	);
	LUT4 #(
		.INIT('hc963)
	) name20946 (
		decrypt_pad,
		\u0_R10_reg[1]/NET0131 ,
		\u0_uk_K_r10_reg[12]/NET0131 ,
		\u0_uk_K_r10_reg[3]/NET0131 ,
		_w26773_
	);
	LUT4 #(
		.INIT('hffc8)
	) name20947 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26774_
	);
	LUT3 #(
		.INIT('h45)
	) name20948 (
		_w26769_,
		_w26772_,
		_w26774_,
		_w26775_
	);
	LUT4 #(
		.INIT('hfd0d)
	) name20949 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26776_
	);
	LUT4 #(
		.INIT('haff3)
	) name20950 (
		_w26770_,
		_w26771_,
		_w26767_,
		_w26773_,
		_w26777_
	);
	LUT3 #(
		.INIT('hd0)
	) name20951 (
		_w26770_,
		_w26776_,
		_w26777_,
		_w26778_
	);
	LUT3 #(
		.INIT('h8a)
	) name20952 (
		_w26766_,
		_w26775_,
		_w26778_,
		_w26779_
	);
	LUT4 #(
		.INIT('h7c3f)
	) name20953 (
		_w26770_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26780_
	);
	LUT2 #(
		.INIT('h1)
	) name20954 (
		_w26771_,
		_w26780_,
		_w26781_
	);
	LUT2 #(
		.INIT('h8)
	) name20955 (
		_w26770_,
		_w26771_,
		_w26782_
	);
	LUT3 #(
		.INIT('h60)
	) name20956 (
		_w26767_,
		_w26768_,
		_w26773_,
		_w26783_
	);
	LUT4 #(
		.INIT('h0008)
	) name20957 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26784_
	);
	LUT4 #(
		.INIT('heef6)
	) name20958 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26785_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name20959 (
		_w26770_,
		_w26771_,
		_w26783_,
		_w26785_,
		_w26786_
	);
	LUT3 #(
		.INIT('h45)
	) name20960 (
		_w26766_,
		_w26781_,
		_w26786_,
		_w26787_
	);
	LUT4 #(
		.INIT('h8000)
	) name20961 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26788_
	);
	LUT3 #(
		.INIT('h47)
	) name20962 (
		_w26771_,
		_w26768_,
		_w26773_,
		_w26789_
	);
	LUT4 #(
		.INIT('h7adf)
	) name20963 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26790_
	);
	LUT2 #(
		.INIT('h1)
	) name20964 (
		_w26770_,
		_w26790_,
		_w26791_
	);
	LUT2 #(
		.INIT('h1)
	) name20965 (
		_w26771_,
		_w26773_,
		_w26792_
	);
	LUT4 #(
		.INIT('h0020)
	) name20966 (
		_w26770_,
		_w26771_,
		_w26767_,
		_w26773_,
		_w26793_
	);
	LUT3 #(
		.INIT('h08)
	) name20967 (
		_w26770_,
		_w26771_,
		_w26773_,
		_w26794_
	);
	LUT3 #(
		.INIT('h13)
	) name20968 (
		_w26769_,
		_w26793_,
		_w26794_,
		_w26795_
	);
	LUT2 #(
		.INIT('h4)
	) name20969 (
		_w26791_,
		_w26795_,
		_w26796_
	);
	LUT4 #(
		.INIT('h5655)
	) name20970 (
		\u0_L10_reg[31]/NET0131 ,
		_w26787_,
		_w26779_,
		_w26796_,
		_w26797_
	);
	LUT4 #(
		.INIT('hc693)
	) name20971 (
		decrypt_pad,
		\u0_R10_reg[26]/NET0131 ,
		\u0_uk_K_r10_reg[16]/NET0131 ,
		\u0_uk_K_r10_reg[21]/NET0131 ,
		_w26798_
	);
	LUT4 #(
		.INIT('hc693)
	) name20972 (
		decrypt_pad,
		\u0_R10_reg[25]/NET0131 ,
		\u0_uk_K_r10_reg[0]/NET0131 ,
		\u0_uk_K_r10_reg[36]/NET0131 ,
		_w26799_
	);
	LUT4 #(
		.INIT('hc963)
	) name20973 (
		decrypt_pad,
		\u0_R10_reg[24]/NET0131 ,
		\u0_uk_K_r10_reg[1]/NET0131 ,
		\u0_uk_K_r10_reg[51]/NET0131 ,
		_w26800_
	);
	LUT4 #(
		.INIT('hc693)
	) name20974 (
		decrypt_pad,
		\u0_R10_reg[29]/NET0131 ,
		\u0_uk_K_r10_reg[28]/NET0131 ,
		\u0_uk_K_r10_reg[9]/NET0131 ,
		_w26801_
	);
	LUT4 #(
		.INIT('h0200)
	) name20975 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w26802_
	);
	LUT4 #(
		.INIT('hadff)
	) name20976 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w26803_
	);
	LUT4 #(
		.INIT('hc693)
	) name20977 (
		decrypt_pad,
		\u0_R10_reg[28]/NET0131 ,
		\u0_uk_K_r10_reg[36]/NET0131 ,
		\u0_uk_K_r10_reg[45]/P0001 ,
		_w26804_
	);
	LUT4 #(
		.INIT('hc963)
	) name20978 (
		decrypt_pad,
		\u0_R10_reg[27]/NET0131 ,
		\u0_uk_K_r10_reg[30]/NET0131 ,
		\u0_uk_K_r10_reg[49]/NET0131 ,
		_w26805_
	);
	LUT4 #(
		.INIT('h006f)
	) name20979 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26805_,
		_w26806_
	);
	LUT3 #(
		.INIT('hb0)
	) name20980 (
		_w26803_,
		_w26804_,
		_w26806_,
		_w26807_
	);
	LUT2 #(
		.INIT('h2)
	) name20981 (
		_w26798_,
		_w26799_,
		_w26808_
	);
	LUT4 #(
		.INIT('h0400)
	) name20982 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w26809_
	);
	LUT4 #(
		.INIT('hfbbf)
	) name20983 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w26810_
	);
	LUT4 #(
		.INIT('h000b)
	) name20984 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w26811_
	);
	LUT3 #(
		.INIT('h08)
	) name20985 (
		_w26805_,
		_w26810_,
		_w26811_,
		_w26812_
	);
	LUT2 #(
		.INIT('h1)
	) name20986 (
		_w26807_,
		_w26812_,
		_w26813_
	);
	LUT2 #(
		.INIT('h8)
	) name20987 (
		_w26800_,
		_w26805_,
		_w26814_
	);
	LUT4 #(
		.INIT('hddad)
	) name20988 (
		_w26800_,
		_w26799_,
		_w26801_,
		_w26805_,
		_w26815_
	);
	LUT2 #(
		.INIT('h1)
	) name20989 (
		_w26798_,
		_w26815_,
		_w26816_
	);
	LUT4 #(
		.INIT('h7f75)
	) name20990 (
		_w26800_,
		_w26798_,
		_w26801_,
		_w26805_,
		_w26817_
	);
	LUT2 #(
		.INIT('h2)
	) name20991 (
		_w26799_,
		_w26817_,
		_w26818_
	);
	LUT4 #(
		.INIT('h0004)
	) name20992 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w26819_
	);
	LUT4 #(
		.INIT('h77fb)
	) name20993 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w26820_
	);
	LUT4 #(
		.INIT('h1000)
	) name20994 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w26821_
	);
	LUT4 #(
		.INIT('h0054)
	) name20995 (
		_w26804_,
		_w26805_,
		_w26820_,
		_w26821_,
		_w26822_
	);
	LUT3 #(
		.INIT('h10)
	) name20996 (
		_w26818_,
		_w26816_,
		_w26822_,
		_w26823_
	);
	LUT3 #(
		.INIT('h9d)
	) name20997 (
		_w26798_,
		_w26799_,
		_w26801_,
		_w26824_
	);
	LUT2 #(
		.INIT('h2)
	) name20998 (
		_w26814_,
		_w26824_,
		_w26825_
	);
	LUT4 #(
		.INIT('h0001)
	) name20999 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w26826_
	);
	LUT3 #(
		.INIT('h02)
	) name21000 (
		_w26804_,
		_w26809_,
		_w26826_,
		_w26827_
	);
	LUT2 #(
		.INIT('h4)
	) name21001 (
		_w26825_,
		_w26827_,
		_w26828_
	);
	LUT4 #(
		.INIT('h6665)
	) name21002 (
		\u0_L10_reg[22]/NET0131 ,
		_w26813_,
		_w26823_,
		_w26828_,
		_w26829_
	);
	LUT4 #(
		.INIT('hc693)
	) name21003 (
		decrypt_pad,
		\u0_R10_reg[24]/NET0131 ,
		\u0_uk_K_r10_reg[29]/NET0131 ,
		\u0_uk_K_r10_reg[38]/NET0131 ,
		_w26830_
	);
	LUT4 #(
		.INIT('hc693)
	) name21004 (
		decrypt_pad,
		\u0_R10_reg[23]/NET0131 ,
		\u0_uk_K_r10_reg[31]/NET0131 ,
		\u0_uk_K_r10_reg[8]/NET0131 ,
		_w26831_
	);
	LUT4 #(
		.INIT('hc693)
	) name21005 (
		decrypt_pad,
		\u0_R10_reg[22]/NET0131 ,
		\u0_uk_K_r10_reg[14]/NET0131 ,
		\u0_uk_K_r10_reg[50]/NET0131 ,
		_w26832_
	);
	LUT4 #(
		.INIT('hc963)
	) name21006 (
		decrypt_pad,
		\u0_R10_reg[20]/NET0131 ,
		\u0_uk_K_r10_reg[44]/NET0131 ,
		\u0_uk_K_r10_reg[8]/NET0131 ,
		_w26833_
	);
	LUT4 #(
		.INIT('hc693)
	) name21007 (
		decrypt_pad,
		\u0_R10_reg[21]/NET0131 ,
		\u0_uk_K_r10_reg[23]/NET0131 ,
		\u0_uk_K_r10_reg[28]/NET0131 ,
		_w26834_
	);
	LUT3 #(
		.INIT('h20)
	) name21008 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26835_
	);
	LUT4 #(
		.INIT('h1400)
	) name21009 (
		_w26831_,
		_w26832_,
		_w26833_,
		_w26834_,
		_w26836_
	);
	LUT2 #(
		.INIT('h1)
	) name21010 (
		_w26831_,
		_w26832_,
		_w26837_
	);
	LUT4 #(
		.INIT('hc963)
	) name21011 (
		decrypt_pad,
		\u0_R10_reg[25]/NET0131 ,
		\u0_uk_K_r10_reg[29]/NET0131 ,
		\u0_uk_K_r10_reg[52]/NET0131 ,
		_w26838_
	);
	LUT4 #(
		.INIT('h0010)
	) name21012 (
		_w26831_,
		_w26832_,
		_w26833_,
		_w26838_,
		_w26839_
	);
	LUT4 #(
		.INIT('h0800)
	) name21013 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26840_
	);
	LUT2 #(
		.INIT('h1)
	) name21014 (
		_w26839_,
		_w26840_,
		_w26841_
	);
	LUT3 #(
		.INIT('ha2)
	) name21015 (
		_w26833_,
		_w26834_,
		_w26838_,
		_w26842_
	);
	LUT3 #(
		.INIT('hcd)
	) name21016 (
		_w26831_,
		_w26832_,
		_w26833_,
		_w26843_
	);
	LUT3 #(
		.INIT('h47)
	) name21017 (
		_w26832_,
		_w26833_,
		_w26838_,
		_w26844_
	);
	LUT2 #(
		.INIT('h2)
	) name21018 (
		_w26831_,
		_w26834_,
		_w26845_
	);
	LUT4 #(
		.INIT('he0ee)
	) name21019 (
		_w26842_,
		_w26843_,
		_w26844_,
		_w26845_,
		_w26846_
	);
	LUT4 #(
		.INIT('h5155)
	) name21020 (
		_w26830_,
		_w26841_,
		_w26836_,
		_w26846_,
		_w26847_
	);
	LUT4 #(
		.INIT('h168a)
	) name21021 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26848_
	);
	LUT2 #(
		.INIT('h1)
	) name21022 (
		_w26831_,
		_w26848_,
		_w26849_
	);
	LUT4 #(
		.INIT('h0004)
	) name21023 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26850_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name21024 (
		_w26831_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26851_
	);
	LUT4 #(
		.INIT('hef00)
	) name21025 (
		_w26835_,
		_w26850_,
		_w26851_,
		_w26830_,
		_w26852_
	);
	LUT3 #(
		.INIT('h04)
	) name21026 (
		_w26833_,
		_w26834_,
		_w26838_,
		_w26853_
	);
	LUT4 #(
		.INIT('h0010)
	) name21027 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26854_
	);
	LUT4 #(
		.INIT('h77ef)
	) name21028 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26855_
	);
	LUT2 #(
		.INIT('h2)
	) name21029 (
		_w26831_,
		_w26855_,
		_w26856_
	);
	LUT3 #(
		.INIT('hf6)
	) name21030 (
		_w26833_,
		_w26834_,
		_w26838_,
		_w26857_
	);
	LUT3 #(
		.INIT('h10)
	) name21031 (
		_w26833_,
		_w26834_,
		_w26838_,
		_w26858_
	);
	LUT4 #(
		.INIT('hdcfe)
	) name21032 (
		_w26831_,
		_w26832_,
		_w26857_,
		_w26858_,
		_w26859_
	);
	LUT4 #(
		.INIT('h0b00)
	) name21033 (
		_w26849_,
		_w26852_,
		_w26856_,
		_w26859_,
		_w26860_
	);
	LUT3 #(
		.INIT('h9a)
	) name21034 (
		\u0_L10_reg[11]/NET0131 ,
		_w26847_,
		_w26860_,
		_w26861_
	);
	LUT4 #(
		.INIT('hfe3c)
	) name21035 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26862_
	);
	LUT4 #(
		.INIT('h8008)
	) name21036 (
		_w26770_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26863_
	);
	LUT4 #(
		.INIT('hf7df)
	) name21037 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26864_
	);
	LUT4 #(
		.INIT('h0e00)
	) name21038 (
		_w26770_,
		_w26862_,
		_w26863_,
		_w26864_,
		_w26865_
	);
	LUT4 #(
		.INIT('h0040)
	) name21039 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26866_
	);
	LUT4 #(
		.INIT('hcc9d)
	) name21040 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26867_
	);
	LUT4 #(
		.INIT('h4041)
	) name21041 (
		_w26770_,
		_w26771_,
		_w26767_,
		_w26773_,
		_w26868_
	);
	LUT4 #(
		.INIT('h0400)
	) name21042 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26869_
	);
	LUT4 #(
		.INIT('h5bff)
	) name21043 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w26870_
	);
	LUT4 #(
		.INIT('h0d00)
	) name21044 (
		_w26770_,
		_w26867_,
		_w26868_,
		_w26870_,
		_w26871_
	);
	LUT3 #(
		.INIT('hed)
	) name21045 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26872_
	);
	LUT2 #(
		.INIT('h8)
	) name21046 (
		_w26770_,
		_w26773_,
		_w26873_
	);
	LUT2 #(
		.INIT('h4)
	) name21047 (
		_w26872_,
		_w26873_,
		_w26874_
	);
	LUT4 #(
		.INIT('h00d8)
	) name21048 (
		_w26766_,
		_w26871_,
		_w26865_,
		_w26874_,
		_w26875_
	);
	LUT2 #(
		.INIT('h9)
	) name21049 (
		\u0_L10_reg[17]/NET0131 ,
		_w26875_,
		_w26876_
	);
	LUT4 #(
		.INIT('hc693)
	) name21050 (
		decrypt_pad,
		\u0_R10_reg[15]/NET0131 ,
		\u0_uk_K_r10_reg[24]/NET0131 ,
		\u0_uk_K_r10_reg[33]/NET0131 ,
		_w26877_
	);
	LUT4 #(
		.INIT('hc963)
	) name21051 (
		decrypt_pad,
		\u0_R10_reg[13]/NET0131 ,
		\u0_uk_K_r10_reg[24]/NET0131 ,
		\u0_uk_K_r10_reg[47]/NET0131 ,
		_w26878_
	);
	LUT2 #(
		.INIT('h8)
	) name21052 (
		_w26877_,
		_w26878_,
		_w26879_
	);
	LUT4 #(
		.INIT('hc693)
	) name21053 (
		decrypt_pad,
		\u0_R10_reg[12]/NET0131 ,
		\u0_uk_K_r10_reg[53]/NET0131 ,
		\u0_uk_K_r10_reg[5]/NET0131 ,
		_w26880_
	);
	LUT4 #(
		.INIT('hc693)
	) name21054 (
		decrypt_pad,
		\u0_R10_reg[17]/NET0131 ,
		\u0_uk_K_r10_reg[12]/NET0131 ,
		\u0_uk_K_r10_reg[46]/NET0131 ,
		_w26881_
	);
	LUT4 #(
		.INIT('hc963)
	) name21055 (
		decrypt_pad,
		\u0_R10_reg[14]/NET0131 ,
		\u0_uk_K_r10_reg[25]/NET0131 ,
		\u0_uk_K_r10_reg[48]/NET0131 ,
		_w26882_
	);
	LUT3 #(
		.INIT('hd8)
	) name21056 (
		_w26880_,
		_w26881_,
		_w26882_,
		_w26883_
	);
	LUT4 #(
		.INIT('hc693)
	) name21057 (
		decrypt_pad,
		\u0_R10_reg[16]/NET0131 ,
		\u0_uk_K_r10_reg[32]/NET0131 ,
		\u0_uk_K_r10_reg[41]/P0001 ,
		_w26884_
	);
	LUT3 #(
		.INIT('h07)
	) name21058 (
		_w26879_,
		_w26883_,
		_w26884_,
		_w26885_
	);
	LUT4 #(
		.INIT('h0002)
	) name21059 (
		_w26877_,
		_w26878_,
		_w26880_,
		_w26881_,
		_w26886_
	);
	LUT4 #(
		.INIT('h0040)
	) name21060 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w26887_
	);
	LUT2 #(
		.INIT('h1)
	) name21061 (
		_w26886_,
		_w26887_,
		_w26888_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name21062 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w26889_
	);
	LUT3 #(
		.INIT('h20)
	) name21063 (
		_w26880_,
		_w26881_,
		_w26882_,
		_w26890_
	);
	LUT4 #(
		.INIT('ha3af)
	) name21064 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w26891_
	);
	LUT3 #(
		.INIT('hc8)
	) name21065 (
		_w26877_,
		_w26889_,
		_w26891_,
		_w26892_
	);
	LUT3 #(
		.INIT('h80)
	) name21066 (
		_w26885_,
		_w26888_,
		_w26892_,
		_w26893_
	);
	LUT4 #(
		.INIT('h0014)
	) name21067 (
		_w26877_,
		_w26878_,
		_w26880_,
		_w26882_,
		_w26894_
	);
	LUT4 #(
		.INIT('h0080)
	) name21068 (
		_w26877_,
		_w26878_,
		_w26880_,
		_w26881_,
		_w26895_
	);
	LUT2 #(
		.INIT('h2)
	) name21069 (
		_w26877_,
		_w26878_,
		_w26896_
	);
	LUT4 #(
		.INIT('h0200)
	) name21070 (
		_w26877_,
		_w26878_,
		_w26880_,
		_w26881_,
		_w26897_
	);
	LUT4 #(
		.INIT('h0002)
	) name21071 (
		_w26884_,
		_w26897_,
		_w26895_,
		_w26894_,
		_w26898_
	);
	LUT4 #(
		.INIT('h0001)
	) name21072 (
		_w26877_,
		_w26878_,
		_w26880_,
		_w26881_,
		_w26899_
	);
	LUT4 #(
		.INIT('h0020)
	) name21073 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w26900_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name21074 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w26901_
	);
	LUT3 #(
		.INIT('h70)
	) name21075 (
		_w26882_,
		_w26899_,
		_w26901_,
		_w26902_
	);
	LUT2 #(
		.INIT('h8)
	) name21076 (
		_w26898_,
		_w26902_,
		_w26903_
	);
	LUT3 #(
		.INIT('h01)
	) name21077 (
		_w26880_,
		_w26881_,
		_w26882_,
		_w26904_
	);
	LUT3 #(
		.INIT('hde)
	) name21078 (
		_w26880_,
		_w26881_,
		_w26882_,
		_w26905_
	);
	LUT2 #(
		.INIT('h2)
	) name21079 (
		_w26896_,
		_w26905_,
		_w26906_
	);
	LUT4 #(
		.INIT('h0008)
	) name21080 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w26907_
	);
	LUT3 #(
		.INIT('h1b)
	) name21081 (
		_w26877_,
		_w26900_,
		_w26907_,
		_w26908_
	);
	LUT2 #(
		.INIT('h4)
	) name21082 (
		_w26906_,
		_w26908_,
		_w26909_
	);
	LUT4 #(
		.INIT('ha955)
	) name21083 (
		\u0_L10_reg[20]/NET0131 ,
		_w26893_,
		_w26903_,
		_w26909_,
		_w26910_
	);
	LUT4 #(
		.INIT('h77dc)
	) name21084 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26911_
	);
	LUT2 #(
		.INIT('h1)
	) name21085 (
		_w26831_,
		_w26911_,
		_w26912_
	);
	LUT4 #(
		.INIT('hcf6f)
	) name21086 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26913_
	);
	LUT2 #(
		.INIT('h2)
	) name21087 (
		_w26831_,
		_w26913_,
		_w26914_
	);
	LUT4 #(
		.INIT('h0102)
	) name21088 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26915_
	);
	LUT3 #(
		.INIT('h01)
	) name21089 (
		_w26839_,
		_w26840_,
		_w26915_,
		_w26916_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name21090 (
		_w26830_,
		_w26914_,
		_w26912_,
		_w26916_,
		_w26917_
	);
	LUT4 #(
		.INIT('h3fd2)
	) name21091 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26918_
	);
	LUT4 #(
		.INIT('hab6f)
	) name21092 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26919_
	);
	LUT4 #(
		.INIT('h0200)
	) name21093 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26920_
	);
	LUT4 #(
		.INIT('h00d8)
	) name21094 (
		_w26831_,
		_w26918_,
		_w26919_,
		_w26920_,
		_w26921_
	);
	LUT4 #(
		.INIT('h2000)
	) name21095 (
		_w26831_,
		_w26832_,
		_w26834_,
		_w26838_,
		_w26922_
	);
	LUT2 #(
		.INIT('h1)
	) name21096 (
		_w26850_,
		_w26922_,
		_w26923_
	);
	LUT3 #(
		.INIT('he0)
	) name21097 (
		_w26830_,
		_w26921_,
		_w26923_,
		_w26924_
	);
	LUT3 #(
		.INIT('h9a)
	) name21098 (
		\u0_L10_reg[29]/NET0131 ,
		_w26917_,
		_w26924_,
		_w26925_
	);
	LUT4 #(
		.INIT('hc963)
	) name21099 (
		decrypt_pad,
		\u0_R10_reg[30]/NET0131 ,
		\u0_uk_K_r10_reg[43]/NET0131 ,
		\u0_uk_K_r10_reg[7]/NET0131 ,
		_w26926_
	);
	LUT4 #(
		.INIT('hc693)
	) name21100 (
		decrypt_pad,
		\u0_R10_reg[29]/NET0131 ,
		\u0_uk_K_r10_reg[37]/NET0131 ,
		\u0_uk_K_r10_reg[42]/NET0131 ,
		_w26927_
	);
	LUT4 #(
		.INIT('hc693)
	) name21101 (
		decrypt_pad,
		\u0_R10_reg[1]/NET0131 ,
		\u0_uk_K_r10_reg[22]/NET0131 ,
		\u0_uk_K_r10_reg[31]/NET0131 ,
		_w26928_
	);
	LUT2 #(
		.INIT('h8)
	) name21102 (
		_w26927_,
		_w26928_,
		_w26929_
	);
	LUT4 #(
		.INIT('hc963)
	) name21103 (
		decrypt_pad,
		\u0_R10_reg[28]/NET0131 ,
		\u0_uk_K_r10_reg[15]/NET0131 ,
		\u0_uk_K_r10_reg[38]/NET0131 ,
		_w26930_
	);
	LUT4 #(
		.INIT('h0080)
	) name21104 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w26931_
	);
	LUT2 #(
		.INIT('h2)
	) name21105 (
		_w26927_,
		_w26928_,
		_w26932_
	);
	LUT4 #(
		.INIT('h0400)
	) name21106 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w26933_
	);
	LUT4 #(
		.INIT('h590c)
	) name21107 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w26934_
	);
	LUT4 #(
		.INIT('hc963)
	) name21108 (
		decrypt_pad,
		\u0_R10_reg[31]/P0001 ,
		\u0_uk_K_r10_reg[0]/NET0131 ,
		\u0_uk_K_r10_reg[50]/NET0131 ,
		_w26935_
	);
	LUT4 #(
		.INIT('h00df)
	) name21109 (
		_w26926_,
		_w26927_,
		_w26930_,
		_w26935_,
		_w26936_
	);
	LUT4 #(
		.INIT('h00de)
	) name21110 (
		_w26926_,
		_w26927_,
		_w26930_,
		_w26935_,
		_w26937_
	);
	LUT4 #(
		.INIT('h5510)
	) name21111 (
		_w26931_,
		_w26934_,
		_w26935_,
		_w26937_,
		_w26938_
	);
	LUT4 #(
		.INIT('hc693)
	) name21112 (
		decrypt_pad,
		\u0_R10_reg[32]/NET0131 ,
		\u0_uk_K_r10_reg[1]/NET0131 ,
		\u0_uk_K_r10_reg[37]/NET0131 ,
		_w26939_
	);
	LUT2 #(
		.INIT('h4)
	) name21113 (
		_w26938_,
		_w26939_,
		_w26940_
	);
	LUT4 #(
		.INIT('h0200)
	) name21114 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w26941_
	);
	LUT4 #(
		.INIT('hfb00)
	) name21115 (
		_w26927_,
		_w26928_,
		_w26930_,
		_w26935_,
		_w26942_
	);
	LUT3 #(
		.INIT('h02)
	) name21116 (
		_w26926_,
		_w26928_,
		_w26930_,
		_w26943_
	);
	LUT3 #(
		.INIT('h07)
	) name21117 (
		_w26927_,
		_w26928_,
		_w26935_,
		_w26944_
	);
	LUT4 #(
		.INIT('h8acf)
	) name21118 (
		_w26943_,
		_w26941_,
		_w26942_,
		_w26944_,
		_w26945_
	);
	LUT4 #(
		.INIT('h8000)
	) name21119 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w26946_
	);
	LUT3 #(
		.INIT('h04)
	) name21120 (
		_w26926_,
		_w26930_,
		_w26935_,
		_w26947_
	);
	LUT3 #(
		.INIT('h01)
	) name21121 (
		_w26933_,
		_w26947_,
		_w26946_,
		_w26948_
	);
	LUT4 #(
		.INIT('h0001)
	) name21122 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w26949_
	);
	LUT4 #(
		.INIT('hfff6)
	) name21123 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w26950_
	);
	LUT4 #(
		.INIT('h0020)
	) name21124 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w26951_
	);
	LUT4 #(
		.INIT('hefd6)
	) name21125 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w26952_
	);
	LUT4 #(
		.INIT('h5f13)
	) name21126 (
		_w26932_,
		_w26935_,
		_w26947_,
		_w26952_,
		_w26953_
	);
	LUT4 #(
		.INIT('hba00)
	) name21127 (
		_w26939_,
		_w26945_,
		_w26948_,
		_w26953_,
		_w26954_
	);
	LUT3 #(
		.INIT('h9a)
	) name21128 (
		\u0_L10_reg[5]/NET0131 ,
		_w26940_,
		_w26954_,
		_w26955_
	);
	LUT3 #(
		.INIT('h32)
	) name21129 (
		_w26837_,
		_w26842_,
		_w26854_,
		_w26956_
	);
	LUT3 #(
		.INIT('h80)
	) name21130 (
		_w26832_,
		_w26834_,
		_w26838_,
		_w26957_
	);
	LUT4 #(
		.INIT('h2000)
	) name21131 (
		_w26831_,
		_w26832_,
		_w26833_,
		_w26838_,
		_w26958_
	);
	LUT3 #(
		.INIT('h02)
	) name21132 (
		_w26830_,
		_w26958_,
		_w26957_,
		_w26959_
	);
	LUT2 #(
		.INIT('h4)
	) name21133 (
		_w26956_,
		_w26959_,
		_w26960_
	);
	LUT3 #(
		.INIT('h10)
	) name21134 (
		_w26832_,
		_w26833_,
		_w26838_,
		_w26961_
	);
	LUT4 #(
		.INIT('haa2a)
	) name21135 (
		_w26831_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26962_
	);
	LUT3 #(
		.INIT('h10)
	) name21136 (
		_w26840_,
		_w26961_,
		_w26962_,
		_w26963_
	);
	LUT4 #(
		.INIT('h5545)
	) name21137 (
		_w26831_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26964_
	);
	LUT2 #(
		.INIT('h4)
	) name21138 (
		_w26920_,
		_w26964_,
		_w26965_
	);
	LUT4 #(
		.INIT('h1000)
	) name21139 (
		_w26831_,
		_w26832_,
		_w26833_,
		_w26838_,
		_w26966_
	);
	LUT3 #(
		.INIT('h01)
	) name21140 (
		_w26850_,
		_w26830_,
		_w26966_,
		_w26967_
	);
	LUT3 #(
		.INIT('he0)
	) name21141 (
		_w26963_,
		_w26965_,
		_w26967_,
		_w26968_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name21142 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w26969_
	);
	LUT4 #(
		.INIT('h4445)
	) name21143 (
		_w26831_,
		_w26832_,
		_w26833_,
		_w26838_,
		_w26970_
	);
	LUT3 #(
		.INIT('hb6)
	) name21144 (
		_w26833_,
		_w26834_,
		_w26838_,
		_w26971_
	);
	LUT2 #(
		.INIT('h8)
	) name21145 (
		_w26831_,
		_w26832_,
		_w26972_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name21146 (
		_w26969_,
		_w26970_,
		_w26971_,
		_w26972_,
		_w26973_
	);
	LUT4 #(
		.INIT('ha955)
	) name21147 (
		\u0_L10_reg[4]/NET0131 ,
		_w26960_,
		_w26968_,
		_w26973_,
		_w26974_
	);
	LUT4 #(
		.INIT('hc963)
	) name21148 (
		decrypt_pad,
		\u0_R10_reg[8]/NET0131 ,
		\u0_uk_K_r10_reg[40]/NET0131 ,
		\u0_uk_K_r10_reg[6]/NET0131 ,
		_w26975_
	);
	LUT4 #(
		.INIT('hc693)
	) name21149 (
		decrypt_pad,
		\u0_R10_reg[6]/NET0131 ,
		\u0_uk_K_r10_reg[46]/NET0131 ,
		\u0_uk_K_r10_reg[55]/NET0131 ,
		_w26976_
	);
	LUT4 #(
		.INIT('hc693)
	) name21150 (
		decrypt_pad,
		\u0_R10_reg[9]/NET0131 ,
		\u0_uk_K_r10_reg[11]/NET0131 ,
		\u0_uk_K_r10_reg[20]/NET0131 ,
		_w26977_
	);
	LUT4 #(
		.INIT('hc963)
	) name21151 (
		decrypt_pad,
		\u0_R10_reg[5]/NET0131 ,
		\u0_uk_K_r10_reg[32]/NET0131 ,
		\u0_uk_K_r10_reg[55]/NET0131 ,
		_w26978_
	);
	LUT4 #(
		.INIT('hc963)
	) name21152 (
		decrypt_pad,
		\u0_R10_reg[7]/NET0131 ,
		\u0_uk_K_r10_reg[17]/NET0131 ,
		\u0_uk_K_r10_reg[40]/NET0131 ,
		_w26979_
	);
	LUT4 #(
		.INIT('h0004)
	) name21153 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26979_,
		_w26980_
	);
	LUT4 #(
		.INIT('hc693)
	) name21154 (
		decrypt_pad,
		\u0_R10_reg[4]/NET0131 ,
		\u0_uk_K_r10_reg[19]/NET0131 ,
		\u0_uk_K_r10_reg[53]/NET0131 ,
		_w26981_
	);
	LUT2 #(
		.INIT('h2)
	) name21155 (
		_w26977_,
		_w26981_,
		_w26982_
	);
	LUT3 #(
		.INIT('h08)
	) name21156 (
		_w26977_,
		_w26978_,
		_w26981_,
		_w26983_
	);
	LUT4 #(
		.INIT('h0080)
	) name21157 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w26984_
	);
	LUT2 #(
		.INIT('h1)
	) name21158 (
		_w26980_,
		_w26984_,
		_w26985_
	);
	LUT4 #(
		.INIT('h0800)
	) name21159 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w26986_
	);
	LUT4 #(
		.INIT('h0103)
	) name21160 (
		_w26979_,
		_w26980_,
		_w26984_,
		_w26986_,
		_w26987_
	);
	LUT2 #(
		.INIT('h8)
	) name21161 (
		_w26977_,
		_w26981_,
		_w26988_
	);
	LUT4 #(
		.INIT('h1014)
	) name21162 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w26989_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name21163 (
		_w26977_,
		_w26978_,
		_w26979_,
		_w26981_,
		_w26990_
	);
	LUT4 #(
		.INIT('h51f3)
	) name21164 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w26991_
	);
	LUT3 #(
		.INIT('h51)
	) name21165 (
		_w26989_,
		_w26990_,
		_w26991_,
		_w26992_
	);
	LUT3 #(
		.INIT('h15)
	) name21166 (
		_w26975_,
		_w26987_,
		_w26992_,
		_w26993_
	);
	LUT4 #(
		.INIT('hf7cc)
	) name21167 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w26994_
	);
	LUT4 #(
		.INIT('h00c4)
	) name21168 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w26995_
	);
	LUT3 #(
		.INIT('h0b)
	) name21169 (
		_w26976_,
		_w26978_,
		_w26979_,
		_w26996_
	);
	LUT4 #(
		.INIT('hf200)
	) name21170 (
		_w26975_,
		_w26994_,
		_w26995_,
		_w26996_,
		_w26997_
	);
	LUT4 #(
		.INIT('h0002)
	) name21171 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w26998_
	);
	LUT4 #(
		.INIT('haffd)
	) name21172 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w26999_
	);
	LUT2 #(
		.INIT('h2)
	) name21173 (
		_w26979_,
		_w26999_,
		_w27000_
	);
	LUT4 #(
		.INIT('h0100)
	) name21174 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27001_
	);
	LUT4 #(
		.INIT('hc040)
	) name21175 (
		_w26976_,
		_w26978_,
		_w26979_,
		_w26981_,
		_w27002_
	);
	LUT4 #(
		.INIT('h4000)
	) name21176 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27003_
	);
	LUT4 #(
		.INIT('haaa8)
	) name21177 (
		_w26975_,
		_w27001_,
		_w27002_,
		_w27003_,
		_w27004_
	);
	LUT3 #(
		.INIT('h01)
	) name21178 (
		_w27000_,
		_w27004_,
		_w26997_,
		_w27005_
	);
	LUT3 #(
		.INIT('h65)
	) name21179 (
		\u0_L10_reg[2]/NET0131 ,
		_w26993_,
		_w27005_,
		_w27006_
	);
	LUT4 #(
		.INIT('h33cb)
	) name21180 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27007_
	);
	LUT4 #(
		.INIT('h0100)
	) name21181 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27008_
	);
	LUT4 #(
		.INIT('h0031)
	) name21182 (
		_w26935_,
		_w26939_,
		_w27007_,
		_w27008_,
		_w27009_
	);
	LUT4 #(
		.INIT('hbf00)
	) name21183 (
		_w26926_,
		_w26927_,
		_w26930_,
		_w26939_,
		_w27010_
	);
	LUT2 #(
		.INIT('h4)
	) name21184 (
		_w26927_,
		_w26935_,
		_w27011_
	);
	LUT4 #(
		.INIT('h0100)
	) name21185 (
		_w26927_,
		_w26928_,
		_w26930_,
		_w26935_,
		_w27012_
	);
	LUT4 #(
		.INIT('h0020)
	) name21186 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26935_,
		_w27013_
	);
	LUT4 #(
		.INIT('h2000)
	) name21187 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27014_
	);
	LUT4 #(
		.INIT('hdff7)
	) name21188 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27015_
	);
	LUT4 #(
		.INIT('h1000)
	) name21189 (
		_w27012_,
		_w27013_,
		_w27010_,
		_w27015_,
		_w27016_
	);
	LUT2 #(
		.INIT('h1)
	) name21190 (
		_w27009_,
		_w27016_,
		_w27017_
	);
	LUT4 #(
		.INIT('h0040)
	) name21191 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27018_
	);
	LUT3 #(
		.INIT('h08)
	) name21192 (
		_w26936_,
		_w26950_,
		_w27018_,
		_w27019_
	);
	LUT4 #(
		.INIT('h0010)
	) name21193 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27020_
	);
	LUT3 #(
		.INIT('h04)
	) name21194 (
		_w26931_,
		_w26935_,
		_w27020_,
		_w27021_
	);
	LUT4 #(
		.INIT('h0004)
	) name21195 (
		_w26927_,
		_w26930_,
		_w26935_,
		_w26939_,
		_w27022_
	);
	LUT3 #(
		.INIT('h0e)
	) name21196 (
		_w27019_,
		_w27021_,
		_w27022_,
		_w27023_
	);
	LUT3 #(
		.INIT('h65)
	) name21197 (
		\u0_L10_reg[15]/P0001 ,
		_w27017_,
		_w27023_,
		_w27024_
	);
	LUT4 #(
		.INIT('h0002)
	) name21198 (
		_w26927_,
		_w26928_,
		_w26930_,
		_w26935_,
		_w27025_
	);
	LUT3 #(
		.INIT('h01)
	) name21199 (
		_w26939_,
		_w26949_,
		_w27025_,
		_w27026_
	);
	LUT3 #(
		.INIT('h40)
	) name21200 (
		_w26926_,
		_w26928_,
		_w26930_,
		_w27027_
	);
	LUT3 #(
		.INIT('h45)
	) name21201 (
		_w26941_,
		_w27011_,
		_w27027_,
		_w27028_
	);
	LUT4 #(
		.INIT('hf5f1)
	) name21202 (
		_w26927_,
		_w26928_,
		_w26930_,
		_w26935_,
		_w27029_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name21203 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27030_
	);
	LUT4 #(
		.INIT('hf531)
	) name21204 (
		_w26926_,
		_w26935_,
		_w27029_,
		_w27030_,
		_w27031_
	);
	LUT3 #(
		.INIT('h80)
	) name21205 (
		_w27026_,
		_w27028_,
		_w27031_,
		_w27032_
	);
	LUT4 #(
		.INIT('h00ef)
	) name21206 (
		_w26926_,
		_w26928_,
		_w26930_,
		_w26935_,
		_w27033_
	);
	LUT4 #(
		.INIT('hf700)
	) name21207 (
		_w26927_,
		_w26928_,
		_w26930_,
		_w26935_,
		_w27034_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21208 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27035_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name21209 (
		_w27014_,
		_w27033_,
		_w27034_,
		_w27035_,
		_w27036_
	);
	LUT4 #(
		.INIT('h0802)
	) name21210 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27037_
	);
	LUT3 #(
		.INIT('h02)
	) name21211 (
		_w26939_,
		_w27020_,
		_w27037_,
		_w27038_
	);
	LUT2 #(
		.INIT('h4)
	) name21212 (
		_w27036_,
		_w27038_,
		_w27039_
	);
	LUT4 #(
		.INIT('h0100)
	) name21213 (
		_w26926_,
		_w26927_,
		_w26930_,
		_w26935_,
		_w27040_
	);
	LUT3 #(
		.INIT('h07)
	) name21214 (
		_w26929_,
		_w26947_,
		_w27040_,
		_w27041_
	);
	LUT4 #(
		.INIT('ha955)
	) name21215 (
		\u0_L10_reg[21]/NET0131 ,
		_w27032_,
		_w27039_,
		_w27041_,
		_w27042_
	);
	LUT4 #(
		.INIT('hc963)
	) name21216 (
		decrypt_pad,
		\u0_R10_reg[20]/NET0131 ,
		\u0_uk_K_r10_reg[22]/NET0131 ,
		\u0_uk_K_r10_reg[45]/P0001 ,
		_w27043_
	);
	LUT4 #(
		.INIT('hc693)
	) name21217 (
		decrypt_pad,
		\u0_R10_reg[19]/NET0131 ,
		\u0_uk_K_r10_reg[2]/NET0131 ,
		\u0_uk_K_r10_reg[7]/NET0131 ,
		_w27044_
	);
	LUT4 #(
		.INIT('hc693)
	) name21218 (
		decrypt_pad,
		\u0_R10_reg[17]/NET0131 ,
		\u0_uk_K_r10_reg[21]/NET0131 ,
		\u0_uk_K_r10_reg[2]/NET0131 ,
		_w27045_
	);
	LUT4 #(
		.INIT('hc693)
	) name21219 (
		decrypt_pad,
		\u0_R10_reg[16]/NET0131 ,
		\u0_uk_K_r10_reg[30]/NET0131 ,
		\u0_uk_K_r10_reg[35]/NET0131 ,
		_w27046_
	);
	LUT4 #(
		.INIT('hc693)
	) name21220 (
		decrypt_pad,
		\u0_R10_reg[18]/NET0131 ,
		\u0_uk_K_r10_reg[15]/NET0131 ,
		\u0_uk_K_r10_reg[51]/NET0131 ,
		_w27047_
	);
	LUT4 #(
		.INIT('hc963)
	) name21221 (
		decrypt_pad,
		\u0_R10_reg[21]/NET0131 ,
		\u0_uk_K_r10_reg[23]/NET0131 ,
		\u0_uk_K_r10_reg[42]/NET0131 ,
		_w27048_
	);
	LUT3 #(
		.INIT('h80)
	) name21222 (
		_w27045_,
		_w27048_,
		_w27046_,
		_w27049_
	);
	LUT4 #(
		.INIT('h3ec4)
	) name21223 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27050_
	);
	LUT3 #(
		.INIT('h40)
	) name21224 (
		_w27045_,
		_w27048_,
		_w27046_,
		_w27051_
	);
	LUT4 #(
		.INIT('hcfbb)
	) name21225 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27052_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name21226 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27053_
	);
	LUT4 #(
		.INIT('hd800)
	) name21227 (
		_w27044_,
		_w27050_,
		_w27052_,
		_w27053_,
		_w27054_
	);
	LUT2 #(
		.INIT('h2)
	) name21228 (
		_w27044_,
		_w27048_,
		_w27055_
	);
	LUT4 #(
		.INIT('hfc77)
	) name21229 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27056_
	);
	LUT3 #(
		.INIT('ha2)
	) name21230 (
		_w27044_,
		_w27045_,
		_w27048_,
		_w27057_
	);
	LUT4 #(
		.INIT('h2223)
	) name21231 (
		_w27044_,
		_w27047_,
		_w27045_,
		_w27046_,
		_w27058_
	);
	LUT4 #(
		.INIT('he0ee)
	) name21232 (
		_w27055_,
		_w27056_,
		_w27057_,
		_w27058_,
		_w27059_
	);
	LUT3 #(
		.INIT('h04)
	) name21233 (
		_w27047_,
		_w27048_,
		_w27046_,
		_w27060_
	);
	LUT4 #(
		.INIT('hf7ed)
	) name21234 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27061_
	);
	LUT2 #(
		.INIT('h4)
	) name21235 (
		_w27044_,
		_w27047_,
		_w27062_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name21236 (
		_w27044_,
		_w27047_,
		_w27045_,
		_w27048_,
		_w27063_
	);
	LUT4 #(
		.INIT('hf531)
	) name21237 (
		_w27044_,
		_w27046_,
		_w27061_,
		_w27063_,
		_w27064_
	);
	LUT4 #(
		.INIT('he200)
	) name21238 (
		_w27059_,
		_w27043_,
		_w27054_,
		_w27064_,
		_w27065_
	);
	LUT2 #(
		.INIT('h9)
	) name21239 (
		\u0_L10_reg[25]/NET0131 ,
		_w27065_,
		_w27066_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name21240 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w27067_
	);
	LUT2 #(
		.INIT('h2)
	) name21241 (
		_w26831_,
		_w27067_,
		_w27068_
	);
	LUT4 #(
		.INIT('h2050)
	) name21242 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w27069_
	);
	LUT4 #(
		.INIT('hfb00)
	) name21243 (
		_w26831_,
		_w26833_,
		_w26834_,
		_w26830_,
		_w27070_
	);
	LUT3 #(
		.INIT('h10)
	) name21244 (
		_w26915_,
		_w27069_,
		_w27070_,
		_w27071_
	);
	LUT4 #(
		.INIT('h4554)
	) name21245 (
		_w26831_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w27072_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name21246 (
		_w26831_,
		_w26832_,
		_w26833_,
		_w26834_,
		_w27073_
	);
	LUT3 #(
		.INIT('h23)
	) name21247 (
		_w26853_,
		_w27072_,
		_w27073_,
		_w27074_
	);
	LUT4 #(
		.INIT('h8000)
	) name21248 (
		_w26832_,
		_w26833_,
		_w26834_,
		_w26838_,
		_w27075_
	);
	LUT2 #(
		.INIT('h1)
	) name21249 (
		_w26830_,
		_w27075_,
		_w27076_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name21250 (
		_w27068_,
		_w27071_,
		_w27074_,
		_w27076_,
		_w27077_
	);
	LUT3 #(
		.INIT('hd7)
	) name21251 (
		_w26833_,
		_w26834_,
		_w26838_,
		_w27078_
	);
	LUT4 #(
		.INIT('hdfce)
	) name21252 (
		_w26831_,
		_w26832_,
		_w26858_,
		_w27078_,
		_w27079_
	);
	LUT3 #(
		.INIT('h65)
	) name21253 (
		\u0_L10_reg[19]/NET0131 ,
		_w27077_,
		_w27079_,
		_w27080_
	);
	LUT4 #(
		.INIT('h404c)
	) name21254 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27081_
	);
	LUT4 #(
		.INIT('h0400)
	) name21255 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27082_
	);
	LUT4 #(
		.INIT('hfad8)
	) name21256 (
		_w26877_,
		_w26904_,
		_w27081_,
		_w27082_,
		_w27083_
	);
	LUT4 #(
		.INIT('h7fd7)
	) name21257 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27084_
	);
	LUT3 #(
		.INIT('h45)
	) name21258 (
		_w26884_,
		_w27083_,
		_w27084_,
		_w27085_
	);
	LUT3 #(
		.INIT('hb0)
	) name21259 (
		_w26880_,
		_w26881_,
		_w26882_,
		_w27086_
	);
	LUT2 #(
		.INIT('h4)
	) name21260 (
		_w26877_,
		_w26878_,
		_w27087_
	);
	LUT4 #(
		.INIT('h4404)
	) name21261 (
		_w26877_,
		_w26878_,
		_w26880_,
		_w26881_,
		_w27088_
	);
	LUT4 #(
		.INIT('h0800)
	) name21262 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27089_
	);
	LUT4 #(
		.INIT('he6ff)
	) name21263 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27090_
	);
	LUT4 #(
		.INIT('h20aa)
	) name21264 (
		_w26884_,
		_w27086_,
		_w27088_,
		_w27090_,
		_w27091_
	);
	LUT4 #(
		.INIT('h6fff)
	) name21265 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27092_
	);
	LUT4 #(
		.INIT('h6dff)
	) name21266 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27093_
	);
	LUT2 #(
		.INIT('h2)
	) name21267 (
		_w26877_,
		_w27093_,
		_w27094_
	);
	LUT4 #(
		.INIT('hafab)
	) name21268 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27095_
	);
	LUT2 #(
		.INIT('h8)
	) name21269 (
		_w26877_,
		_w26884_,
		_w27096_
	);
	LUT2 #(
		.INIT('h4)
	) name21270 (
		_w27095_,
		_w27096_,
		_w27097_
	);
	LUT4 #(
		.INIT('h135f)
	) name21271 (
		_w26882_,
		_w26890_,
		_w26899_,
		_w27087_,
		_w27098_
	);
	LUT4 #(
		.INIT('h0100)
	) name21272 (
		_w27094_,
		_w27097_,
		_w27091_,
		_w27098_,
		_w27099_
	);
	LUT3 #(
		.INIT('h65)
	) name21273 (
		\u0_L10_reg[1]/NET0131 ,
		_w27085_,
		_w27099_,
		_w27100_
	);
	LUT4 #(
		.INIT('hfbef)
	) name21274 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w27101_
	);
	LUT4 #(
		.INIT('h0288)
	) name21275 (
		_w26770_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w27102_
	);
	LUT4 #(
		.INIT('h0032)
	) name21276 (
		_w26770_,
		_w26788_,
		_w27101_,
		_w27102_,
		_w27103_
	);
	LUT2 #(
		.INIT('h1)
	) name21277 (
		_w26782_,
		_w27103_,
		_w27104_
	);
	LUT4 #(
		.INIT('h3800)
	) name21278 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w27105_
	);
	LUT3 #(
		.INIT('h14)
	) name21279 (
		_w26767_,
		_w26768_,
		_w26773_,
		_w27106_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name21280 (
		_w26770_,
		_w26784_,
		_w27105_,
		_w27106_,
		_w27107_
	);
	LUT4 #(
		.INIT('h002a)
	) name21281 (
		_w26766_,
		_w26769_,
		_w26794_,
		_w26866_,
		_w27108_
	);
	LUT4 #(
		.INIT('h1554)
	) name21282 (
		_w26766_,
		_w26771_,
		_w26768_,
		_w26773_,
		_w27109_
	);
	LUT4 #(
		.INIT('h4440)
	) name21283 (
		_w26770_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w27110_
	);
	LUT2 #(
		.INIT('h2)
	) name21284 (
		_w26770_,
		_w26767_,
		_w27111_
	);
	LUT4 #(
		.INIT('h8caf)
	) name21285 (
		_w26792_,
		_w26789_,
		_w27110_,
		_w27111_,
		_w27112_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name21286 (
		_w27107_,
		_w27108_,
		_w27109_,
		_w27112_,
		_w27113_
	);
	LUT3 #(
		.INIT('ha9)
	) name21287 (
		\u0_L10_reg[23]/NET0131 ,
		_w27104_,
		_w27113_,
		_w27114_
	);
	LUT4 #(
		.INIT('hff2e)
	) name21288 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27115_
	);
	LUT3 #(
		.INIT('h02)
	) name21289 (
		_w26976_,
		_w26978_,
		_w26981_,
		_w27116_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name21290 (
		_w26976_,
		_w26978_,
		_w26979_,
		_w26981_,
		_w27117_
	);
	LUT4 #(
		.INIT('h0ef3)
	) name21291 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27118_
	);
	LUT4 #(
		.INIT('h7277)
	) name21292 (
		_w26979_,
		_w27115_,
		_w27116_,
		_w27118_,
		_w27119_
	);
	LUT4 #(
		.INIT('h0802)
	) name21293 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27120_
	);
	LUT4 #(
		.INIT('h2000)
	) name21294 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27121_
	);
	LUT3 #(
		.INIT('h01)
	) name21295 (
		_w26975_,
		_w27121_,
		_w27120_,
		_w27122_
	);
	LUT2 #(
		.INIT('h4)
	) name21296 (
		_w27119_,
		_w27122_,
		_w27123_
	);
	LUT3 #(
		.INIT('h90)
	) name21297 (
		_w26977_,
		_w26978_,
		_w26981_,
		_w27124_
	);
	LUT4 #(
		.INIT('h0020)
	) name21298 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27125_
	);
	LUT3 #(
		.INIT('h02)
	) name21299 (
		_w26979_,
		_w27125_,
		_w27124_,
		_w27126_
	);
	LUT4 #(
		.INIT('hdf2e)
	) name21300 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27127_
	);
	LUT2 #(
		.INIT('h8)
	) name21301 (
		_w27117_,
		_w27127_,
		_w27128_
	);
	LUT2 #(
		.INIT('h8)
	) name21302 (
		_w26979_,
		_w26981_,
		_w27129_
	);
	LUT4 #(
		.INIT('h0dff)
	) name21303 (
		_w26977_,
		_w26978_,
		_w26979_,
		_w26981_,
		_w27130_
	);
	LUT4 #(
		.INIT('h0008)
	) name21304 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27131_
	);
	LUT4 #(
		.INIT('h00a8)
	) name21305 (
		_w26975_,
		_w26976_,
		_w27130_,
		_w27131_,
		_w27132_
	);
	LUT3 #(
		.INIT('he0)
	) name21306 (
		_w27126_,
		_w27128_,
		_w27132_,
		_w27133_
	);
	LUT3 #(
		.INIT('ha9)
	) name21307 (
		\u0_L10_reg[28]/NET0131 ,
		_w27123_,
		_w27133_,
		_w27134_
	);
	LUT4 #(
		.INIT('hcf2f)
	) name21308 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27135_
	);
	LUT4 #(
		.INIT('h0100)
	) name21309 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27136_
	);
	LUT4 #(
		.INIT('h3eff)
	) name21310 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27137_
	);
	LUT4 #(
		.INIT('hf7b9)
	) name21311 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27138_
	);
	LUT4 #(
		.INIT('hd800)
	) name21312 (
		_w27044_,
		_w27137_,
		_w27135_,
		_w27138_,
		_w27139_
	);
	LUT4 #(
		.INIT('h0200)
	) name21313 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27140_
	);
	LUT4 #(
		.INIT('h0020)
	) name21314 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27141_
	);
	LUT4 #(
		.INIT('hf7b7)
	) name21315 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27142_
	);
	LUT4 #(
		.INIT('he4ee)
	) name21316 (
		_w27044_,
		_w27140_,
		_w27141_,
		_w27142_,
		_w27143_
	);
	LUT4 #(
		.INIT('h0028)
	) name21317 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27144_
	);
	LUT4 #(
		.INIT('h0001)
	) name21318 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27145_
	);
	LUT4 #(
		.INIT('hcffe)
	) name21319 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27146_
	);
	LUT2 #(
		.INIT('h1)
	) name21320 (
		_w27044_,
		_w27047_,
		_w27147_
	);
	LUT3 #(
		.INIT('h10)
	) name21321 (
		_w27044_,
		_w27047_,
		_w27046_,
		_w27148_
	);
	LUT4 #(
		.INIT('h000d)
	) name21322 (
		_w27044_,
		_w27146_,
		_w27144_,
		_w27148_,
		_w27149_
	);
	LUT4 #(
		.INIT('h3120)
	) name21323 (
		_w27043_,
		_w27143_,
		_w27149_,
		_w27139_,
		_w27150_
	);
	LUT2 #(
		.INIT('h9)
	) name21324 (
		\u0_L10_reg[8]/NET0131 ,
		_w27150_,
		_w27151_
	);
	LUT4 #(
		.INIT('h5f5e)
	) name21325 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27152_
	);
	LUT2 #(
		.INIT('h2)
	) name21326 (
		_w26805_,
		_w27152_,
		_w27153_
	);
	LUT3 #(
		.INIT('hd9)
	) name21327 (
		_w26800_,
		_w26801_,
		_w26805_,
		_w27154_
	);
	LUT2 #(
		.INIT('h2)
	) name21328 (
		_w26808_,
		_w27154_,
		_w27155_
	);
	LUT4 #(
		.INIT('hefbf)
	) name21329 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27156_
	);
	LUT3 #(
		.INIT('h40)
	) name21330 (
		_w26802_,
		_w26804_,
		_w27156_,
		_w27157_
	);
	LUT3 #(
		.INIT('h10)
	) name21331 (
		_w27153_,
		_w27155_,
		_w27157_,
		_w27158_
	);
	LUT4 #(
		.INIT('h41eb)
	) name21332 (
		_w26800_,
		_w26799_,
		_w26801_,
		_w26805_,
		_w27159_
	);
	LUT3 #(
		.INIT('h09)
	) name21333 (
		_w26799_,
		_w26801_,
		_w26805_,
		_w27160_
	);
	LUT3 #(
		.INIT('h04)
	) name21334 (
		_w26800_,
		_w26799_,
		_w26801_,
		_w27161_
	);
	LUT4 #(
		.INIT('hddd8)
	) name21335 (
		_w26798_,
		_w27159_,
		_w27161_,
		_w27160_,
		_w27162_
	);
	LUT3 #(
		.INIT('h02)
	) name21336 (
		_w26800_,
		_w26798_,
		_w26801_,
		_w27163_
	);
	LUT4 #(
		.INIT('h2d7d)
	) name21337 (
		_w26800_,
		_w26798_,
		_w26801_,
		_w26805_,
		_w27164_
	);
	LUT3 #(
		.INIT('h32)
	) name21338 (
		_w26799_,
		_w26804_,
		_w27164_,
		_w27165_
	);
	LUT2 #(
		.INIT('h4)
	) name21339 (
		_w27162_,
		_w27165_,
		_w27166_
	);
	LUT3 #(
		.INIT('ha9)
	) name21340 (
		\u0_L10_reg[12]/NET0131 ,
		_w27158_,
		_w27166_,
		_w27167_
	);
	LUT4 #(
		.INIT('hfdbd)
	) name21341 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27168_
	);
	LUT4 #(
		.INIT('hf3db)
	) name21342 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27169_
	);
	LUT4 #(
		.INIT('hc480)
	) name21343 (
		_w26877_,
		_w27092_,
		_w27168_,
		_w27169_,
		_w27170_
	);
	LUT2 #(
		.INIT('h2)
	) name21344 (
		_w26884_,
		_w27170_,
		_w27171_
	);
	LUT4 #(
		.INIT('hdd01)
	) name21345 (
		_w26877_,
		_w26878_,
		_w26881_,
		_w26882_,
		_w27172_
	);
	LUT4 #(
		.INIT('h0020)
	) name21346 (
		_w26877_,
		_w26878_,
		_w26881_,
		_w26882_,
		_w27173_
	);
	LUT3 #(
		.INIT('h02)
	) name21347 (
		_w26880_,
		_w27173_,
		_w27172_,
		_w27174_
	);
	LUT4 #(
		.INIT('h0020)
	) name21348 (
		_w26877_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27175_
	);
	LUT3 #(
		.INIT('h02)
	) name21349 (
		_w26889_,
		_w26899_,
		_w27175_,
		_w27176_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name21350 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w27177_
	);
	LUT4 #(
		.INIT('h0800)
	) name21351 (
		_w26877_,
		_w26878_,
		_w26880_,
		_w26882_,
		_w27178_
	);
	LUT4 #(
		.INIT('h0072)
	) name21352 (
		_w26877_,
		_w26907_,
		_w27177_,
		_w27178_,
		_w27179_
	);
	LUT4 #(
		.INIT('hba00)
	) name21353 (
		_w26884_,
		_w27174_,
		_w27176_,
		_w27179_,
		_w27180_
	);
	LUT3 #(
		.INIT('h65)
	) name21354 (
		\u0_L10_reg[10]/NET0131 ,
		_w27171_,
		_w27180_,
		_w27181_
	);
	LUT4 #(
		.INIT('h9fff)
	) name21355 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27182_
	);
	LUT4 #(
		.INIT('hfec7)
	) name21356 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27183_
	);
	LUT4 #(
		.INIT('h0313)
	) name21357 (
		_w26975_,
		_w26979_,
		_w27182_,
		_w27183_,
		_w27184_
	);
	LUT3 #(
		.INIT('h12)
	) name21358 (
		_w26977_,
		_w26978_,
		_w26981_,
		_w27185_
	);
	LUT4 #(
		.INIT('he0f0)
	) name21359 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27186_
	);
	LUT3 #(
		.INIT('h02)
	) name21360 (
		_w26979_,
		_w27186_,
		_w27185_,
		_w27187_
	);
	LUT3 #(
		.INIT('h54)
	) name21361 (
		_w26976_,
		_w26978_,
		_w26979_,
		_w27188_
	);
	LUT2 #(
		.INIT('h8)
	) name21362 (
		_w26982_,
		_w27188_,
		_w27189_
	);
	LUT3 #(
		.INIT('h8a)
	) name21363 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w27190_
	);
	LUT3 #(
		.INIT('h15)
	) name21364 (
		_w26975_,
		_w27129_,
		_w27190_,
		_w27191_
	);
	LUT3 #(
		.INIT('h10)
	) name21365 (
		_w27189_,
		_w27187_,
		_w27191_,
		_w27192_
	);
	LUT3 #(
		.INIT('h02)
	) name21366 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w27193_
	);
	LUT3 #(
		.INIT('h08)
	) name21367 (
		_w26976_,
		_w26977_,
		_w26981_,
		_w27194_
	);
	LUT4 #(
		.INIT('hfe00)
	) name21368 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26979_,
		_w27195_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name21369 (
		_w26990_,
		_w27193_,
		_w27194_,
		_w27195_,
		_w27196_
	);
	LUT4 #(
		.INIT('h0010)
	) name21370 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27197_
	);
	LUT3 #(
		.INIT('h08)
	) name21371 (
		_w26975_,
		_w27182_,
		_w27197_,
		_w27198_
	);
	LUT3 #(
		.INIT('h20)
	) name21372 (
		_w26985_,
		_w27196_,
		_w27198_,
		_w27199_
	);
	LUT4 #(
		.INIT('h999a)
	) name21373 (
		\u0_L10_reg[13]/NET0131 ,
		_w27184_,
		_w27192_,
		_w27199_,
		_w27200_
	);
	LUT3 #(
		.INIT('h04)
	) name21374 (
		_w27045_,
		_w27048_,
		_w27046_,
		_w27201_
	);
	LUT4 #(
		.INIT('ha34f)
	) name21375 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27202_
	);
	LUT2 #(
		.INIT('h2)
	) name21376 (
		_w27044_,
		_w27202_,
		_w27203_
	);
	LUT3 #(
		.INIT('hf6)
	) name21377 (
		_w27045_,
		_w27048_,
		_w27046_,
		_w27204_
	);
	LUT2 #(
		.INIT('h2)
	) name21378 (
		_w27147_,
		_w27204_,
		_w27205_
	);
	LUT4 #(
		.INIT('h1200)
	) name21379 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27206_
	);
	LUT4 #(
		.INIT('h0400)
	) name21380 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27207_
	);
	LUT4 #(
		.INIT('h0007)
	) name21381 (
		_w27062_,
		_w27049_,
		_w27207_,
		_w27206_,
		_w27208_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name21382 (
		_w27043_,
		_w27205_,
		_w27203_,
		_w27208_,
		_w27209_
	);
	LUT4 #(
		.INIT('h2004)
	) name21383 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27210_
	);
	LUT4 #(
		.INIT('haa8a)
	) name21384 (
		_w27044_,
		_w27047_,
		_w27045_,
		_w27046_,
		_w27211_
	);
	LUT4 #(
		.INIT('h5ffc)
	) name21385 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27212_
	);
	LUT2 #(
		.INIT('h8)
	) name21386 (
		_w27211_,
		_w27212_,
		_w27213_
	);
	LUT4 #(
		.INIT('h5515)
	) name21387 (
		_w27044_,
		_w27047_,
		_w27045_,
		_w27048_,
		_w27214_
	);
	LUT4 #(
		.INIT('h4000)
	) name21388 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27215_
	);
	LUT4 #(
		.INIT('hbeff)
	) name21389 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27216_
	);
	LUT3 #(
		.INIT('h40)
	) name21390 (
		_w27201_,
		_w27214_,
		_w27216_,
		_w27217_
	);
	LUT4 #(
		.INIT('h4445)
	) name21391 (
		_w27043_,
		_w27210_,
		_w27213_,
		_w27217_,
		_w27218_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name21392 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27219_
	);
	LUT3 #(
		.INIT('hb1)
	) name21393 (
		_w27044_,
		_w27144_,
		_w27219_,
		_w27220_
	);
	LUT4 #(
		.INIT('h5655)
	) name21394 (
		\u0_L10_reg[14]/NET0131 ,
		_w27218_,
		_w27209_,
		_w27220_,
		_w27221_
	);
	LUT4 #(
		.INIT('h8228)
	) name21395 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w27222_
	);
	LUT3 #(
		.INIT('h43)
	) name21396 (
		_w26767_,
		_w26768_,
		_w26773_,
		_w27223_
	);
	LUT2 #(
		.INIT('h2)
	) name21397 (
		_w26770_,
		_w26771_,
		_w27224_
	);
	LUT4 #(
		.INIT('h0015)
	) name21398 (
		_w26869_,
		_w27223_,
		_w27224_,
		_w27222_,
		_w27225_
	);
	LUT2 #(
		.INIT('h2)
	) name21399 (
		_w26766_,
		_w27225_,
		_w27226_
	);
	LUT3 #(
		.INIT('h40)
	) name21400 (
		_w26771_,
		_w26767_,
		_w26773_,
		_w27227_
	);
	LUT3 #(
		.INIT('h28)
	) name21401 (
		_w26770_,
		_w26768_,
		_w26773_,
		_w27228_
	);
	LUT4 #(
		.INIT('h4000)
	) name21402 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w27229_
	);
	LUT3 #(
		.INIT('h0b)
	) name21403 (
		_w27227_,
		_w27228_,
		_w27229_,
		_w27230_
	);
	LUT4 #(
		.INIT('h1005)
	) name21404 (
		_w26770_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w27231_
	);
	LUT4 #(
		.INIT('h0082)
	) name21405 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w27232_
	);
	LUT2 #(
		.INIT('h1)
	) name21406 (
		_w27231_,
		_w27232_,
		_w27233_
	);
	LUT4 #(
		.INIT('h9fff)
	) name21407 (
		_w26771_,
		_w26767_,
		_w26768_,
		_w26773_,
		_w27234_
	);
	LUT2 #(
		.INIT('h1)
	) name21408 (
		_w26770_,
		_w27234_,
		_w27235_
	);
	LUT4 #(
		.INIT('h00ea)
	) name21409 (
		_w26766_,
		_w27230_,
		_w27233_,
		_w27235_,
		_w27236_
	);
	LUT3 #(
		.INIT('h65)
	) name21410 (
		\u0_L10_reg[9]/NET0131 ,
		_w27226_,
		_w27236_,
		_w27237_
	);
	LUT4 #(
		.INIT('hf32e)
	) name21411 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27238_
	);
	LUT2 #(
		.INIT('h1)
	) name21412 (
		_w26935_,
		_w27238_,
		_w27239_
	);
	LUT4 #(
		.INIT('hef6f)
	) name21413 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27240_
	);
	LUT2 #(
		.INIT('h6)
	) name21414 (
		_w26928_,
		_w26930_,
		_w27241_
	);
	LUT4 #(
		.INIT('hc400)
	) name21415 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26935_,
		_w27242_
	);
	LUT4 #(
		.INIT('h4500)
	) name21416 (
		_w26941_,
		_w27241_,
		_w27242_,
		_w27240_,
		_w27243_
	);
	LUT3 #(
		.INIT('h8a)
	) name21417 (
		_w26939_,
		_w27239_,
		_w27243_,
		_w27244_
	);
	LUT4 #(
		.INIT('hb0b8)
	) name21418 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27245_
	);
	LUT4 #(
		.INIT('hfb00)
	) name21419 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26935_,
		_w27246_
	);
	LUT4 #(
		.INIT('h4544)
	) name21420 (
		_w26939_,
		_w26951_,
		_w27245_,
		_w27246_,
		_w27247_
	);
	LUT4 #(
		.INIT('heff7)
	) name21421 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26930_,
		_w27248_
	);
	LUT2 #(
		.INIT('h1)
	) name21422 (
		_w26935_,
		_w27248_,
		_w27249_
	);
	LUT4 #(
		.INIT('h0080)
	) name21423 (
		_w26926_,
		_w26928_,
		_w26930_,
		_w26935_,
		_w27250_
	);
	LUT3 #(
		.INIT('h54)
	) name21424 (
		_w26939_,
		_w27025_,
		_w27250_,
		_w27251_
	);
	LUT4 #(
		.INIT('h0200)
	) name21425 (
		_w26926_,
		_w26927_,
		_w26928_,
		_w26935_,
		_w27252_
	);
	LUT3 #(
		.INIT('h07)
	) name21426 (
		_w26932_,
		_w26947_,
		_w27252_,
		_w27253_
	);
	LUT4 #(
		.INIT('h0100)
	) name21427 (
		_w27247_,
		_w27249_,
		_w27251_,
		_w27253_,
		_w27254_
	);
	LUT3 #(
		.INIT('h65)
	) name21428 (
		\u0_L10_reg[27]/NET0131 ,
		_w27244_,
		_w27254_,
		_w27255_
	);
	LUT3 #(
		.INIT('h21)
	) name21429 (
		_w26800_,
		_w26798_,
		_w26801_,
		_w27256_
	);
	LUT4 #(
		.INIT('hf6ad)
	) name21430 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27257_
	);
	LUT2 #(
		.INIT('h1)
	) name21431 (
		_w26805_,
		_w27257_,
		_w27258_
	);
	LUT2 #(
		.INIT('h2)
	) name21432 (
		_w26798_,
		_w26801_,
		_w27259_
	);
	LUT3 #(
		.INIT('ha8)
	) name21433 (
		_w26800_,
		_w26799_,
		_w26805_,
		_w27260_
	);
	LUT4 #(
		.INIT('hcffa)
	) name21434 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27261_
	);
	LUT4 #(
		.INIT('h3f15)
	) name21435 (
		_w26805_,
		_w27259_,
		_w27260_,
		_w27261_,
		_w27262_
	);
	LUT3 #(
		.INIT('h8a)
	) name21436 (
		_w26804_,
		_w27258_,
		_w27262_,
		_w27263_
	);
	LUT3 #(
		.INIT('hb5)
	) name21437 (
		_w26798_,
		_w26799_,
		_w26801_,
		_w27264_
	);
	LUT2 #(
		.INIT('h8)
	) name21438 (
		_w27260_,
		_w27264_,
		_w27265_
	);
	LUT3 #(
		.INIT('ha2)
	) name21439 (
		_w26810_,
		_w27160_,
		_w27163_,
		_w27266_
	);
	LUT4 #(
		.INIT('h9fbf)
	) name21440 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27267_
	);
	LUT3 #(
		.INIT('h72)
	) name21441 (
		_w26805_,
		_w26809_,
		_w27267_,
		_w27268_
	);
	LUT4 #(
		.INIT('hba00)
	) name21442 (
		_w26804_,
		_w27265_,
		_w27266_,
		_w27268_,
		_w27269_
	);
	LUT3 #(
		.INIT('h65)
	) name21443 (
		\u0_L10_reg[32]/NET0131 ,
		_w27263_,
		_w27269_,
		_w27270_
	);
	LUT4 #(
		.INIT('hc693)
	) name21444 (
		decrypt_pad,
		\u0_R10_reg[11]/NET0131 ,
		\u0_uk_K_r10_reg[26]/NET0131 ,
		\u0_uk_K_r10_reg[3]/NET0131 ,
		_w27271_
	);
	LUT4 #(
		.INIT('hc963)
	) name21445 (
		decrypt_pad,
		\u0_R10_reg[12]/NET0131 ,
		\u0_uk_K_r10_reg[18]/NET0131 ,
		\u0_uk_K_r10_reg[41]/P0001 ,
		_w27272_
	);
	LUT4 #(
		.INIT('hc693)
	) name21446 (
		decrypt_pad,
		\u0_R10_reg[13]/NET0131 ,
		\u0_uk_K_r10_reg[54]/NET0131 ,
		\u0_uk_K_r10_reg[6]/NET0131 ,
		_w27273_
	);
	LUT4 #(
		.INIT('hc693)
	) name21447 (
		decrypt_pad,
		\u0_R10_reg[9]/NET0131 ,
		\u0_uk_K_r10_reg[17]/NET0131 ,
		\u0_uk_K_r10_reg[26]/NET0131 ,
		_w27274_
	);
	LUT4 #(
		.INIT('hc693)
	) name21448 (
		decrypt_pad,
		\u0_R10_reg[8]/NET0131 ,
		\u0_uk_K_r10_reg[20]/NET0131 ,
		\u0_uk_K_r10_reg[54]/NET0131 ,
		_w27275_
	);
	LUT4 #(
		.INIT('hc693)
	) name21449 (
		decrypt_pad,
		\u0_R10_reg[10]/NET0131 ,
		\u0_uk_K_r10_reg[25]/NET0131 ,
		\u0_uk_K_r10_reg[34]/NET0131 ,
		_w27276_
	);
	LUT4 #(
		.INIT('h95b5)
	) name21450 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27277_
	);
	LUT2 #(
		.INIT('h1)
	) name21451 (
		_w27273_,
		_w27275_,
		_w27278_
	);
	LUT4 #(
		.INIT('h0001)
	) name21452 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27279_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name21453 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27280_
	);
	LUT4 #(
		.INIT('h08cc)
	) name21454 (
		_w27272_,
		_w27271_,
		_w27277_,
		_w27280_,
		_w27281_
	);
	LUT2 #(
		.INIT('h8)
	) name21455 (
		_w27273_,
		_w27275_,
		_w27282_
	);
	LUT2 #(
		.INIT('h6)
	) name21456 (
		_w27273_,
		_w27275_,
		_w27283_
	);
	LUT4 #(
		.INIT('h000d)
	) name21457 (
		_w27271_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27284_
	);
	LUT4 #(
		.INIT('h0020)
	) name21458 (
		_w27271_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27285_
	);
	LUT4 #(
		.INIT('h4000)
	) name21459 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27286_
	);
	LUT4 #(
		.INIT('h0103)
	) name21460 (
		_w27283_,
		_w27285_,
		_w27286_,
		_w27284_,
		_w27287_
	);
	LUT3 #(
		.INIT('h20)
	) name21461 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27288_
	);
	LUT4 #(
		.INIT('h2000)
	) name21462 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27289_
	);
	LUT4 #(
		.INIT('h9990)
	) name21463 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27290_
	);
	LUT4 #(
		.INIT('h0990)
	) name21464 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27291_
	);
	LUT3 #(
		.INIT('h0b)
	) name21465 (
		_w27271_,
		_w27289_,
		_w27291_,
		_w27292_
	);
	LUT3 #(
		.INIT('h80)
	) name21466 (
		_w27272_,
		_w27274_,
		_w27276_,
		_w27293_
	);
	LUT3 #(
		.INIT('h80)
	) name21467 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27294_
	);
	LUT4 #(
		.INIT('h7b5b)
	) name21468 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27295_
	);
	LUT2 #(
		.INIT('h2)
	) name21469 (
		_w27272_,
		_w27271_,
		_w27296_
	);
	LUT4 #(
		.INIT('h7077)
	) name21470 (
		_w27278_,
		_w27293_,
		_w27295_,
		_w27296_,
		_w27297_
	);
	LUT4 #(
		.INIT('hea00)
	) name21471 (
		_w27272_,
		_w27287_,
		_w27292_,
		_w27297_,
		_w27298_
	);
	LUT3 #(
		.INIT('h65)
	) name21472 (
		\u0_L10_reg[6]/NET0131 ,
		_w27281_,
		_w27298_,
		_w27299_
	);
	LUT3 #(
		.INIT('h02)
	) name21473 (
		_w27044_,
		_w27141_,
		_w27136_,
		_w27300_
	);
	LUT4 #(
		.INIT('h2000)
	) name21474 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27301_
	);
	LUT4 #(
		.INIT('h0001)
	) name21475 (
		_w27044_,
		_w27145_,
		_w27207_,
		_w27301_,
		_w27302_
	);
	LUT2 #(
		.INIT('h1)
	) name21476 (
		_w27300_,
		_w27302_,
		_w27303_
	);
	LUT4 #(
		.INIT('h1510)
	) name21477 (
		_w27044_,
		_w27047_,
		_w27048_,
		_w27046_,
		_w27304_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name21478 (
		_w27044_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27305_
	);
	LUT4 #(
		.INIT('h8acf)
	) name21479 (
		_w27060_,
		_w27051_,
		_w27304_,
		_w27305_,
		_w27306_
	);
	LUT4 #(
		.INIT('h2022)
	) name21480 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27307_
	);
	LUT2 #(
		.INIT('h1)
	) name21481 (
		_w27043_,
		_w27307_,
		_w27308_
	);
	LUT4 #(
		.INIT('haff3)
	) name21482 (
		_w27047_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27309_
	);
	LUT2 #(
		.INIT('h2)
	) name21483 (
		_w27044_,
		_w27309_,
		_w27310_
	);
	LUT4 #(
		.INIT('h0040)
	) name21484 (
		_w27044_,
		_w27045_,
		_w27048_,
		_w27046_,
		_w27311_
	);
	LUT4 #(
		.INIT('h0002)
	) name21485 (
		_w27043_,
		_w27140_,
		_w27215_,
		_w27311_,
		_w27312_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name21486 (
		_w27306_,
		_w27308_,
		_w27310_,
		_w27312_,
		_w27313_
	);
	LUT3 #(
		.INIT('h56)
	) name21487 (
		\u0_L10_reg[3]/NET0131 ,
		_w27303_,
		_w27313_,
		_w27314_
	);
	LUT4 #(
		.INIT('hae16)
	) name21488 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27315_
	);
	LUT2 #(
		.INIT('h1)
	) name21489 (
		_w26805_,
		_w27315_,
		_w27316_
	);
	LUT4 #(
		.INIT('h4880)
	) name21490 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27317_
	);
	LUT4 #(
		.INIT('h2210)
	) name21491 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27318_
	);
	LUT4 #(
		.INIT('h002a)
	) name21492 (
		_w26804_,
		_w26805_,
		_w27318_,
		_w27317_,
		_w27319_
	);
	LUT4 #(
		.INIT('h4080)
	) name21493 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27320_
	);
	LUT4 #(
		.INIT('hdf00)
	) name21494 (
		_w26800_,
		_w26799_,
		_w26801_,
		_w26805_,
		_w27321_
	);
	LUT4 #(
		.INIT('h5455)
	) name21495 (
		_w26804_,
		_w27256_,
		_w27320_,
		_w27321_,
		_w27322_
	);
	LUT3 #(
		.INIT('h0b)
	) name21496 (
		_w27316_,
		_w27319_,
		_w27322_,
		_w27323_
	);
	LUT2 #(
		.INIT('h2)
	) name21497 (
		_w26805_,
		_w26819_,
		_w27324_
	);
	LUT4 #(
		.INIT('hddeb)
	) name21498 (
		_w26800_,
		_w26798_,
		_w26799_,
		_w26801_,
		_w27325_
	);
	LUT4 #(
		.INIT('h0302)
	) name21499 (
		_w26804_,
		_w26805_,
		_w27317_,
		_w27325_,
		_w27326_
	);
	LUT2 #(
		.INIT('h1)
	) name21500 (
		_w27324_,
		_w27326_,
		_w27327_
	);
	LUT3 #(
		.INIT('h56)
	) name21501 (
		\u0_L10_reg[7]/NET0131 ,
		_w27323_,
		_w27327_,
		_w27328_
	);
	LUT3 #(
		.INIT('h1d)
	) name21502 (
		_w26976_,
		_w26978_,
		_w26979_,
		_w27329_
	);
	LUT3 #(
		.INIT('h0b)
	) name21503 (
		_w26976_,
		_w26978_,
		_w26981_,
		_w27330_
	);
	LUT4 #(
		.INIT('hdefe)
	) name21504 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w26981_,
		_w27331_
	);
	LUT4 #(
		.INIT('h3500)
	) name21505 (
		_w26988_,
		_w27330_,
		_w27329_,
		_w27331_,
		_w27332_
	);
	LUT2 #(
		.INIT('h1)
	) name21506 (
		_w26975_,
		_w27332_,
		_w27333_
	);
	LUT4 #(
		.INIT('h4060)
	) name21507 (
		_w26977_,
		_w26978_,
		_w26979_,
		_w26981_,
		_w27334_
	);
	LUT3 #(
		.INIT('ha8)
	) name21508 (
		_w26975_,
		_w26998_,
		_w27334_,
		_w27335_
	);
	LUT3 #(
		.INIT('hb8)
	) name21509 (
		_w26976_,
		_w26977_,
		_w26978_,
		_w27336_
	);
	LUT2 #(
		.INIT('h8)
	) name21510 (
		_w26975_,
		_w26981_,
		_w27337_
	);
	LUT4 #(
		.INIT('h4544)
	) name21511 (
		_w26979_,
		_w26983_,
		_w27336_,
		_w27337_,
		_w27338_
	);
	LUT4 #(
		.INIT('h80b0)
	) name21512 (
		_w26976_,
		_w26977_,
		_w26979_,
		_w26981_,
		_w27339_
	);
	LUT2 #(
		.INIT('h4)
	) name21513 (
		_w27330_,
		_w27339_,
		_w27340_
	);
	LUT3 #(
		.INIT('h01)
	) name21514 (
		_w27338_,
		_w27335_,
		_w27340_,
		_w27341_
	);
	LUT3 #(
		.INIT('h65)
	) name21515 (
		\u0_L10_reg[18]/NET0131 ,
		_w27333_,
		_w27341_,
		_w27342_
	);
	LUT4 #(
		.INIT('h3dc3)
	) name21516 (
		_w27271_,
		_w27273_,
		_w27275_,
		_w27274_,
		_w27343_
	);
	LUT4 #(
		.INIT('h0110)
	) name21517 (
		_w27271_,
		_w27273_,
		_w27275_,
		_w27276_,
		_w27344_
	);
	LUT4 #(
		.INIT('h0074)
	) name21518 (
		_w27288_,
		_w27276_,
		_w27343_,
		_w27344_,
		_w27345_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name21519 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27346_
	);
	LUT4 #(
		.INIT('h2880)
	) name21520 (
		_w27271_,
		_w27273_,
		_w27275_,
		_w27274_,
		_w27347_
	);
	LUT4 #(
		.INIT('h0032)
	) name21521 (
		_w27271_,
		_w27279_,
		_w27346_,
		_w27347_,
		_w27348_
	);
	LUT4 #(
		.INIT('hbeff)
	) name21522 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27349_
	);
	LUT4 #(
		.INIT('h0400)
	) name21523 (
		_w27271_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27350_
	);
	LUT3 #(
		.INIT('h0d)
	) name21524 (
		_w27271_,
		_w27349_,
		_w27350_,
		_w27351_
	);
	LUT4 #(
		.INIT('he400)
	) name21525 (
		_w27272_,
		_w27348_,
		_w27345_,
		_w27351_,
		_w27352_
	);
	LUT2 #(
		.INIT('h9)
	) name21526 (
		\u0_L10_reg[16]/NET0131 ,
		_w27352_,
		_w27353_
	);
	LUT2 #(
		.INIT('h4)
	) name21527 (
		_w27271_,
		_w27290_,
		_w27354_
	);
	LUT4 #(
		.INIT('h1dff)
	) name21528 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27355_
	);
	LUT2 #(
		.INIT('h2)
	) name21529 (
		_w27271_,
		_w27355_,
		_w27356_
	);
	LUT2 #(
		.INIT('h2)
	) name21530 (
		_w27271_,
		_w27276_,
		_w27357_
	);
	LUT3 #(
		.INIT('h0d)
	) name21531 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27358_
	);
	LUT4 #(
		.INIT('h0777)
	) name21532 (
		_w27283_,
		_w27284_,
		_w27357_,
		_w27358_,
		_w27359_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name21533 (
		_w27272_,
		_w27356_,
		_w27354_,
		_w27359_,
		_w27360_
	);
	LUT4 #(
		.INIT('he2cd)
	) name21534 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27361_
	);
	LUT4 #(
		.INIT('h0400)
	) name21535 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27362_
	);
	LUT4 #(
		.INIT('h5504)
	) name21536 (
		_w27272_,
		_w27271_,
		_w27361_,
		_w27362_,
		_w27363_
	);
	LUT4 #(
		.INIT('h0009)
	) name21537 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27364_
	);
	LUT4 #(
		.INIT('h9db6)
	) name21538 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27365_
	);
	LUT2 #(
		.INIT('h1)
	) name21539 (
		_w27272_,
		_w27271_,
		_w27366_
	);
	LUT2 #(
		.INIT('h4)
	) name21540 (
		_w27365_,
		_w27366_,
		_w27367_
	);
	LUT3 #(
		.INIT('hdb)
	) name21541 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27368_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name21542 (
		_w27271_,
		_w27276_,
		_w27294_,
		_w27368_,
		_w27369_
	);
	LUT3 #(
		.INIT('h10)
	) name21543 (
		_w27363_,
		_w27367_,
		_w27369_,
		_w27370_
	);
	LUT3 #(
		.INIT('h65)
	) name21544 (
		\u0_L10_reg[24]/NET0131 ,
		_w27360_,
		_w27370_,
		_w27371_
	);
	LUT4 #(
		.INIT('h0200)
	) name21545 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27372_
	);
	LUT3 #(
		.INIT('h01)
	) name21546 (
		_w27272_,
		_w27364_,
		_w27372_,
		_w27373_
	);
	LUT2 #(
		.INIT('h8)
	) name21547 (
		_w27275_,
		_w27276_,
		_w27374_
	);
	LUT4 #(
		.INIT('h73af)
	) name21548 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27375_
	);
	LUT4 #(
		.INIT('hdf53)
	) name21549 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27376_
	);
	LUT3 #(
		.INIT('hd8)
	) name21550 (
		_w27271_,
		_w27375_,
		_w27376_,
		_w27377_
	);
	LUT4 #(
		.INIT('heed9)
	) name21551 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27378_
	);
	LUT4 #(
		.INIT('h23ef)
	) name21552 (
		_w27273_,
		_w27275_,
		_w27274_,
		_w27276_,
		_w27379_
	);
	LUT4 #(
		.INIT('ha820)
	) name21553 (
		_w27272_,
		_w27271_,
		_w27379_,
		_w27378_,
		_w27380_
	);
	LUT3 #(
		.INIT('h07)
	) name21554 (
		_w27373_,
		_w27377_,
		_w27380_,
		_w27381_
	);
	LUT3 #(
		.INIT('h08)
	) name21555 (
		_w27271_,
		_w27273_,
		_w27274_,
		_w27382_
	);
	LUT2 #(
		.INIT('h8)
	) name21556 (
		_w27374_,
		_w27382_,
		_w27383_
	);
	LUT4 #(
		.INIT('h1000)
	) name21557 (
		_w27271_,
		_w27273_,
		_w27274_,
		_w27276_,
		_w27384_
	);
	LUT3 #(
		.INIT('h0b)
	) name21558 (
		_w27282_,
		_w27293_,
		_w27384_,
		_w27385_
	);
	LUT2 #(
		.INIT('h4)
	) name21559 (
		_w27383_,
		_w27385_,
		_w27386_
	);
	LUT3 #(
		.INIT('h9a)
	) name21560 (
		\u0_L10_reg[30]/NET0131 ,
		_w27381_,
		_w27386_,
		_w27387_
	);
	LUT4 #(
		.INIT('hc963)
	) name21561 (
		decrypt_pad,
		\u0_R9_reg[27]/NET0131 ,
		\u0_uk_K_r9_reg[16]/NET0131 ,
		\u0_uk_K_r9_reg[8]/NET0131 ,
		_w27388_
	);
	LUT4 #(
		.INIT('hc693)
	) name21562 (
		decrypt_pad,
		\u0_R9_reg[26]/NET0131 ,
		\u0_uk_K_r9_reg[30]/NET0131 ,
		\u0_uk_K_r9_reg[7]/NET0131 ,
		_w27389_
	);
	LUT4 #(
		.INIT('hc693)
	) name21563 (
		decrypt_pad,
		\u0_R9_reg[24]/NET0131 ,
		\u0_uk_K_r9_reg[38]/NET0131 ,
		\u0_uk_K_r9_reg[42]/NET0131 ,
		_w27390_
	);
	LUT4 #(
		.INIT('hc693)
	) name21564 (
		decrypt_pad,
		\u0_R9_reg[25]/NET0131 ,
		\u0_uk_K_r9_reg[14]/NET0131 ,
		\u0_uk_K_r9_reg[22]/NET0131 ,
		_w27391_
	);
	LUT4 #(
		.INIT('hc693)
	) name21565 (
		decrypt_pad,
		\u0_R9_reg[29]/NET0131 ,
		\u0_uk_K_r9_reg[42]/NET0131 ,
		\u0_uk_K_r9_reg[50]/NET0131 ,
		_w27392_
	);
	LUT4 #(
		.INIT('h0002)
	) name21566 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27393_
	);
	LUT2 #(
		.INIT('h6)
	) name21567 (
		_w27389_,
		_w27390_,
		_w27394_
	);
	LUT4 #(
		.INIT('h5a2d)
	) name21568 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27395_
	);
	LUT2 #(
		.INIT('h8)
	) name21569 (
		_w27388_,
		_w27390_,
		_w27396_
	);
	LUT4 #(
		.INIT('h0200)
	) name21570 (
		_w27388_,
		_w27389_,
		_w27391_,
		_w27390_,
		_w27397_
	);
	LUT4 #(
		.INIT('h8400)
	) name21571 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27398_
	);
	LUT4 #(
		.INIT('h000e)
	) name21572 (
		_w27388_,
		_w27395_,
		_w27397_,
		_w27398_,
		_w27399_
	);
	LUT4 #(
		.INIT('hc963)
	) name21573 (
		decrypt_pad,
		\u0_R9_reg[28]/NET0131 ,
		\u0_uk_K_r9_reg[31]/P0001 ,
		\u0_uk_K_r9_reg[50]/NET0131 ,
		_w27400_
	);
	LUT2 #(
		.INIT('h1)
	) name21574 (
		_w27399_,
		_w27400_,
		_w27401_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name21575 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27402_
	);
	LUT4 #(
		.INIT('h1400)
	) name21576 (
		_w27388_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27403_
	);
	LUT2 #(
		.INIT('h4)
	) name21577 (
		_w27402_,
		_w27403_,
		_w27404_
	);
	LUT3 #(
		.INIT('h9d)
	) name21578 (
		_w27389_,
		_w27391_,
		_w27392_,
		_w27405_
	);
	LUT4 #(
		.INIT('h0200)
	) name21579 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27406_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name21580 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27407_
	);
	LUT3 #(
		.INIT('hd0)
	) name21581 (
		_w27396_,
		_w27405_,
		_w27407_,
		_w27408_
	);
	LUT4 #(
		.INIT('h0208)
	) name21582 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27409_
	);
	LUT4 #(
		.INIT('hfdc6)
	) name21583 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27410_
	);
	LUT4 #(
		.INIT('h4010)
	) name21584 (
		_w27388_,
		_w27389_,
		_w27391_,
		_w27390_,
		_w27411_
	);
	LUT3 #(
		.INIT('h0d)
	) name21585 (
		_w27388_,
		_w27410_,
		_w27411_,
		_w27412_
	);
	LUT4 #(
		.INIT('h7500)
	) name21586 (
		_w27400_,
		_w27404_,
		_w27408_,
		_w27412_,
		_w27413_
	);
	LUT3 #(
		.INIT('h65)
	) name21587 (
		\u0_L9_reg[22]/NET0131 ,
		_w27401_,
		_w27413_,
		_w27414_
	);
	LUT4 #(
		.INIT('hc693)
	) name21588 (
		decrypt_pad,
		\u0_R9_reg[4]/NET0131 ,
		\u0_uk_K_r9_reg[19]/NET0131 ,
		\u0_uk_K_r9_reg[25]/NET0131 ,
		_w27415_
	);
	LUT4 #(
		.INIT('hc693)
	) name21589 (
		decrypt_pad,
		\u0_R9_reg[3]/NET0131 ,
		\u0_uk_K_r9_reg[41]/NET0131 ,
		\u0_uk_K_r9_reg[47]/NET0131 ,
		_w27416_
	);
	LUT4 #(
		.INIT('hc693)
	) name21590 (
		decrypt_pad,
		\u0_R9_reg[1]/NET0131 ,
		\u0_uk_K_r9_reg[17]/NET0131 ,
		\u0_uk_K_r9_reg[55]/NET0131 ,
		_w27417_
	);
	LUT4 #(
		.INIT('hc693)
	) name21591 (
		decrypt_pad,
		\u0_R9_reg[5]/NET0131 ,
		\u0_uk_K_r9_reg[47]/NET0131 ,
		\u0_uk_K_r9_reg[53]/NET0131 ,
		_w27418_
	);
	LUT4 #(
		.INIT('hc963)
	) name21592 (
		decrypt_pad,
		\u0_R9_reg[2]/NET0131 ,
		\u0_uk_K_r9_reg[13]/NET0131 ,
		\u0_uk_K_r9_reg[32]/NET0131 ,
		_w27419_
	);
	LUT4 #(
		.INIT('hc963)
	) name21593 (
		decrypt_pad,
		\u0_R9_reg[32]/NET0131 ,
		\u0_uk_K_r9_reg[34]/NET0131 ,
		\u0_uk_K_r9_reg[53]/NET0131 ,
		_w27420_
	);
	LUT4 #(
		.INIT('hf0dd)
	) name21594 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27421_
	);
	LUT2 #(
		.INIT('h2)
	) name21595 (
		_w27416_,
		_w27421_,
		_w27422_
	);
	LUT4 #(
		.INIT('hafac)
	) name21596 (
		_w27416_,
		_w27419_,
		_w27417_,
		_w27418_,
		_w27423_
	);
	LUT2 #(
		.INIT('h2)
	) name21597 (
		_w27416_,
		_w27419_,
		_w27424_
	);
	LUT3 #(
		.INIT('hd0)
	) name21598 (
		_w27416_,
		_w27419_,
		_w27417_,
		_w27425_
	);
	LUT3 #(
		.INIT('h32)
	) name21599 (
		_w27419_,
		_w27420_,
		_w27418_,
		_w27426_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name21600 (
		_w27420_,
		_w27423_,
		_w27425_,
		_w27426_,
		_w27427_
	);
	LUT3 #(
		.INIT('h8a)
	) name21601 (
		_w27415_,
		_w27422_,
		_w27427_,
		_w27428_
	);
	LUT4 #(
		.INIT('hefe6)
	) name21602 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27429_
	);
	LUT2 #(
		.INIT('h1)
	) name21603 (
		_w27416_,
		_w27429_,
		_w27430_
	);
	LUT2 #(
		.INIT('h1)
	) name21604 (
		_w27420_,
		_w27418_,
		_w27431_
	);
	LUT3 #(
		.INIT('h48)
	) name21605 (
		_w27420_,
		_w27417_,
		_w27418_,
		_w27432_
	);
	LUT4 #(
		.INIT('h73cf)
	) name21606 (
		_w27416_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27433_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name21607 (
		_w27416_,
		_w27419_,
		_w27432_,
		_w27433_,
		_w27434_
	);
	LUT3 #(
		.INIT('h45)
	) name21608 (
		_w27415_,
		_w27430_,
		_w27434_,
		_w27435_
	);
	LUT4 #(
		.INIT('h7daf)
	) name21609 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27436_
	);
	LUT2 #(
		.INIT('h1)
	) name21610 (
		_w27416_,
		_w27436_,
		_w27437_
	);
	LUT4 #(
		.INIT('h0020)
	) name21611 (
		_w27416_,
		_w27419_,
		_w27420_,
		_w27417_,
		_w27438_
	);
	LUT3 #(
		.INIT('h08)
	) name21612 (
		_w27416_,
		_w27419_,
		_w27417_,
		_w27439_
	);
	LUT3 #(
		.INIT('h15)
	) name21613 (
		_w27438_,
		_w27431_,
		_w27439_,
		_w27440_
	);
	LUT2 #(
		.INIT('h4)
	) name21614 (
		_w27437_,
		_w27440_,
		_w27441_
	);
	LUT4 #(
		.INIT('h5655)
	) name21615 (
		\u0_L9_reg[31]/NET0131 ,
		_w27435_,
		_w27428_,
		_w27441_,
		_w27442_
	);
	LUT4 #(
		.INIT('hc693)
	) name21616 (
		decrypt_pad,
		\u0_R9_reg[24]/NET0131 ,
		\u0_uk_K_r9_reg[43]/NET0131 ,
		\u0_uk_K_r9_reg[51]/NET0131 ,
		_w27443_
	);
	LUT4 #(
		.INIT('hc693)
	) name21617 (
		decrypt_pad,
		\u0_R9_reg[23]/NET0131 ,
		\u0_uk_K_r9_reg[45]/NET0131 ,
		\u0_uk_K_r9_reg[49]/NET0131 ,
		_w27444_
	);
	LUT4 #(
		.INIT('hc963)
	) name21618 (
		decrypt_pad,
		\u0_R9_reg[21]/NET0131 ,
		\u0_uk_K_r9_reg[14]/NET0131 ,
		\u0_uk_K_r9_reg[37]/NET0131 ,
		_w27445_
	);
	LUT4 #(
		.INIT('hc693)
	) name21619 (
		decrypt_pad,
		\u0_R9_reg[22]/NET0131 ,
		\u0_uk_K_r9_reg[28]/NET0131 ,
		\u0_uk_K_r9_reg[36]/NET0131 ,
		_w27446_
	);
	LUT4 #(
		.INIT('hc693)
	) name21620 (
		decrypt_pad,
		\u0_R9_reg[20]/NET0131 ,
		\u0_uk_K_r9_reg[22]/NET0131 ,
		\u0_uk_K_r9_reg[30]/NET0131 ,
		_w27447_
	);
	LUT4 #(
		.INIT('hc963)
	) name21621 (
		decrypt_pad,
		\u0_R9_reg[25]/NET0131 ,
		\u0_uk_K_r9_reg[15]/NET0131 ,
		\u0_uk_K_r9_reg[7]/NET0131 ,
		_w27448_
	);
	LUT3 #(
		.INIT('hd0)
	) name21622 (
		_w27445_,
		_w27448_,
		_w27447_,
		_w27449_
	);
	LUT4 #(
		.INIT('h3e77)
	) name21623 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27450_
	);
	LUT2 #(
		.INIT('h2)
	) name21624 (
		_w27444_,
		_w27450_,
		_w27451_
	);
	LUT4 #(
		.INIT('ha088)
	) name21625 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27452_
	);
	LUT4 #(
		.INIT('h5515)
	) name21626 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27453_
	);
	LUT3 #(
		.INIT('h01)
	) name21627 (
		_w27444_,
		_w27453_,
		_w27452_,
		_w27454_
	);
	LUT2 #(
		.INIT('h1)
	) name21628 (
		_w27446_,
		_w27444_,
		_w27455_
	);
	LUT4 #(
		.INIT('h1000)
	) name21629 (
		_w27446_,
		_w27444_,
		_w27448_,
		_w27447_,
		_w27456_
	);
	LUT2 #(
		.INIT('h4)
	) name21630 (
		_w27445_,
		_w27456_,
		_w27457_
	);
	LUT4 #(
		.INIT('haaa8)
	) name21631 (
		_w27443_,
		_w27454_,
		_w27451_,
		_w27457_,
		_w27458_
	);
	LUT4 #(
		.INIT('h0408)
	) name21632 (
		_w27446_,
		_w27445_,
		_w27444_,
		_w27447_,
		_w27459_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name21633 (
		_w27446_,
		_w27445_,
		_w27444_,
		_w27448_,
		_w27460_
	);
	LUT4 #(
		.INIT('hef00)
	) name21634 (
		_w27446_,
		_w27445_,
		_w27444_,
		_w27447_,
		_w27461_
	);
	LUT2 #(
		.INIT('h4)
	) name21635 (
		_w27460_,
		_w27461_,
		_w27462_
	);
	LUT4 #(
		.INIT('h2000)
	) name21636 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27463_
	);
	LUT3 #(
		.INIT('h04)
	) name21637 (
		_w27446_,
		_w27444_,
		_w27447_,
		_w27464_
	);
	LUT4 #(
		.INIT('h0040)
	) name21638 (
		_w27445_,
		_w27444_,
		_w27448_,
		_w27447_,
		_w27465_
	);
	LUT3 #(
		.INIT('h01)
	) name21639 (
		_w27463_,
		_w27464_,
		_w27465_,
		_w27466_
	);
	LUT4 #(
		.INIT('h00ef)
	) name21640 (
		_w27462_,
		_w27459_,
		_w27466_,
		_w27443_,
		_w27467_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name21641 (
		_w27445_,
		_w27444_,
		_w27448_,
		_w27447_,
		_w27468_
	);
	LUT2 #(
		.INIT('h1)
	) name21642 (
		_w27446_,
		_w27468_,
		_w27469_
	);
	LUT4 #(
		.INIT('h0004)
	) name21643 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27470_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name21644 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27471_
	);
	LUT4 #(
		.INIT('h0001)
	) name21645 (
		_w27446_,
		_w27444_,
		_w27448_,
		_w27447_,
		_w27472_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name21646 (
		_w27445_,
		_w27444_,
		_w27471_,
		_w27472_,
		_w27473_
	);
	LUT2 #(
		.INIT('h4)
	) name21647 (
		_w27469_,
		_w27473_,
		_w27474_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name21648 (
		\u0_L9_reg[11]/NET0131 ,
		_w27467_,
		_w27458_,
		_w27474_,
		_w27475_
	);
	LUT4 #(
		.INIT('hc693)
	) name21649 (
		decrypt_pad,
		\u0_R9_reg[12]/NET0131 ,
		\u0_uk_K_r9_reg[10]/NET0131 ,
		\u0_uk_K_r9_reg[48]/NET0131 ,
		_w27476_
	);
	LUT4 #(
		.INIT('hc963)
	) name21650 (
		decrypt_pad,
		\u0_R9_reg[13]/NET0131 ,
		\u0_uk_K_r9_reg[10]/NET0131 ,
		\u0_uk_K_r9_reg[4]/NET0131 ,
		_w27477_
	);
	LUT4 #(
		.INIT('hc693)
	) name21651 (
		decrypt_pad,
		\u0_R9_reg[17]/NET0131 ,
		\u0_uk_K_r9_reg[26]/NET0131 ,
		\u0_uk_K_r9_reg[32]/NET0131 ,
		_w27478_
	);
	LUT2 #(
		.INIT('h4)
	) name21652 (
		_w27476_,
		_w27478_,
		_w27479_
	);
	LUT4 #(
		.INIT('hc693)
	) name21653 (
		decrypt_pad,
		\u0_R9_reg[15]/NET0131 ,
		\u0_uk_K_r9_reg[13]/NET0131 ,
		\u0_uk_K_r9_reg[19]/NET0131 ,
		_w27480_
	);
	LUT4 #(
		.INIT('h7e00)
	) name21654 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27480_,
		_w27481_
	);
	LUT4 #(
		.INIT('hc963)
	) name21655 (
		decrypt_pad,
		\u0_R9_reg[14]/NET0131 ,
		\u0_uk_K_r9_reg[11]/NET0131 ,
		\u0_uk_K_r9_reg[5]/NET0131 ,
		_w27482_
	);
	LUT3 #(
		.INIT('h20)
	) name21656 (
		_w27476_,
		_w27478_,
		_w27482_,
		_w27483_
	);
	LUT3 #(
		.INIT('h0b)
	) name21657 (
		_w27477_,
		_w27478_,
		_w27480_,
		_w27484_
	);
	LUT3 #(
		.INIT('h45)
	) name21658 (
		_w27481_,
		_w27483_,
		_w27484_,
		_w27485_
	);
	LUT3 #(
		.INIT('h04)
	) name21659 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27486_
	);
	LUT4 #(
		.INIT('h0400)
	) name21660 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27487_
	);
	LUT3 #(
		.INIT('h01)
	) name21661 (
		_w27476_,
		_w27478_,
		_w27482_,
		_w27488_
	);
	LUT4 #(
		.INIT('h0001)
	) name21662 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27489_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name21663 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27490_
	);
	LUT4 #(
		.INIT('h0020)
	) name21664 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27491_
	);
	LUT4 #(
		.INIT('hc963)
	) name21665 (
		decrypt_pad,
		\u0_R9_reg[16]/NET0131 ,
		\u0_uk_K_r9_reg[27]/P0001 ,
		\u0_uk_K_r9_reg[46]/NET0131 ,
		_w27492_
	);
	LUT3 #(
		.INIT('h80)
	) name21666 (
		_w27477_,
		_w27482_,
		_w27480_,
		_w27493_
	);
	LUT4 #(
		.INIT('h4000)
	) name21667 (
		_w27476_,
		_w27477_,
		_w27482_,
		_w27480_,
		_w27494_
	);
	LUT4 #(
		.INIT('h0002)
	) name21668 (
		_w27490_,
		_w27492_,
		_w27494_,
		_w27491_,
		_w27495_
	);
	LUT4 #(
		.INIT('h0006)
	) name21669 (
		_w27476_,
		_w27477_,
		_w27482_,
		_w27480_,
		_w27496_
	);
	LUT4 #(
		.INIT('h1000)
	) name21670 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27480_,
		_w27497_
	);
	LUT4 #(
		.INIT('h8000)
	) name21671 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27498_
	);
	LUT4 #(
		.INIT('h0002)
	) name21672 (
		_w27492_,
		_w27497_,
		_w27496_,
		_w27498_,
		_w27499_
	);
	LUT4 #(
		.INIT('h0100)
	) name21673 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27500_
	);
	LUT3 #(
		.INIT('h20)
	) name21674 (
		_w27476_,
		_w27478_,
		_w27480_,
		_w27501_
	);
	LUT4 #(
		.INIT('h0800)
	) name21675 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27480_,
		_w27502_
	);
	LUT2 #(
		.INIT('h2)
	) name21676 (
		_w27478_,
		_w27482_,
		_w27503_
	);
	LUT4 #(
		.INIT('h0040)
	) name21677 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27504_
	);
	LUT2 #(
		.INIT('h1)
	) name21678 (
		_w27502_,
		_w27504_,
		_w27505_
	);
	LUT4 #(
		.INIT('h000b)
	) name21679 (
		_w27480_,
		_w27500_,
		_w27502_,
		_w27504_,
		_w27506_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name21680 (
		_w27485_,
		_w27495_,
		_w27499_,
		_w27506_,
		_w27507_
	);
	LUT4 #(
		.INIT('h0200)
	) name21681 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27508_
	);
	LUT4 #(
		.INIT('hfcb8)
	) name21682 (
		_w27489_,
		_w27480_,
		_w27504_,
		_w27508_,
		_w27509_
	);
	LUT2 #(
		.INIT('h2)
	) name21683 (
		_w27477_,
		_w27482_,
		_w27510_
	);
	LUT2 #(
		.INIT('h8)
	) name21684 (
		_w27501_,
		_w27510_,
		_w27511_
	);
	LUT2 #(
		.INIT('h1)
	) name21685 (
		_w27509_,
		_w27511_,
		_w27512_
	);
	LUT3 #(
		.INIT('h65)
	) name21686 (
		\u0_L9_reg[20]/NET0131 ,
		_w27507_,
		_w27512_,
		_w27513_
	);
	LUT4 #(
		.INIT('hc963)
	) name21687 (
		decrypt_pad,
		\u0_R9_reg[28]/NET0131 ,
		\u0_uk_K_r9_reg[1]/NET0131 ,
		\u0_uk_K_r9_reg[52]/NET0131 ,
		_w27514_
	);
	LUT4 #(
		.INIT('hc693)
	) name21688 (
		decrypt_pad,
		\u0_R9_reg[30]/NET0131 ,
		\u0_uk_K_r9_reg[21]/NET0131 ,
		\u0_uk_K_r9_reg[29]/NET0131 ,
		_w27515_
	);
	LUT4 #(
		.INIT('hc963)
	) name21689 (
		decrypt_pad,
		\u0_R9_reg[29]/NET0131 ,
		\u0_uk_K_r9_reg[28]/NET0131 ,
		\u0_uk_K_r9_reg[51]/NET0131 ,
		_w27516_
	);
	LUT4 #(
		.INIT('hc693)
	) name21690 (
		decrypt_pad,
		\u0_R9_reg[1]/NET0131 ,
		\u0_uk_K_r9_reg[36]/NET0131 ,
		\u0_uk_K_r9_reg[44]/NET0131 ,
		_w27517_
	);
	LUT4 #(
		.INIT('hc963)
	) name21691 (
		decrypt_pad,
		\u0_R9_reg[31]/P0001 ,
		\u0_uk_K_r9_reg[45]/NET0131 ,
		\u0_uk_K_r9_reg[9]/NET0131 ,
		_w27518_
	);
	LUT2 #(
		.INIT('h1)
	) name21692 (
		_w27515_,
		_w27518_,
		_w27519_
	);
	LUT4 #(
		.INIT('h7d4c)
	) name21693 (
		_w27516_,
		_w27515_,
		_w27517_,
		_w27518_,
		_w27520_
	);
	LUT2 #(
		.INIT('h2)
	) name21694 (
		_w27514_,
		_w27520_,
		_w27521_
	);
	LUT4 #(
		.INIT('h0020)
	) name21695 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27522_
	);
	LUT4 #(
		.INIT('heedf)
	) name21696 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27523_
	);
	LUT3 #(
		.INIT('h0b)
	) name21697 (
		_w27514_,
		_w27515_,
		_w27517_,
		_w27524_
	);
	LUT3 #(
		.INIT('h0b)
	) name21698 (
		_w27516_,
		_w27517_,
		_w27518_,
		_w27525_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name21699 (
		_w27523_,
		_w27518_,
		_w27524_,
		_w27525_,
		_w27526_
	);
	LUT4 #(
		.INIT('hc693)
	) name21700 (
		decrypt_pad,
		\u0_R9_reg[32]/NET0131 ,
		\u0_uk_K_r9_reg[15]/NET0131 ,
		\u0_uk_K_r9_reg[23]/P0001 ,
		_w27527_
	);
	LUT3 #(
		.INIT('h0b)
	) name21701 (
		_w27521_,
		_w27526_,
		_w27527_,
		_w27528_
	);
	LUT4 #(
		.INIT('h0008)
	) name21702 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27529_
	);
	LUT4 #(
		.INIT('hf531)
	) name21703 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27530_
	);
	LUT3 #(
		.INIT('h02)
	) name21704 (
		_w27518_,
		_w27530_,
		_w27529_,
		_w27531_
	);
	LUT4 #(
		.INIT('h4000)
	) name21705 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27532_
	);
	LUT4 #(
		.INIT('h0001)
	) name21706 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27518_,
		_w27533_
	);
	LUT2 #(
		.INIT('h1)
	) name21707 (
		_w27532_,
		_w27533_,
		_w27534_
	);
	LUT3 #(
		.INIT('h8a)
	) name21708 (
		_w27527_,
		_w27531_,
		_w27534_,
		_w27535_
	);
	LUT4 #(
		.INIT('h0240)
	) name21709 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27536_
	);
	LUT4 #(
		.INIT('h0001)
	) name21710 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27537_
	);
	LUT4 #(
		.INIT('h1000)
	) name21711 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27538_
	);
	LUT4 #(
		.INIT('hedbe)
	) name21712 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27539_
	);
	LUT2 #(
		.INIT('h2)
	) name21713 (
		_w27518_,
		_w27539_,
		_w27540_
	);
	LUT3 #(
		.INIT('h08)
	) name21714 (
		_w27514_,
		_w27516_,
		_w27517_,
		_w27541_
	);
	LUT3 #(
		.INIT('h20)
	) name21715 (
		_w27514_,
		_w27516_,
		_w27527_,
		_w27542_
	);
	LUT4 #(
		.INIT('hcdef)
	) name21716 (
		_w27515_,
		_w27518_,
		_w27541_,
		_w27542_,
		_w27543_
	);
	LUT2 #(
		.INIT('h4)
	) name21717 (
		_w27540_,
		_w27543_,
		_w27544_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name21718 (
		\u0_L9_reg[5]/NET0131 ,
		_w27528_,
		_w27535_,
		_w27544_,
		_w27545_
	);
	LUT3 #(
		.INIT('h02)
	) name21719 (
		_w27480_,
		_w27491_,
		_w27504_,
		_w27546_
	);
	LUT4 #(
		.INIT('hecfc)
	) name21720 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27547_
	);
	LUT2 #(
		.INIT('h1)
	) name21721 (
		_w27492_,
		_w27547_,
		_w27548_
	);
	LUT4 #(
		.INIT('h0002)
	) name21722 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27549_
	);
	LUT4 #(
		.INIT('h0084)
	) name21723 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27550_
	);
	LUT3 #(
		.INIT('h01)
	) name21724 (
		_w27480_,
		_w27550_,
		_w27549_,
		_w27551_
	);
	LUT3 #(
		.INIT('h45)
	) name21725 (
		_w27546_,
		_w27548_,
		_w27551_,
		_w27552_
	);
	LUT4 #(
		.INIT('h0100)
	) name21726 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27480_,
		_w27553_
	);
	LUT4 #(
		.INIT('h0800)
	) name21727 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27554_
	);
	LUT4 #(
		.INIT('h0004)
	) name21728 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27555_
	);
	LUT4 #(
		.INIT('h0002)
	) name21729 (
		_w27492_,
		_w27555_,
		_w27554_,
		_w27553_,
		_w27556_
	);
	LUT4 #(
		.INIT('h5f4f)
	) name21730 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27557_
	);
	LUT3 #(
		.INIT('h0d)
	) name21731 (
		_w27476_,
		_w27482_,
		_w27480_,
		_w27558_
	);
	LUT4 #(
		.INIT('hafbf)
	) name21732 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27480_,
		_w27559_
	);
	LUT4 #(
		.INIT('hcf45)
	) name21733 (
		_w27482_,
		_w27557_,
		_w27558_,
		_w27559_,
		_w27560_
	);
	LUT4 #(
		.INIT('h00fd)
	) name21734 (
		_w27476_,
		_w27477_,
		_w27482_,
		_w27492_,
		_w27561_
	);
	LUT3 #(
		.INIT('hb0)
	) name21735 (
		_w27479_,
		_w27493_,
		_w27561_,
		_w27562_
	);
	LUT4 #(
		.INIT('h153f)
	) name21736 (
		_w27505_,
		_w27556_,
		_w27560_,
		_w27562_,
		_w27563_
	);
	LUT3 #(
		.INIT('h56)
	) name21737 (
		\u0_L9_reg[26]/NET0131 ,
		_w27552_,
		_w27563_,
		_w27564_
	);
	LUT4 #(
		.INIT('hc963)
	) name21738 (
		decrypt_pad,
		\u0_R9_reg[7]/NET0131 ,
		\u0_uk_K_r9_reg[3]/NET0131 ,
		\u0_uk_K_r9_reg[54]/NET0131 ,
		_w27565_
	);
	LUT4 #(
		.INIT('hc693)
	) name21739 (
		decrypt_pad,
		\u0_R9_reg[5]/NET0131 ,
		\u0_uk_K_r9_reg[12]/NET0131 ,
		\u0_uk_K_r9_reg[18]/NET0131 ,
		_w27566_
	);
	LUT4 #(
		.INIT('hc693)
	) name21740 (
		decrypt_pad,
		\u0_R9_reg[9]/NET0131 ,
		\u0_uk_K_r9_reg[25]/NET0131 ,
		\u0_uk_K_r9_reg[6]/NET0131 ,
		_w27567_
	);
	LUT4 #(
		.INIT('hc693)
	) name21741 (
		decrypt_pad,
		\u0_R9_reg[4]/NET0131 ,
		\u0_uk_K_r9_reg[33]/NET0131 ,
		\u0_uk_K_r9_reg[39]/NET0131 ,
		_w27568_
	);
	LUT4 #(
		.INIT('hc693)
	) name21742 (
		decrypt_pad,
		\u0_R9_reg[6]/NET0131 ,
		\u0_uk_K_r9_reg[3]/NET0131 ,
		\u0_uk_K_r9_reg[41]/NET0131 ,
		_w27569_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name21743 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27570_
	);
	LUT3 #(
		.INIT('h10)
	) name21744 (
		_w27566_,
		_w27568_,
		_w27569_,
		_w27571_
	);
	LUT4 #(
		.INIT('h00ef)
	) name21745 (
		_w27566_,
		_w27568_,
		_w27569_,
		_w27565_,
		_w27572_
	);
	LUT4 #(
		.INIT('h5b4b)
	) name21746 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27573_
	);
	LUT4 #(
		.INIT('h7277)
	) name21747 (
		_w27565_,
		_w27570_,
		_w27571_,
		_w27573_,
		_w27574_
	);
	LUT2 #(
		.INIT('h8)
	) name21748 (
		_w27567_,
		_w27568_,
		_w27575_
	);
	LUT4 #(
		.INIT('h4100)
	) name21749 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27576_
	);
	LUT4 #(
		.INIT('h2000)
	) name21750 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27577_
	);
	LUT4 #(
		.INIT('hc693)
	) name21751 (
		decrypt_pad,
		\u0_R9_reg[8]/NET0131 ,
		\u0_uk_K_r9_reg[20]/NET0131 ,
		\u0_uk_K_r9_reg[26]/NET0131 ,
		_w27578_
	);
	LUT3 #(
		.INIT('h01)
	) name21752 (
		_w27577_,
		_w27576_,
		_w27578_,
		_w27579_
	);
	LUT2 #(
		.INIT('h4)
	) name21753 (
		_w27574_,
		_w27579_,
		_w27580_
	);
	LUT3 #(
		.INIT('hd0)
	) name21754 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27581_
	);
	LUT3 #(
		.INIT('h90)
	) name21755 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27582_
	);
	LUT4 #(
		.INIT('h0200)
	) name21756 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27583_
	);
	LUT3 #(
		.INIT('h02)
	) name21757 (
		_w27565_,
		_w27583_,
		_w27582_,
		_w27584_
	);
	LUT4 #(
		.INIT('hd7f4)
	) name21758 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27585_
	);
	LUT2 #(
		.INIT('h8)
	) name21759 (
		_w27572_,
		_w27585_,
		_w27586_
	);
	LUT4 #(
		.INIT('h0400)
	) name21760 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27587_
	);
	LUT3 #(
		.INIT('h0b)
	) name21761 (
		_w27566_,
		_w27567_,
		_w27565_,
		_w27588_
	);
	LUT2 #(
		.INIT('h2)
	) name21762 (
		_w27568_,
		_w27569_,
		_w27589_
	);
	LUT4 #(
		.INIT('h008a)
	) name21763 (
		_w27578_,
		_w27588_,
		_w27589_,
		_w27587_,
		_w27590_
	);
	LUT3 #(
		.INIT('he0)
	) name21764 (
		_w27584_,
		_w27586_,
		_w27590_,
		_w27591_
	);
	LUT3 #(
		.INIT('ha9)
	) name21765 (
		\u0_L9_reg[28]/NET0131 ,
		_w27580_,
		_w27591_,
		_w27592_
	);
	LUT4 #(
		.INIT('h3cf6)
	) name21766 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27593_
	);
	LUT4 #(
		.INIT('h5044)
	) name21767 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27594_
	);
	LUT4 #(
		.INIT('ha7bb)
	) name21768 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27595_
	);
	LUT4 #(
		.INIT('h0020)
	) name21769 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27596_
	);
	LUT4 #(
		.INIT('h00e4)
	) name21770 (
		_w27444_,
		_w27595_,
		_w27593_,
		_w27596_,
		_w27597_
	);
	LUT2 #(
		.INIT('h1)
	) name21771 (
		_w27443_,
		_w27597_,
		_w27598_
	);
	LUT4 #(
		.INIT('hf73b)
	) name21772 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27599_
	);
	LUT2 #(
		.INIT('h2)
	) name21773 (
		_w27444_,
		_w27599_,
		_w27600_
	);
	LUT3 #(
		.INIT('h28)
	) name21774 (
		_w27446_,
		_w27448_,
		_w27447_,
		_w27601_
	);
	LUT4 #(
		.INIT('hc0d0)
	) name21775 (
		_w27446_,
		_w27445_,
		_w27444_,
		_w27448_,
		_w27602_
	);
	LUT3 #(
		.INIT('h01)
	) name21776 (
		_w27594_,
		_w27602_,
		_w27601_,
		_w27603_
	);
	LUT4 #(
		.INIT('h0100)
	) name21777 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27604_
	);
	LUT4 #(
		.INIT('h4000)
	) name21778 (
		_w27446_,
		_w27445_,
		_w27444_,
		_w27448_,
		_w27605_
	);
	LUT2 #(
		.INIT('h1)
	) name21779 (
		_w27604_,
		_w27605_,
		_w27606_
	);
	LUT4 #(
		.INIT('h5700)
	) name21780 (
		_w27443_,
		_w27600_,
		_w27603_,
		_w27606_,
		_w27607_
	);
	LUT3 #(
		.INIT('h9a)
	) name21781 (
		\u0_L9_reg[29]/NET0131 ,
		_w27598_,
		_w27607_,
		_w27608_
	);
	LUT4 #(
		.INIT('h0a02)
	) name21782 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27609_
	);
	LUT3 #(
		.INIT('h01)
	) name21783 (
		_w27480_,
		_w27504_,
		_w27609_,
		_w27610_
	);
	LUT3 #(
		.INIT('h04)
	) name21784 (
		_w27486_,
		_w27480_,
		_w27491_,
		_w27611_
	);
	LUT4 #(
		.INIT('h6fff)
	) name21785 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27612_
	);
	LUT4 #(
		.INIT('h02aa)
	) name21786 (
		_w27492_,
		_w27610_,
		_w27611_,
		_w27612_,
		_w27613_
	);
	LUT4 #(
		.INIT('h0001)
	) name21787 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27480_,
		_w27614_
	);
	LUT3 #(
		.INIT('h08)
	) name21788 (
		_w27476_,
		_w27477_,
		_w27482_,
		_w27615_
	);
	LUT4 #(
		.INIT('h0008)
	) name21789 (
		_w27476_,
		_w27478_,
		_w27482_,
		_w27480_,
		_w27616_
	);
	LUT3 #(
		.INIT('h01)
	) name21790 (
		_w27614_,
		_w27615_,
		_w27616_,
		_w27617_
	);
	LUT4 #(
		.INIT('h0400)
	) name21791 (
		_w27476_,
		_w27478_,
		_w27482_,
		_w27480_,
		_w27618_
	);
	LUT3 #(
		.INIT('h20)
	) name21792 (
		_w27476_,
		_w27477_,
		_w27480_,
		_w27619_
	);
	LUT3 #(
		.INIT('h23)
	) name21793 (
		_w27503_,
		_w27618_,
		_w27619_,
		_w27620_
	);
	LUT4 #(
		.INIT('h1333)
	) name21794 (
		_w27490_,
		_w27492_,
		_w27617_,
		_w27620_,
		_w27621_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name21795 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27622_
	);
	LUT2 #(
		.INIT('h1)
	) name21796 (
		_w27480_,
		_w27622_,
		_w27623_
	);
	LUT3 #(
		.INIT('h15)
	) name21797 (
		_w27494_,
		_w27501_,
		_w27510_,
		_w27624_
	);
	LUT2 #(
		.INIT('h4)
	) name21798 (
		_w27623_,
		_w27624_,
		_w27625_
	);
	LUT4 #(
		.INIT('h5655)
	) name21799 (
		\u0_L9_reg[10]/NET0131 ,
		_w27621_,
		_w27613_,
		_w27625_,
		_w27626_
	);
	LUT4 #(
		.INIT('hc693)
	) name21800 (
		decrypt_pad,
		\u0_R9_reg[20]/NET0131 ,
		\u0_uk_K_r9_reg[0]/P0001 ,
		\u0_uk_K_r9_reg[8]/NET0131 ,
		_w27627_
	);
	LUT4 #(
		.INIT('hc693)
	) name21801 (
		decrypt_pad,
		\u0_R9_reg[19]/NET0131 ,
		\u0_uk_K_r9_reg[16]/NET0131 ,
		\u0_uk_K_r9_reg[52]/NET0131 ,
		_w27628_
	);
	LUT4 #(
		.INIT('hc693)
	) name21802 (
		decrypt_pad,
		\u0_R9_reg[17]/NET0131 ,
		\u0_uk_K_r9_reg[35]/NET0131 ,
		\u0_uk_K_r9_reg[43]/NET0131 ,
		_w27629_
	);
	LUT4 #(
		.INIT('hc963)
	) name21803 (
		decrypt_pad,
		\u0_R9_reg[16]/NET0131 ,
		\u0_uk_K_r9_reg[21]/NET0131 ,
		\u0_uk_K_r9_reg[44]/NET0131 ,
		_w27630_
	);
	LUT4 #(
		.INIT('hc693)
	) name21804 (
		decrypt_pad,
		\u0_R9_reg[21]/NET0131 ,
		\u0_uk_K_r9_reg[1]/NET0131 ,
		\u0_uk_K_r9_reg[9]/NET0131 ,
		_w27631_
	);
	LUT2 #(
		.INIT('h2)
	) name21805 (
		_w27630_,
		_w27631_,
		_w27632_
	);
	LUT4 #(
		.INIT('hc693)
	) name21806 (
		decrypt_pad,
		\u0_R9_reg[18]/NET0131 ,
		\u0_uk_K_r9_reg[29]/NET0131 ,
		\u0_uk_K_r9_reg[37]/NET0131 ,
		_w27633_
	);
	LUT4 #(
		.INIT('h938f)
	) name21807 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27634_
	);
	LUT2 #(
		.INIT('h2)
	) name21808 (
		_w27628_,
		_w27634_,
		_w27635_
	);
	LUT3 #(
		.INIT('hbe)
	) name21809 (
		_w27630_,
		_w27631_,
		_w27629_,
		_w27636_
	);
	LUT2 #(
		.INIT('h1)
	) name21810 (
		_w27633_,
		_w27628_,
		_w27637_
	);
	LUT2 #(
		.INIT('h4)
	) name21811 (
		_w27636_,
		_w27637_,
		_w27638_
	);
	LUT3 #(
		.INIT('h80)
	) name21812 (
		_w27630_,
		_w27631_,
		_w27629_,
		_w27639_
	);
	LUT2 #(
		.INIT('h2)
	) name21813 (
		_w27633_,
		_w27628_,
		_w27640_
	);
	LUT4 #(
		.INIT('h0400)
	) name21814 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27641_
	);
	LUT4 #(
		.INIT('h0008)
	) name21815 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27642_
	);
	LUT4 #(
		.INIT('hfbb7)
	) name21816 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27643_
	);
	LUT3 #(
		.INIT('h70)
	) name21817 (
		_w27639_,
		_w27640_,
		_w27643_,
		_w27644_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name21818 (
		_w27627_,
		_w27635_,
		_w27638_,
		_w27644_,
		_w27645_
	);
	LUT4 #(
		.INIT('h7f00)
	) name21819 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27628_,
		_w27646_
	);
	LUT4 #(
		.INIT('heefc)
	) name21820 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27647_
	);
	LUT2 #(
		.INIT('h8)
	) name21821 (
		_w27646_,
		_w27647_,
		_w27648_
	);
	LUT3 #(
		.INIT('h04)
	) name21822 (
		_w27630_,
		_w27631_,
		_w27629_,
		_w27649_
	);
	LUT4 #(
		.INIT('h00df)
	) name21823 (
		_w27633_,
		_w27631_,
		_w27629_,
		_w27628_,
		_w27650_
	);
	LUT4 #(
		.INIT('h0004)
	) name21824 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27651_
	);
	LUT4 #(
		.INIT('h4000)
	) name21825 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27652_
	);
	LUT4 #(
		.INIT('hbffb)
	) name21826 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27653_
	);
	LUT3 #(
		.INIT('h40)
	) name21827 (
		_w27649_,
		_w27650_,
		_w27653_,
		_w27654_
	);
	LUT4 #(
		.INIT('h0080)
	) name21828 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27655_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name21829 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27656_
	);
	LUT4 #(
		.INIT('h001f)
	) name21830 (
		_w27648_,
		_w27654_,
		_w27656_,
		_w27627_,
		_w27657_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name21831 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27658_
	);
	LUT4 #(
		.INIT('h0020)
	) name21832 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27659_
	);
	LUT4 #(
		.INIT('hfddf)
	) name21833 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27660_
	);
	LUT3 #(
		.INIT('hd8)
	) name21834 (
		_w27628_,
		_w27658_,
		_w27660_,
		_w27661_
	);
	LUT4 #(
		.INIT('h5655)
	) name21835 (
		\u0_L9_reg[14]/NET0131 ,
		_w27657_,
		_w27645_,
		_w27661_,
		_w27662_
	);
	LUT4 #(
		.INIT('h7773)
	) name21836 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27663_
	);
	LUT4 #(
		.INIT('h6673)
	) name21837 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27664_
	);
	LUT4 #(
		.INIT('h0002)
	) name21838 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27665_
	);
	LUT4 #(
		.INIT('h3302)
	) name21839 (
		_w27518_,
		_w27527_,
		_w27664_,
		_w27665_,
		_w27666_
	);
	LUT4 #(
		.INIT('h0040)
	) name21840 (
		_w27516_,
		_w27515_,
		_w27517_,
		_w27518_,
		_w27667_
	);
	LUT4 #(
		.INIT('hf7b7)
	) name21841 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27668_
	);
	LUT4 #(
		.INIT('h0100)
	) name21842 (
		_w27514_,
		_w27516_,
		_w27517_,
		_w27518_,
		_w27669_
	);
	LUT4 #(
		.INIT('h2000)
	) name21843 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27670_
	);
	LUT4 #(
		.INIT('h0100)
	) name21844 (
		_w27669_,
		_w27667_,
		_w27670_,
		_w27668_,
		_w27671_
	);
	LUT3 #(
		.INIT('h02)
	) name21845 (
		_w27514_,
		_w27516_,
		_w27527_,
		_w27672_
	);
	LUT4 #(
		.INIT('hfbbf)
	) name21846 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27673_
	);
	LUT4 #(
		.INIT('h00df)
	) name21847 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27518_,
		_w27674_
	);
	LUT4 #(
		.INIT('h1000)
	) name21848 (
		_w27537_,
		_w27672_,
		_w27674_,
		_w27673_,
		_w27675_
	);
	LUT4 #(
		.INIT('h0100)
	) name21849 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27676_
	);
	LUT3 #(
		.INIT('h02)
	) name21850 (
		_w27518_,
		_w27532_,
		_w27676_,
		_w27677_
	);
	LUT4 #(
		.INIT('hddd0)
	) name21851 (
		_w27527_,
		_w27671_,
		_w27675_,
		_w27677_,
		_w27678_
	);
	LUT3 #(
		.INIT('h65)
	) name21852 (
		\u0_L9_reg[15]/P0001 ,
		_w27666_,
		_w27678_,
		_w27679_
	);
	LUT4 #(
		.INIT('h0004)
	) name21853 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27680_
	);
	LUT4 #(
		.INIT('h00bf)
	) name21854 (
		_w27388_,
		_w27389_,
		_w27390_,
		_w27400_,
		_w27681_
	);
	LUT3 #(
		.INIT('h41)
	) name21855 (
		_w27388_,
		_w27391_,
		_w27392_,
		_w27682_
	);
	LUT4 #(
		.INIT('h0100)
	) name21856 (
		_w27393_,
		_w27680_,
		_w27682_,
		_w27681_,
		_w27683_
	);
	LUT3 #(
		.INIT('h08)
	) name21857 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27684_
	);
	LUT4 #(
		.INIT('h2800)
	) name21858 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27685_
	);
	LUT3 #(
		.INIT('h04)
	) name21859 (
		_w27389_,
		_w27390_,
		_w27392_,
		_w27686_
	);
	LUT4 #(
		.INIT('hf5cf)
	) name21860 (
		_w27388_,
		_w27389_,
		_w27390_,
		_w27392_,
		_w27687_
	);
	LUT3 #(
		.INIT('h32)
	) name21861 (
		_w27391_,
		_w27685_,
		_w27687_,
		_w27688_
	);
	LUT2 #(
		.INIT('h8)
	) name21862 (
		_w27683_,
		_w27688_,
		_w27689_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name21863 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27690_
	);
	LUT2 #(
		.INIT('h2)
	) name21864 (
		_w27388_,
		_w27690_,
		_w27691_
	);
	LUT4 #(
		.INIT('h1400)
	) name21865 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27692_
	);
	LUT4 #(
		.INIT('h0028)
	) name21866 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27693_
	);
	LUT4 #(
		.INIT('h008c)
	) name21867 (
		_w27388_,
		_w27400_,
		_w27406_,
		_w27693_,
		_w27694_
	);
	LUT3 #(
		.INIT('h10)
	) name21868 (
		_w27692_,
		_w27691_,
		_w27694_,
		_w27695_
	);
	LUT3 #(
		.INIT('ha9)
	) name21869 (
		\u0_L9_reg[12]/NET0131 ,
		_w27689_,
		_w27695_,
		_w27696_
	);
	LUT4 #(
		.INIT('hc6cd)
	) name21870 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27697_
	);
	LUT2 #(
		.INIT('h2)
	) name21871 (
		_w27492_,
		_w27697_,
		_w27698_
	);
	LUT3 #(
		.INIT('h40)
	) name21872 (
		_w27487_,
		_w27480_,
		_w27612_,
		_w27699_
	);
	LUT4 #(
		.INIT('hae3b)
	) name21873 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27700_
	);
	LUT2 #(
		.INIT('h2)
	) name21874 (
		_w27492_,
		_w27700_,
		_w27701_
	);
	LUT3 #(
		.INIT('h01)
	) name21875 (
		_w27480_,
		_w27500_,
		_w27554_,
		_w27702_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name21876 (
		_w27698_,
		_w27699_,
		_w27701_,
		_w27702_,
		_w27703_
	);
	LUT4 #(
		.INIT('h202a)
	) name21877 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27704_
	);
	LUT4 #(
		.INIT('hfbc8)
	) name21878 (
		_w27488_,
		_w27480_,
		_w27508_,
		_w27704_,
		_w27705_
	);
	LUT4 #(
		.INIT('h7fb7)
	) name21879 (
		_w27476_,
		_w27477_,
		_w27478_,
		_w27482_,
		_w27706_
	);
	LUT3 #(
		.INIT('h45)
	) name21880 (
		_w27492_,
		_w27705_,
		_w27706_,
		_w27707_
	);
	LUT3 #(
		.INIT('h56)
	) name21881 (
		\u0_L9_reg[1]/NET0131 ,
		_w27703_,
		_w27707_,
		_w27708_
	);
	LUT4 #(
		.INIT('h080a)
	) name21882 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27709_
	);
	LUT3 #(
		.INIT('h01)
	) name21883 (
		_w27518_,
		_w27670_,
		_w27709_,
		_w27710_
	);
	LUT4 #(
		.INIT('h8381)
	) name21884 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27711_
	);
	LUT4 #(
		.INIT('hbf00)
	) name21885 (
		_w27514_,
		_w27516_,
		_w27517_,
		_w27518_,
		_w27712_
	);
	LUT2 #(
		.INIT('h4)
	) name21886 (
		_w27711_,
		_w27712_,
		_w27713_
	);
	LUT4 #(
		.INIT('h0090)
	) name21887 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27714_
	);
	LUT3 #(
		.INIT('h02)
	) name21888 (
		_w27527_,
		_w27676_,
		_w27714_,
		_w27715_
	);
	LUT3 #(
		.INIT('he0)
	) name21889 (
		_w27710_,
		_w27713_,
		_w27715_,
		_w27716_
	);
	LUT4 #(
		.INIT('hde56)
	) name21890 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27717_
	);
	LUT2 #(
		.INIT('h2)
	) name21891 (
		_w27518_,
		_w27717_,
		_w27718_
	);
	LUT4 #(
		.INIT('h00bf)
	) name21892 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27527_,
		_w27719_
	);
	LUT2 #(
		.INIT('h4)
	) name21893 (
		_w27522_,
		_w27719_,
		_w27720_
	);
	LUT2 #(
		.INIT('h8)
	) name21894 (
		_w27514_,
		_w27517_,
		_w27721_
	);
	LUT3 #(
		.INIT('hdc)
	) name21895 (
		_w27516_,
		_w27515_,
		_w27518_,
		_w27722_
	);
	LUT2 #(
		.INIT('h2)
	) name21896 (
		_w27721_,
		_w27722_,
		_w27723_
	);
	LUT2 #(
		.INIT('h1)
	) name21897 (
		_w27514_,
		_w27518_,
		_w27724_
	);
	LUT3 #(
		.INIT('h35)
	) name21898 (
		_w27516_,
		_w27515_,
		_w27517_,
		_w27725_
	);
	LUT3 #(
		.INIT('h51)
	) name21899 (
		_w27537_,
		_w27724_,
		_w27725_,
		_w27726_
	);
	LUT4 #(
		.INIT('h1000)
	) name21900 (
		_w27718_,
		_w27723_,
		_w27720_,
		_w27726_,
		_w27727_
	);
	LUT3 #(
		.INIT('ha9)
	) name21901 (
		\u0_L9_reg[21]/NET0131 ,
		_w27716_,
		_w27727_,
		_w27728_
	);
	LUT4 #(
		.INIT('h3dc8)
	) name21902 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27729_
	);
	LUT4 #(
		.INIT('hee3f)
	) name21903 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27730_
	);
	LUT4 #(
		.INIT('ha7ff)
	) name21904 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27731_
	);
	LUT4 #(
		.INIT('hd800)
	) name21905 (
		_w27628_,
		_w27729_,
		_w27730_,
		_w27731_,
		_w27732_
	);
	LUT2 #(
		.INIT('h2)
	) name21906 (
		_w27627_,
		_w27732_,
		_w27733_
	);
	LUT4 #(
		.INIT('hddf3)
	) name21907 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27734_
	);
	LUT2 #(
		.INIT('h1)
	) name21908 (
		_w27628_,
		_w27734_,
		_w27735_
	);
	LUT4 #(
		.INIT('h1000)
	) name21909 (
		_w27633_,
		_w27631_,
		_w27629_,
		_w27628_,
		_w27736_
	);
	LUT4 #(
		.INIT('h0001)
	) name21910 (
		_w27633_,
		_w27630_,
		_w27629_,
		_w27628_,
		_w27737_
	);
	LUT4 #(
		.INIT('h2000)
	) name21911 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27738_
	);
	LUT3 #(
		.INIT('h01)
	) name21912 (
		_w27737_,
		_w27738_,
		_w27736_,
		_w27739_
	);
	LUT4 #(
		.INIT('hf7ed)
	) name21913 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27740_
	);
	LUT4 #(
		.INIT('h0008)
	) name21914 (
		_w27633_,
		_w27630_,
		_w27629_,
		_w27628_,
		_w27741_
	);
	LUT4 #(
		.INIT('h0031)
	) name21915 (
		_w27628_,
		_w27652_,
		_w27740_,
		_w27741_,
		_w27742_
	);
	LUT4 #(
		.INIT('hba00)
	) name21916 (
		_w27627_,
		_w27735_,
		_w27739_,
		_w27742_,
		_w27743_
	);
	LUT3 #(
		.INIT('h65)
	) name21917 (
		\u0_L9_reg[25]/NET0131 ,
		_w27733_,
		_w27743_,
		_w27744_
	);
	LUT4 #(
		.INIT('hf3ec)
	) name21918 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27745_
	);
	LUT3 #(
		.INIT('h7d)
	) name21919 (
		_w27420_,
		_w27417_,
		_w27418_,
		_w27746_
	);
	LUT4 #(
		.INIT('hfd7f)
	) name21920 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27747_
	);
	LUT4 #(
		.INIT('he400)
	) name21921 (
		_w27416_,
		_w27745_,
		_w27746_,
		_w27747_,
		_w27748_
	);
	LUT4 #(
		.INIT('h4555)
	) name21922 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27749_
	);
	LUT4 #(
		.INIT('haa8a)
	) name21923 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27750_
	);
	LUT3 #(
		.INIT('h02)
	) name21924 (
		_w27416_,
		_w27750_,
		_w27749_,
		_w27751_
	);
	LUT4 #(
		.INIT('h0400)
	) name21925 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27752_
	);
	LUT4 #(
		.INIT('hc9cd)
	) name21926 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27753_
	);
	LUT4 #(
		.INIT('h4041)
	) name21927 (
		_w27416_,
		_w27419_,
		_w27420_,
		_w27417_,
		_w27754_
	);
	LUT4 #(
		.INIT('h0040)
	) name21928 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27755_
	);
	LUT4 #(
		.INIT('h5fbf)
	) name21929 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27756_
	);
	LUT4 #(
		.INIT('h0d00)
	) name21930 (
		_w27416_,
		_w27753_,
		_w27754_,
		_w27756_,
		_w27757_
	);
	LUT4 #(
		.INIT('h0e04)
	) name21931 (
		_w27415_,
		_w27748_,
		_w27751_,
		_w27757_,
		_w27758_
	);
	LUT2 #(
		.INIT('h9)
	) name21932 (
		\u0_L9_reg[17]/NET0131 ,
		_w27758_,
		_w27759_
	);
	LUT4 #(
		.INIT('h0026)
	) name21933 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27760_
	);
	LUT3 #(
		.INIT('h40)
	) name21934 (
		_w27566_,
		_w27569_,
		_w27565_,
		_w27761_
	);
	LUT3 #(
		.INIT('h13)
	) name21935 (
		_w27575_,
		_w27760_,
		_w27761_,
		_w27762_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name21936 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27763_
	);
	LUT4 #(
		.INIT('h00bf)
	) name21937 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27565_,
		_w27764_
	);
	LUT2 #(
		.INIT('h2)
	) name21938 (
		_w27567_,
		_w27569_,
		_w27765_
	);
	LUT4 #(
		.INIT('h0004)
	) name21939 (
		_w27566_,
		_w27567_,
		_w27569_,
		_w27565_,
		_w27766_
	);
	LUT4 #(
		.INIT('h0800)
	) name21940 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27767_
	);
	LUT4 #(
		.INIT('h000b)
	) name21941 (
		_w27763_,
		_w27764_,
		_w27766_,
		_w27767_,
		_w27768_
	);
	LUT3 #(
		.INIT('h15)
	) name21942 (
		_w27578_,
		_w27762_,
		_w27768_,
		_w27769_
	);
	LUT4 #(
		.INIT('hbc6e)
	) name21943 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27770_
	);
	LUT4 #(
		.INIT('h0804)
	) name21944 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27771_
	);
	LUT4 #(
		.INIT('h0051)
	) name21945 (
		_w27565_,
		_w27578_,
		_w27770_,
		_w27771_,
		_w27772_
	);
	LUT4 #(
		.INIT('h5f45)
	) name21946 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27773_
	);
	LUT3 #(
		.INIT('h10)
	) name21947 (
		_w27566_,
		_w27567_,
		_w27569_,
		_w27774_
	);
	LUT4 #(
		.INIT('h0100)
	) name21948 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27775_
	);
	LUT4 #(
		.INIT('hf700)
	) name21949 (
		_w27566_,
		_w27568_,
		_w27569_,
		_w27565_,
		_w27776_
	);
	LUT4 #(
		.INIT('h0d00)
	) name21950 (
		_w27578_,
		_w27773_,
		_w27775_,
		_w27776_,
		_w27777_
	);
	LUT2 #(
		.INIT('h1)
	) name21951 (
		_w27772_,
		_w27777_,
		_w27778_
	);
	LUT3 #(
		.INIT('h56)
	) name21952 (
		\u0_L9_reg[2]/NET0131 ,
		_w27769_,
		_w27778_,
		_w27779_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name21953 (
		_w27445_,
		_w27444_,
		_w27448_,
		_w27447_,
		_w27780_
	);
	LUT4 #(
		.INIT('hdfaf)
	) name21954 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27781_
	);
	LUT4 #(
		.INIT('h3331)
	) name21955 (
		_w27445_,
		_w27444_,
		_w27448_,
		_w27447_,
		_w27782_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name21956 (
		_w27596_,
		_w27780_,
		_w27781_,
		_w27782_,
		_w27783_
	);
	LUT3 #(
		.INIT('h01)
	) name21957 (
		_w27443_,
		_w27456_,
		_w27604_,
		_w27784_
	);
	LUT3 #(
		.INIT('h15)
	) name21958 (
		_w27446_,
		_w27448_,
		_w27447_,
		_w27785_
	);
	LUT4 #(
		.INIT('hd850)
	) name21959 (
		_w27446_,
		_w27445_,
		_w27444_,
		_w27448_,
		_w27786_
	);
	LUT2 #(
		.INIT('h4)
	) name21960 (
		_w27785_,
		_w27786_,
		_w27787_
	);
	LUT4 #(
		.INIT('h2202)
	) name21961 (
		_w27443_,
		_w27470_,
		_w27455_,
		_w27449_,
		_w27788_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name21962 (
		_w27783_,
		_w27784_,
		_w27787_,
		_w27788_,
		_w27789_
	);
	LUT4 #(
		.INIT('h1233)
	) name21963 (
		_w27445_,
		_w27444_,
		_w27448_,
		_w27447_,
		_w27790_
	);
	LUT4 #(
		.INIT('hc448)
	) name21964 (
		_w27445_,
		_w27444_,
		_w27448_,
		_w27447_,
		_w27791_
	);
	LUT4 #(
		.INIT('h3331)
	) name21965 (
		_w27446_,
		_w27472_,
		_w27791_,
		_w27790_,
		_w27792_
	);
	LUT3 #(
		.INIT('h65)
	) name21966 (
		\u0_L9_reg[4]/NET0131 ,
		_w27789_,
		_w27792_,
		_w27793_
	);
	LUT4 #(
		.INIT('hfcc7)
	) name21967 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27794_
	);
	LUT2 #(
		.INIT('h1)
	) name21968 (
		_w27416_,
		_w27794_,
		_w27795_
	);
	LUT3 #(
		.INIT('ha8)
	) name21969 (
		_w27416_,
		_w27419_,
		_w27418_,
		_w27796_
	);
	LUT2 #(
		.INIT('h8)
	) name21970 (
		_w27432_,
		_w27796_,
		_w27797_
	);
	LUT3 #(
		.INIT('h07)
	) name21971 (
		_w27431_,
		_w27439_,
		_w27752_,
		_w27798_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name21972 (
		_w27415_,
		_w27795_,
		_w27797_,
		_w27798_,
		_w27799_
	);
	LUT4 #(
		.INIT('h373f)
	) name21973 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27800_
	);
	LUT2 #(
		.INIT('h1)
	) name21974 (
		_w27416_,
		_w27800_,
		_w27801_
	);
	LUT4 #(
		.INIT('h0020)
	) name21975 (
		_w27416_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27802_
	);
	LUT4 #(
		.INIT('h0800)
	) name21976 (
		_w27416_,
		_w27419_,
		_w27420_,
		_w27418_,
		_w27803_
	);
	LUT3 #(
		.INIT('h7e)
	) name21977 (
		_w27419_,
		_w27417_,
		_w27418_,
		_w27804_
	);
	LUT3 #(
		.INIT('h10)
	) name21978 (
		_w27802_,
		_w27803_,
		_w27804_,
		_w27805_
	);
	LUT3 #(
		.INIT('hd9)
	) name21979 (
		_w27420_,
		_w27417_,
		_w27418_,
		_w27806_
	);
	LUT4 #(
		.INIT('h7ebf)
	) name21980 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w27807_
	);
	LUT4 #(
		.INIT('hfda8)
	) name21981 (
		_w27416_,
		_w27419_,
		_w27806_,
		_w27807_,
		_w27808_
	);
	LUT4 #(
		.INIT('hba00)
	) name21982 (
		_w27415_,
		_w27801_,
		_w27805_,
		_w27808_,
		_w27809_
	);
	LUT3 #(
		.INIT('h9a)
	) name21983 (
		\u0_L9_reg[23]/NET0131 ,
		_w27799_,
		_w27809_,
		_w27810_
	);
	LUT4 #(
		.INIT('hba76)
	) name21984 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27811_
	);
	LUT2 #(
		.INIT('h1)
	) name21985 (
		_w27518_,
		_w27811_,
		_w27812_
	);
	LUT3 #(
		.INIT('hd0)
	) name21986 (
		_w27514_,
		_w27517_,
		_w27518_,
		_w27813_
	);
	LUT4 #(
		.INIT('hbcdf)
	) name21987 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27814_
	);
	LUT3 #(
		.INIT('hb0)
	) name21988 (
		_w27663_,
		_w27813_,
		_w27814_,
		_w27815_
	);
	LUT3 #(
		.INIT('h8a)
	) name21989 (
		_w27527_,
		_w27812_,
		_w27815_,
		_w27816_
	);
	LUT4 #(
		.INIT('hfd00)
	) name21990 (
		_w27516_,
		_w27515_,
		_w27517_,
		_w27518_,
		_w27817_
	);
	LUT4 #(
		.INIT('h0cbf)
	) name21991 (
		_w27514_,
		_w27516_,
		_w27515_,
		_w27517_,
		_w27818_
	);
	LUT2 #(
		.INIT('h8)
	) name21992 (
		_w27817_,
		_w27818_,
		_w27819_
	);
	LUT4 #(
		.INIT('h0080)
	) name21993 (
		_w27514_,
		_w27515_,
		_w27517_,
		_w27518_,
		_w27820_
	);
	LUT4 #(
		.INIT('h0004)
	) name21994 (
		_w27514_,
		_w27516_,
		_w27517_,
		_w27518_,
		_w27821_
	);
	LUT3 #(
		.INIT('h01)
	) name21995 (
		_w27538_,
		_w27821_,
		_w27820_,
		_w27822_
	);
	LUT3 #(
		.INIT('h45)
	) name21996 (
		_w27527_,
		_w27819_,
		_w27822_,
		_w27823_
	);
	LUT2 #(
		.INIT('h4)
	) name21997 (
		_w27518_,
		_w27536_,
		_w27824_
	);
	LUT4 #(
		.INIT('h0400)
	) name21998 (
		_w27516_,
		_w27515_,
		_w27517_,
		_w27518_,
		_w27825_
	);
	LUT3 #(
		.INIT('h07)
	) name21999 (
		_w27519_,
		_w27541_,
		_w27825_,
		_w27826_
	);
	LUT2 #(
		.INIT('h4)
	) name22000 (
		_w27824_,
		_w27826_,
		_w27827_
	);
	LUT4 #(
		.INIT('h5655)
	) name22001 (
		\u0_L9_reg[27]/NET0131 ,
		_w27816_,
		_w27823_,
		_w27827_,
		_w27828_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name22002 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27829_
	);
	LUT4 #(
		.INIT('hf9ed)
	) name22003 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27830_
	);
	LUT4 #(
		.INIT('h0515)
	) name22004 (
		_w27565_,
		_w27578_,
		_w27829_,
		_w27830_,
		_w27831_
	);
	LUT4 #(
		.INIT('h2e9e)
	) name22005 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27832_
	);
	LUT2 #(
		.INIT('h2)
	) name22006 (
		_w27565_,
		_w27832_,
		_w27833_
	);
	LUT3 #(
		.INIT('h32)
	) name22007 (
		_w27566_,
		_w27568_,
		_w27565_,
		_w27834_
	);
	LUT3 #(
		.INIT('h15)
	) name22008 (
		_w27578_,
		_w27765_,
		_w27834_,
		_w27835_
	);
	LUT2 #(
		.INIT('h4)
	) name22009 (
		_w27833_,
		_w27835_,
		_w27836_
	);
	LUT3 #(
		.INIT('h20)
	) name22010 (
		_w27567_,
		_w27568_,
		_w27569_,
		_w27837_
	);
	LUT4 #(
		.INIT('hfe00)
	) name22011 (
		_w27566_,
		_w27567_,
		_w27569_,
		_w27565_,
		_w27838_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name22012 (
		_w27764_,
		_w27774_,
		_w27837_,
		_w27838_,
		_w27839_
	);
	LUT4 #(
		.INIT('h0002)
	) name22013 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27840_
	);
	LUT4 #(
		.INIT('h0002)
	) name22014 (
		_w27578_,
		_w27766_,
		_w27767_,
		_w27840_,
		_w27841_
	);
	LUT3 #(
		.INIT('h20)
	) name22015 (
		_w27829_,
		_w27839_,
		_w27841_,
		_w27842_
	);
	LUT4 #(
		.INIT('h999a)
	) name22016 (
		\u0_L9_reg[13]/NET0131 ,
		_w27831_,
		_w27836_,
		_w27842_,
		_w27843_
	);
	LUT4 #(
		.INIT('h0ee2)
	) name22017 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27844_
	);
	LUT4 #(
		.INIT('hd001)
	) name22018 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27845_
	);
	LUT3 #(
		.INIT('h01)
	) name22019 (
		_w27388_,
		_w27845_,
		_w27844_,
		_w27846_
	);
	LUT4 #(
		.INIT('h0080)
	) name22020 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27847_
	);
	LUT4 #(
		.INIT('hbb5c)
	) name22021 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27848_
	);
	LUT3 #(
		.INIT('h31)
	) name22022 (
		_w27388_,
		_w27847_,
		_w27848_,
		_w27849_
	);
	LUT3 #(
		.INIT('h8a)
	) name22023 (
		_w27400_,
		_w27846_,
		_w27849_,
		_w27850_
	);
	LUT4 #(
		.INIT('hcfaf)
	) name22024 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27851_
	);
	LUT3 #(
		.INIT('h31)
	) name22025 (
		_w27388_,
		_w27409_,
		_w27851_,
		_w27852_
	);
	LUT4 #(
		.INIT('h8040)
	) name22026 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27853_
	);
	LUT3 #(
		.INIT('h0b)
	) name22027 (
		_w27686_,
		_w27682_,
		_w27853_,
		_w27854_
	);
	LUT4 #(
		.INIT('h4404)
	) name22028 (
		_w27388_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27855_
	);
	LUT4 #(
		.INIT('h135f)
	) name22029 (
		_w27388_,
		_w27394_,
		_w27406_,
		_w27855_,
		_w27856_
	);
	LUT4 #(
		.INIT('hea00)
	) name22030 (
		_w27400_,
		_w27852_,
		_w27854_,
		_w27856_,
		_w27857_
	);
	LUT3 #(
		.INIT('h65)
	) name22031 (
		\u0_L9_reg[32]/NET0131 ,
		_w27850_,
		_w27857_,
		_w27858_
	);
	LUT4 #(
		.INIT('hc693)
	) name22032 (
		decrypt_pad,
		\u0_R9_reg[11]/P0001 ,
		\u0_uk_K_r9_reg[40]/NET0131 ,
		\u0_uk_K_r9_reg[46]/NET0131 ,
		_w27859_
	);
	LUT4 #(
		.INIT('hc963)
	) name22033 (
		decrypt_pad,
		\u0_R9_reg[12]/NET0131 ,
		\u0_uk_K_r9_reg[4]/NET0131 ,
		\u0_uk_K_r9_reg[55]/NET0131 ,
		_w27860_
	);
	LUT4 #(
		.INIT('hc693)
	) name22034 (
		decrypt_pad,
		\u0_R9_reg[13]/NET0131 ,
		\u0_uk_K_r9_reg[11]/NET0131 ,
		\u0_uk_K_r9_reg[17]/NET0131 ,
		_w27861_
	);
	LUT4 #(
		.INIT('hc963)
	) name22035 (
		decrypt_pad,
		\u0_R9_reg[9]/NET0131 ,
		\u0_uk_K_r9_reg[12]/NET0131 ,
		\u0_uk_K_r9_reg[6]/NET0131 ,
		_w27862_
	);
	LUT4 #(
		.INIT('hc963)
	) name22036 (
		decrypt_pad,
		\u0_R9_reg[10]/NET0131 ,
		\u0_uk_K_r9_reg[20]/NET0131 ,
		\u0_uk_K_r9_reg[39]/NET0131 ,
		_w27863_
	);
	LUT4 #(
		.INIT('hc693)
	) name22037 (
		decrypt_pad,
		\u0_R9_reg[8]/NET0131 ,
		\u0_uk_K_r9_reg[34]/NET0131 ,
		\u0_uk_K_r9_reg[40]/NET0131 ,
		_w27864_
	);
	LUT4 #(
		.INIT('h95b5)
	) name22038 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27865_
	);
	LUT2 #(
		.INIT('h1)
	) name22039 (
		_w27861_,
		_w27864_,
		_w27866_
	);
	LUT2 #(
		.INIT('h1)
	) name22040 (
		_w27862_,
		_w27863_,
		_w27867_
	);
	LUT4 #(
		.INIT('h0001)
	) name22041 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27868_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name22042 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27869_
	);
	LUT4 #(
		.INIT('h08cc)
	) name22043 (
		_w27860_,
		_w27859_,
		_w27865_,
		_w27869_,
		_w27870_
	);
	LUT2 #(
		.INIT('h8)
	) name22044 (
		_w27861_,
		_w27864_,
		_w27871_
	);
	LUT2 #(
		.INIT('h6)
	) name22045 (
		_w27861_,
		_w27864_,
		_w27872_
	);
	LUT4 #(
		.INIT('h0990)
	) name22046 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27873_
	);
	LUT4 #(
		.INIT('h2000)
	) name22047 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27874_
	);
	LUT2 #(
		.INIT('h4)
	) name22048 (
		_w27864_,
		_w27859_,
		_w27875_
	);
	LUT4 #(
		.INIT('h0400)
	) name22049 (
		_w27864_,
		_w27862_,
		_w27863_,
		_w27859_,
		_w27876_
	);
	LUT3 #(
		.INIT('h0b)
	) name22050 (
		_w27859_,
		_w27874_,
		_w27876_,
		_w27877_
	);
	LUT4 #(
		.INIT('h4000)
	) name22051 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27878_
	);
	LUT4 #(
		.INIT('h0203)
	) name22052 (
		_w27864_,
		_w27862_,
		_w27863_,
		_w27859_,
		_w27879_
	);
	LUT3 #(
		.INIT('h13)
	) name22053 (
		_w27872_,
		_w27878_,
		_w27879_,
		_w27880_
	);
	LUT4 #(
		.INIT('h4555)
	) name22054 (
		_w27860_,
		_w27873_,
		_w27877_,
		_w27880_,
		_w27881_
	);
	LUT3 #(
		.INIT('h80)
	) name22055 (
		_w27862_,
		_w27863_,
		_w27860_,
		_w27882_
	);
	LUT3 #(
		.INIT('h51)
	) name22056 (
		_w27864_,
		_w27862_,
		_w27863_,
		_w27883_
	);
	LUT2 #(
		.INIT('h2)
	) name22057 (
		_w27860_,
		_w27859_,
		_w27884_
	);
	LUT4 #(
		.INIT('h0090)
	) name22058 (
		_w27861_,
		_w27862_,
		_w27860_,
		_w27859_,
		_w27885_
	);
	LUT4 #(
		.INIT('h7077)
	) name22059 (
		_w27866_,
		_w27882_,
		_w27883_,
		_w27885_,
		_w27886_
	);
	LUT4 #(
		.INIT('h5655)
	) name22060 (
		\u0_L9_reg[6]/NET0131 ,
		_w27881_,
		_w27870_,
		_w27886_,
		_w27887_
	);
	LUT2 #(
		.INIT('h2)
	) name22061 (
		_w27388_,
		_w27400_,
		_w27888_
	);
	LUT3 #(
		.INIT('h28)
	) name22062 (
		_w27391_,
		_w27390_,
		_w27392_,
		_w27889_
	);
	LUT4 #(
		.INIT('h877a)
	) name22063 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27890_
	);
	LUT2 #(
		.INIT('h2)
	) name22064 (
		_w27888_,
		_w27890_,
		_w27891_
	);
	LUT4 #(
		.INIT('h2880)
	) name22065 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27892_
	);
	LUT4 #(
		.INIT('h5004)
	) name22066 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27893_
	);
	LUT2 #(
		.INIT('h4)
	) name22067 (
		_w27388_,
		_w27400_,
		_w27894_
	);
	LUT2 #(
		.INIT('h9)
	) name22068 (
		_w27388_,
		_w27400_,
		_w27895_
	);
	LUT3 #(
		.INIT('h10)
	) name22069 (
		_w27892_,
		_w27893_,
		_w27895_,
		_w27896_
	);
	LUT4 #(
		.INIT('h21a1)
	) name22070 (
		_w27389_,
		_w27391_,
		_w27390_,
		_w27392_,
		_w27897_
	);
	LUT4 #(
		.INIT('h0010)
	) name22071 (
		_w27684_,
		_w27889_,
		_w27894_,
		_w27897_,
		_w27898_
	);
	LUT4 #(
		.INIT('h00ab)
	) name22072 (
		_w27393_,
		_w27891_,
		_w27896_,
		_w27898_,
		_w27899_
	);
	LUT2 #(
		.INIT('h6)
	) name22073 (
		\u0_L9_reg[7]/NET0131 ,
		_w27899_,
		_w27900_
	);
	LUT3 #(
		.INIT('h02)
	) name22074 (
		_w27628_,
		_w27651_,
		_w27639_,
		_w27901_
	);
	LUT4 #(
		.INIT('h3010)
	) name22075 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27902_
	);
	LUT4 #(
		.INIT('h00f7)
	) name22076 (
		_w27630_,
		_w27631_,
		_w27629_,
		_w27628_,
		_w27903_
	);
	LUT2 #(
		.INIT('h4)
	) name22077 (
		_w27902_,
		_w27903_,
		_w27904_
	);
	LUT4 #(
		.INIT('he6fd)
	) name22078 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27905_
	);
	LUT4 #(
		.INIT('h0155)
	) name22079 (
		_w27627_,
		_w27901_,
		_w27904_,
		_w27905_,
		_w27906_
	);
	LUT4 #(
		.INIT('h0001)
	) name22080 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27907_
	);
	LUT4 #(
		.INIT('hff3e)
	) name22081 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27908_
	);
	LUT3 #(
		.INIT('h04)
	) name22082 (
		_w27633_,
		_w27630_,
		_w27628_,
		_w27909_
	);
	LUT4 #(
		.INIT('h00c4)
	) name22083 (
		_w27628_,
		_w27660_,
		_w27908_,
		_w27909_,
		_w27910_
	);
	LUT4 #(
		.INIT('he5df)
	) name22084 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27911_
	);
	LUT4 #(
		.INIT('haf23)
	) name22085 (
		_w27631_,
		_w27628_,
		_w27741_,
		_w27911_,
		_w27912_
	);
	LUT3 #(
		.INIT('hd0)
	) name22086 (
		_w27627_,
		_w27910_,
		_w27912_,
		_w27913_
	);
	LUT3 #(
		.INIT('h65)
	) name22087 (
		\u0_L9_reg[8]/NET0131 ,
		_w27906_,
		_w27913_,
		_w27914_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name22088 (
		_w27446_,
		_w27445_,
		_w27444_,
		_w27447_,
		_w27915_
	);
	LUT3 #(
		.INIT('h0d)
	) name22089 (
		_w27445_,
		_w27448_,
		_w27447_,
		_w27916_
	);
	LUT4 #(
		.INIT('h8000)
	) name22090 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27917_
	);
	LUT4 #(
		.INIT('h0021)
	) name22091 (
		_w27445_,
		_w27444_,
		_w27448_,
		_w27447_,
		_w27918_
	);
	LUT4 #(
		.INIT('h0301)
	) name22092 (
		_w27915_,
		_w27917_,
		_w27918_,
		_w27916_,
		_w27919_
	);
	LUT4 #(
		.INIT('h4300)
	) name22093 (
		_w27446_,
		_w27445_,
		_w27444_,
		_w27447_,
		_w27920_
	);
	LUT4 #(
		.INIT('h0082)
	) name22094 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27921_
	);
	LUT4 #(
		.INIT('h0414)
	) name22095 (
		_w27446_,
		_w27445_,
		_w27448_,
		_w27447_,
		_w27922_
	);
	LUT4 #(
		.INIT('h0001)
	) name22096 (
		_w27465_,
		_w27921_,
		_w27922_,
		_w27920_,
		_w27923_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name22097 (
		_w27446_,
		_w27445_,
		_w27468_,
		_w27456_,
		_w27924_
	);
	LUT4 #(
		.INIT('hd800)
	) name22098 (
		_w27443_,
		_w27923_,
		_w27919_,
		_w27924_,
		_w27925_
	);
	LUT2 #(
		.INIT('h9)
	) name22099 (
		\u0_L9_reg[19]/P0001 ,
		_w27925_,
		_w27926_
	);
	LUT3 #(
		.INIT('h80)
	) name22100 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27927_
	);
	LUT4 #(
		.INIT('h6979)
	) name22101 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27859_,
		_w27928_
	);
	LUT3 #(
		.INIT('h04)
	) name22102 (
		_w27861_,
		_w27864_,
		_w27863_,
		_w27929_
	);
	LUT4 #(
		.INIT('h0014)
	) name22103 (
		_w27861_,
		_w27864_,
		_w27863_,
		_w27859_,
		_w27930_
	);
	LUT4 #(
		.INIT('h0302)
	) name22104 (
		_w27863_,
		_w27874_,
		_w27930_,
		_w27928_,
		_w27931_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name22105 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27932_
	);
	LUT4 #(
		.INIT('h6800)
	) name22106 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27859_,
		_w27933_
	);
	LUT4 #(
		.INIT('h0032)
	) name22107 (
		_w27859_,
		_w27868_,
		_w27932_,
		_w27933_,
		_w27934_
	);
	LUT4 #(
		.INIT('h0020)
	) name22108 (
		_w27864_,
		_w27862_,
		_w27863_,
		_w27859_,
		_w27935_
	);
	LUT4 #(
		.INIT('hbeff)
	) name22109 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27936_
	);
	LUT3 #(
		.INIT('h31)
	) name22110 (
		_w27859_,
		_w27935_,
		_w27936_,
		_w27937_
	);
	LUT4 #(
		.INIT('hd800)
	) name22111 (
		_w27860_,
		_w27931_,
		_w27934_,
		_w27937_,
		_w27938_
	);
	LUT2 #(
		.INIT('h9)
	) name22112 (
		\u0_L9_reg[16]/NET0131 ,
		_w27938_,
		_w27939_
	);
	LUT4 #(
		.INIT('h0400)
	) name22113 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27940_
	);
	LUT4 #(
		.INIT('he2cd)
	) name22114 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27941_
	);
	LUT4 #(
		.INIT('h5054)
	) name22115 (
		_w27860_,
		_w27859_,
		_w27940_,
		_w27941_,
		_w27942_
	);
	LUT4 #(
		.INIT('h1df2)
	) name22116 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27943_
	);
	LUT2 #(
		.INIT('h2)
	) name22117 (
		_w27859_,
		_w27943_,
		_w27944_
	);
	LUT4 #(
		.INIT('hfe3e)
	) name22118 (
		_w27859_,
		_w27872_,
		_w27867_,
		_w27875_,
		_w27945_
	);
	LUT3 #(
		.INIT('h8a)
	) name22119 (
		_w27860_,
		_w27944_,
		_w27945_,
		_w27946_
	);
	LUT4 #(
		.INIT('h9db6)
	) name22120 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27947_
	);
	LUT2 #(
		.INIT('h1)
	) name22121 (
		_w27860_,
		_w27859_,
		_w27948_
	);
	LUT2 #(
		.INIT('h4)
	) name22122 (
		_w27947_,
		_w27948_,
		_w27949_
	);
	LUT2 #(
		.INIT('h8)
	) name22123 (
		_w27861_,
		_w27876_,
		_w27950_
	);
	LUT2 #(
		.INIT('h4)
	) name22124 (
		_w27862_,
		_w27859_,
		_w27951_
	);
	LUT2 #(
		.INIT('h2)
	) name22125 (
		_w27863_,
		_w27859_,
		_w27952_
	);
	LUT4 #(
		.INIT('h135f)
	) name22126 (
		_w27929_,
		_w27927_,
		_w27951_,
		_w27952_,
		_w27953_
	);
	LUT3 #(
		.INIT('h10)
	) name22127 (
		_w27949_,
		_w27950_,
		_w27953_,
		_w27954_
	);
	LUT4 #(
		.INIT('h5655)
	) name22128 (
		\u0_L9_reg[24]/NET0131 ,
		_w27946_,
		_w27942_,
		_w27954_,
		_w27955_
	);
	LUT4 #(
		.INIT('h23af)
	) name22129 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27956_
	);
	LUT4 #(
		.INIT('hbf00)
	) name22130 (
		_w27861_,
		_w27862_,
		_w27863_,
		_w27859_,
		_w27957_
	);
	LUT3 #(
		.INIT('h0e)
	) name22131 (
		_w27864_,
		_w27862_,
		_w27859_,
		_w27958_
	);
	LUT4 #(
		.INIT('hfdf6)
	) name22132 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27959_
	);
	LUT4 #(
		.INIT('h2700)
	) name22133 (
		_w27956_,
		_w27958_,
		_w27957_,
		_w27959_,
		_w27960_
	);
	LUT2 #(
		.INIT('h1)
	) name22134 (
		_w27860_,
		_w27960_,
		_w27961_
	);
	LUT4 #(
		.INIT('h1200)
	) name22135 (
		_w27861_,
		_w27864_,
		_w27863_,
		_w27859_,
		_w27962_
	);
	LUT4 #(
		.INIT('haa80)
	) name22136 (
		_w27860_,
		_w27929_,
		_w27951_,
		_w27962_,
		_w27963_
	);
	LUT4 #(
		.INIT('h23ef)
	) name22137 (
		_w27861_,
		_w27864_,
		_w27862_,
		_w27863_,
		_w27964_
	);
	LUT2 #(
		.INIT('h2)
	) name22138 (
		_w27884_,
		_w27964_,
		_w27965_
	);
	LUT3 #(
		.INIT('h80)
	) name22139 (
		_w27861_,
		_w27864_,
		_w27863_,
		_w27966_
	);
	LUT2 #(
		.INIT('h8)
	) name22140 (
		_w27951_,
		_w27966_,
		_w27967_
	);
	LUT4 #(
		.INIT('h0040)
	) name22141 (
		_w27861_,
		_w27862_,
		_w27863_,
		_w27859_,
		_w27968_
	);
	LUT3 #(
		.INIT('h0d)
	) name22142 (
		_w27882_,
		_w27871_,
		_w27968_,
		_w27969_
	);
	LUT4 #(
		.INIT('h0100)
	) name22143 (
		_w27963_,
		_w27965_,
		_w27967_,
		_w27969_,
		_w27970_
	);
	LUT3 #(
		.INIT('h9a)
	) name22144 (
		\u0_L9_reg[30]/NET0131 ,
		_w27961_,
		_w27970_,
		_w27971_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name22145 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27972_
	);
	LUT2 #(
		.INIT('h2)
	) name22146 (
		_w27628_,
		_w27972_,
		_w27973_
	);
	LUT4 #(
		.INIT('h0040)
	) name22147 (
		_w27630_,
		_w27631_,
		_w27629_,
		_w27628_,
		_w27974_
	);
	LUT4 #(
		.INIT('h0004)
	) name22148 (
		_w27652_,
		_w27627_,
		_w27642_,
		_w27974_,
		_w27975_
	);
	LUT4 #(
		.INIT('he3ef)
	) name22149 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27976_
	);
	LUT2 #(
		.INIT('h2)
	) name22150 (
		_w27628_,
		_w27976_,
		_w27977_
	);
	LUT4 #(
		.INIT('h5010)
	) name22151 (
		_w27633_,
		_w27630_,
		_w27631_,
		_w27629_,
		_w27978_
	);
	LUT3 #(
		.INIT('hd0)
	) name22152 (
		_w27633_,
		_w27629_,
		_w27628_,
		_w27979_
	);
	LUT4 #(
		.INIT('h5554)
	) name22153 (
		_w27627_,
		_w27632_,
		_w27979_,
		_w27978_,
		_w27980_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name22154 (
		_w27973_,
		_w27975_,
		_w27977_,
		_w27980_,
		_w27981_
	);
	LUT3 #(
		.INIT('h02)
	) name22155 (
		_w27628_,
		_w27651_,
		_w27659_,
		_w27982_
	);
	LUT4 #(
		.INIT('h0001)
	) name22156 (
		_w27628_,
		_w27655_,
		_w27641_,
		_w27907_,
		_w27983_
	);
	LUT2 #(
		.INIT('h1)
	) name22157 (
		_w27982_,
		_w27983_,
		_w27984_
	);
	LUT3 #(
		.INIT('h56)
	) name22158 (
		\u0_L9_reg[3]/NET0131 ,
		_w27981_,
		_w27984_,
		_w27985_
	);
	LUT4 #(
		.INIT('h2600)
	) name22159 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27565_,
		_w27986_
	);
	LUT3 #(
		.INIT('h07)
	) name22160 (
		_w27567_,
		_w27569_,
		_w27565_,
		_w27987_
	);
	LUT4 #(
		.INIT('h0103)
	) name22161 (
		_w27581_,
		_w27775_,
		_w27986_,
		_w27987_,
		_w27988_
	);
	LUT4 #(
		.INIT('h0121)
	) name22162 (
		_w27566_,
		_w27568_,
		_w27569_,
		_w27565_,
		_w27989_
	);
	LUT3 #(
		.INIT('h1b)
	) name22163 (
		_w27566_,
		_w27569_,
		_w27565_,
		_w27990_
	);
	LUT4 #(
		.INIT('hdfee)
	) name22164 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27991_
	);
	LUT4 #(
		.INIT('h0d00)
	) name22165 (
		_w27575_,
		_w27990_,
		_w27989_,
		_w27991_,
		_w27992_
	);
	LUT4 #(
		.INIT('h0008)
	) name22166 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27565_,
		_w27993_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name22167 (
		_w27566_,
		_w27567_,
		_w27568_,
		_w27569_,
		_w27994_
	);
	LUT3 #(
		.INIT('h31)
	) name22168 (
		_w27565_,
		_w27993_,
		_w27994_,
		_w27995_
	);
	LUT4 #(
		.INIT('he400)
	) name22169 (
		_w27578_,
		_w27992_,
		_w27988_,
		_w27995_,
		_w27996_
	);
	LUT2 #(
		.INIT('h9)
	) name22170 (
		\u0_L9_reg[18]/NET0131 ,
		_w27996_,
		_w27997_
	);
	LUT4 #(
		.INIT('hc963)
	) name22171 (
		decrypt_pad,
		\u0_R8_reg[4]/NET0131 ,
		\u0_uk_K_r8_reg[11]/NET0131 ,
		\u0_uk_K_r8_reg[33]/NET0131 ,
		_w27998_
	);
	LUT4 #(
		.INIT('hc693)
	) name22172 (
		decrypt_pad,
		\u0_R8_reg[32]/NET0131 ,
		\u0_uk_K_r8_reg[10]/NET0131 ,
		\u0_uk_K_r8_reg[20]/NET0131 ,
		_w27999_
	);
	LUT4 #(
		.INIT('hc963)
	) name22173 (
		decrypt_pad,
		\u0_R8_reg[5]/NET0131 ,
		\u0_uk_K_r8_reg[39]/NET0131 ,
		\u0_uk_K_r8_reg[4]/NET0131 ,
		_w28000_
	);
	LUT2 #(
		.INIT('h1)
	) name22174 (
		_w27999_,
		_w28000_,
		_w28001_
	);
	LUT4 #(
		.INIT('hc963)
	) name22175 (
		decrypt_pad,
		\u0_R8_reg[3]/NET0131 ,
		\u0_uk_K_r8_reg[33]/NET0131 ,
		\u0_uk_K_r8_reg[55]/NET0131 ,
		_w28002_
	);
	LUT4 #(
		.INIT('hc963)
	) name22176 (
		decrypt_pad,
		\u0_R8_reg[2]/NET0131 ,
		\u0_uk_K_r8_reg[24]/NET0131 ,
		\u0_uk_K_r8_reg[46]/NET0131 ,
		_w28003_
	);
	LUT3 #(
		.INIT('h02)
	) name22177 (
		_w28002_,
		_w28003_,
		_w27999_,
		_w28004_
	);
	LUT4 #(
		.INIT('hc963)
	) name22178 (
		decrypt_pad,
		\u0_R8_reg[1]/NET0131 ,
		\u0_uk_K_r8_reg[41]/NET0131 ,
		\u0_uk_K_r8_reg[6]/NET0131 ,
		_w28005_
	);
	LUT4 #(
		.INIT('hffc8)
	) name22179 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28006_
	);
	LUT3 #(
		.INIT('h45)
	) name22180 (
		_w28001_,
		_w28004_,
		_w28006_,
		_w28007_
	);
	LUT4 #(
		.INIT('hfd0d)
	) name22181 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28008_
	);
	LUT4 #(
		.INIT('haff3)
	) name22182 (
		_w28002_,
		_w28003_,
		_w27999_,
		_w28005_,
		_w28009_
	);
	LUT3 #(
		.INIT('hd0)
	) name22183 (
		_w28002_,
		_w28008_,
		_w28009_,
		_w28010_
	);
	LUT3 #(
		.INIT('h8a)
	) name22184 (
		_w27998_,
		_w28007_,
		_w28010_,
		_w28011_
	);
	LUT4 #(
		.INIT('h7c3f)
	) name22185 (
		_w28002_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28012_
	);
	LUT2 #(
		.INIT('h1)
	) name22186 (
		_w28003_,
		_w28012_,
		_w28013_
	);
	LUT2 #(
		.INIT('h8)
	) name22187 (
		_w28002_,
		_w28003_,
		_w28014_
	);
	LUT3 #(
		.INIT('h60)
	) name22188 (
		_w27999_,
		_w28000_,
		_w28005_,
		_w28015_
	);
	LUT4 #(
		.INIT('h0008)
	) name22189 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28016_
	);
	LUT4 #(
		.INIT('heef6)
	) name22190 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28017_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name22191 (
		_w28002_,
		_w28003_,
		_w28015_,
		_w28017_,
		_w28018_
	);
	LUT3 #(
		.INIT('h45)
	) name22192 (
		_w27998_,
		_w28013_,
		_w28018_,
		_w28019_
	);
	LUT4 #(
		.INIT('h8000)
	) name22193 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28020_
	);
	LUT3 #(
		.INIT('h47)
	) name22194 (
		_w28003_,
		_w28000_,
		_w28005_,
		_w28021_
	);
	LUT4 #(
		.INIT('h7adf)
	) name22195 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28022_
	);
	LUT2 #(
		.INIT('h1)
	) name22196 (
		_w28002_,
		_w28022_,
		_w28023_
	);
	LUT2 #(
		.INIT('h1)
	) name22197 (
		_w28003_,
		_w28005_,
		_w28024_
	);
	LUT4 #(
		.INIT('h0020)
	) name22198 (
		_w28002_,
		_w28003_,
		_w27999_,
		_w28005_,
		_w28025_
	);
	LUT3 #(
		.INIT('h08)
	) name22199 (
		_w28002_,
		_w28003_,
		_w28005_,
		_w28026_
	);
	LUT3 #(
		.INIT('h13)
	) name22200 (
		_w28001_,
		_w28025_,
		_w28026_,
		_w28027_
	);
	LUT2 #(
		.INIT('h4)
	) name22201 (
		_w28023_,
		_w28027_,
		_w28028_
	);
	LUT4 #(
		.INIT('h5655)
	) name22202 (
		\u0_L8_reg[31]/NET0131 ,
		_w28019_,
		_w28011_,
		_w28028_,
		_w28029_
	);
	LUT4 #(
		.INIT('hc693)
	) name22203 (
		decrypt_pad,
		\u0_R8_reg[24]/NET0131 ,
		\u0_uk_K_r8_reg[2]/NET0131 ,
		\u0_uk_K_r8_reg[37]/P0001 ,
		_w28030_
	);
	LUT4 #(
		.INIT('hc693)
	) name22204 (
		decrypt_pad,
		\u0_R8_reg[23]/NET0131 ,
		\u0_uk_K_r8_reg[0]/NET0131 ,
		\u0_uk_K_r8_reg[35]/NET0131 ,
		_w28031_
	);
	LUT4 #(
		.INIT('hc963)
	) name22205 (
		decrypt_pad,
		\u0_R8_reg[20]/NET0131 ,
		\u0_uk_K_r8_reg[16]/NET0131 ,
		\u0_uk_K_r8_reg[36]/NET0131 ,
		_w28032_
	);
	LUT4 #(
		.INIT('hc963)
	) name22206 (
		decrypt_pad,
		\u0_R8_reg[21]/NET0131 ,
		\u0_uk_K_r8_reg[0]/NET0131 ,
		\u0_uk_K_r8_reg[51]/NET0131 ,
		_w28033_
	);
	LUT4 #(
		.INIT('hc963)
	) name22207 (
		decrypt_pad,
		\u0_R8_reg[25]/NET0131 ,
		\u0_uk_K_r8_reg[1]/NET0131 ,
		\u0_uk_K_r8_reg[21]/NET0131 ,
		_w28034_
	);
	LUT4 #(
		.INIT('hc963)
	) name22208 (
		decrypt_pad,
		\u0_R8_reg[22]/NET0131 ,
		\u0_uk_K_r8_reg[22]/NET0131 ,
		\u0_uk_K_r8_reg[42]/NET0131 ,
		_w28035_
	);
	LUT4 #(
		.INIT('h0002)
	) name22209 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28036_
	);
	LUT4 #(
		.INIT('h27fd)
	) name22210 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28037_
	);
	LUT2 #(
		.INIT('h2)
	) name22211 (
		_w28031_,
		_w28037_,
		_w28038_
	);
	LUT2 #(
		.INIT('h1)
	) name22212 (
		_w28031_,
		_w28035_,
		_w28039_
	);
	LUT4 #(
		.INIT('h0008)
	) name22213 (
		_w28032_,
		_w28034_,
		_w28031_,
		_w28035_,
		_w28040_
	);
	LUT3 #(
		.INIT('hbc)
	) name22214 (
		_w28032_,
		_w28035_,
		_w28033_,
		_w28041_
	);
	LUT4 #(
		.INIT('h0704)
	) name22215 (
		_w28032_,
		_w28034_,
		_w28031_,
		_w28035_,
		_w28042_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name22216 (
		_w28033_,
		_w28040_,
		_w28041_,
		_w28042_,
		_w28043_
	);
	LUT3 #(
		.INIT('h8a)
	) name22217 (
		_w28030_,
		_w28038_,
		_w28043_,
		_w28044_
	);
	LUT4 #(
		.INIT('h0080)
	) name22218 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28045_
	);
	LUT2 #(
		.INIT('h2)
	) name22219 (
		_w28032_,
		_w28034_,
		_w28046_
	);
	LUT3 #(
		.INIT('hce)
	) name22220 (
		_w28031_,
		_w28035_,
		_w28033_,
		_w28047_
	);
	LUT4 #(
		.INIT('h0040)
	) name22221 (
		_w28032_,
		_w28034_,
		_w28031_,
		_w28033_,
		_w28048_
	);
	LUT4 #(
		.INIT('h000d)
	) name22222 (
		_w28046_,
		_w28047_,
		_w28048_,
		_w28045_,
		_w28049_
	);
	LUT4 #(
		.INIT('he97b)
	) name22223 (
		_w28032_,
		_w28031_,
		_w28035_,
		_w28033_,
		_w28050_
	);
	LUT3 #(
		.INIT('h15)
	) name22224 (
		_w28030_,
		_w28049_,
		_w28050_,
		_w28051_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name22225 (
		_w28032_,
		_w28034_,
		_w28031_,
		_w28033_,
		_w28052_
	);
	LUT2 #(
		.INIT('h1)
	) name22226 (
		_w28035_,
		_w28052_,
		_w28053_
	);
	LUT3 #(
		.INIT('h0e)
	) name22227 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28054_
	);
	LUT3 #(
		.INIT('h70)
	) name22228 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28055_
	);
	LUT3 #(
		.INIT('ha8)
	) name22229 (
		_w28031_,
		_w28035_,
		_w28033_,
		_w28056_
	);
	LUT3 #(
		.INIT('h10)
	) name22230 (
		_w28055_,
		_w28054_,
		_w28056_,
		_w28057_
	);
	LUT3 #(
		.INIT('h01)
	) name22231 (
		_w28032_,
		_w28034_,
		_w28033_,
		_w28058_
	);
	LUT2 #(
		.INIT('h8)
	) name22232 (
		_w28039_,
		_w28058_,
		_w28059_
	);
	LUT3 #(
		.INIT('h01)
	) name22233 (
		_w28057_,
		_w28053_,
		_w28059_,
		_w28060_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name22234 (
		\u0_L8_reg[11]/NET0131 ,
		_w28051_,
		_w28044_,
		_w28060_,
		_w28061_
	);
	LUT4 #(
		.INIT('hc963)
	) name22235 (
		decrypt_pad,
		\u0_R8_reg[28]/NET0131 ,
		\u0_uk_K_r8_reg[44]/NET0131 ,
		\u0_uk_K_r8_reg[9]/P0001 ,
		_w28062_
	);
	LUT4 #(
		.INIT('hc693)
	) name22236 (
		decrypt_pad,
		\u0_R8_reg[27]/NET0131 ,
		\u0_uk_K_r8_reg[22]/NET0131 ,
		\u0_uk_K_r8_reg[2]/NET0131 ,
		_w28063_
	);
	LUT4 #(
		.INIT('hc963)
	) name22237 (
		decrypt_pad,
		\u0_R8_reg[24]/NET0131 ,
		\u0_uk_K_r8_reg[28]/NET0131 ,
		\u0_uk_K_r8_reg[52]/NET0131 ,
		_w28064_
	);
	LUT4 #(
		.INIT('hc693)
	) name22238 (
		decrypt_pad,
		\u0_R8_reg[25]/NET0131 ,
		\u0_uk_K_r8_reg[28]/NET0131 ,
		\u0_uk_K_r8_reg[8]/NET0131 ,
		_w28065_
	);
	LUT4 #(
		.INIT('hc693)
	) name22239 (
		decrypt_pad,
		\u0_R8_reg[29]/NET0131 ,
		\u0_uk_K_r8_reg[1]/NET0131 ,
		\u0_uk_K_r8_reg[36]/NET0131 ,
		_w28066_
	);
	LUT4 #(
		.INIT('hc693)
	) name22240 (
		decrypt_pad,
		\u0_R8_reg[26]/NET0131 ,
		\u0_uk_K_r8_reg[44]/NET0131 ,
		\u0_uk_K_r8_reg[52]/NET0131 ,
		_w28067_
	);
	LUT4 #(
		.INIT('h0004)
	) name22241 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28068_
	);
	LUT4 #(
		.INIT('h775b)
	) name22242 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28069_
	);
	LUT2 #(
		.INIT('h1)
	) name22243 (
		_w28063_,
		_w28069_,
		_w28070_
	);
	LUT2 #(
		.INIT('h1)
	) name22244 (
		_w28067_,
		_w28065_,
		_w28071_
	);
	LUT3 #(
		.INIT('h8a)
	) name22245 (
		_w28064_,
		_w28063_,
		_w28066_,
		_w28072_
	);
	LUT2 #(
		.INIT('h6)
	) name22246 (
		_w28064_,
		_w28067_,
		_w28073_
	);
	LUT4 #(
		.INIT('h9000)
	) name22247 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28074_
	);
	LUT4 #(
		.INIT('h0100)
	) name22248 (
		_w28064_,
		_w28067_,
		_w28063_,
		_w28066_,
		_w28075_
	);
	LUT4 #(
		.INIT('h0111)
	) name22249 (
		_w28074_,
		_w28075_,
		_w28071_,
		_w28072_,
		_w28076_
	);
	LUT3 #(
		.INIT('h45)
	) name22250 (
		_w28062_,
		_w28070_,
		_w28076_,
		_w28077_
	);
	LUT2 #(
		.INIT('h6)
	) name22251 (
		_w28067_,
		_w28065_,
		_w28078_
	);
	LUT4 #(
		.INIT('h8808)
	) name22252 (
		_w28064_,
		_w28063_,
		_w28065_,
		_w28066_,
		_w28079_
	);
	LUT2 #(
		.INIT('h8)
	) name22253 (
		_w28078_,
		_w28079_,
		_w28080_
	);
	LUT4 #(
		.INIT('h0401)
	) name22254 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28081_
	);
	LUT2 #(
		.INIT('h6)
	) name22255 (
		_w28064_,
		_w28065_,
		_w28082_
	);
	LUT4 #(
		.INIT('h0700)
	) name22256 (
		_w28064_,
		_w28067_,
		_w28063_,
		_w28066_,
		_w28083_
	);
	LUT3 #(
		.INIT('h15)
	) name22257 (
		_w28081_,
		_w28082_,
		_w28083_,
		_w28084_
	);
	LUT4 #(
		.INIT('h0900)
	) name22258 (
		_w28064_,
		_w28067_,
		_w28063_,
		_w28065_,
		_w28085_
	);
	LUT2 #(
		.INIT('h4)
	) name22259 (
		_w28065_,
		_w28066_,
		_w28086_
	);
	LUT4 #(
		.INIT('h0440)
	) name22260 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28087_
	);
	LUT4 #(
		.INIT('hfbb4)
	) name22261 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28088_
	);
	LUT3 #(
		.INIT('h31)
	) name22262 (
		_w28063_,
		_w28085_,
		_w28088_,
		_w28089_
	);
	LUT4 #(
		.INIT('h7500)
	) name22263 (
		_w28062_,
		_w28080_,
		_w28084_,
		_w28089_,
		_w28090_
	);
	LUT3 #(
		.INIT('h65)
	) name22264 (
		\u0_L8_reg[22]/NET0131 ,
		_w28077_,
		_w28090_,
		_w28091_
	);
	LUT4 #(
		.INIT('hfe3c)
	) name22265 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28092_
	);
	LUT4 #(
		.INIT('h8008)
	) name22266 (
		_w28002_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28093_
	);
	LUT4 #(
		.INIT('hf7df)
	) name22267 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28094_
	);
	LUT4 #(
		.INIT('h0e00)
	) name22268 (
		_w28002_,
		_w28092_,
		_w28093_,
		_w28094_,
		_w28095_
	);
	LUT4 #(
		.INIT('h0040)
	) name22269 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28096_
	);
	LUT4 #(
		.INIT('hcc9d)
	) name22270 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28097_
	);
	LUT4 #(
		.INIT('h4041)
	) name22271 (
		_w28002_,
		_w28003_,
		_w27999_,
		_w28005_,
		_w28098_
	);
	LUT4 #(
		.INIT('h0400)
	) name22272 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28099_
	);
	LUT4 #(
		.INIT('h5bff)
	) name22273 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28100_
	);
	LUT4 #(
		.INIT('h0d00)
	) name22274 (
		_w28002_,
		_w28097_,
		_w28098_,
		_w28100_,
		_w28101_
	);
	LUT3 #(
		.INIT('hed)
	) name22275 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28102_
	);
	LUT2 #(
		.INIT('h8)
	) name22276 (
		_w28002_,
		_w28005_,
		_w28103_
	);
	LUT2 #(
		.INIT('h4)
	) name22277 (
		_w28102_,
		_w28103_,
		_w28104_
	);
	LUT4 #(
		.INIT('h00d8)
	) name22278 (
		_w27998_,
		_w28101_,
		_w28095_,
		_w28104_,
		_w28105_
	);
	LUT2 #(
		.INIT('h9)
	) name22279 (
		\u0_L8_reg[17]/NET0131 ,
		_w28105_,
		_w28106_
	);
	LUT4 #(
		.INIT('hc693)
	) name22280 (
		decrypt_pad,
		\u0_R8_reg[13]/NET0131 ,
		\u0_uk_K_r8_reg[18]/NET0131 ,
		\u0_uk_K_r8_reg[53]/NET0131 ,
		_w28107_
	);
	LUT4 #(
		.INIT('hc693)
	) name22281 (
		decrypt_pad,
		\u0_R8_reg[15]/NET0131 ,
		\u0_uk_K_r8_reg[27]/NET0131 ,
		\u0_uk_K_r8_reg[5]/NET0131 ,
		_w28108_
	);
	LUT4 #(
		.INIT('hc963)
	) name22282 (
		decrypt_pad,
		\u0_R8_reg[17]/NET0131 ,
		\u0_uk_K_r8_reg[18]/NET0131 ,
		\u0_uk_K_r8_reg[40]/NET0131 ,
		_w28109_
	);
	LUT4 #(
		.INIT('hc693)
	) name22283 (
		decrypt_pad,
		\u0_R8_reg[12]/NET0131 ,
		\u0_uk_K_r8_reg[24]/NET0131 ,
		\u0_uk_K_r8_reg[34]/NET0131 ,
		_w28110_
	);
	LUT2 #(
		.INIT('h2)
	) name22284 (
		_w28109_,
		_w28110_,
		_w28111_
	);
	LUT4 #(
		.INIT('h0200)
	) name22285 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28108_,
		_w28112_
	);
	LUT4 #(
		.INIT('hc963)
	) name22286 (
		decrypt_pad,
		\u0_R8_reg[16]/NET0131 ,
		\u0_uk_K_r8_reg[13]/P0001 ,
		\u0_uk_K_r8_reg[3]/NET0131 ,
		_w28113_
	);
	LUT4 #(
		.INIT('hc693)
	) name22287 (
		decrypt_pad,
		\u0_R8_reg[14]/NET0131 ,
		\u0_uk_K_r8_reg[19]/NET0131 ,
		\u0_uk_K_r8_reg[54]/NET0131 ,
		_w28114_
	);
	LUT2 #(
		.INIT('h2)
	) name22288 (
		_w28107_,
		_w28110_,
		_w28115_
	);
	LUT4 #(
		.INIT('h0006)
	) name22289 (
		_w28107_,
		_w28110_,
		_w28114_,
		_w28108_,
		_w28116_
	);
	LUT4 #(
		.INIT('h8000)
	) name22290 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28117_
	);
	LUT4 #(
		.INIT('h0100)
	) name22291 (
		_w28112_,
		_w28116_,
		_w28117_,
		_w28113_,
		_w28118_
	);
	LUT4 #(
		.INIT('h4000)
	) name22292 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28108_,
		_w28119_
	);
	LUT3 #(
		.INIT('h08)
	) name22293 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28120_
	);
	LUT4 #(
		.INIT('h0008)
	) name22294 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28121_
	);
	LUT2 #(
		.INIT('h1)
	) name22295 (
		_w28119_,
		_w28121_,
		_w28122_
	);
	LUT4 #(
		.INIT('h0001)
	) name22296 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28108_,
		_w28123_
	);
	LUT4 #(
		.INIT('h0123)
	) name22297 (
		_w28114_,
		_w28119_,
		_w28120_,
		_w28123_,
		_w28124_
	);
	LUT2 #(
		.INIT('h8)
	) name22298 (
		_w28118_,
		_w28124_,
		_w28125_
	);
	LUT4 #(
		.INIT('h0100)
	) name22299 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28108_,
		_w28126_
	);
	LUT4 #(
		.INIT('h8000)
	) name22300 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28108_,
		_w28127_
	);
	LUT3 #(
		.INIT('h01)
	) name22301 (
		_w28113_,
		_w28126_,
		_w28127_,
		_w28128_
	);
	LUT3 #(
		.INIT('h80)
	) name22302 (
		_w28107_,
		_w28114_,
		_w28108_,
		_w28129_
	);
	LUT4 #(
		.INIT('h2000)
	) name22303 (
		_w28107_,
		_w28110_,
		_w28114_,
		_w28108_,
		_w28130_
	);
	LUT4 #(
		.INIT('h0020)
	) name22304 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28131_
	);
	LUT2 #(
		.INIT('h1)
	) name22305 (
		_w28130_,
		_w28131_,
		_w28132_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name22306 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28133_
	);
	LUT4 #(
		.INIT('h8ddd)
	) name22307 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28134_
	);
	LUT3 #(
		.INIT('hc8)
	) name22308 (
		_w28108_,
		_w28133_,
		_w28134_,
		_w28135_
	);
	LUT3 #(
		.INIT('h80)
	) name22309 (
		_w28128_,
		_w28132_,
		_w28135_,
		_w28136_
	);
	LUT4 #(
		.INIT('heffe)
	) name22310 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28137_
	);
	LUT2 #(
		.INIT('h4)
	) name22311 (
		_w28137_,
		_w28108_,
		_w28138_
	);
	LUT3 #(
		.INIT('h02)
	) name22312 (
		_w28109_,
		_w28114_,
		_w28108_,
		_w28139_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name22313 (
		_w28114_,
		_w28119_,
		_w28115_,
		_w28139_,
		_w28140_
	);
	LUT2 #(
		.INIT('h4)
	) name22314 (
		_w28138_,
		_w28140_,
		_w28141_
	);
	LUT4 #(
		.INIT('ha955)
	) name22315 (
		\u0_L8_reg[20]/NET0131 ,
		_w28125_,
		_w28136_,
		_w28141_,
		_w28142_
	);
	LUT4 #(
		.INIT('h67dc)
	) name22316 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28143_
	);
	LUT4 #(
		.INIT('h0d08)
	) name22317 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28144_
	);
	LUT4 #(
		.INIT('hd2f7)
	) name22318 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28145_
	);
	LUT4 #(
		.INIT('h0040)
	) name22319 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28146_
	);
	LUT4 #(
		.INIT('h00e4)
	) name22320 (
		_w28031_,
		_w28145_,
		_w28143_,
		_w28146_,
		_w28147_
	);
	LUT2 #(
		.INIT('h1)
	) name22321 (
		_w28030_,
		_w28147_,
		_w28148_
	);
	LUT4 #(
		.INIT('h9aff)
	) name22322 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28149_
	);
	LUT2 #(
		.INIT('h2)
	) name22323 (
		_w28031_,
		_w28149_,
		_w28150_
	);
	LUT3 #(
		.INIT('h60)
	) name22324 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28151_
	);
	LUT4 #(
		.INIT('hcc04)
	) name22325 (
		_w28034_,
		_w28031_,
		_w28035_,
		_w28033_,
		_w28152_
	);
	LUT3 #(
		.INIT('h01)
	) name22326 (
		_w28144_,
		_w28152_,
		_w28151_,
		_w28153_
	);
	LUT4 #(
		.INIT('h0800)
	) name22327 (
		_w28034_,
		_w28031_,
		_w28035_,
		_w28033_,
		_w28154_
	);
	LUT2 #(
		.INIT('h1)
	) name22328 (
		_w28036_,
		_w28154_,
		_w28155_
	);
	LUT4 #(
		.INIT('h5700)
	) name22329 (
		_w28030_,
		_w28150_,
		_w28153_,
		_w28155_,
		_w28156_
	);
	LUT3 #(
		.INIT('h9a)
	) name22330 (
		\u0_L8_reg[29]/NET0131 ,
		_w28148_,
		_w28156_,
		_w28157_
	);
	LUT4 #(
		.INIT('hc693)
	) name22331 (
		decrypt_pad,
		\u0_R8_reg[7]/NET0131 ,
		\u0_uk_K_r8_reg[11]/NET0131 ,
		\u0_uk_K_r8_reg[46]/NET0131 ,
		_w28158_
	);
	LUT4 #(
		.INIT('hc963)
	) name22332 (
		decrypt_pad,
		\u0_R8_reg[9]/NET0131 ,
		\u0_uk_K_r8_reg[17]/NET0131 ,
		\u0_uk_K_r8_reg[39]/NET0131 ,
		_w28159_
	);
	LUT4 #(
		.INIT('hc963)
	) name22333 (
		decrypt_pad,
		\u0_R8_reg[4]/NET0131 ,
		\u0_uk_K_r8_reg[25]/NET0131 ,
		\u0_uk_K_r8_reg[47]/NET0131 ,
		_w28160_
	);
	LUT4 #(
		.INIT('hc693)
	) name22334 (
		decrypt_pad,
		\u0_R8_reg[5]/NET0131 ,
		\u0_uk_K_r8_reg[26]/NET0131 ,
		\u0_uk_K_r8_reg[4]/NET0131 ,
		_w28161_
	);
	LUT4 #(
		.INIT('hc693)
	) name22335 (
		decrypt_pad,
		\u0_R8_reg[6]/NET0131 ,
		\u0_uk_K_r8_reg[17]/NET0131 ,
		\u0_uk_K_r8_reg[27]/NET0131 ,
		_w28162_
	);
	LUT4 #(
		.INIT('h2002)
	) name22336 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28163_
	);
	LUT4 #(
		.INIT('hc963)
	) name22337 (
		decrypt_pad,
		\u0_R8_reg[8]/NET0131 ,
		\u0_uk_K_r8_reg[12]/NET0131 ,
		\u0_uk_K_r8_reg[34]/NET0131 ,
		_w28164_
	);
	LUT3 #(
		.INIT('h3b)
	) name22338 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28165_
	);
	LUT4 #(
		.INIT('h39fd)
	) name22339 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28166_
	);
	LUT4 #(
		.INIT('h5051)
	) name22340 (
		_w28158_,
		_w28164_,
		_w28163_,
		_w28166_,
		_w28167_
	);
	LUT4 #(
		.INIT('h0b7b)
	) name22341 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28158_,
		_w28168_
	);
	LUT2 #(
		.INIT('h1)
	) name22342 (
		_w28168_,
		_w28162_,
		_w28169_
	);
	LUT3 #(
		.INIT('h54)
	) name22343 (
		_w28160_,
		_w28161_,
		_w28158_,
		_w28170_
	);
	LUT4 #(
		.INIT('hc001)
	) name22344 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28158_,
		_w28171_
	);
	LUT4 #(
		.INIT('h0d00)
	) name22345 (
		_w28159_,
		_w28160_,
		_w28158_,
		_w28162_,
		_w28172_
	);
	LUT3 #(
		.INIT('h15)
	) name22346 (
		_w28171_,
		_w28165_,
		_w28172_,
		_w28173_
	);
	LUT3 #(
		.INIT('hb0)
	) name22347 (
		_w28169_,
		_w28173_,
		_w28164_,
		_w28174_
	);
	LUT4 #(
		.INIT('h0052)
	) name22348 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28175_
	);
	LUT2 #(
		.INIT('h2)
	) name22349 (
		_w28159_,
		_w28162_,
		_w28176_
	);
	LUT4 #(
		.INIT('h0002)
	) name22350 (
		_w28159_,
		_w28161_,
		_w28158_,
		_w28162_,
		_w28177_
	);
	LUT4 #(
		.INIT('h2000)
	) name22351 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28178_
	);
	LUT4 #(
		.INIT('h5554)
	) name22352 (
		_w28164_,
		_w28175_,
		_w28177_,
		_w28178_,
		_w28179_
	);
	LUT4 #(
		.INIT('h0800)
	) name22353 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28180_
	);
	LUT4 #(
		.INIT('h0100)
	) name22354 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28181_
	);
	LUT4 #(
		.INIT('hfe3f)
	) name22355 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28182_
	);
	LUT4 #(
		.INIT('h20aa)
	) name22356 (
		_w28158_,
		_w28164_,
		_w28180_,
		_w28182_,
		_w28183_
	);
	LUT2 #(
		.INIT('h1)
	) name22357 (
		_w28179_,
		_w28183_,
		_w28184_
	);
	LUT4 #(
		.INIT('h5655)
	) name22358 (
		\u0_L8_reg[2]/NET0131 ,
		_w28174_,
		_w28167_,
		_w28184_,
		_w28185_
	);
	LUT4 #(
		.INIT('hd97b)
	) name22359 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28186_
	);
	LUT2 #(
		.INIT('h2)
	) name22360 (
		_w28031_,
		_w28186_,
		_w28187_
	);
	LUT4 #(
		.INIT('heebf)
	) name22361 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28188_
	);
	LUT4 #(
		.INIT('h0302)
	) name22362 (
		_w28031_,
		_w28036_,
		_w28040_,
		_w28188_,
		_w28189_
	);
	LUT3 #(
		.INIT('h45)
	) name22363 (
		_w28030_,
		_w28187_,
		_w28189_,
		_w28190_
	);
	LUT3 #(
		.INIT('h10)
	) name22364 (
		_w28034_,
		_w28035_,
		_w28033_,
		_w28191_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name22365 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28192_
	);
	LUT4 #(
		.INIT('h0080)
	) name22366 (
		_w28032_,
		_w28034_,
		_w28031_,
		_w28035_,
		_w28193_
	);
	LUT4 #(
		.INIT('hc100)
	) name22367 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28194_
	);
	LUT4 #(
		.INIT('h0032)
	) name22368 (
		_w28031_,
		_w28193_,
		_w28192_,
		_w28194_,
		_w28195_
	);
	LUT4 #(
		.INIT('h70d0)
	) name22369 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28196_
	);
	LUT4 #(
		.INIT('h0f01)
	) name22370 (
		_w28032_,
		_w28034_,
		_w28031_,
		_w28035_,
		_w28197_
	);
	LUT3 #(
		.INIT('hbe)
	) name22371 (
		_w28032_,
		_w28034_,
		_w28033_,
		_w28198_
	);
	LUT3 #(
		.INIT('h9e)
	) name22372 (
		_w28032_,
		_w28034_,
		_w28033_,
		_w28199_
	);
	LUT2 #(
		.INIT('h8)
	) name22373 (
		_w28031_,
		_w28035_,
		_w28200_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name22374 (
		_w28196_,
		_w28197_,
		_w28199_,
		_w28200_,
		_w28201_
	);
	LUT3 #(
		.INIT('hd0)
	) name22375 (
		_w28030_,
		_w28195_,
		_w28201_,
		_w28202_
	);
	LUT3 #(
		.INIT('h65)
	) name22376 (
		\u0_L8_reg[4]/NET0131 ,
		_w28190_,
		_w28202_,
		_w28203_
	);
	LUT4 #(
		.INIT('hc693)
	) name22377 (
		decrypt_pad,
		\u0_R8_reg[32]/NET0131 ,
		\u0_uk_K_r8_reg[29]/NET0131 ,
		\u0_uk_K_r8_reg[9]/P0001 ,
		_w28204_
	);
	LUT4 #(
		.INIT('hc963)
	) name22378 (
		decrypt_pad,
		\u0_R8_reg[1]/NET0131 ,
		\u0_uk_K_r8_reg[30]/NET0131 ,
		\u0_uk_K_r8_reg[50]/NET0131 ,
		_w28205_
	);
	LUT4 #(
		.INIT('hc963)
	) name22379 (
		decrypt_pad,
		\u0_R8_reg[30]/NET0131 ,
		\u0_uk_K_r8_reg[15]/NET0131 ,
		\u0_uk_K_r8_reg[35]/NET0131 ,
		_w28206_
	);
	LUT4 #(
		.INIT('hc963)
	) name22380 (
		decrypt_pad,
		\u0_R8_reg[29]/NET0131 ,
		\u0_uk_K_r8_reg[14]/NET0131 ,
		\u0_uk_K_r8_reg[38]/NET0131 ,
		_w28207_
	);
	LUT4 #(
		.INIT('hc963)
	) name22381 (
		decrypt_pad,
		\u0_R8_reg[28]/NET0131 ,
		\u0_uk_K_r8_reg[42]/NET0131 ,
		\u0_uk_K_r8_reg[7]/NET0131 ,
		_w28208_
	);
	LUT4 #(
		.INIT('hfcdf)
	) name22382 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28209_
	);
	LUT4 #(
		.INIT('hc693)
	) name22383 (
		decrypt_pad,
		\u0_R8_reg[31]/P0001 ,
		\u0_uk_K_r8_reg[23]/NET0131 ,
		\u0_uk_K_r8_reg[31]/NET0131 ,
		_w28210_
	);
	LUT2 #(
		.INIT('h4)
	) name22384 (
		_w28209_,
		_w28210_,
		_w28211_
	);
	LUT3 #(
		.INIT('h0d)
	) name22385 (
		_w28206_,
		_w28208_,
		_w28205_,
		_w28212_
	);
	LUT3 #(
		.INIT('h0b)
	) name22386 (
		_w28207_,
		_w28205_,
		_w28210_,
		_w28213_
	);
	LUT2 #(
		.INIT('h4)
	) name22387 (
		_w28212_,
		_w28213_,
		_w28214_
	);
	LUT4 #(
		.INIT('h8000)
	) name22388 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28215_
	);
	LUT3 #(
		.INIT('h04)
	) name22389 (
		_w28206_,
		_w28208_,
		_w28210_,
		_w28216_
	);
	LUT4 #(
		.INIT('h0040)
	) name22390 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28217_
	);
	LUT3 #(
		.INIT('h01)
	) name22391 (
		_w28215_,
		_w28216_,
		_w28217_,
		_w28218_
	);
	LUT4 #(
		.INIT('h5455)
	) name22392 (
		_w28204_,
		_w28211_,
		_w28214_,
		_w28218_,
		_w28219_
	);
	LUT4 #(
		.INIT('h0200)
	) name22393 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28220_
	);
	LUT4 #(
		.INIT('h0001)
	) name22394 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28221_
	);
	LUT4 #(
		.INIT('haf23)
	) name22395 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28222_
	);
	LUT4 #(
		.INIT('h1008)
	) name22396 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28223_
	);
	LUT4 #(
		.INIT('hedf6)
	) name22397 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28224_
	);
	LUT2 #(
		.INIT('h2)
	) name22398 (
		_w28210_,
		_w28224_,
		_w28225_
	);
	LUT3 #(
		.INIT('h02)
	) name22399 (
		_w28210_,
		_w28217_,
		_w28222_,
		_w28226_
	);
	LUT4 #(
		.INIT('h0800)
	) name22400 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28227_
	);
	LUT4 #(
		.INIT('h0001)
	) name22401 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28210_,
		_w28228_
	);
	LUT2 #(
		.INIT('h1)
	) name22402 (
		_w28227_,
		_w28228_,
		_w28229_
	);
	LUT3 #(
		.INIT('h20)
	) name22403 (
		_w28204_,
		_w28207_,
		_w28208_,
		_w28230_
	);
	LUT4 #(
		.INIT('hcdcf)
	) name22404 (
		_w28206_,
		_w28210_,
		_w28217_,
		_w28230_,
		_w28231_
	);
	LUT4 #(
		.INIT('h7500)
	) name22405 (
		_w28204_,
		_w28226_,
		_w28229_,
		_w28231_,
		_w28232_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name22406 (
		\u0_L8_reg[5]/NET0131 ,
		_w28219_,
		_w28225_,
		_w28232_,
		_w28233_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name22407 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28234_
	);
	LUT4 #(
		.INIT('h0200)
	) name22408 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28235_
	);
	LUT4 #(
		.INIT('hedeb)
	) name22409 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28236_
	);
	LUT4 #(
		.INIT('h0515)
	) name22410 (
		_w28158_,
		_w28164_,
		_w28234_,
		_w28236_,
		_w28237_
	);
	LUT4 #(
		.INIT('hf6b6)
	) name22411 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28238_
	);
	LUT2 #(
		.INIT('h2)
	) name22412 (
		_w28158_,
		_w28238_,
		_w28239_
	);
	LUT2 #(
		.INIT('h8)
	) name22413 (
		_w28170_,
		_w28176_,
		_w28240_
	);
	LUT2 #(
		.INIT('h8)
	) name22414 (
		_w28160_,
		_w28158_,
		_w28241_
	);
	LUT3 #(
		.INIT('hb0)
	) name22415 (
		_w28159_,
		_w28161_,
		_w28162_,
		_w28242_
	);
	LUT3 #(
		.INIT('h15)
	) name22416 (
		_w28164_,
		_w28241_,
		_w28242_,
		_w28243_
	);
	LUT3 #(
		.INIT('h10)
	) name22417 (
		_w28239_,
		_w28240_,
		_w28243_,
		_w28244_
	);
	LUT3 #(
		.INIT('h01)
	) name22418 (
		_w28159_,
		_w28161_,
		_w28162_,
		_w28245_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name22419 (
		_w28159_,
		_w28160_,
		_w28158_,
		_w28162_,
		_w28246_
	);
	LUT3 #(
		.INIT('h08)
	) name22420 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28247_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name22421 (
		_w28159_,
		_w28161_,
		_w28158_,
		_w28162_,
		_w28248_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name22422 (
		_w28245_,
		_w28246_,
		_w28247_,
		_w28248_,
		_w28249_
	);
	LUT4 #(
		.INIT('h0010)
	) name22423 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28250_
	);
	LUT4 #(
		.INIT('h0002)
	) name22424 (
		_w28164_,
		_w28177_,
		_w28178_,
		_w28250_,
		_w28251_
	);
	LUT3 #(
		.INIT('h20)
	) name22425 (
		_w28234_,
		_w28249_,
		_w28251_,
		_w28252_
	);
	LUT4 #(
		.INIT('h999a)
	) name22426 (
		\u0_L8_reg[13]/NET0131 ,
		_w28237_,
		_w28244_,
		_w28252_,
		_w28253_
	);
	LUT4 #(
		.INIT('hc963)
	) name22427 (
		decrypt_pad,
		\u0_R8_reg[18]/NET0131 ,
		\u0_uk_K_r8_reg[23]/NET0131 ,
		\u0_uk_K_r8_reg[43]/NET0131 ,
		_w28254_
	);
	LUT4 #(
		.INIT('hc693)
	) name22428 (
		decrypt_pad,
		\u0_R8_reg[19]/NET0131 ,
		\u0_uk_K_r8_reg[30]/NET0131 ,
		\u0_uk_K_r8_reg[38]/NET0131 ,
		_w28255_
	);
	LUT2 #(
		.INIT('h1)
	) name22429 (
		_w28254_,
		_w28255_,
		_w28256_
	);
	LUT4 #(
		.INIT('hc963)
	) name22430 (
		decrypt_pad,
		\u0_R8_reg[17]/NET0131 ,
		\u0_uk_K_r8_reg[29]/NET0131 ,
		\u0_uk_K_r8_reg[49]/NET0131 ,
		_w28257_
	);
	LUT4 #(
		.INIT('hc693)
	) name22431 (
		decrypt_pad,
		\u0_R8_reg[21]/NET0131 ,
		\u0_uk_K_r8_reg[15]/NET0131 ,
		\u0_uk_K_r8_reg[50]/NET0131 ,
		_w28258_
	);
	LUT4 #(
		.INIT('hc693)
	) name22432 (
		decrypt_pad,
		\u0_R8_reg[16]/NET0131 ,
		\u0_uk_K_r8_reg[31]/NET0131 ,
		\u0_uk_K_r8_reg[7]/NET0131 ,
		_w28259_
	);
	LUT3 #(
		.INIT('hf6)
	) name22433 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28260_
	);
	LUT2 #(
		.INIT('h2)
	) name22434 (
		_w28256_,
		_w28260_,
		_w28261_
	);
	LUT4 #(
		.INIT('h0040)
	) name22435 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28262_
	);
	LUT3 #(
		.INIT('ha2)
	) name22436 (
		_w28257_,
		_w28254_,
		_w28255_,
		_w28263_
	);
	LUT4 #(
		.INIT('h80a0)
	) name22437 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28264_
	);
	LUT3 #(
		.INIT('h45)
	) name22438 (
		_w28262_,
		_w28263_,
		_w28264_,
		_w28265_
	);
	LUT3 #(
		.INIT('h02)
	) name22439 (
		_w28257_,
		_w28259_,
		_w28254_,
		_w28266_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name22440 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28267_
	);
	LUT4 #(
		.INIT('hea00)
	) name22441 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28255_,
		_w28268_
	);
	LUT4 #(
		.INIT('h1000)
	) name22442 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28269_
	);
	LUT4 #(
		.INIT('hc693)
	) name22443 (
		decrypt_pad,
		\u0_R8_reg[20]/NET0131 ,
		\u0_uk_K_r8_reg[14]/NET0131 ,
		\u0_uk_K_r8_reg[49]/NET0131 ,
		_w28270_
	);
	LUT4 #(
		.INIT('h0700)
	) name22444 (
		_w28267_,
		_w28268_,
		_w28269_,
		_w28270_,
		_w28271_
	);
	LUT3 #(
		.INIT('h40)
	) name22445 (
		_w28261_,
		_w28265_,
		_w28271_,
		_w28272_
	);
	LUT3 #(
		.INIT('h02)
	) name22446 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28273_
	);
	LUT4 #(
		.INIT('h00bf)
	) name22447 (
		_w28258_,
		_w28257_,
		_w28254_,
		_w28255_,
		_w28274_
	);
	LUT4 #(
		.INIT('h0080)
	) name22448 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28275_
	);
	LUT4 #(
		.INIT('h0010)
	) name22449 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28276_
	);
	LUT4 #(
		.INIT('hff6f)
	) name22450 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28277_
	);
	LUT3 #(
		.INIT('h40)
	) name22451 (
		_w28273_,
		_w28274_,
		_w28277_,
		_w28278_
	);
	LUT4 #(
		.INIT('hfe00)
	) name22452 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28255_,
		_w28279_
	);
	LUT2 #(
		.INIT('h8)
	) name22453 (
		_w28267_,
		_w28279_,
		_w28280_
	);
	LUT4 #(
		.INIT('h0004)
	) name22454 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28281_
	);
	LUT4 #(
		.INIT('h2000)
	) name22455 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28282_
	);
	LUT3 #(
		.INIT('h01)
	) name22456 (
		_w28270_,
		_w28282_,
		_w28281_,
		_w28283_
	);
	LUT3 #(
		.INIT('he0)
	) name22457 (
		_w28278_,
		_w28280_,
		_w28283_,
		_w28284_
	);
	LUT4 #(
		.INIT('hfebf)
	) name22458 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28285_
	);
	LUT4 #(
		.INIT('h0200)
	) name22459 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28286_
	);
	LUT4 #(
		.INIT('hf9ff)
	) name22460 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28287_
	);
	LUT3 #(
		.INIT('hd8)
	) name22461 (
		_w28255_,
		_w28285_,
		_w28287_,
		_w28288_
	);
	LUT4 #(
		.INIT('ha955)
	) name22462 (
		\u0_L8_reg[14]/NET0131 ,
		_w28272_,
		_w28284_,
		_w28288_,
		_w28289_
	);
	LUT4 #(
		.INIT('heffa)
	) name22463 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28290_
	);
	LUT4 #(
		.INIT('hdf8f)
	) name22464 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28291_
	);
	LUT4 #(
		.INIT('h7fb7)
	) name22465 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28292_
	);
	LUT4 #(
		.INIT('hd800)
	) name22466 (
		_w28108_,
		_w28290_,
		_w28291_,
		_w28292_,
		_w28293_
	);
	LUT2 #(
		.INIT('h1)
	) name22467 (
		_w28113_,
		_w28293_,
		_w28294_
	);
	LUT4 #(
		.INIT('hf773)
	) name22468 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28295_
	);
	LUT4 #(
		.INIT('h4000)
	) name22469 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28296_
	);
	LUT4 #(
		.INIT('hbcff)
	) name22470 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28297_
	);
	LUT4 #(
		.INIT('h04cc)
	) name22471 (
		_w28108_,
		_w28113_,
		_w28295_,
		_w28297_,
		_w28298_
	);
	LUT4 #(
		.INIT('h7dff)
	) name22472 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28299_
	);
	LUT4 #(
		.INIT('h79ff)
	) name22473 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28300_
	);
	LUT2 #(
		.INIT('h2)
	) name22474 (
		_w28108_,
		_w28300_,
		_w28301_
	);
	LUT2 #(
		.INIT('h4)
	) name22475 (
		_w28108_,
		_w28296_,
		_w28302_
	);
	LUT4 #(
		.INIT('hddcd)
	) name22476 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28303_
	);
	LUT2 #(
		.INIT('h8)
	) name22477 (
		_w28108_,
		_w28113_,
		_w28304_
	);
	LUT4 #(
		.INIT('h7077)
	) name22478 (
		_w28114_,
		_w28123_,
		_w28303_,
		_w28304_,
		_w28305_
	);
	LUT4 #(
		.INIT('h0100)
	) name22479 (
		_w28301_,
		_w28302_,
		_w28298_,
		_w28305_,
		_w28306_
	);
	LUT3 #(
		.INIT('h65)
	) name22480 (
		\u0_L8_reg[1]/NET0131 ,
		_w28294_,
		_w28306_,
		_w28307_
	);
	LUT4 #(
		.INIT('hafe7)
	) name22481 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28308_
	);
	LUT4 #(
		.INIT('hfbdb)
	) name22482 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28309_
	);
	LUT4 #(
		.INIT('hc480)
	) name22483 (
		_w28108_,
		_w28299_,
		_w28309_,
		_w28308_,
		_w28310_
	);
	LUT2 #(
		.INIT('h2)
	) name22484 (
		_w28113_,
		_w28310_,
		_w28311_
	);
	LUT4 #(
		.INIT('hc2f1)
	) name22485 (
		_w28109_,
		_w28107_,
		_w28114_,
		_w28108_,
		_w28312_
	);
	LUT2 #(
		.INIT('h2)
	) name22486 (
		_w28110_,
		_w28312_,
		_w28313_
	);
	LUT4 #(
		.INIT('h0200)
	) name22487 (
		_w28109_,
		_w28110_,
		_w28114_,
		_w28108_,
		_w28314_
	);
	LUT3 #(
		.INIT('h04)
	) name22488 (
		_w28123_,
		_w28133_,
		_w28314_,
		_w28315_
	);
	LUT3 #(
		.INIT('h45)
	) name22489 (
		_w28113_,
		_w28313_,
		_w28315_,
		_w28316_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name22490 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28317_
	);
	LUT2 #(
		.INIT('h1)
	) name22491 (
		_w28108_,
		_w28317_,
		_w28318_
	);
	LUT3 #(
		.INIT('h0b)
	) name22492 (
		_w28114_,
		_w28119_,
		_w28130_,
		_w28319_
	);
	LUT2 #(
		.INIT('h4)
	) name22493 (
		_w28318_,
		_w28319_,
		_w28320_
	);
	LUT4 #(
		.INIT('h5655)
	) name22494 (
		\u0_L8_reg[10]/NET0131 ,
		_w28316_,
		_w28311_,
		_w28320_,
		_w28321_
	);
	LUT3 #(
		.INIT('hb0)
	) name22495 (
		_w28064_,
		_w28067_,
		_w28063_,
		_w28322_
	);
	LUT3 #(
		.INIT('h10)
	) name22496 (
		_w28086_,
		_w28082_,
		_w28322_,
		_w28323_
	);
	LUT4 #(
		.INIT('h0400)
	) name22497 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28324_
	);
	LUT4 #(
		.INIT('h1248)
	) name22498 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28325_
	);
	LUT4 #(
		.INIT('h080c)
	) name22499 (
		_w28063_,
		_w28062_,
		_w28325_,
		_w28324_,
		_w28326_
	);
	LUT2 #(
		.INIT('h4)
	) name22500 (
		_w28323_,
		_w28326_,
		_w28327_
	);
	LUT2 #(
		.INIT('h4)
	) name22501 (
		_w28064_,
		_w28066_,
		_w28328_
	);
	LUT4 #(
		.INIT('h0814)
	) name22502 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28329_
	);
	LUT4 #(
		.INIT('h0770)
	) name22503 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28330_
	);
	LUT2 #(
		.INIT('h1)
	) name22504 (
		_w28063_,
		_w28330_,
		_w28331_
	);
	LUT3 #(
		.INIT('h53)
	) name22505 (
		_w28067_,
		_w28063_,
		_w28065_,
		_w28332_
	);
	LUT4 #(
		.INIT('h0002)
	) name22506 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28333_
	);
	LUT4 #(
		.INIT('h0051)
	) name22507 (
		_w28062_,
		_w28328_,
		_w28332_,
		_w28333_,
		_w28334_
	);
	LUT3 #(
		.INIT('h10)
	) name22508 (
		_w28331_,
		_w28329_,
		_w28334_,
		_w28335_
	);
	LUT3 #(
		.INIT('ha9)
	) name22509 (
		\u0_L8_reg[12]/NET0131 ,
		_w28327_,
		_w28335_,
		_w28336_
	);
	LUT4 #(
		.INIT('h0100)
	) name22510 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28210_,
		_w28337_
	);
	LUT2 #(
		.INIT('h1)
	) name22511 (
		_w28204_,
		_w28337_,
		_w28338_
	);
	LUT4 #(
		.INIT('hf2fe)
	) name22512 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28339_
	);
	LUT3 #(
		.INIT('h80)
	) name22513 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28340_
	);
	LUT4 #(
		.INIT('hef00)
	) name22514 (
		_w28206_,
		_w28207_,
		_w28205_,
		_w28210_,
		_w28341_
	);
	LUT3 #(
		.INIT('h40)
	) name22515 (
		_w28340_,
		_w28339_,
		_w28341_,
		_w28342_
	);
	LUT4 #(
		.INIT('h2000)
	) name22516 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28343_
	);
	LUT4 #(
		.INIT('h00fb)
	) name22517 (
		_w28206_,
		_w28208_,
		_w28205_,
		_w28210_,
		_w28344_
	);
	LUT2 #(
		.INIT('h4)
	) name22518 (
		_w28343_,
		_w28344_,
		_w28345_
	);
	LUT4 #(
		.INIT('h0100)
	) name22519 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28346_
	);
	LUT4 #(
		.INIT('hfe7d)
	) name22520 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28347_
	);
	LUT4 #(
		.INIT('h0155)
	) name22521 (
		_w28338_,
		_w28342_,
		_w28345_,
		_w28347_,
		_w28348_
	);
	LUT4 #(
		.INIT('h0040)
	) name22522 (
		_w28206_,
		_w28208_,
		_w28205_,
		_w28210_,
		_w28349_
	);
	LUT2 #(
		.INIT('h8)
	) name22523 (
		_w28207_,
		_w28349_,
		_w28350_
	);
	LUT4 #(
		.INIT('hffde)
	) name22524 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28351_
	);
	LUT2 #(
		.INIT('h4)
	) name22525 (
		_w28349_,
		_w28351_,
		_w28352_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name22526 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28353_
	);
	LUT2 #(
		.INIT('h2)
	) name22527 (
		_w28210_,
		_w28353_,
		_w28354_
	);
	LUT4 #(
		.INIT('hb7f7)
	) name22528 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28355_
	);
	LUT4 #(
		.INIT('h0020)
	) name22529 (
		_w28206_,
		_w28208_,
		_w28205_,
		_w28210_,
		_w28356_
	);
	LUT4 #(
		.INIT('h0002)
	) name22530 (
		_w28207_,
		_w28208_,
		_w28205_,
		_w28210_,
		_w28357_
	);
	LUT3 #(
		.INIT('h10)
	) name22531 (
		_w28356_,
		_w28357_,
		_w28355_,
		_w28358_
	);
	LUT4 #(
		.INIT('h4555)
	) name22532 (
		_w28204_,
		_w28354_,
		_w28358_,
		_w28352_,
		_w28359_
	);
	LUT4 #(
		.INIT('h5556)
	) name22533 (
		\u0_L8_reg[21]/NET0131 ,
		_w28348_,
		_w28350_,
		_w28359_,
		_w28360_
	);
	LUT4 #(
		.INIT('h3c3b)
	) name22534 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28361_
	);
	LUT4 #(
		.INIT('h0010)
	) name22535 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28362_
	);
	LUT4 #(
		.INIT('h5504)
	) name22536 (
		_w28204_,
		_w28210_,
		_w28361_,
		_w28362_,
		_w28363_
	);
	LUT4 #(
		.INIT('h0020)
	) name22537 (
		_w28206_,
		_w28207_,
		_w28205_,
		_w28210_,
		_w28364_
	);
	LUT4 #(
		.INIT('hbfb7)
	) name22538 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28365_
	);
	LUT4 #(
		.INIT('h0100)
	) name22539 (
		_w28207_,
		_w28208_,
		_w28205_,
		_w28210_,
		_w28366_
	);
	LUT4 #(
		.INIT('h0100)
	) name22540 (
		_w28343_,
		_w28366_,
		_w28364_,
		_w28365_,
		_w28367_
	);
	LUT3 #(
		.INIT('h10)
	) name22541 (
		_w28204_,
		_w28207_,
		_w28208_,
		_w28368_
	);
	LUT4 #(
		.INIT('hfbf7)
	) name22542 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28369_
	);
	LUT4 #(
		.INIT('h00df)
	) name22543 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28210_,
		_w28370_
	);
	LUT4 #(
		.INIT('h1000)
	) name22544 (
		_w28221_,
		_w28368_,
		_w28370_,
		_w28369_,
		_w28371_
	);
	LUT3 #(
		.INIT('h02)
	) name22545 (
		_w28210_,
		_w28227_,
		_w28346_,
		_w28372_
	);
	LUT4 #(
		.INIT('hddd0)
	) name22546 (
		_w28204_,
		_w28367_,
		_w28371_,
		_w28372_,
		_w28373_
	);
	LUT3 #(
		.INIT('h65)
	) name22547 (
		\u0_L8_reg[15]/P0001 ,
		_w28363_,
		_w28373_,
		_w28374_
	);
	LUT4 #(
		.INIT('h4e55)
	) name22548 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28375_
	);
	LUT4 #(
		.INIT('h8000)
	) name22549 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28376_
	);
	LUT4 #(
		.INIT('h0e04)
	) name22550 (
		_w28031_,
		_w28198_,
		_w28376_,
		_w28375_,
		_w28377_
	);
	LUT2 #(
		.INIT('h1)
	) name22551 (
		_w28030_,
		_w28377_,
		_w28378_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name22552 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28379_
	);
	LUT2 #(
		.INIT('h2)
	) name22553 (
		_w28031_,
		_w28379_,
		_w28380_
	);
	LUT4 #(
		.INIT('h4010)
	) name22554 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28381_
	);
	LUT4 #(
		.INIT('h0004)
	) name22555 (
		_w28032_,
		_w28034_,
		_w28035_,
		_w28033_,
		_w28382_
	);
	LUT3 #(
		.INIT('h02)
	) name22556 (
		_w28032_,
		_w28031_,
		_w28033_,
		_w28383_
	);
	LUT4 #(
		.INIT('h0001)
	) name22557 (
		_w28191_,
		_w28381_,
		_w28382_,
		_w28383_,
		_w28384_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name22558 (
		_w28035_,
		_w28033_,
		_w28052_,
		_w28040_,
		_w28385_
	);
	LUT4 #(
		.INIT('h7500)
	) name22559 (
		_w28030_,
		_w28380_,
		_w28384_,
		_w28385_,
		_w28386_
	);
	LUT3 #(
		.INIT('h65)
	) name22560 (
		\u0_L8_reg[19]/NET0131 ,
		_w28378_,
		_w28386_,
		_w28387_
	);
	LUT4 #(
		.INIT('hfbef)
	) name22561 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28388_
	);
	LUT4 #(
		.INIT('h0288)
	) name22562 (
		_w28002_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28389_
	);
	LUT4 #(
		.INIT('h0032)
	) name22563 (
		_w28002_,
		_w28020_,
		_w28388_,
		_w28389_,
		_w28390_
	);
	LUT2 #(
		.INIT('h1)
	) name22564 (
		_w28014_,
		_w28390_,
		_w28391_
	);
	LUT4 #(
		.INIT('h3800)
	) name22565 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28392_
	);
	LUT3 #(
		.INIT('h14)
	) name22566 (
		_w27999_,
		_w28000_,
		_w28005_,
		_w28393_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name22567 (
		_w28002_,
		_w28016_,
		_w28392_,
		_w28393_,
		_w28394_
	);
	LUT4 #(
		.INIT('h002a)
	) name22568 (
		_w27998_,
		_w28001_,
		_w28026_,
		_w28096_,
		_w28395_
	);
	LUT4 #(
		.INIT('h1554)
	) name22569 (
		_w27998_,
		_w28003_,
		_w28000_,
		_w28005_,
		_w28396_
	);
	LUT4 #(
		.INIT('h4440)
	) name22570 (
		_w28002_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28397_
	);
	LUT2 #(
		.INIT('h2)
	) name22571 (
		_w28002_,
		_w27999_,
		_w28398_
	);
	LUT4 #(
		.INIT('h8caf)
	) name22572 (
		_w28024_,
		_w28021_,
		_w28397_,
		_w28398_,
		_w28399_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name22573 (
		_w28394_,
		_w28395_,
		_w28396_,
		_w28399_,
		_w28400_
	);
	LUT3 #(
		.INIT('ha9)
	) name22574 (
		\u0_L8_reg[23]/NET0131 ,
		_w28391_,
		_w28400_,
		_w28401_
	);
	LUT4 #(
		.INIT('hecee)
	) name22575 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28402_
	);
	LUT4 #(
		.INIT('h0094)
	) name22576 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28403_
	);
	LUT4 #(
		.INIT('h0504)
	) name22577 (
		_w28108_,
		_w28113_,
		_w28403_,
		_w28402_,
		_w28404_
	);
	LUT3 #(
		.INIT('h02)
	) name22578 (
		_w28108_,
		_w28121_,
		_w28131_,
		_w28405_
	);
	LUT2 #(
		.INIT('h1)
	) name22579 (
		_w28404_,
		_w28405_,
		_w28406_
	);
	LUT4 #(
		.INIT('h4004)
	) name22580 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28407_
	);
	LUT3 #(
		.INIT('h02)
	) name22581 (
		_w28113_,
		_w28126_,
		_w28407_,
		_w28408_
	);
	LUT4 #(
		.INIT('h5ffd)
	) name22582 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28114_,
		_w28409_
	);
	LUT4 #(
		.INIT('hf5f7)
	) name22583 (
		_w28109_,
		_w28107_,
		_w28110_,
		_w28108_,
		_w28410_
	);
	LUT4 #(
		.INIT('hfc54)
	) name22584 (
		_w28114_,
		_w28108_,
		_w28409_,
		_w28410_,
		_w28411_
	);
	LUT4 #(
		.INIT('h00fb)
	) name22585 (
		_w28107_,
		_w28110_,
		_w28114_,
		_w28113_,
		_w28412_
	);
	LUT3 #(
		.INIT('hb0)
	) name22586 (
		_w28111_,
		_w28129_,
		_w28412_,
		_w28413_
	);
	LUT4 #(
		.INIT('h153f)
	) name22587 (
		_w28122_,
		_w28408_,
		_w28411_,
		_w28413_,
		_w28414_
	);
	LUT3 #(
		.INIT('h56)
	) name22588 (
		\u0_L8_reg[26]/NET0131 ,
		_w28406_,
		_w28414_,
		_w28415_
	);
	LUT4 #(
		.INIT('h6b7b)
	) name22589 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28416_
	);
	LUT2 #(
		.INIT('h2)
	) name22590 (
		_w28158_,
		_w28416_,
		_w28417_
	);
	LUT4 #(
		.INIT('hdfce)
	) name22591 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28418_
	);
	LUT2 #(
		.INIT('h1)
	) name22592 (
		_w28158_,
		_w28418_,
		_w28419_
	);
	LUT4 #(
		.INIT('h33f7)
	) name22593 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28158_,
		_w28420_
	);
	LUT3 #(
		.INIT('h32)
	) name22594 (
		_w28162_,
		_w28235_,
		_w28420_,
		_w28421_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name22595 (
		_w28164_,
		_w28419_,
		_w28417_,
		_w28421_,
		_w28422_
	);
	LUT4 #(
		.INIT('h3d39)
	) name22596 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28423_
	);
	LUT4 #(
		.INIT('hb6ff)
	) name22597 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28424_
	);
	LUT4 #(
		.INIT('hd800)
	) name22598 (
		_w28158_,
		_w28418_,
		_w28423_,
		_w28424_,
		_w28425_
	);
	LUT4 #(
		.INIT('hbcff)
	) name22599 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28426_
	);
	LUT2 #(
		.INIT('h1)
	) name22600 (
		_w28158_,
		_w28426_,
		_w28427_
	);
	LUT3 #(
		.INIT('h0e)
	) name22601 (
		_w28164_,
		_w28425_,
		_w28427_,
		_w28428_
	);
	LUT3 #(
		.INIT('h65)
	) name22602 (
		\u0_L8_reg[28]/NET0131 ,
		_w28422_,
		_w28428_,
		_w28429_
	);
	LUT4 #(
		.INIT('h7f6f)
	) name22603 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28430_
	);
	LUT2 #(
		.INIT('h2)
	) name22604 (
		_w28255_,
		_w28430_,
		_w28431_
	);
	LUT4 #(
		.INIT('hbeff)
	) name22605 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28432_
	);
	LUT3 #(
		.INIT('h20)
	) name22606 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28433_
	);
	LUT4 #(
		.INIT('hd7d5)
	) name22607 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28434_
	);
	LUT4 #(
		.INIT('h3200)
	) name22608 (
		_w28255_,
		_w28266_,
		_w28434_,
		_w28432_,
		_w28435_
	);
	LUT3 #(
		.INIT('h45)
	) name22609 (
		_w28270_,
		_w28431_,
		_w28435_,
		_w28436_
	);
	LUT4 #(
		.INIT('h0001)
	) name22610 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28437_
	);
	LUT4 #(
		.INIT('hdfde)
	) name22611 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28438_
	);
	LUT3 #(
		.INIT('h02)
	) name22612 (
		_w28259_,
		_w28254_,
		_w28255_,
		_w28439_
	);
	LUT4 #(
		.INIT('h00c4)
	) name22613 (
		_w28255_,
		_w28287_,
		_w28438_,
		_w28439_,
		_w28440_
	);
	LUT4 #(
		.INIT('hb9f7)
	) name22614 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28441_
	);
	LUT3 #(
		.INIT('hb1)
	) name22615 (
		_w28255_,
		_w28269_,
		_w28441_,
		_w28442_
	);
	LUT3 #(
		.INIT('hd0)
	) name22616 (
		_w28270_,
		_w28440_,
		_w28442_,
		_w28443_
	);
	LUT3 #(
		.INIT('h65)
	) name22617 (
		\u0_L8_reg[8]/NET0131 ,
		_w28436_,
		_w28443_,
		_w28444_
	);
	LUT4 #(
		.INIT('hf23e)
	) name22618 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28445_
	);
	LUT4 #(
		.INIT('h3ffb)
	) name22619 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28446_
	);
	LUT4 #(
		.INIT('he6df)
	) name22620 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28205_,
		_w28447_
	);
	LUT4 #(
		.INIT('hd800)
	) name22621 (
		_w28210_,
		_w28446_,
		_w28445_,
		_w28447_,
		_w28448_
	);
	LUT2 #(
		.INIT('h2)
	) name22622 (
		_w28204_,
		_w28448_,
		_w28449_
	);
	LUT4 #(
		.INIT('hf700)
	) name22623 (
		_w28206_,
		_w28207_,
		_w28208_,
		_w28210_,
		_w28450_
	);
	LUT3 #(
		.INIT('h4b)
	) name22624 (
		_w28206_,
		_w28207_,
		_w28205_,
		_w28451_
	);
	LUT2 #(
		.INIT('h8)
	) name22625 (
		_w28450_,
		_w28451_,
		_w28452_
	);
	LUT4 #(
		.INIT('h0080)
	) name22626 (
		_w28206_,
		_w28208_,
		_w28205_,
		_w28210_,
		_w28453_
	);
	LUT3 #(
		.INIT('h01)
	) name22627 (
		_w28220_,
		_w28357_,
		_w28453_,
		_w28454_
	);
	LUT4 #(
		.INIT('h0200)
	) name22628 (
		_w28206_,
		_w28207_,
		_w28205_,
		_w28210_,
		_w28455_
	);
	LUT4 #(
		.INIT('h00ab)
	) name22629 (
		_w28210_,
		_w28217_,
		_w28223_,
		_w28455_,
		_w28456_
	);
	LUT4 #(
		.INIT('hba00)
	) name22630 (
		_w28204_,
		_w28452_,
		_w28454_,
		_w28456_,
		_w28457_
	);
	LUT3 #(
		.INIT('h65)
	) name22631 (
		\u0_L8_reg[27]/NET0131 ,
		_w28449_,
		_w28457_,
		_w28458_
	);
	LUT4 #(
		.INIT('h0102)
	) name22632 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28459_
	);
	LUT3 #(
		.INIT('h04)
	) name22633 (
		_w28064_,
		_w28065_,
		_w28066_,
		_w28460_
	);
	LUT4 #(
		.INIT('h0800)
	) name22634 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28461_
	);
	LUT4 #(
		.INIT('h0001)
	) name22635 (
		_w28063_,
		_w28459_,
		_w28461_,
		_w28460_,
		_w28462_
	);
	LUT3 #(
		.INIT('h02)
	) name22636 (
		_w28064_,
		_w28067_,
		_w28066_,
		_w28463_
	);
	LUT4 #(
		.INIT('h308d)
	) name22637 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28464_
	);
	LUT3 #(
		.INIT('h02)
	) name22638 (
		_w28063_,
		_w28324_,
		_w28464_,
		_w28465_
	);
	LUT4 #(
		.INIT('h0080)
	) name22639 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28466_
	);
	LUT2 #(
		.INIT('h2)
	) name22640 (
		_w28062_,
		_w28466_,
		_w28467_
	);
	LUT3 #(
		.INIT('he0)
	) name22641 (
		_w28462_,
		_w28465_,
		_w28467_,
		_w28468_
	);
	LUT4 #(
		.INIT('h8020)
	) name22642 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28469_
	);
	LUT3 #(
		.INIT('h01)
	) name22643 (
		_w28062_,
		_w28087_,
		_w28469_,
		_w28470_
	);
	LUT3 #(
		.INIT('h20)
	) name22644 (
		_w28064_,
		_w28065_,
		_w28066_,
		_w28471_
	);
	LUT3 #(
		.INIT('h41)
	) name22645 (
		_w28063_,
		_w28065_,
		_w28066_,
		_w28472_
	);
	LUT4 #(
		.INIT('h4457)
	) name22646 (
		_w28063_,
		_w28463_,
		_w28471_,
		_w28472_,
		_w28473_
	);
	LUT2 #(
		.INIT('h8)
	) name22647 (
		_w28470_,
		_w28473_,
		_w28474_
	);
	LUT4 #(
		.INIT('h3010)
	) name22648 (
		_w28064_,
		_w28063_,
		_w28065_,
		_w28066_,
		_w28475_
	);
	LUT2 #(
		.INIT('h8)
	) name22649 (
		_w28073_,
		_w28475_,
		_w28476_
	);
	LUT4 #(
		.INIT('h55a9)
	) name22650 (
		\u0_L8_reg[32]/NET0131 ,
		_w28468_,
		_w28474_,
		_w28476_,
		_w28477_
	);
	LUT3 #(
		.INIT('hb0)
	) name22651 (
		_w28257_,
		_w28254_,
		_w28255_,
		_w28478_
	);
	LUT4 #(
		.INIT('h50da)
	) name22652 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28479_
	);
	LUT2 #(
		.INIT('h1)
	) name22653 (
		_w28478_,
		_w28479_,
		_w28480_
	);
	LUT4 #(
		.INIT('hbfb5)
	) name22654 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28481_
	);
	LUT3 #(
		.INIT('h31)
	) name22655 (
		_w28255_,
		_w28270_,
		_w28481_,
		_w28482_
	);
	LUT4 #(
		.INIT('hfb5b)
	) name22656 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w28483_
	);
	LUT2 #(
		.INIT('h2)
	) name22657 (
		_w28255_,
		_w28483_,
		_w28484_
	);
	LUT4 #(
		.INIT('h0008)
	) name22658 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28255_,
		_w28485_
	);
	LUT4 #(
		.INIT('h0004)
	) name22659 (
		_w28269_,
		_w28270_,
		_w28275_,
		_w28485_,
		_w28486_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name22660 (
		_w28480_,
		_w28482_,
		_w28484_,
		_w28486_,
		_w28487_
	);
	LUT4 #(
		.INIT('h0001)
	) name22661 (
		_w28262_,
		_w28255_,
		_w28282_,
		_w28437_,
		_w28488_
	);
	LUT3 #(
		.INIT('h02)
	) name22662 (
		_w28255_,
		_w28276_,
		_w28286_,
		_w28489_
	);
	LUT2 #(
		.INIT('h1)
	) name22663 (
		_w28488_,
		_w28489_,
		_w28490_
	);
	LUT3 #(
		.INIT('h56)
	) name22664 (
		\u0_L8_reg[3]/NET0131 ,
		_w28487_,
		_w28490_,
		_w28491_
	);
	LUT4 #(
		.INIT('hc963)
	) name22665 (
		decrypt_pad,
		\u0_R8_reg[11]/NET0131 ,
		\u0_uk_K_r8_reg[32]/NET0131 ,
		\u0_uk_K_r8_reg[54]/NET0131 ,
		_w28492_
	);
	LUT4 #(
		.INIT('hc693)
	) name22666 (
		decrypt_pad,
		\u0_R8_reg[12]/NET0131 ,
		\u0_uk_K_r8_reg[12]/NET0131 ,
		\u0_uk_K_r8_reg[47]/NET0131 ,
		_w28493_
	);
	LUT4 #(
		.INIT('hc693)
	) name22667 (
		decrypt_pad,
		\u0_R8_reg[13]/NET0131 ,
		\u0_uk_K_r8_reg[25]/NET0131 ,
		\u0_uk_K_r8_reg[3]/NET0131 ,
		_w28494_
	);
	LUT4 #(
		.INIT('hc693)
	) name22668 (
		decrypt_pad,
		\u0_R8_reg[9]/NET0131 ,
		\u0_uk_K_r8_reg[20]/NET0131 ,
		\u0_uk_K_r8_reg[55]/NET0131 ,
		_w28495_
	);
	LUT4 #(
		.INIT('hc963)
	) name22669 (
		decrypt_pad,
		\u0_R8_reg[8]/NET0131 ,
		\u0_uk_K_r8_reg[26]/NET0131 ,
		\u0_uk_K_r8_reg[48]/NET0131 ,
		_w28496_
	);
	LUT4 #(
		.INIT('hc693)
	) name22670 (
		decrypt_pad,
		\u0_R8_reg[10]/NET0131 ,
		\u0_uk_K_r8_reg[53]/NET0131 ,
		\u0_uk_K_r8_reg[6]/NET0131 ,
		_w28497_
	);
	LUT4 #(
		.INIT('h95b5)
	) name22671 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28498_
	);
	LUT2 #(
		.INIT('h1)
	) name22672 (
		_w28494_,
		_w28496_,
		_w28499_
	);
	LUT4 #(
		.INIT('h0001)
	) name22673 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28500_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name22674 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28501_
	);
	LUT4 #(
		.INIT('h08cc)
	) name22675 (
		_w28493_,
		_w28492_,
		_w28498_,
		_w28501_,
		_w28502_
	);
	LUT2 #(
		.INIT('h8)
	) name22676 (
		_w28494_,
		_w28496_,
		_w28503_
	);
	LUT2 #(
		.INIT('h6)
	) name22677 (
		_w28494_,
		_w28496_,
		_w28504_
	);
	LUT4 #(
		.INIT('h000d)
	) name22678 (
		_w28492_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28505_
	);
	LUT4 #(
		.INIT('h0020)
	) name22679 (
		_w28492_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28506_
	);
	LUT4 #(
		.INIT('h4000)
	) name22680 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28507_
	);
	LUT4 #(
		.INIT('h0103)
	) name22681 (
		_w28504_,
		_w28506_,
		_w28507_,
		_w28505_,
		_w28508_
	);
	LUT3 #(
		.INIT('h20)
	) name22682 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28509_
	);
	LUT4 #(
		.INIT('h2000)
	) name22683 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28510_
	);
	LUT4 #(
		.INIT('h9990)
	) name22684 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28511_
	);
	LUT4 #(
		.INIT('h0990)
	) name22685 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28512_
	);
	LUT3 #(
		.INIT('h0b)
	) name22686 (
		_w28492_,
		_w28510_,
		_w28512_,
		_w28513_
	);
	LUT3 #(
		.INIT('h80)
	) name22687 (
		_w28493_,
		_w28495_,
		_w28497_,
		_w28514_
	);
	LUT3 #(
		.INIT('h80)
	) name22688 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28515_
	);
	LUT4 #(
		.INIT('h7b5b)
	) name22689 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28516_
	);
	LUT2 #(
		.INIT('h2)
	) name22690 (
		_w28493_,
		_w28492_,
		_w28517_
	);
	LUT4 #(
		.INIT('h7077)
	) name22691 (
		_w28499_,
		_w28514_,
		_w28516_,
		_w28517_,
		_w28518_
	);
	LUT4 #(
		.INIT('hea00)
	) name22692 (
		_w28493_,
		_w28508_,
		_w28513_,
		_w28518_,
		_w28519_
	);
	LUT3 #(
		.INIT('h65)
	) name22693 (
		\u0_L8_reg[6]/NET0131 ,
		_w28502_,
		_w28519_,
		_w28520_
	);
	LUT2 #(
		.INIT('h2)
	) name22694 (
		_w28063_,
		_w28062_,
		_w28521_
	);
	LUT4 #(
		.INIT('h4080)
	) name22695 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28522_
	);
	LUT4 #(
		.INIT('h956e)
	) name22696 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28523_
	);
	LUT2 #(
		.INIT('h2)
	) name22697 (
		_w28521_,
		_w28523_,
		_w28524_
	);
	LUT4 #(
		.INIT('h2210)
	) name22698 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28525_
	);
	LUT2 #(
		.INIT('h4)
	) name22699 (
		_w28063_,
		_w28062_,
		_w28526_
	);
	LUT2 #(
		.INIT('h9)
	) name22700 (
		_w28063_,
		_w28062_,
		_w28527_
	);
	LUT4 #(
		.INIT('h0100)
	) name22701 (
		_w28461_,
		_w28522_,
		_w28525_,
		_w28527_,
		_w28528_
	);
	LUT3 #(
		.INIT('h48)
	) name22702 (
		_w28064_,
		_w28065_,
		_w28066_,
		_w28529_
	);
	LUT3 #(
		.INIT('h41)
	) name22703 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28530_
	);
	LUT4 #(
		.INIT('h0888)
	) name22704 (
		_w28064_,
		_w28067_,
		_w28065_,
		_w28066_,
		_w28531_
	);
	LUT4 #(
		.INIT('h0002)
	) name22705 (
		_w28526_,
		_w28531_,
		_w28530_,
		_w28529_,
		_w28532_
	);
	LUT4 #(
		.INIT('h00ab)
	) name22706 (
		_w28068_,
		_w28524_,
		_w28528_,
		_w28532_,
		_w28533_
	);
	LUT2 #(
		.INIT('h6)
	) name22707 (
		\u0_L8_reg[7]/NET0131 ,
		_w28533_,
		_w28534_
	);
	LUT4 #(
		.INIT('h8228)
	) name22708 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28535_
	);
	LUT3 #(
		.INIT('h43)
	) name22709 (
		_w27999_,
		_w28000_,
		_w28005_,
		_w28536_
	);
	LUT2 #(
		.INIT('h2)
	) name22710 (
		_w28002_,
		_w28003_,
		_w28537_
	);
	LUT4 #(
		.INIT('h0015)
	) name22711 (
		_w28099_,
		_w28536_,
		_w28537_,
		_w28535_,
		_w28538_
	);
	LUT2 #(
		.INIT('h2)
	) name22712 (
		_w27998_,
		_w28538_,
		_w28539_
	);
	LUT3 #(
		.INIT('h40)
	) name22713 (
		_w28003_,
		_w27999_,
		_w28005_,
		_w28540_
	);
	LUT3 #(
		.INIT('h28)
	) name22714 (
		_w28002_,
		_w28000_,
		_w28005_,
		_w28541_
	);
	LUT4 #(
		.INIT('h4000)
	) name22715 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28542_
	);
	LUT3 #(
		.INIT('h0b)
	) name22716 (
		_w28540_,
		_w28541_,
		_w28542_,
		_w28543_
	);
	LUT4 #(
		.INIT('h1005)
	) name22717 (
		_w28002_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28544_
	);
	LUT4 #(
		.INIT('h0082)
	) name22718 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28545_
	);
	LUT2 #(
		.INIT('h1)
	) name22719 (
		_w28544_,
		_w28545_,
		_w28546_
	);
	LUT4 #(
		.INIT('h9fff)
	) name22720 (
		_w28003_,
		_w27999_,
		_w28000_,
		_w28005_,
		_w28547_
	);
	LUT2 #(
		.INIT('h1)
	) name22721 (
		_w28002_,
		_w28547_,
		_w28548_
	);
	LUT4 #(
		.INIT('h00ea)
	) name22722 (
		_w27998_,
		_w28543_,
		_w28546_,
		_w28548_,
		_w28549_
	);
	LUT3 #(
		.INIT('h65)
	) name22723 (
		\u0_L8_reg[9]/NET0131 ,
		_w28539_,
		_w28549_,
		_w28550_
	);
	LUT4 #(
		.INIT('h3dc3)
	) name22724 (
		_w28492_,
		_w28494_,
		_w28496_,
		_w28495_,
		_w28551_
	);
	LUT4 #(
		.INIT('h0110)
	) name22725 (
		_w28492_,
		_w28494_,
		_w28496_,
		_w28497_,
		_w28552_
	);
	LUT4 #(
		.INIT('h0074)
	) name22726 (
		_w28509_,
		_w28497_,
		_w28551_,
		_w28552_,
		_w28553_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name22727 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28554_
	);
	LUT4 #(
		.INIT('h2880)
	) name22728 (
		_w28492_,
		_w28494_,
		_w28496_,
		_w28495_,
		_w28555_
	);
	LUT4 #(
		.INIT('h0032)
	) name22729 (
		_w28492_,
		_w28500_,
		_w28554_,
		_w28555_,
		_w28556_
	);
	LUT4 #(
		.INIT('hbeff)
	) name22730 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28557_
	);
	LUT4 #(
		.INIT('h0400)
	) name22731 (
		_w28492_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28558_
	);
	LUT3 #(
		.INIT('h0d)
	) name22732 (
		_w28492_,
		_w28557_,
		_w28558_,
		_w28559_
	);
	LUT4 #(
		.INIT('he400)
	) name22733 (
		_w28493_,
		_w28556_,
		_w28553_,
		_w28559_,
		_w28560_
	);
	LUT2 #(
		.INIT('h9)
	) name22734 (
		\u0_L8_reg[16]/NET0131 ,
		_w28560_,
		_w28561_
	);
	LUT2 #(
		.INIT('h4)
	) name22735 (
		_w28492_,
		_w28511_,
		_w28562_
	);
	LUT4 #(
		.INIT('h1dff)
	) name22736 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28563_
	);
	LUT2 #(
		.INIT('h2)
	) name22737 (
		_w28492_,
		_w28563_,
		_w28564_
	);
	LUT2 #(
		.INIT('h2)
	) name22738 (
		_w28492_,
		_w28497_,
		_w28565_
	);
	LUT3 #(
		.INIT('h0d)
	) name22739 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28566_
	);
	LUT4 #(
		.INIT('h0777)
	) name22740 (
		_w28504_,
		_w28505_,
		_w28565_,
		_w28566_,
		_w28567_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name22741 (
		_w28493_,
		_w28564_,
		_w28562_,
		_w28567_,
		_w28568_
	);
	LUT4 #(
		.INIT('he2cd)
	) name22742 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28569_
	);
	LUT4 #(
		.INIT('h0400)
	) name22743 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28570_
	);
	LUT4 #(
		.INIT('h5504)
	) name22744 (
		_w28493_,
		_w28492_,
		_w28569_,
		_w28570_,
		_w28571_
	);
	LUT4 #(
		.INIT('h0009)
	) name22745 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28572_
	);
	LUT4 #(
		.INIT('h9db6)
	) name22746 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28573_
	);
	LUT2 #(
		.INIT('h1)
	) name22747 (
		_w28493_,
		_w28492_,
		_w28574_
	);
	LUT2 #(
		.INIT('h4)
	) name22748 (
		_w28573_,
		_w28574_,
		_w28575_
	);
	LUT3 #(
		.INIT('hdb)
	) name22749 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28576_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name22750 (
		_w28492_,
		_w28497_,
		_w28515_,
		_w28576_,
		_w28577_
	);
	LUT3 #(
		.INIT('h10)
	) name22751 (
		_w28571_,
		_w28575_,
		_w28577_,
		_w28578_
	);
	LUT3 #(
		.INIT('h65)
	) name22752 (
		\u0_L8_reg[24]/NET0131 ,
		_w28568_,
		_w28578_,
		_w28579_
	);
	LUT4 #(
		.INIT('h0200)
	) name22753 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28580_
	);
	LUT3 #(
		.INIT('h01)
	) name22754 (
		_w28493_,
		_w28572_,
		_w28580_,
		_w28581_
	);
	LUT2 #(
		.INIT('h8)
	) name22755 (
		_w28496_,
		_w28497_,
		_w28582_
	);
	LUT4 #(
		.INIT('h73af)
	) name22756 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28583_
	);
	LUT4 #(
		.INIT('hdf53)
	) name22757 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28584_
	);
	LUT3 #(
		.INIT('hd8)
	) name22758 (
		_w28492_,
		_w28583_,
		_w28584_,
		_w28585_
	);
	LUT4 #(
		.INIT('heed9)
	) name22759 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28586_
	);
	LUT4 #(
		.INIT('h23ef)
	) name22760 (
		_w28494_,
		_w28496_,
		_w28495_,
		_w28497_,
		_w28587_
	);
	LUT4 #(
		.INIT('ha820)
	) name22761 (
		_w28493_,
		_w28492_,
		_w28587_,
		_w28586_,
		_w28588_
	);
	LUT3 #(
		.INIT('h07)
	) name22762 (
		_w28581_,
		_w28585_,
		_w28588_,
		_w28589_
	);
	LUT3 #(
		.INIT('h08)
	) name22763 (
		_w28492_,
		_w28494_,
		_w28495_,
		_w28590_
	);
	LUT2 #(
		.INIT('h8)
	) name22764 (
		_w28582_,
		_w28590_,
		_w28591_
	);
	LUT4 #(
		.INIT('h1000)
	) name22765 (
		_w28492_,
		_w28494_,
		_w28495_,
		_w28497_,
		_w28592_
	);
	LUT3 #(
		.INIT('h0b)
	) name22766 (
		_w28503_,
		_w28514_,
		_w28592_,
		_w28593_
	);
	LUT2 #(
		.INIT('h4)
	) name22767 (
		_w28591_,
		_w28593_,
		_w28594_
	);
	LUT3 #(
		.INIT('h9a)
	) name22768 (
		\u0_L8_reg[30]/NET0131 ,
		_w28589_,
		_w28594_,
		_w28595_
	);
	LUT4 #(
		.INIT('h5200)
	) name22769 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28158_,
		_w28596_
	);
	LUT4 #(
		.INIT('hfb73)
	) name22770 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28597_
	);
	LUT4 #(
		.INIT('h0032)
	) name22771 (
		_w28158_,
		_w28181_,
		_w28597_,
		_w28596_,
		_w28598_
	);
	LUT4 #(
		.INIT('h8000)
	) name22772 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28158_,
		_w28599_
	);
	LUT4 #(
		.INIT('hbffa)
	) name22773 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28600_
	);
	LUT4 #(
		.INIT('h0411)
	) name22774 (
		_w28160_,
		_w28161_,
		_w28158_,
		_w28162_,
		_w28601_
	);
	LUT4 #(
		.INIT('h0100)
	) name22775 (
		_w28180_,
		_w28599_,
		_w28601_,
		_w28600_,
		_w28602_
	);
	LUT4 #(
		.INIT('h0020)
	) name22776 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28158_,
		_w28603_
	);
	LUT4 #(
		.INIT('h77ef)
	) name22777 (
		_w28159_,
		_w28160_,
		_w28161_,
		_w28162_,
		_w28604_
	);
	LUT3 #(
		.INIT('h31)
	) name22778 (
		_w28158_,
		_w28603_,
		_w28604_,
		_w28605_
	);
	LUT4 #(
		.INIT('hd800)
	) name22779 (
		_w28164_,
		_w28598_,
		_w28602_,
		_w28605_,
		_w28606_
	);
	LUT2 #(
		.INIT('h9)
	) name22780 (
		\u0_L8_reg[18]/NET0131 ,
		_w28606_,
		_w28607_
	);
	LUT4 #(
		.INIT('hc693)
	) name22781 (
		decrypt_pad,
		\u0_R7_reg[28]/NET0131 ,
		\u0_uk_K_r7_reg[23]/P0001 ,
		\u0_uk_K_r7_reg[30]/P0001 ,
		_w28608_
	);
	LUT4 #(
		.INIT('hc693)
	) name22782 (
		decrypt_pad,
		\u0_R7_reg[27]/NET0131 ,
		\u0_uk_K_r7_reg[36]/NET0131 ,
		\u0_uk_K_r7_reg[43]/NET0131 ,
		_w28609_
	);
	LUT4 #(
		.INIT('hc693)
	) name22783 (
		decrypt_pad,
		\u0_R7_reg[26]/NET0131 ,
		\u0_uk_K_r7_reg[31]/NET0131 ,
		\u0_uk_K_r7_reg[38]/NET0131 ,
		_w28610_
	);
	LUT4 #(
		.INIT('hc963)
	) name22784 (
		decrypt_pad,
		\u0_R7_reg[24]/NET0131 ,
		\u0_uk_K_r7_reg[14]/NET0131 ,
		\u0_uk_K_r7_reg[7]/NET0131 ,
		_w28611_
	);
	LUT2 #(
		.INIT('h9)
	) name22785 (
		_w28610_,
		_w28611_,
		_w28612_
	);
	LUT4 #(
		.INIT('hc693)
	) name22786 (
		decrypt_pad,
		\u0_R7_reg[29]/NET0131 ,
		\u0_uk_K_r7_reg[15]/NET0131 ,
		\u0_uk_K_r7_reg[22]/NET0131 ,
		_w28613_
	);
	LUT4 #(
		.INIT('hc693)
	) name22787 (
		decrypt_pad,
		\u0_R7_reg[25]/NET0131 ,
		\u0_uk_K_r7_reg[42]/NET0131 ,
		\u0_uk_K_r7_reg[49]/NET0131 ,
		_w28614_
	);
	LUT4 #(
		.INIT('h0002)
	) name22788 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28615_
	);
	LUT4 #(
		.INIT('h6369)
	) name22789 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28616_
	);
	LUT4 #(
		.INIT('h9000)
	) name22790 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28617_
	);
	LUT3 #(
		.INIT('h04)
	) name22791 (
		_w28610_,
		_w28611_,
		_w28614_,
		_w28618_
	);
	LUT4 #(
		.INIT('h1054)
	) name22792 (
		_w28617_,
		_w28609_,
		_w28616_,
		_w28618_,
		_w28619_
	);
	LUT2 #(
		.INIT('h1)
	) name22793 (
		_w28608_,
		_w28619_,
		_w28620_
	);
	LUT3 #(
		.INIT('h0b)
	) name22794 (
		_w28610_,
		_w28611_,
		_w28614_,
		_w28621_
	);
	LUT4 #(
		.INIT('h20a0)
	) name22795 (
		_w28608_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28622_
	);
	LUT4 #(
		.INIT('h3031)
	) name22796 (
		_w28612_,
		_w28609_,
		_w28621_,
		_w28622_,
		_w28623_
	);
	LUT4 #(
		.INIT('h0200)
	) name22797 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28624_
	);
	LUT4 #(
		.INIT('h0020)
	) name22798 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28625_
	);
	LUT4 #(
		.INIT('hffd2)
	) name22799 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28626_
	);
	LUT3 #(
		.INIT('h20)
	) name22800 (
		_w28609_,
		_w28624_,
		_w28626_,
		_w28627_
	);
	LUT3 #(
		.INIT('h40)
	) name22801 (
		_w28610_,
		_w28613_,
		_w28614_,
		_w28628_
	);
	LUT3 #(
		.INIT('hb5)
	) name22802 (
		_w28610_,
		_w28613_,
		_w28614_,
		_w28629_
	);
	LUT2 #(
		.INIT('h8)
	) name22803 (
		_w28611_,
		_w28609_,
		_w28630_
	);
	LUT4 #(
		.INIT('hffde)
	) name22804 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28631_
	);
	LUT4 #(
		.INIT('h20aa)
	) name22805 (
		_w28608_,
		_w28629_,
		_w28630_,
		_w28631_,
		_w28632_
	);
	LUT3 #(
		.INIT('h0e)
	) name22806 (
		_w28623_,
		_w28627_,
		_w28632_,
		_w28633_
	);
	LUT3 #(
		.INIT('h65)
	) name22807 (
		\u0_L7_reg[22]/NET0131 ,
		_w28620_,
		_w28633_,
		_w28634_
	);
	LUT4 #(
		.INIT('hc693)
	) name22808 (
		decrypt_pad,
		\u0_R7_reg[32]/NET0131 ,
		\u0_uk_K_r7_reg[24]/NET0131 ,
		\u0_uk_K_r7_reg[6]/NET0131 ,
		_w28635_
	);
	LUT4 #(
		.INIT('hc693)
	) name22809 (
		decrypt_pad,
		\u0_R7_reg[5]/NET0131 ,
		\u0_uk_K_r7_reg[18]/NET0131 ,
		\u0_uk_K_r7_reg[25]/NET0131 ,
		_w28636_
	);
	LUT2 #(
		.INIT('h4)
	) name22810 (
		_w28635_,
		_w28636_,
		_w28637_
	);
	LUT4 #(
		.INIT('hc693)
	) name22811 (
		decrypt_pad,
		\u0_R7_reg[3]/NET0131 ,
		\u0_uk_K_r7_reg[12]/NET0131 ,
		\u0_uk_K_r7_reg[19]/NET0131 ,
		_w28638_
	);
	LUT4 #(
		.INIT('hc963)
	) name22812 (
		decrypt_pad,
		\u0_R7_reg[2]/NET0131 ,
		\u0_uk_K_r7_reg[10]/NET0131 ,
		\u0_uk_K_r7_reg[3]/NET0131 ,
		_w28639_
	);
	LUT2 #(
		.INIT('h2)
	) name22813 (
		_w28638_,
		_w28639_,
		_w28640_
	);
	LUT4 #(
		.INIT('hc693)
	) name22814 (
		decrypt_pad,
		\u0_R7_reg[1]/NET0131 ,
		\u0_uk_K_r7_reg[20]/NET0131 ,
		\u0_uk_K_r7_reg[27]/NET0131 ,
		_w28641_
	);
	LUT3 #(
		.INIT('hd0)
	) name22815 (
		_w28638_,
		_w28639_,
		_w28641_,
		_w28642_
	);
	LUT4 #(
		.INIT('hc693)
	) name22816 (
		decrypt_pad,
		\u0_R7_reg[4]/NET0131 ,
		\u0_uk_K_r7_reg[47]/NET0131 ,
		\u0_uk_K_r7_reg[54]/NET0131 ,
		_w28643_
	);
	LUT4 #(
		.INIT('h0004)
	) name22817 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28644_
	);
	LUT4 #(
		.INIT('h00c4)
	) name22818 (
		_w28637_,
		_w28643_,
		_w28642_,
		_w28644_,
		_w28645_
	);
	LUT3 #(
		.INIT('h0d)
	) name22819 (
		_w28639_,
		_w28635_,
		_w28636_,
		_w28646_
	);
	LUT3 #(
		.INIT('h2a)
	) name22820 (
		_w28638_,
		_w28641_,
		_w28636_,
		_w28647_
	);
	LUT4 #(
		.INIT('h500c)
	) name22821 (
		_w28638_,
		_w28639_,
		_w28635_,
		_w28641_,
		_w28648_
	);
	LUT3 #(
		.INIT('h0b)
	) name22822 (
		_w28646_,
		_w28647_,
		_w28648_,
		_w28649_
	);
	LUT4 #(
		.INIT('h73cf)
	) name22823 (
		_w28638_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28650_
	);
	LUT2 #(
		.INIT('h1)
	) name22824 (
		_w28639_,
		_w28650_,
		_w28651_
	);
	LUT2 #(
		.INIT('h6)
	) name22825 (
		_w28635_,
		_w28636_,
		_w28652_
	);
	LUT3 #(
		.INIT('h80)
	) name22826 (
		_w28638_,
		_w28639_,
		_w28641_,
		_w28653_
	);
	LUT3 #(
		.INIT('h15)
	) name22827 (
		_w28643_,
		_w28652_,
		_w28653_,
		_w28654_
	);
	LUT4 #(
		.INIT('h7077)
	) name22828 (
		_w28645_,
		_w28649_,
		_w28651_,
		_w28654_,
		_w28655_
	);
	LUT2 #(
		.INIT('h9)
	) name22829 (
		_w28639_,
		_w28635_,
		_w28656_
	);
	LUT4 #(
		.INIT('h0047)
	) name22830 (
		_w28639_,
		_w28641_,
		_w28636_,
		_w28643_,
		_w28657_
	);
	LUT4 #(
		.INIT('h7daf)
	) name22831 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28658_
	);
	LUT4 #(
		.INIT('h4055)
	) name22832 (
		_w28638_,
		_w28656_,
		_w28657_,
		_w28658_,
		_w28659_
	);
	LUT4 #(
		.INIT('h0020)
	) name22833 (
		_w28638_,
		_w28639_,
		_w28635_,
		_w28641_,
		_w28660_
	);
	LUT3 #(
		.INIT('h02)
	) name22834 (
		_w28639_,
		_w28641_,
		_w28636_,
		_w28661_
	);
	LUT2 #(
		.INIT('h2)
	) name22835 (
		_w28638_,
		_w28635_,
		_w28662_
	);
	LUT3 #(
		.INIT('h15)
	) name22836 (
		_w28660_,
		_w28661_,
		_w28662_,
		_w28663_
	);
	LUT2 #(
		.INIT('h4)
	) name22837 (
		_w28659_,
		_w28663_,
		_w28664_
	);
	LUT3 #(
		.INIT('h65)
	) name22838 (
		\u0_L7_reg[31]/NET0131 ,
		_w28655_,
		_w28664_,
		_w28665_
	);
	LUT4 #(
		.INIT('hc693)
	) name22839 (
		decrypt_pad,
		\u0_R7_reg[23]/NET0131 ,
		\u0_uk_K_r7_reg[14]/NET0131 ,
		\u0_uk_K_r7_reg[21]/NET0131 ,
		_w28666_
	);
	LUT4 #(
		.INIT('hc693)
	) name22840 (
		decrypt_pad,
		\u0_R7_reg[25]/NET0131 ,
		\u0_uk_K_r7_reg[35]/NET0131 ,
		\u0_uk_K_r7_reg[42]/NET0131 ,
		_w28667_
	);
	LUT4 #(
		.INIT('hc963)
	) name22841 (
		decrypt_pad,
		\u0_R7_reg[20]/NET0131 ,
		\u0_uk_K_r7_reg[2]/NET0131 ,
		\u0_uk_K_r7_reg[50]/NET0131 ,
		_w28668_
	);
	LUT4 #(
		.INIT('hc693)
	) name22842 (
		decrypt_pad,
		\u0_R7_reg[22]/NET0131 ,
		\u0_uk_K_r7_reg[1]/NET0131 ,
		\u0_uk_K_r7_reg[8]/NET0131 ,
		_w28669_
	);
	LUT3 #(
		.INIT('h80)
	) name22843 (
		_w28667_,
		_w28668_,
		_w28669_,
		_w28670_
	);
	LUT4 #(
		.INIT('hc693)
	) name22844 (
		decrypt_pad,
		\u0_R7_reg[21]/NET0131 ,
		\u0_uk_K_r7_reg[38]/NET0131 ,
		\u0_uk_K_r7_reg[45]/NET0131 ,
		_w28671_
	);
	LUT4 #(
		.INIT('hfdcc)
	) name22845 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28672_
	);
	LUT4 #(
		.INIT('hc693)
	) name22846 (
		decrypt_pad,
		\u0_R7_reg[24]/NET0131 ,
		\u0_uk_K_r7_reg[16]/NET0131 ,
		\u0_uk_K_r7_reg[23]/P0001 ,
		_w28673_
	);
	LUT4 #(
		.INIT('h0010)
	) name22847 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28674_
	);
	LUT2 #(
		.INIT('h2)
	) name22848 (
		_w28673_,
		_w28674_,
		_w28675_
	);
	LUT4 #(
		.INIT('h3032)
	) name22849 (
		_w28673_,
		_w28670_,
		_w28672_,
		_w28674_,
		_w28676_
	);
	LUT2 #(
		.INIT('h2)
	) name22850 (
		_w28666_,
		_w28676_,
		_w28677_
	);
	LUT4 #(
		.INIT('h0004)
	) name22851 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28678_
	);
	LUT3 #(
		.INIT('h40)
	) name22852 (
		_w28668_,
		_w28671_,
		_w28669_,
		_w28679_
	);
	LUT4 #(
		.INIT('h4f7b)
	) name22853 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28680_
	);
	LUT2 #(
		.INIT('h2)
	) name22854 (
		_w28666_,
		_w28680_,
		_w28681_
	);
	LUT3 #(
		.INIT('h07)
	) name22855 (
		_w28667_,
		_w28671_,
		_w28669_,
		_w28682_
	);
	LUT3 #(
		.INIT('h15)
	) name22856 (
		_w28666_,
		_w28667_,
		_w28668_,
		_w28683_
	);
	LUT3 #(
		.INIT('h10)
	) name22857 (
		_w28679_,
		_w28682_,
		_w28683_,
		_w28684_
	);
	LUT3 #(
		.INIT('h08)
	) name22858 (
		_w28667_,
		_w28668_,
		_w28669_,
		_w28685_
	);
	LUT2 #(
		.INIT('h1)
	) name22859 (
		_w28666_,
		_w28671_,
		_w28686_
	);
	LUT2 #(
		.INIT('h8)
	) name22860 (
		_w28685_,
		_w28686_,
		_w28687_
	);
	LUT3 #(
		.INIT('h2a)
	) name22861 (
		_w28673_,
		_w28685_,
		_w28686_,
		_w28688_
	);
	LUT3 #(
		.INIT('h10)
	) name22862 (
		_w28681_,
		_w28684_,
		_w28688_,
		_w28689_
	);
	LUT4 #(
		.INIT('h1040)
	) name22863 (
		_w28666_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28690_
	);
	LUT2 #(
		.INIT('h1)
	) name22864 (
		_w28673_,
		_w28690_,
		_w28691_
	);
	LUT4 #(
		.INIT('hf5cf)
	) name22865 (
		_w28666_,
		_w28667_,
		_w28671_,
		_w28669_,
		_w28692_
	);
	LUT2 #(
		.INIT('h1)
	) name22866 (
		_w28666_,
		_w28669_,
		_w28693_
	);
	LUT4 #(
		.INIT('h0010)
	) name22867 (
		_w28666_,
		_w28667_,
		_w28668_,
		_w28669_,
		_w28694_
	);
	LUT4 #(
		.INIT('h0800)
	) name22868 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28695_
	);
	LUT4 #(
		.INIT('h000d)
	) name22869 (
		_w28668_,
		_w28692_,
		_w28694_,
		_w28695_,
		_w28696_
	);
	LUT2 #(
		.INIT('h8)
	) name22870 (
		_w28691_,
		_w28696_,
		_w28697_
	);
	LUT3 #(
		.INIT('h01)
	) name22871 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28698_
	);
	LUT4 #(
		.INIT('h4555)
	) name22872 (
		_w28666_,
		_w28667_,
		_w28668_,
		_w28671_,
		_w28699_
	);
	LUT4 #(
		.INIT('h0002)
	) name22873 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28700_
	);
	LUT3 #(
		.INIT('h32)
	) name22874 (
		_w28693_,
		_w28699_,
		_w28700_,
		_w28701_
	);
	LUT4 #(
		.INIT('h7075)
	) name22875 (
		_w28693_,
		_w28698_,
		_w28699_,
		_w28700_,
		_w28702_
	);
	LUT4 #(
		.INIT('h0e00)
	) name22876 (
		_w28689_,
		_w28697_,
		_w28677_,
		_w28702_,
		_w28703_
	);
	LUT2 #(
		.INIT('h6)
	) name22877 (
		\u0_L7_reg[11]/NET0131 ,
		_w28703_,
		_w28704_
	);
	LUT4 #(
		.INIT('hc693)
	) name22878 (
		decrypt_pad,
		\u0_R7_reg[31]/P0001 ,
		\u0_uk_K_r7_reg[37]/NET0131 ,
		\u0_uk_K_r7_reg[44]/NET0131 ,
		_w28705_
	);
	LUT4 #(
		.INIT('hc693)
	) name22879 (
		decrypt_pad,
		\u0_R7_reg[28]/NET0131 ,
		\u0_uk_K_r7_reg[21]/NET0131 ,
		\u0_uk_K_r7_reg[28]/NET0131 ,
		_w28706_
	);
	LUT4 #(
		.INIT('hc963)
	) name22880 (
		decrypt_pad,
		\u0_R7_reg[30]/NET0131 ,
		\u0_uk_K_r7_reg[1]/NET0131 ,
		\u0_uk_K_r7_reg[49]/NET0131 ,
		_w28707_
	);
	LUT4 #(
		.INIT('hc963)
	) name22881 (
		decrypt_pad,
		\u0_R7_reg[1]/NET0131 ,
		\u0_uk_K_r7_reg[16]/NET0131 ,
		\u0_uk_K_r7_reg[9]/NET0131 ,
		_w28708_
	);
	LUT4 #(
		.INIT('hc963)
	) name22882 (
		decrypt_pad,
		\u0_R7_reg[29]/NET0131 ,
		\u0_uk_K_r7_reg[0]/NET0131 ,
		\u0_uk_K_r7_reg[52]/NET0131 ,
		_w28709_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name22883 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28710_
	);
	LUT4 #(
		.INIT('h0200)
	) name22884 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28711_
	);
	LUT4 #(
		.INIT('hc693)
	) name22885 (
		decrypt_pad,
		\u0_R7_reg[32]/NET0131 ,
		\u0_uk_K_r7_reg[43]/NET0131 ,
		\u0_uk_K_r7_reg[50]/NET0131 ,
		_w28712_
	);
	LUT3 #(
		.INIT('h01)
	) name22886 (
		_w28706_,
		_w28707_,
		_w28709_,
		_w28713_
	);
	LUT4 #(
		.INIT('h0001)
	) name22887 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28714_
	);
	LUT4 #(
		.INIT('h0040)
	) name22888 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28715_
	);
	LUT4 #(
		.INIT('hefb6)
	) name22889 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28716_
	);
	LUT4 #(
		.INIT('hef00)
	) name22890 (
		_w28711_,
		_w28710_,
		_w28712_,
		_w28716_,
		_w28717_
	);
	LUT2 #(
		.INIT('h2)
	) name22891 (
		_w28705_,
		_w28717_,
		_w28718_
	);
	LUT4 #(
		.INIT('hff9b)
	) name22892 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28719_
	);
	LUT3 #(
		.INIT('h20)
	) name22893 (
		_w28705_,
		_w28711_,
		_w28719_,
		_w28720_
	);
	LUT4 #(
		.INIT('hdc10)
	) name22894 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28721_
	);
	LUT3 #(
		.INIT('h51)
	) name22895 (
		_w28705_,
		_w28706_,
		_w28707_,
		_w28722_
	);
	LUT2 #(
		.INIT('h4)
	) name22896 (
		_w28721_,
		_w28722_,
		_w28723_
	);
	LUT4 #(
		.INIT('h8000)
	) name22897 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28724_
	);
	LUT2 #(
		.INIT('h1)
	) name22898 (
		_w28712_,
		_w28724_,
		_w28725_
	);
	LUT4 #(
		.INIT('hfd5a)
	) name22899 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28726_
	);
	LUT3 #(
		.INIT('h40)
	) name22900 (
		_w28706_,
		_w28708_,
		_w28709_,
		_w28727_
	);
	LUT4 #(
		.INIT('h4000)
	) name22901 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28728_
	);
	LUT4 #(
		.INIT('h0c08)
	) name22902 (
		_w28705_,
		_w28712_,
		_w28728_,
		_w28726_,
		_w28729_
	);
	LUT4 #(
		.INIT('h001f)
	) name22903 (
		_w28720_,
		_w28723_,
		_w28725_,
		_w28729_,
		_w28730_
	);
	LUT3 #(
		.INIT('ha9)
	) name22904 (
		\u0_L7_reg[5]/NET0131 ,
		_w28718_,
		_w28730_,
		_w28731_
	);
	LUT2 #(
		.INIT('h2)
	) name22905 (
		_w28705_,
		_w28706_,
		_w28732_
	);
	LUT3 #(
		.INIT('h08)
	) name22906 (
		_w28708_,
		_w28707_,
		_w28709_,
		_w28733_
	);
	LUT2 #(
		.INIT('h4)
	) name22907 (
		_w28732_,
		_w28733_,
		_w28734_
	);
	LUT3 #(
		.INIT('h20)
	) name22908 (
		_w28706_,
		_w28707_,
		_w28709_,
		_w28735_
	);
	LUT4 #(
		.INIT('hdf00)
	) name22909 (
		_w28706_,
		_w28707_,
		_w28709_,
		_w28712_,
		_w28736_
	);
	LUT4 #(
		.INIT('h1000)
	) name22910 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28737_
	);
	LUT4 #(
		.INIT('h0002)
	) name22911 (
		_w28705_,
		_w28706_,
		_w28708_,
		_w28709_,
		_w28738_
	);
	LUT3 #(
		.INIT('h10)
	) name22912 (
		_w28737_,
		_w28738_,
		_w28736_,
		_w28739_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name22913 (
		_w28705_,
		_w28706_,
		_w28708_,
		_w28709_,
		_w28740_
	);
	LUT4 #(
		.INIT('h10bb)
	) name22914 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28741_
	);
	LUT4 #(
		.INIT('h0002)
	) name22915 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28742_
	);
	LUT4 #(
		.INIT('h1101)
	) name22916 (
		_w28712_,
		_w28742_,
		_w28740_,
		_w28741_,
		_w28743_
	);
	LUT3 #(
		.INIT('h0b)
	) name22917 (
		_w28734_,
		_w28739_,
		_w28743_,
		_w28744_
	);
	LUT4 #(
		.INIT('h0004)
	) name22918 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28745_
	);
	LUT3 #(
		.INIT('h02)
	) name22919 (
		_w28705_,
		_w28728_,
		_w28745_,
		_w28746_
	);
	LUT4 #(
		.INIT('h080a)
	) name22920 (
		_w28706_,
		_w28707_,
		_w28709_,
		_w28712_,
		_w28747_
	);
	LUT4 #(
		.INIT('h0400)
	) name22921 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28748_
	);
	LUT4 #(
		.INIT('h0001)
	) name22922 (
		_w28705_,
		_w28737_,
		_w28747_,
		_w28748_,
		_w28749_
	);
	LUT3 #(
		.INIT('h23)
	) name22923 (
		_w28714_,
		_w28746_,
		_w28749_,
		_w28750_
	);
	LUT3 #(
		.INIT('h56)
	) name22924 (
		\u0_L7_reg[15]/P0001 ,
		_w28744_,
		_w28750_,
		_w28751_
	);
	LUT4 #(
		.INIT('hc963)
	) name22925 (
		decrypt_pad,
		\u0_R7_reg[17]/NET0131 ,
		\u0_uk_K_r7_reg[4]/NET0131 ,
		\u0_uk_K_r7_reg[54]/NET0131 ,
		_w28752_
	);
	LUT4 #(
		.INIT('hc693)
	) name22926 (
		decrypt_pad,
		\u0_R7_reg[14]/NET0131 ,
		\u0_uk_K_r7_reg[33]/NET0131 ,
		\u0_uk_K_r7_reg[40]/NET0131 ,
		_w28753_
	);
	LUT4 #(
		.INIT('hc693)
	) name22927 (
		decrypt_pad,
		\u0_R7_reg[13]/NET0131 ,
		\u0_uk_K_r7_reg[32]/NET0131 ,
		\u0_uk_K_r7_reg[39]/NET0131 ,
		_w28754_
	);
	LUT4 #(
		.INIT('hc693)
	) name22928 (
		decrypt_pad,
		\u0_R7_reg[12]/NET0131 ,
		\u0_uk_K_r7_reg[13]/NET0131 ,
		\u0_uk_K_r7_reg[20]/NET0131 ,
		_w28755_
	);
	LUT2 #(
		.INIT('h4)
	) name22929 (
		_w28755_,
		_w28753_,
		_w28756_
	);
	LUT4 #(
		.INIT('hc693)
	) name22930 (
		decrypt_pad,
		\u0_R7_reg[15]/NET0131 ,
		\u0_uk_K_r7_reg[41]/NET0131 ,
		\u0_uk_K_r7_reg[48]/NET0131 ,
		_w28757_
	);
	LUT4 #(
		.INIT('h44cf)
	) name22931 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28757_,
		_w28758_
	);
	LUT2 #(
		.INIT('h2)
	) name22932 (
		_w28752_,
		_w28758_,
		_w28759_
	);
	LUT2 #(
		.INIT('h8)
	) name22933 (
		_w28754_,
		_w28752_,
		_w28760_
	);
	LUT2 #(
		.INIT('h4)
	) name22934 (
		_w28754_,
		_w28757_,
		_w28761_
	);
	LUT4 #(
		.INIT('h4044)
	) name22935 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28757_,
		_w28762_
	);
	LUT2 #(
		.INIT('h4)
	) name22936 (
		_w28760_,
		_w28762_,
		_w28763_
	);
	LUT3 #(
		.INIT('h20)
	) name22937 (
		_w28755_,
		_w28754_,
		_w28757_,
		_w28764_
	);
	LUT3 #(
		.INIT('h01)
	) name22938 (
		_w28754_,
		_w28757_,
		_w28752_,
		_w28765_
	);
	LUT4 #(
		.INIT('hc693)
	) name22939 (
		decrypt_pad,
		\u0_R7_reg[16]/NET0131 ,
		\u0_uk_K_r7_reg[17]/NET0131 ,
		\u0_uk_K_r7_reg[24]/NET0131 ,
		_w28766_
	);
	LUT3 #(
		.INIT('ha2)
	) name22940 (
		_w28766_,
		_w28755_,
		_w28753_,
		_w28767_
	);
	LUT3 #(
		.INIT('h10)
	) name22941 (
		_w28765_,
		_w28764_,
		_w28767_,
		_w28768_
	);
	LUT3 #(
		.INIT('h10)
	) name22942 (
		_w28759_,
		_w28763_,
		_w28768_,
		_w28769_
	);
	LUT4 #(
		.INIT('h0004)
	) name22943 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28757_,
		_w28770_
	);
	LUT3 #(
		.INIT('h02)
	) name22944 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28771_
	);
	LUT3 #(
		.INIT('h01)
	) name22945 (
		_w28771_,
		_w28770_,
		_w28765_,
		_w28772_
	);
	LUT4 #(
		.INIT('h0080)
	) name22946 (
		_w28755_,
		_w28754_,
		_w28757_,
		_w28752_,
		_w28773_
	);
	LUT2 #(
		.INIT('h4)
	) name22947 (
		_w28753_,
		_w28752_,
		_w28774_
	);
	LUT4 #(
		.INIT('h1000)
	) name22948 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28775_
	);
	LUT2 #(
		.INIT('h4)
	) name22949 (
		_w28755_,
		_w28752_,
		_w28776_
	);
	LUT3 #(
		.INIT('h80)
	) name22950 (
		_w28753_,
		_w28754_,
		_w28757_,
		_w28777_
	);
	LUT4 #(
		.INIT('h1011)
	) name22951 (
		_w28773_,
		_w28775_,
		_w28776_,
		_w28777_,
		_w28778_
	);
	LUT4 #(
		.INIT('hdfed)
	) name22952 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28779_
	);
	LUT3 #(
		.INIT('hed)
	) name22953 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28780_
	);
	LUT4 #(
		.INIT('hfa72)
	) name22954 (
		_w28757_,
		_w28752_,
		_w28779_,
		_w28780_,
		_w28781_
	);
	LUT4 #(
		.INIT('hea00)
	) name22955 (
		_w28766_,
		_w28772_,
		_w28778_,
		_w28781_,
		_w28782_
	);
	LUT3 #(
		.INIT('h65)
	) name22956 (
		\u0_L7_reg[26]/NET0131 ,
		_w28769_,
		_w28782_,
		_w28783_
	);
	LUT3 #(
		.INIT('h8c)
	) name22957 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28784_
	);
	LUT4 #(
		.INIT('h0080)
	) name22958 (
		_w28666_,
		_w28667_,
		_w28668_,
		_w28669_,
		_w28785_
	);
	LUT3 #(
		.INIT('h80)
	) name22959 (
		_w28667_,
		_w28671_,
		_w28669_,
		_w28786_
	);
	LUT4 #(
		.INIT('h0031)
	) name22960 (
		_w28693_,
		_w28785_,
		_w28784_,
		_w28786_,
		_w28787_
	);
	LUT2 #(
		.INIT('h8)
	) name22961 (
		_w28675_,
		_w28787_,
		_w28788_
	);
	LUT4 #(
		.INIT('h0200)
	) name22962 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28789_
	);
	LUT4 #(
		.INIT('hef67)
	) name22963 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28790_
	);
	LUT3 #(
		.INIT('h10)
	) name22964 (
		_w28666_,
		_w28789_,
		_w28790_,
		_w28791_
	);
	LUT3 #(
		.INIT('h02)
	) name22965 (
		_w28667_,
		_w28668_,
		_w28669_,
		_w28792_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name22966 (
		_w28666_,
		_w28667_,
		_w28668_,
		_w28671_,
		_w28793_
	);
	LUT3 #(
		.INIT('h10)
	) name22967 (
		_w28695_,
		_w28792_,
		_w28793_,
		_w28794_
	);
	LUT2 #(
		.INIT('h1)
	) name22968 (
		_w28673_,
		_w28678_,
		_w28795_
	);
	LUT3 #(
		.INIT('he0)
	) name22969 (
		_w28791_,
		_w28794_,
		_w28795_,
		_w28796_
	);
	LUT3 #(
		.INIT('h9e)
	) name22970 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28797_
	);
	LUT4 #(
		.INIT('h7bee)
	) name22971 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28798_
	);
	LUT4 #(
		.INIT('hf7a2)
	) name22972 (
		_w28666_,
		_w28669_,
		_w28797_,
		_w28798_,
		_w28799_
	);
	LUT4 #(
		.INIT('ha955)
	) name22973 (
		\u0_L7_reg[4]/NET0131 ,
		_w28788_,
		_w28796_,
		_w28799_,
		_w28800_
	);
	LUT4 #(
		.INIT('h0a22)
	) name22974 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28801_
	);
	LUT3 #(
		.INIT('h08)
	) name22975 (
		_w28755_,
		_w28753_,
		_w28752_,
		_w28802_
	);
	LUT4 #(
		.INIT('h0008)
	) name22976 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28803_
	);
	LUT3 #(
		.INIT('h01)
	) name22977 (
		_w28755_,
		_w28753_,
		_w28752_,
		_w28804_
	);
	LUT4 #(
		.INIT('heee4)
	) name22978 (
		_w28757_,
		_w28801_,
		_w28804_,
		_w28803_,
		_w28805_
	);
	LUT4 #(
		.INIT('h8000)
	) name22979 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28806_
	);
	LUT4 #(
		.INIT('h6fdf)
	) name22980 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28807_
	);
	LUT3 #(
		.INIT('h45)
	) name22981 (
		_w28766_,
		_w28805_,
		_w28807_,
		_w28808_
	);
	LUT4 #(
		.INIT('h00ef)
	) name22982 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28809_
	);
	LUT4 #(
		.INIT('h0070)
	) name22983 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28757_,
		_w28810_
	);
	LUT4 #(
		.INIT('h0080)
	) name22984 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28811_
	);
	LUT4 #(
		.INIT('hfb7b)
	) name22985 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28812_
	);
	LUT4 #(
		.INIT('h20aa)
	) name22986 (
		_w28766_,
		_w28809_,
		_w28810_,
		_w28812_,
		_w28813_
	);
	LUT4 #(
		.INIT('h0040)
	) name22987 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28814_
	);
	LUT4 #(
		.INIT('h7bff)
	) name22988 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28815_
	);
	LUT4 #(
		.INIT('h7bbf)
	) name22989 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28816_
	);
	LUT2 #(
		.INIT('h2)
	) name22990 (
		_w28757_,
		_w28816_,
		_w28817_
	);
	LUT2 #(
		.INIT('h4)
	) name22991 (
		_w28757_,
		_w28811_,
		_w28818_
	);
	LUT3 #(
		.INIT('h20)
	) name22992 (
		_w28766_,
		_w28754_,
		_w28757_,
		_w28819_
	);
	LUT3 #(
		.INIT('hf2)
	) name22993 (
		_w28755_,
		_w28753_,
		_w28752_,
		_w28820_
	);
	LUT4 #(
		.INIT('h0777)
	) name22994 (
		_w28756_,
		_w28765_,
		_w28819_,
		_w28820_,
		_w28821_
	);
	LUT4 #(
		.INIT('h0100)
	) name22995 (
		_w28817_,
		_w28818_,
		_w28813_,
		_w28821_,
		_w28822_
	);
	LUT3 #(
		.INIT('h65)
	) name22996 (
		\u0_L7_reg[1]/NET0131 ,
		_w28808_,
		_w28822_,
		_w28823_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name22997 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28824_
	);
	LUT3 #(
		.INIT('h41)
	) name22998 (
		_w28638_,
		_w28635_,
		_w28636_,
		_w28825_
	);
	LUT4 #(
		.INIT('h8008)
	) name22999 (
		_w28638_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28826_
	);
	LUT4 #(
		.INIT('h0080)
	) name23000 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28827_
	);
	LUT4 #(
		.INIT('hfd7f)
	) name23001 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28828_
	);
	LUT4 #(
		.INIT('h4500)
	) name23002 (
		_w28826_,
		_w28824_,
		_w28825_,
		_w28828_,
		_w28829_
	);
	LUT4 #(
		.INIT('h0400)
	) name23003 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28830_
	);
	LUT4 #(
		.INIT('hc9cd)
	) name23004 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28831_
	);
	LUT4 #(
		.INIT('h4041)
	) name23005 (
		_w28638_,
		_w28639_,
		_w28635_,
		_w28641_,
		_w28832_
	);
	LUT4 #(
		.INIT('h0040)
	) name23006 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28833_
	);
	LUT4 #(
		.INIT('h5fbf)
	) name23007 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w28834_
	);
	LUT4 #(
		.INIT('h0d00)
	) name23008 (
		_w28638_,
		_w28831_,
		_w28832_,
		_w28834_,
		_w28835_
	);
	LUT3 #(
		.INIT('hb7)
	) name23009 (
		_w28639_,
		_w28641_,
		_w28636_,
		_w28836_
	);
	LUT2 #(
		.INIT('h2)
	) name23010 (
		_w28662_,
		_w28836_,
		_w28837_
	);
	LUT4 #(
		.INIT('h0d08)
	) name23011 (
		_w28643_,
		_w28835_,
		_w28837_,
		_w28829_,
		_w28838_
	);
	LUT2 #(
		.INIT('h9)
	) name23012 (
		\u0_L7_reg[17]/NET0131 ,
		_w28838_,
		_w28839_
	);
	LUT4 #(
		.INIT('hc693)
	) name23013 (
		decrypt_pad,
		\u0_R7_reg[8]/NET0131 ,
		\u0_uk_K_r7_reg[48]/NET0131 ,
		\u0_uk_K_r7_reg[55]/P0001 ,
		_w28840_
	);
	LUT4 #(
		.INIT('hc963)
	) name23014 (
		decrypt_pad,
		\u0_R7_reg[6]/NET0131 ,
		\u0_uk_K_r7_reg[13]/NET0131 ,
		\u0_uk_K_r7_reg[6]/NET0131 ,
		_w28841_
	);
	LUT4 #(
		.INIT('hc963)
	) name23015 (
		decrypt_pad,
		\u0_R7_reg[9]/NET0131 ,
		\u0_uk_K_r7_reg[3]/NET0131 ,
		\u0_uk_K_r7_reg[53]/NET0131 ,
		_w28842_
	);
	LUT4 #(
		.INIT('hc693)
	) name23016 (
		decrypt_pad,
		\u0_R7_reg[5]/NET0131 ,
		\u0_uk_K_r7_reg[40]/NET0131 ,
		\u0_uk_K_r7_reg[47]/NET0131 ,
		_w28843_
	);
	LUT4 #(
		.INIT('hc693)
	) name23017 (
		decrypt_pad,
		\u0_R7_reg[7]/NET0131 ,
		\u0_uk_K_r7_reg[25]/NET0131 ,
		\u0_uk_K_r7_reg[32]/NET0131 ,
		_w28844_
	);
	LUT4 #(
		.INIT('h0004)
	) name23018 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28844_,
		_w28845_
	);
	LUT4 #(
		.INIT('hc963)
	) name23019 (
		decrypt_pad,
		\u0_R7_reg[4]/NET0131 ,
		\u0_uk_K_r7_reg[11]/NET0131 ,
		\u0_uk_K_r7_reg[4]/NET0131 ,
		_w28846_
	);
	LUT2 #(
		.INIT('h2)
	) name23020 (
		_w28842_,
		_w28846_,
		_w28847_
	);
	LUT3 #(
		.INIT('h08)
	) name23021 (
		_w28842_,
		_w28843_,
		_w28846_,
		_w28848_
	);
	LUT4 #(
		.INIT('h0080)
	) name23022 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28849_
	);
	LUT2 #(
		.INIT('h1)
	) name23023 (
		_w28845_,
		_w28849_,
		_w28850_
	);
	LUT4 #(
		.INIT('h0800)
	) name23024 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28851_
	);
	LUT4 #(
		.INIT('h0103)
	) name23025 (
		_w28844_,
		_w28845_,
		_w28849_,
		_w28851_,
		_w28852_
	);
	LUT2 #(
		.INIT('h8)
	) name23026 (
		_w28842_,
		_w28846_,
		_w28853_
	);
	LUT4 #(
		.INIT('h1014)
	) name23027 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28854_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name23028 (
		_w28842_,
		_w28843_,
		_w28844_,
		_w28846_,
		_w28855_
	);
	LUT4 #(
		.INIT('h51f3)
	) name23029 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28856_
	);
	LUT3 #(
		.INIT('h51)
	) name23030 (
		_w28854_,
		_w28855_,
		_w28856_,
		_w28857_
	);
	LUT3 #(
		.INIT('h15)
	) name23031 (
		_w28840_,
		_w28852_,
		_w28857_,
		_w28858_
	);
	LUT4 #(
		.INIT('hf7cc)
	) name23032 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28859_
	);
	LUT4 #(
		.INIT('h00c4)
	) name23033 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28860_
	);
	LUT3 #(
		.INIT('h0b)
	) name23034 (
		_w28841_,
		_w28843_,
		_w28844_,
		_w28861_
	);
	LUT4 #(
		.INIT('hf200)
	) name23035 (
		_w28840_,
		_w28859_,
		_w28860_,
		_w28861_,
		_w28862_
	);
	LUT4 #(
		.INIT('h0002)
	) name23036 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28863_
	);
	LUT4 #(
		.INIT('haffd)
	) name23037 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28864_
	);
	LUT2 #(
		.INIT('h2)
	) name23038 (
		_w28844_,
		_w28864_,
		_w28865_
	);
	LUT4 #(
		.INIT('h0100)
	) name23039 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28866_
	);
	LUT4 #(
		.INIT('hc040)
	) name23040 (
		_w28841_,
		_w28843_,
		_w28844_,
		_w28846_,
		_w28867_
	);
	LUT4 #(
		.INIT('h4000)
	) name23041 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28868_
	);
	LUT4 #(
		.INIT('haaa8)
	) name23042 (
		_w28840_,
		_w28866_,
		_w28867_,
		_w28868_,
		_w28869_
	);
	LUT3 #(
		.INIT('h01)
	) name23043 (
		_w28865_,
		_w28869_,
		_w28862_,
		_w28870_
	);
	LUT3 #(
		.INIT('h65)
	) name23044 (
		\u0_L7_reg[2]/NET0131 ,
		_w28858_,
		_w28870_,
		_w28871_
	);
	LUT4 #(
		.INIT('h0282)
	) name23045 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28872_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name23046 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28873_
	);
	LUT4 #(
		.INIT('hd8fa)
	) name23047 (
		_w28705_,
		_w28727_,
		_w28872_,
		_w28873_,
		_w28874_
	);
	LUT4 #(
		.INIT('h2010)
	) name23048 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28875_
	);
	LUT3 #(
		.INIT('h02)
	) name23049 (
		_w28712_,
		_w28745_,
		_w28875_,
		_w28876_
	);
	LUT2 #(
		.INIT('h4)
	) name23050 (
		_w28874_,
		_w28876_,
		_w28877_
	);
	LUT2 #(
		.INIT('h2)
	) name23051 (
		_w28705_,
		_w28709_,
		_w28878_
	);
	LUT3 #(
		.INIT('h08)
	) name23052 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28879_
	);
	LUT2 #(
		.INIT('h4)
	) name23053 (
		_w28878_,
		_w28879_,
		_w28880_
	);
	LUT4 #(
		.INIT('h5040)
	) name23054 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28881_
	);
	LUT4 #(
		.INIT('h0100)
	) name23055 (
		_w28705_,
		_w28706_,
		_w28708_,
		_w28709_,
		_w28882_
	);
	LUT4 #(
		.INIT('h1011)
	) name23056 (
		_w28712_,
		_w28882_,
		_w28878_,
		_w28881_,
		_w28883_
	);
	LUT4 #(
		.INIT('h0021)
	) name23057 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28884_
	);
	LUT4 #(
		.INIT('hdd5f)
	) name23058 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w28885_
	);
	LUT3 #(
		.INIT('h31)
	) name23059 (
		_w28705_,
		_w28884_,
		_w28885_,
		_w28886_
	);
	LUT3 #(
		.INIT('h40)
	) name23060 (
		_w28880_,
		_w28883_,
		_w28886_,
		_w28887_
	);
	LUT2 #(
		.INIT('h4)
	) name23061 (
		_w28705_,
		_w28708_,
		_w28888_
	);
	LUT4 #(
		.INIT('h0002)
	) name23062 (
		_w28705_,
		_w28706_,
		_w28707_,
		_w28709_,
		_w28889_
	);
	LUT3 #(
		.INIT('h07)
	) name23063 (
		_w28735_,
		_w28888_,
		_w28889_,
		_w28890_
	);
	LUT4 #(
		.INIT('ha955)
	) name23064 (
		\u0_L7_reg[21]/NET0131 ,
		_w28877_,
		_w28887_,
		_w28890_,
		_w28891_
	);
	LUT4 #(
		.INIT('h9fcf)
	) name23065 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28892_
	);
	LUT2 #(
		.INIT('h2)
	) name23066 (
		_w28666_,
		_w28892_,
		_w28893_
	);
	LUT4 #(
		.INIT('h66fe)
	) name23067 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28894_
	);
	LUT2 #(
		.INIT('h1)
	) name23068 (
		_w28666_,
		_w28894_,
		_w28895_
	);
	LUT4 #(
		.INIT('hfefd)
	) name23069 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28896_
	);
	LUT3 #(
		.INIT('h10)
	) name23070 (
		_w28694_,
		_w28695_,
		_w28896_,
		_w28897_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name23071 (
		_w28673_,
		_w28893_,
		_w28895_,
		_w28897_,
		_w28898_
	);
	LUT4 #(
		.INIT('h697a)
	) name23072 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28899_
	);
	LUT4 #(
		.INIT('h0054)
	) name23073 (
		_w28673_,
		_w28666_,
		_w28789_,
		_w28899_,
		_w28900_
	);
	LUT4 #(
		.INIT('hbf47)
	) name23074 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w28901_
	);
	LUT2 #(
		.INIT('h1)
	) name23075 (
		_w28673_,
		_w28666_,
		_w28902_
	);
	LUT4 #(
		.INIT('h0080)
	) name23076 (
		_w28666_,
		_w28667_,
		_w28671_,
		_w28669_,
		_w28903_
	);
	LUT4 #(
		.INIT('h1011)
	) name23077 (
		_w28678_,
		_w28903_,
		_w28901_,
		_w28902_,
		_w28904_
	);
	LUT2 #(
		.INIT('h4)
	) name23078 (
		_w28900_,
		_w28904_,
		_w28905_
	);
	LUT3 #(
		.INIT('h9a)
	) name23079 (
		\u0_L7_reg[29]/NET0131 ,
		_w28898_,
		_w28905_,
		_w28906_
	);
	LUT4 #(
		.INIT('hc693)
	) name23080 (
		decrypt_pad,
		\u0_R7_reg[20]/NET0131 ,
		\u0_uk_K_r7_reg[28]/NET0131 ,
		\u0_uk_K_r7_reg[35]/NET0131 ,
		_w28907_
	);
	LUT4 #(
		.INIT('hc693)
	) name23081 (
		decrypt_pad,
		\u0_R7_reg[19]/NET0131 ,
		\u0_uk_K_r7_reg[44]/NET0131 ,
		\u0_uk_K_r7_reg[51]/NET0131 ,
		_w28908_
	);
	LUT4 #(
		.INIT('hc963)
	) name23082 (
		decrypt_pad,
		\u0_R7_reg[17]/NET0131 ,
		\u0_uk_K_r7_reg[15]/NET0131 ,
		\u0_uk_K_r7_reg[8]/NET0131 ,
		_w28909_
	);
	LUT4 #(
		.INIT('hc693)
	) name23083 (
		decrypt_pad,
		\u0_R7_reg[16]/NET0131 ,
		\u0_uk_K_r7_reg[45]/NET0131 ,
		\u0_uk_K_r7_reg[52]/NET0131 ,
		_w28910_
	);
	LUT4 #(
		.INIT('hc693)
	) name23084 (
		decrypt_pad,
		\u0_R7_reg[21]/NET0131 ,
		\u0_uk_K_r7_reg[29]/NET0131 ,
		\u0_uk_K_r7_reg[36]/NET0131 ,
		_w28911_
	);
	LUT2 #(
		.INIT('h2)
	) name23085 (
		_w28910_,
		_w28911_,
		_w28912_
	);
	LUT4 #(
		.INIT('hc693)
	) name23086 (
		decrypt_pad,
		\u0_R7_reg[18]/NET0131 ,
		\u0_uk_K_r7_reg[2]/NET0131 ,
		\u0_uk_K_r7_reg[9]/NET0131 ,
		_w28913_
	);
	LUT4 #(
		.INIT('h938f)
	) name23087 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28914_
	);
	LUT2 #(
		.INIT('h2)
	) name23088 (
		_w28908_,
		_w28914_,
		_w28915_
	);
	LUT3 #(
		.INIT('hbe)
	) name23089 (
		_w28910_,
		_w28911_,
		_w28909_,
		_w28916_
	);
	LUT2 #(
		.INIT('h1)
	) name23090 (
		_w28913_,
		_w28908_,
		_w28917_
	);
	LUT2 #(
		.INIT('h4)
	) name23091 (
		_w28916_,
		_w28917_,
		_w28918_
	);
	LUT3 #(
		.INIT('h80)
	) name23092 (
		_w28910_,
		_w28911_,
		_w28909_,
		_w28919_
	);
	LUT2 #(
		.INIT('h2)
	) name23093 (
		_w28913_,
		_w28908_,
		_w28920_
	);
	LUT4 #(
		.INIT('h0400)
	) name23094 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28921_
	);
	LUT4 #(
		.INIT('h0008)
	) name23095 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28922_
	);
	LUT4 #(
		.INIT('hfbb7)
	) name23096 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28923_
	);
	LUT3 #(
		.INIT('h70)
	) name23097 (
		_w28919_,
		_w28920_,
		_w28923_,
		_w28924_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name23098 (
		_w28907_,
		_w28915_,
		_w28918_,
		_w28924_,
		_w28925_
	);
	LUT4 #(
		.INIT('h7f00)
	) name23099 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28908_,
		_w28926_
	);
	LUT4 #(
		.INIT('heefc)
	) name23100 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28927_
	);
	LUT2 #(
		.INIT('h8)
	) name23101 (
		_w28926_,
		_w28927_,
		_w28928_
	);
	LUT3 #(
		.INIT('h04)
	) name23102 (
		_w28910_,
		_w28911_,
		_w28909_,
		_w28929_
	);
	LUT4 #(
		.INIT('h00df)
	) name23103 (
		_w28913_,
		_w28911_,
		_w28909_,
		_w28908_,
		_w28930_
	);
	LUT4 #(
		.INIT('h0004)
	) name23104 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28931_
	);
	LUT4 #(
		.INIT('h4000)
	) name23105 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28932_
	);
	LUT4 #(
		.INIT('hbffb)
	) name23106 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28933_
	);
	LUT3 #(
		.INIT('h40)
	) name23107 (
		_w28929_,
		_w28930_,
		_w28933_,
		_w28934_
	);
	LUT4 #(
		.INIT('h0080)
	) name23108 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28935_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name23109 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28936_
	);
	LUT4 #(
		.INIT('h001f)
	) name23110 (
		_w28928_,
		_w28934_,
		_w28936_,
		_w28907_,
		_w28937_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name23111 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28938_
	);
	LUT4 #(
		.INIT('h0020)
	) name23112 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28939_
	);
	LUT4 #(
		.INIT('hfddf)
	) name23113 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28940_
	);
	LUT3 #(
		.INIT('hd8)
	) name23114 (
		_w28908_,
		_w28938_,
		_w28940_,
		_w28941_
	);
	LUT4 #(
		.INIT('h5655)
	) name23115 (
		\u0_L7_reg[14]/NET0131 ,
		_w28937_,
		_w28925_,
		_w28941_,
		_w28942_
	);
	LUT4 #(
		.INIT('hff2e)
	) name23116 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28943_
	);
	LUT3 #(
		.INIT('h02)
	) name23117 (
		_w28841_,
		_w28843_,
		_w28846_,
		_w28944_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name23118 (
		_w28841_,
		_w28843_,
		_w28844_,
		_w28846_,
		_w28945_
	);
	LUT4 #(
		.INIT('h0ef3)
	) name23119 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28946_
	);
	LUT4 #(
		.INIT('h7277)
	) name23120 (
		_w28844_,
		_w28943_,
		_w28944_,
		_w28946_,
		_w28947_
	);
	LUT4 #(
		.INIT('h0802)
	) name23121 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28948_
	);
	LUT4 #(
		.INIT('h2000)
	) name23122 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28949_
	);
	LUT3 #(
		.INIT('h01)
	) name23123 (
		_w28840_,
		_w28949_,
		_w28948_,
		_w28950_
	);
	LUT2 #(
		.INIT('h4)
	) name23124 (
		_w28947_,
		_w28950_,
		_w28951_
	);
	LUT3 #(
		.INIT('h90)
	) name23125 (
		_w28842_,
		_w28843_,
		_w28846_,
		_w28952_
	);
	LUT4 #(
		.INIT('h0020)
	) name23126 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28953_
	);
	LUT3 #(
		.INIT('h02)
	) name23127 (
		_w28844_,
		_w28953_,
		_w28952_,
		_w28954_
	);
	LUT4 #(
		.INIT('hdf2e)
	) name23128 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28955_
	);
	LUT2 #(
		.INIT('h8)
	) name23129 (
		_w28945_,
		_w28955_,
		_w28956_
	);
	LUT2 #(
		.INIT('h8)
	) name23130 (
		_w28844_,
		_w28846_,
		_w28957_
	);
	LUT4 #(
		.INIT('h0dff)
	) name23131 (
		_w28842_,
		_w28843_,
		_w28844_,
		_w28846_,
		_w28958_
	);
	LUT4 #(
		.INIT('h0008)
	) name23132 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w28959_
	);
	LUT4 #(
		.INIT('h00a8)
	) name23133 (
		_w28840_,
		_w28841_,
		_w28958_,
		_w28959_,
		_w28960_
	);
	LUT3 #(
		.INIT('he0)
	) name23134 (
		_w28954_,
		_w28956_,
		_w28960_,
		_w28961_
	);
	LUT3 #(
		.INIT('ha9)
	) name23135 (
		\u0_L7_reg[28]/NET0131 ,
		_w28951_,
		_w28961_,
		_w28962_
	);
	LUT2 #(
		.INIT('h1)
	) name23136 (
		_w28614_,
		_w28609_,
		_w28963_
	);
	LUT4 #(
		.INIT('h2030)
	) name23137 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28964_
	);
	LUT2 #(
		.INIT('h4)
	) name23138 (
		_w28963_,
		_w28964_,
		_w28965_
	);
	LUT4 #(
		.INIT('h0080)
	) name23139 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28966_
	);
	LUT3 #(
		.INIT('h01)
	) name23140 (
		_w28608_,
		_w28615_,
		_w28966_,
		_w28967_
	);
	LUT4 #(
		.INIT('h0104)
	) name23141 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28968_
	);
	LUT4 #(
		.INIT('h0770)
	) name23142 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28969_
	);
	LUT3 #(
		.INIT('h32)
	) name23143 (
		_w28609_,
		_w28968_,
		_w28969_,
		_w28970_
	);
	LUT3 #(
		.INIT('h40)
	) name23144 (
		_w28965_,
		_w28967_,
		_w28970_,
		_w28971_
	);
	LUT4 #(
		.INIT('h33fe)
	) name23145 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28972_
	);
	LUT2 #(
		.INIT('h2)
	) name23146 (
		_w28609_,
		_w28972_,
		_w28973_
	);
	LUT4 #(
		.INIT('hedb7)
	) name23147 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w28974_
	);
	LUT4 #(
		.INIT('h8a00)
	) name23148 (
		_w28608_,
		_w28609_,
		_w28625_,
		_w28974_,
		_w28975_
	);
	LUT2 #(
		.INIT('h4)
	) name23149 (
		_w28973_,
		_w28975_,
		_w28976_
	);
	LUT3 #(
		.INIT('ha9)
	) name23150 (
		\u0_L7_reg[12]/NET0131 ,
		_w28971_,
		_w28976_,
		_w28977_
	);
	LUT2 #(
		.INIT('h8)
	) name23151 (
		_w28753_,
		_w28757_,
		_w28978_
	);
	LUT4 #(
		.INIT('hafee)
	) name23152 (
		_w28755_,
		_w28754_,
		_w28757_,
		_w28752_,
		_w28979_
	);
	LUT2 #(
		.INIT('h1)
	) name23153 (
		_w28978_,
		_w28979_,
		_w28980_
	);
	LUT4 #(
		.INIT('h2220)
	) name23154 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28981_
	);
	LUT2 #(
		.INIT('h4)
	) name23155 (
		_w28761_,
		_w28981_,
		_w28982_
	);
	LUT3 #(
		.INIT('h0b)
	) name23156 (
		_w28774_,
		_w28764_,
		_w28814_,
		_w28983_
	);
	LUT4 #(
		.INIT('h5455)
	) name23157 (
		_w28766_,
		_w28980_,
		_w28982_,
		_w28983_,
		_w28984_
	);
	LUT4 #(
		.INIT('hef75)
	) name23158 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28985_
	);
	LUT4 #(
		.INIT('h0200)
	) name23159 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28986_
	);
	LUT4 #(
		.INIT('hfdaf)
	) name23160 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28987_
	);
	LUT4 #(
		.INIT('hc480)
	) name23161 (
		_w28757_,
		_w28815_,
		_w28987_,
		_w28985_,
		_w28988_
	);
	LUT4 #(
		.INIT('h0001)
	) name23162 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28989_
	);
	LUT4 #(
		.INIT('h7bfe)
	) name23163 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28752_,
		_w28990_
	);
	LUT2 #(
		.INIT('h1)
	) name23164 (
		_w28757_,
		_w28990_,
		_w28991_
	);
	LUT4 #(
		.INIT('h4000)
	) name23165 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28757_,
		_w28992_
	);
	LUT3 #(
		.INIT('h0b)
	) name23166 (
		_w28753_,
		_w28773_,
		_w28992_,
		_w28993_
	);
	LUT4 #(
		.INIT('h0d00)
	) name23167 (
		_w28766_,
		_w28988_,
		_w28991_,
		_w28993_,
		_w28994_
	);
	LUT3 #(
		.INIT('h65)
	) name23168 (
		\u0_L7_reg[10]/NET0131 ,
		_w28984_,
		_w28994_,
		_w28995_
	);
	LUT4 #(
		.INIT('h3dc8)
	) name23169 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28996_
	);
	LUT4 #(
		.INIT('hee3f)
	) name23170 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28997_
	);
	LUT4 #(
		.INIT('ha7ff)
	) name23171 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w28998_
	);
	LUT4 #(
		.INIT('hd800)
	) name23172 (
		_w28908_,
		_w28996_,
		_w28997_,
		_w28998_,
		_w28999_
	);
	LUT2 #(
		.INIT('h2)
	) name23173 (
		_w28907_,
		_w28999_,
		_w29000_
	);
	LUT4 #(
		.INIT('hddf3)
	) name23174 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29001_
	);
	LUT2 #(
		.INIT('h1)
	) name23175 (
		_w28908_,
		_w29001_,
		_w29002_
	);
	LUT4 #(
		.INIT('h1000)
	) name23176 (
		_w28913_,
		_w28911_,
		_w28909_,
		_w28908_,
		_w29003_
	);
	LUT4 #(
		.INIT('h0001)
	) name23177 (
		_w28913_,
		_w28910_,
		_w28909_,
		_w28908_,
		_w29004_
	);
	LUT4 #(
		.INIT('h2000)
	) name23178 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29005_
	);
	LUT3 #(
		.INIT('h01)
	) name23179 (
		_w29004_,
		_w29005_,
		_w29003_,
		_w29006_
	);
	LUT4 #(
		.INIT('hf7ed)
	) name23180 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29007_
	);
	LUT4 #(
		.INIT('h0008)
	) name23181 (
		_w28913_,
		_w28910_,
		_w28909_,
		_w28908_,
		_w29008_
	);
	LUT4 #(
		.INIT('h0031)
	) name23182 (
		_w28908_,
		_w28932_,
		_w29007_,
		_w29008_,
		_w29009_
	);
	LUT4 #(
		.INIT('hba00)
	) name23183 (
		_w28907_,
		_w29002_,
		_w29006_,
		_w29009_,
		_w29010_
	);
	LUT3 #(
		.INIT('h65)
	) name23184 (
		\u0_L7_reg[25]/NET0131 ,
		_w29000_,
		_w29010_,
		_w29011_
	);
	LUT4 #(
		.INIT('h0401)
	) name23185 (
		_w28666_,
		_w28667_,
		_w28668_,
		_w28671_,
		_w29012_
	);
	LUT4 #(
		.INIT('h23e3)
	) name23186 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w29013_
	);
	LUT4 #(
		.INIT('h8000)
	) name23187 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w29014_
	);
	LUT4 #(
		.INIT('h0051)
	) name23188 (
		_w28673_,
		_w28666_,
		_w29013_,
		_w29014_,
		_w29015_
	);
	LUT3 #(
		.INIT('h04)
	) name23189 (
		_w28666_,
		_w28668_,
		_w28671_,
		_w29016_
	);
	LUT4 #(
		.INIT('haa8a)
	) name23190 (
		_w28673_,
		_w28667_,
		_w28671_,
		_w28669_,
		_w29017_
	);
	LUT3 #(
		.INIT('h10)
	) name23191 (
		_w28700_,
		_w29016_,
		_w29017_,
		_w29018_
	);
	LUT4 #(
		.INIT('hfd3d)
	) name23192 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w29019_
	);
	LUT4 #(
		.INIT('h2100)
	) name23193 (
		_w28667_,
		_w28668_,
		_w28671_,
		_w28669_,
		_w29020_
	);
	LUT3 #(
		.INIT('h0d)
	) name23194 (
		_w28666_,
		_w29019_,
		_w29020_,
		_w29021_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name23195 (
		_w29012_,
		_w29015_,
		_w29018_,
		_w29021_,
		_w29022_
	);
	LUT2 #(
		.INIT('h1)
	) name23196 (
		_w28687_,
		_w28701_,
		_w29023_
	);
	LUT3 #(
		.INIT('h65)
	) name23197 (
		\u0_L7_reg[19]/NET0131 ,
		_w29022_,
		_w29023_,
		_w29024_
	);
	LUT4 #(
		.INIT('hd3cc)
	) name23198 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w29025_
	);
	LUT2 #(
		.INIT('h2)
	) name23199 (
		_w28705_,
		_w29025_,
		_w29026_
	);
	LUT4 #(
		.INIT('h4000)
	) name23200 (
		_w28705_,
		_w28706_,
		_w28708_,
		_w28707_,
		_w29027_
	);
	LUT3 #(
		.INIT('h01)
	) name23201 (
		_w28715_,
		_w28882_,
		_w29027_,
		_w29028_
	);
	LUT3 #(
		.INIT('h45)
	) name23202 (
		_w28712_,
		_w29026_,
		_w29028_,
		_w29029_
	);
	LUT4 #(
		.INIT('h8900)
	) name23203 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w29030_
	);
	LUT3 #(
		.INIT('h60)
	) name23204 (
		_w28706_,
		_w28708_,
		_w28709_,
		_w29031_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name23205 (
		_w28705_,
		_w28713_,
		_w29030_,
		_w29031_,
		_w29032_
	);
	LUT4 #(
		.INIT('hbfd3)
	) name23206 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w29033_
	);
	LUT4 #(
		.INIT('h0020)
	) name23207 (
		_w28705_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w29034_
	);
	LUT4 #(
		.INIT('hedf7)
	) name23208 (
		_w28706_,
		_w28708_,
		_w28707_,
		_w28709_,
		_w29035_
	);
	LUT3 #(
		.INIT('h32)
	) name23209 (
		_w28705_,
		_w29034_,
		_w29035_,
		_w29036_
	);
	LUT4 #(
		.INIT('h7500)
	) name23210 (
		_w28712_,
		_w29032_,
		_w29033_,
		_w29036_,
		_w29037_
	);
	LUT3 #(
		.INIT('h65)
	) name23211 (
		\u0_L7_reg[27]/NET0131 ,
		_w29029_,
		_w29037_,
		_w29038_
	);
	LUT4 #(
		.INIT('hc1e6)
	) name23212 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w29039_
	);
	LUT2 #(
		.INIT('h1)
	) name23213 (
		_w28609_,
		_w29039_,
		_w29040_
	);
	LUT4 #(
		.INIT('h2800)
	) name23214 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w29041_
	);
	LUT4 #(
		.INIT('hd77f)
	) name23215 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w29042_
	);
	LUT3 #(
		.INIT('h41)
	) name23216 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w29043_
	);
	LUT4 #(
		.INIT('h4140)
	) name23217 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w29044_
	);
	LUT4 #(
		.INIT('h2a00)
	) name23218 (
		_w28608_,
		_w28609_,
		_w29044_,
		_w29042_,
		_w29045_
	);
	LUT4 #(
		.INIT('hf700)
	) name23219 (
		_w28611_,
		_w28613_,
		_w28614_,
		_w28609_,
		_w29046_
	);
	LUT4 #(
		.INIT('h5455)
	) name23220 (
		_w28608_,
		_w29043_,
		_w29041_,
		_w29046_,
		_w29047_
	);
	LUT3 #(
		.INIT('h0b)
	) name23221 (
		_w29040_,
		_w29045_,
		_w29047_,
		_w29048_
	);
	LUT2 #(
		.INIT('h1)
	) name23222 (
		_w28609_,
		_w29042_,
		_w29049_
	);
	LUT2 #(
		.INIT('h2)
	) name23223 (
		_w28608_,
		_w28609_,
		_w29050_
	);
	LUT4 #(
		.INIT('h00dc)
	) name23224 (
		_w28609_,
		_w28615_,
		_w29044_,
		_w29050_,
		_w29051_
	);
	LUT2 #(
		.INIT('h1)
	) name23225 (
		_w29049_,
		_w29051_,
		_w29052_
	);
	LUT3 #(
		.INIT('h65)
	) name23226 (
		\u0_L7_reg[7]/NET0131 ,
		_w29048_,
		_w29052_,
		_w29053_
	);
	LUT3 #(
		.INIT('h02)
	) name23227 (
		_w28908_,
		_w28931_,
		_w28919_,
		_w29054_
	);
	LUT4 #(
		.INIT('h3010)
	) name23228 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29055_
	);
	LUT4 #(
		.INIT('h00f7)
	) name23229 (
		_w28910_,
		_w28911_,
		_w28909_,
		_w28908_,
		_w29056_
	);
	LUT2 #(
		.INIT('h4)
	) name23230 (
		_w29055_,
		_w29056_,
		_w29057_
	);
	LUT4 #(
		.INIT('he6fd)
	) name23231 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29058_
	);
	LUT4 #(
		.INIT('h0155)
	) name23232 (
		_w28907_,
		_w29054_,
		_w29057_,
		_w29058_,
		_w29059_
	);
	LUT4 #(
		.INIT('h0001)
	) name23233 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29060_
	);
	LUT4 #(
		.INIT('hff3e)
	) name23234 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29061_
	);
	LUT3 #(
		.INIT('h04)
	) name23235 (
		_w28913_,
		_w28910_,
		_w28908_,
		_w29062_
	);
	LUT4 #(
		.INIT('h00c4)
	) name23236 (
		_w28908_,
		_w28940_,
		_w29061_,
		_w29062_,
		_w29063_
	);
	LUT4 #(
		.INIT('he5df)
	) name23237 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29064_
	);
	LUT4 #(
		.INIT('haf23)
	) name23238 (
		_w28911_,
		_w28908_,
		_w29008_,
		_w29064_,
		_w29065_
	);
	LUT3 #(
		.INIT('hd0)
	) name23239 (
		_w28907_,
		_w29063_,
		_w29065_,
		_w29066_
	);
	LUT3 #(
		.INIT('h65)
	) name23240 (
		\u0_L7_reg[8]/NET0131 ,
		_w29059_,
		_w29066_,
		_w29067_
	);
	LUT4 #(
		.INIT('hbf00)
	) name23241 (
		_w28610_,
		_w28613_,
		_w28614_,
		_w28609_,
		_w29068_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name23242 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w29069_
	);
	LUT2 #(
		.INIT('h8)
	) name23243 (
		_w29068_,
		_w29069_,
		_w29070_
	);
	LUT4 #(
		.INIT('h0014)
	) name23244 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w29071_
	);
	LUT4 #(
		.INIT('h00ef)
	) name23245 (
		_w28611_,
		_w28613_,
		_w28614_,
		_w28609_,
		_w29072_
	);
	LUT3 #(
		.INIT('h10)
	) name23246 (
		_w28966_,
		_w29071_,
		_w29072_,
		_w29073_
	);
	LUT2 #(
		.INIT('h2)
	) name23247 (
		_w28610_,
		_w28613_,
		_w29074_
	);
	LUT4 #(
		.INIT('h0800)
	) name23248 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w29075_
	);
	LUT4 #(
		.INIT('haa02)
	) name23249 (
		_w28608_,
		_w29070_,
		_w29073_,
		_w29075_,
		_w29076_
	);
	LUT4 #(
		.INIT('h6200)
	) name23250 (
		_w28610_,
		_w28611_,
		_w28613_,
		_w28614_,
		_w29077_
	);
	LUT2 #(
		.INIT('h6)
	) name23251 (
		_w28613_,
		_w28614_,
		_w29078_
	);
	LUT4 #(
		.INIT('h5545)
	) name23252 (
		_w28608_,
		_w28610_,
		_w28611_,
		_w28614_,
		_w29079_
	);
	LUT4 #(
		.INIT('h4544)
	) name23253 (
		_w28609_,
		_w29077_,
		_w29078_,
		_w29079_,
		_w29080_
	);
	LUT2 #(
		.INIT('h2)
	) name23254 (
		_w28625_,
		_w29050_,
		_w29081_
	);
	LUT3 #(
		.INIT('ha8)
	) name23255 (
		_w28611_,
		_w28614_,
		_w28609_,
		_w29082_
	);
	LUT4 #(
		.INIT('h5455)
	) name23256 (
		_w28624_,
		_w28628_,
		_w29074_,
		_w29082_,
		_w29083_
	);
	LUT4 #(
		.INIT('h0032)
	) name23257 (
		_w28608_,
		_w29081_,
		_w29083_,
		_w29080_,
		_w29084_
	);
	LUT3 #(
		.INIT('h65)
	) name23258 (
		\u0_L7_reg[32]/NET0131 ,
		_w29076_,
		_w29084_,
		_w29085_
	);
	LUT4 #(
		.INIT('h007e)
	) name23259 (
		_w28639_,
		_w28641_,
		_w28636_,
		_w28643_,
		_w29086_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name23260 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w29087_
	);
	LUT2 #(
		.INIT('h2)
	) name23261 (
		_w29086_,
		_w29087_,
		_w29088_
	);
	LUT3 #(
		.INIT('h07)
	) name23262 (
		_w28661_,
		_w28662_,
		_w28830_,
		_w29089_
	);
	LUT4 #(
		.INIT('h0008)
	) name23263 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w29090_
	);
	LUT4 #(
		.INIT('heb00)
	) name23264 (
		_w28635_,
		_w28641_,
		_w28636_,
		_w28643_,
		_w29091_
	);
	LUT2 #(
		.INIT('h4)
	) name23265 (
		_w29090_,
		_w29091_,
		_w29092_
	);
	LUT4 #(
		.INIT('h8100)
	) name23266 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w29093_
	);
	LUT3 #(
		.INIT('h01)
	) name23267 (
		_w28638_,
		_w28833_,
		_w29093_,
		_w29094_
	);
	LUT4 #(
		.INIT('hea00)
	) name23268 (
		_w29088_,
		_w29089_,
		_w29092_,
		_w29094_,
		_w29095_
	);
	LUT4 #(
		.INIT('hbf00)
	) name23269 (
		_w28635_,
		_w28641_,
		_w28636_,
		_w28643_,
		_w29096_
	);
	LUT2 #(
		.INIT('h4)
	) name23270 (
		_w28827_,
		_w29096_,
		_w29097_
	);
	LUT4 #(
		.INIT('hddcf)
	) name23271 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w29098_
	);
	LUT2 #(
		.INIT('h8)
	) name23272 (
		_w29086_,
		_w29098_,
		_w29099_
	);
	LUT4 #(
		.INIT('h0414)
	) name23273 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w29100_
	);
	LUT2 #(
		.INIT('h2)
	) name23274 (
		_w28638_,
		_w29100_,
		_w29101_
	);
	LUT4 #(
		.INIT('hf800)
	) name23275 (
		_w29089_,
		_w29097_,
		_w29099_,
		_w29101_,
		_w29102_
	);
	LUT3 #(
		.INIT('h56)
	) name23276 (
		\u0_L7_reg[23]/NET0131 ,
		_w29095_,
		_w29102_,
		_w29103_
	);
	LUT4 #(
		.INIT('h9fff)
	) name23277 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w29104_
	);
	LUT4 #(
		.INIT('hfec7)
	) name23278 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w29105_
	);
	LUT4 #(
		.INIT('h0313)
	) name23279 (
		_w28840_,
		_w28844_,
		_w29104_,
		_w29105_,
		_w29106_
	);
	LUT3 #(
		.INIT('h12)
	) name23280 (
		_w28842_,
		_w28843_,
		_w28846_,
		_w29107_
	);
	LUT4 #(
		.INIT('he0f0)
	) name23281 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w29108_
	);
	LUT3 #(
		.INIT('h02)
	) name23282 (
		_w28844_,
		_w29108_,
		_w29107_,
		_w29109_
	);
	LUT3 #(
		.INIT('h54)
	) name23283 (
		_w28841_,
		_w28843_,
		_w28844_,
		_w29110_
	);
	LUT2 #(
		.INIT('h8)
	) name23284 (
		_w28847_,
		_w29110_,
		_w29111_
	);
	LUT3 #(
		.INIT('h8a)
	) name23285 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w29112_
	);
	LUT3 #(
		.INIT('h15)
	) name23286 (
		_w28840_,
		_w28957_,
		_w29112_,
		_w29113_
	);
	LUT3 #(
		.INIT('h10)
	) name23287 (
		_w29111_,
		_w29109_,
		_w29113_,
		_w29114_
	);
	LUT3 #(
		.INIT('h02)
	) name23288 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w29115_
	);
	LUT3 #(
		.INIT('h08)
	) name23289 (
		_w28841_,
		_w28842_,
		_w28846_,
		_w29116_
	);
	LUT4 #(
		.INIT('hfe00)
	) name23290 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28844_,
		_w29117_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name23291 (
		_w28855_,
		_w29115_,
		_w29116_,
		_w29117_,
		_w29118_
	);
	LUT4 #(
		.INIT('h0010)
	) name23292 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w29119_
	);
	LUT3 #(
		.INIT('h08)
	) name23293 (
		_w28840_,
		_w29104_,
		_w29119_,
		_w29120_
	);
	LUT3 #(
		.INIT('h20)
	) name23294 (
		_w28850_,
		_w29118_,
		_w29120_,
		_w29121_
	);
	LUT4 #(
		.INIT('h999a)
	) name23295 (
		\u0_L7_reg[13]/NET0131 ,
		_w29106_,
		_w29114_,
		_w29121_,
		_w29122_
	);
	LUT4 #(
		.INIT('hc693)
	) name23296 (
		decrypt_pad,
		\u0_R7_reg[11]/P0001 ,
		\u0_uk_K_r7_reg[11]/NET0131 ,
		\u0_uk_K_r7_reg[18]/NET0131 ,
		_w29123_
	);
	LUT4 #(
		.INIT('hc693)
	) name23297 (
		decrypt_pad,
		\u0_R7_reg[12]/NET0131 ,
		\u0_uk_K_r7_reg[26]/P0001 ,
		\u0_uk_K_r7_reg[33]/NET0131 ,
		_w29124_
	);
	LUT4 #(
		.INIT('hc693)
	) name23298 (
		decrypt_pad,
		\u0_R7_reg[13]/NET0131 ,
		\u0_uk_K_r7_reg[39]/NET0131 ,
		\u0_uk_K_r7_reg[46]/NET0131 ,
		_w29125_
	);
	LUT4 #(
		.INIT('hc693)
	) name23299 (
		decrypt_pad,
		\u0_R7_reg[9]/NET0131 ,
		\u0_uk_K_r7_reg[34]/NET0131 ,
		\u0_uk_K_r7_reg[41]/NET0131 ,
		_w29126_
	);
	LUT4 #(
		.INIT('hc693)
	) name23300 (
		decrypt_pad,
		\u0_R7_reg[10]/NET0131 ,
		\u0_uk_K_r7_reg[10]/NET0131 ,
		\u0_uk_K_r7_reg[17]/NET0131 ,
		_w29127_
	);
	LUT4 #(
		.INIT('hc963)
	) name23301 (
		decrypt_pad,
		\u0_R7_reg[8]/NET0131 ,
		\u0_uk_K_r7_reg[12]/NET0131 ,
		\u0_uk_K_r7_reg[5]/NET0131 ,
		_w29128_
	);
	LUT2 #(
		.INIT('h2)
	) name23302 (
		_w29125_,
		_w29128_,
		_w29129_
	);
	LUT4 #(
		.INIT('h95b5)
	) name23303 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29130_
	);
	LUT2 #(
		.INIT('h1)
	) name23304 (
		_w29125_,
		_w29128_,
		_w29131_
	);
	LUT4 #(
		.INIT('h0001)
	) name23305 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29132_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name23306 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29133_
	);
	LUT4 #(
		.INIT('h08cc)
	) name23307 (
		_w29124_,
		_w29123_,
		_w29130_,
		_w29133_,
		_w29134_
	);
	LUT2 #(
		.INIT('h6)
	) name23308 (
		_w29126_,
		_w29127_,
		_w29135_
	);
	LUT2 #(
		.INIT('h8)
	) name23309 (
		_w29125_,
		_w29128_,
		_w29136_
	);
	LUT3 #(
		.INIT('h46)
	) name23310 (
		_w29125_,
		_w29128_,
		_w29123_,
		_w29137_
	);
	LUT2 #(
		.INIT('h1)
	) name23311 (
		_w29135_,
		_w29137_,
		_w29138_
	);
	LUT3 #(
		.INIT('h40)
	) name23312 (
		_w29128_,
		_w29126_,
		_w29123_,
		_w29139_
	);
	LUT4 #(
		.INIT('h0660)
	) name23313 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29140_
	);
	LUT3 #(
		.INIT('h45)
	) name23314 (
		_w29124_,
		_w29139_,
		_w29140_,
		_w29141_
	);
	LUT3 #(
		.INIT('h80)
	) name23315 (
		_w29126_,
		_w29127_,
		_w29124_,
		_w29142_
	);
	LUT3 #(
		.INIT('h51)
	) name23316 (
		_w29128_,
		_w29126_,
		_w29127_,
		_w29143_
	);
	LUT4 #(
		.INIT('h0090)
	) name23317 (
		_w29125_,
		_w29126_,
		_w29124_,
		_w29123_,
		_w29144_
	);
	LUT4 #(
		.INIT('h7077)
	) name23318 (
		_w29131_,
		_w29142_,
		_w29143_,
		_w29144_,
		_w29145_
	);
	LUT4 #(
		.INIT('h4500)
	) name23319 (
		_w29134_,
		_w29138_,
		_w29141_,
		_w29145_,
		_w29146_
	);
	LUT2 #(
		.INIT('h9)
	) name23320 (
		\u0_L7_reg[6]/NET0131 ,
		_w29146_,
		_w29147_
	);
	LUT3 #(
		.INIT('h01)
	) name23321 (
		_w29126_,
		_w29127_,
		_w29123_,
		_w29148_
	);
	LUT4 #(
		.INIT('h000d)
	) name23322 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29149_
	);
	LUT3 #(
		.INIT('h09)
	) name23323 (
		_w29125_,
		_w29128_,
		_w29123_,
		_w29150_
	);
	LUT3 #(
		.INIT('h54)
	) name23324 (
		_w29148_,
		_w29149_,
		_w29150_,
		_w29151_
	);
	LUT4 #(
		.INIT('h1dff)
	) name23325 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29152_
	);
	LUT2 #(
		.INIT('h2)
	) name23326 (
		_w29123_,
		_w29152_,
		_w29153_
	);
	LUT4 #(
		.INIT('h0004)
	) name23327 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29154_
	);
	LUT3 #(
		.INIT('h07)
	) name23328 (
		_w29129_,
		_w29148_,
		_w29154_,
		_w29155_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name23329 (
		_w29124_,
		_w29153_,
		_w29151_,
		_w29155_,
		_w29156_
	);
	LUT3 #(
		.INIT('h20)
	) name23330 (
		_w29128_,
		_w29126_,
		_w29127_,
		_w29157_
	);
	LUT4 #(
		.INIT('h0400)
	) name23331 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29158_
	);
	LUT3 #(
		.INIT('h10)
	) name23332 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29159_
	);
	LUT4 #(
		.INIT('he2cd)
	) name23333 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29160_
	);
	LUT4 #(
		.INIT('h5054)
	) name23334 (
		_w29124_,
		_w29123_,
		_w29158_,
		_w29160_,
		_w29161_
	);
	LUT4 #(
		.INIT('h0009)
	) name23335 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29162_
	);
	LUT4 #(
		.INIT('h9db6)
	) name23336 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29163_
	);
	LUT2 #(
		.INIT('h1)
	) name23337 (
		_w29124_,
		_w29123_,
		_w29164_
	);
	LUT2 #(
		.INIT('h4)
	) name23338 (
		_w29163_,
		_w29164_,
		_w29165_
	);
	LUT4 #(
		.INIT('hffdb)
	) name23339 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29166_
	);
	LUT3 #(
		.INIT('h80)
	) name23340 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29167_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name23341 (
		_w29127_,
		_w29123_,
		_w29166_,
		_w29167_,
		_w29168_
	);
	LUT3 #(
		.INIT('h10)
	) name23342 (
		_w29161_,
		_w29165_,
		_w29168_,
		_w29169_
	);
	LUT3 #(
		.INIT('h65)
	) name23343 (
		\u0_L7_reg[24]/NET0131 ,
		_w29156_,
		_w29169_,
		_w29170_
	);
	LUT4 #(
		.INIT('hf04f)
	) name23344 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w29171_
	);
	LUT2 #(
		.INIT('h2)
	) name23345 (
		_w28638_,
		_w29171_,
		_w29172_
	);
	LUT4 #(
		.INIT('h4802)
	) name23346 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w29173_
	);
	LUT3 #(
		.INIT('h43)
	) name23347 (
		_w28635_,
		_w28641_,
		_w28636_,
		_w29174_
	);
	LUT4 #(
		.INIT('h1005)
	) name23348 (
		_w28638_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w29175_
	);
	LUT3 #(
		.INIT('h01)
	) name23349 (
		_w28643_,
		_w29175_,
		_w29173_,
		_w29176_
	);
	LUT4 #(
		.INIT('h8228)
	) name23350 (
		_w28639_,
		_w28635_,
		_w28641_,
		_w28636_,
		_w29177_
	);
	LUT4 #(
		.INIT('h040c)
	) name23351 (
		_w28640_,
		_w28643_,
		_w28833_,
		_w29174_,
		_w29178_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name23352 (
		_w29172_,
		_w29176_,
		_w29177_,
		_w29178_,
		_w29179_
	);
	LUT3 #(
		.INIT('h40)
	) name23353 (
		_w28638_,
		_w28641_,
		_w28636_,
		_w29180_
	);
	LUT2 #(
		.INIT('h4)
	) name23354 (
		_w28656_,
		_w29180_,
		_w29181_
	);
	LUT3 #(
		.INIT('h56)
	) name23355 (
		\u0_L7_reg[9]/NET0131 ,
		_w29179_,
		_w29181_,
		_w29182_
	);
	LUT4 #(
		.INIT('hed00)
	) name23356 (
		_w29125_,
		_w29128_,
		_w29127_,
		_w29123_,
		_w29183_
	);
	LUT3 #(
		.INIT('h07)
	) name23357 (
		_w29128_,
		_w29127_,
		_w29123_,
		_w29184_
	);
	LUT4 #(
		.INIT('h8acf)
	) name23358 (
		_w29159_,
		_w29154_,
		_w29183_,
		_w29184_,
		_w29185_
	);
	LUT2 #(
		.INIT('h2)
	) name23359 (
		_w29124_,
		_w29185_,
		_w29186_
	);
	LUT3 #(
		.INIT('h04)
	) name23360 (
		_w29125_,
		_w29126_,
		_w29127_,
		_w29187_
	);
	LUT4 #(
		.INIT('h8c00)
	) name23361 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29188_
	);
	LUT3 #(
		.INIT('h02)
	) name23362 (
		_w29123_,
		_w29188_,
		_w29187_,
		_w29189_
	);
	LUT4 #(
		.INIT('h008c)
	) name23363 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29190_
	);
	LUT3 #(
		.INIT('h20)
	) name23364 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29191_
	);
	LUT4 #(
		.INIT('h00df)
	) name23365 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29123_,
		_w29192_
	);
	LUT2 #(
		.INIT('h4)
	) name23366 (
		_w29190_,
		_w29192_,
		_w29193_
	);
	LUT4 #(
		.INIT('h0200)
	) name23367 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29194_
	);
	LUT3 #(
		.INIT('h01)
	) name23368 (
		_w29124_,
		_w29162_,
		_w29194_,
		_w29195_
	);
	LUT3 #(
		.INIT('he0)
	) name23369 (
		_w29189_,
		_w29193_,
		_w29195_,
		_w29196_
	);
	LUT2 #(
		.INIT('h8)
	) name23370 (
		_w29125_,
		_w29123_,
		_w29197_
	);
	LUT2 #(
		.INIT('h8)
	) name23371 (
		_w29157_,
		_w29197_,
		_w29198_
	);
	LUT4 #(
		.INIT('h0040)
	) name23372 (
		_w29125_,
		_w29126_,
		_w29127_,
		_w29123_,
		_w29199_
	);
	LUT3 #(
		.INIT('h0d)
	) name23373 (
		_w29142_,
		_w29136_,
		_w29199_,
		_w29200_
	);
	LUT2 #(
		.INIT('h4)
	) name23374 (
		_w29198_,
		_w29200_,
		_w29201_
	);
	LUT4 #(
		.INIT('h56aa)
	) name23375 (
		\u0_L7_reg[30]/NET0131 ,
		_w29186_,
		_w29196_,
		_w29201_,
		_w29202_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name23376 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29203_
	);
	LUT2 #(
		.INIT('h2)
	) name23377 (
		_w28908_,
		_w29203_,
		_w29204_
	);
	LUT4 #(
		.INIT('h0040)
	) name23378 (
		_w28910_,
		_w28911_,
		_w28909_,
		_w28908_,
		_w29205_
	);
	LUT4 #(
		.INIT('h0004)
	) name23379 (
		_w28932_,
		_w28907_,
		_w28922_,
		_w29205_,
		_w29206_
	);
	LUT4 #(
		.INIT('he3ef)
	) name23380 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29207_
	);
	LUT2 #(
		.INIT('h2)
	) name23381 (
		_w28908_,
		_w29207_,
		_w29208_
	);
	LUT4 #(
		.INIT('h5010)
	) name23382 (
		_w28913_,
		_w28910_,
		_w28911_,
		_w28909_,
		_w29209_
	);
	LUT3 #(
		.INIT('hd0)
	) name23383 (
		_w28913_,
		_w28909_,
		_w28908_,
		_w29210_
	);
	LUT4 #(
		.INIT('h5554)
	) name23384 (
		_w28907_,
		_w28912_,
		_w29210_,
		_w29209_,
		_w29211_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name23385 (
		_w29204_,
		_w29206_,
		_w29208_,
		_w29211_,
		_w29212_
	);
	LUT3 #(
		.INIT('h02)
	) name23386 (
		_w28908_,
		_w28931_,
		_w28939_,
		_w29213_
	);
	LUT4 #(
		.INIT('h0001)
	) name23387 (
		_w28908_,
		_w28935_,
		_w28921_,
		_w29060_,
		_w29214_
	);
	LUT2 #(
		.INIT('h1)
	) name23388 (
		_w29213_,
		_w29214_,
		_w29215_
	);
	LUT3 #(
		.INIT('h56)
	) name23389 (
		\u0_L7_reg[3]/NET0131 ,
		_w29212_,
		_w29215_,
		_w29216_
	);
	LUT4 #(
		.INIT('h6979)
	) name23390 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29123_,
		_w29217_
	);
	LUT4 #(
		.INIT('h0014)
	) name23391 (
		_w29125_,
		_w29128_,
		_w29127_,
		_w29123_,
		_w29218_
	);
	LUT4 #(
		.INIT('h0072)
	) name23392 (
		_w29127_,
		_w29191_,
		_w29217_,
		_w29218_,
		_w29219_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name23393 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29220_
	);
	LUT4 #(
		.INIT('h6800)
	) name23394 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29123_,
		_w29221_
	);
	LUT4 #(
		.INIT('h0032)
	) name23395 (
		_w29123_,
		_w29132_,
		_w29220_,
		_w29221_,
		_w29222_
	);
	LUT4 #(
		.INIT('hbeff)
	) name23396 (
		_w29125_,
		_w29128_,
		_w29126_,
		_w29127_,
		_w29223_
	);
	LUT4 #(
		.INIT('h0020)
	) name23397 (
		_w29128_,
		_w29126_,
		_w29127_,
		_w29123_,
		_w29224_
	);
	LUT3 #(
		.INIT('h0d)
	) name23398 (
		_w29123_,
		_w29223_,
		_w29224_,
		_w29225_
	);
	LUT4 #(
		.INIT('hd800)
	) name23399 (
		_w29124_,
		_w29219_,
		_w29222_,
		_w29225_,
		_w29226_
	);
	LUT2 #(
		.INIT('h9)
	) name23400 (
		\u0_L7_reg[16]/NET0131 ,
		_w29226_,
		_w29227_
	);
	LUT3 #(
		.INIT('h1d)
	) name23401 (
		_w28841_,
		_w28843_,
		_w28844_,
		_w29228_
	);
	LUT3 #(
		.INIT('h0b)
	) name23402 (
		_w28841_,
		_w28843_,
		_w28846_,
		_w29229_
	);
	LUT4 #(
		.INIT('hdefe)
	) name23403 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w28846_,
		_w29230_
	);
	LUT4 #(
		.INIT('h3500)
	) name23404 (
		_w28853_,
		_w29229_,
		_w29228_,
		_w29230_,
		_w29231_
	);
	LUT2 #(
		.INIT('h1)
	) name23405 (
		_w28840_,
		_w29231_,
		_w29232_
	);
	LUT4 #(
		.INIT('h4060)
	) name23406 (
		_w28842_,
		_w28843_,
		_w28844_,
		_w28846_,
		_w29233_
	);
	LUT3 #(
		.INIT('ha8)
	) name23407 (
		_w28840_,
		_w28863_,
		_w29233_,
		_w29234_
	);
	LUT3 #(
		.INIT('hb8)
	) name23408 (
		_w28841_,
		_w28842_,
		_w28843_,
		_w29235_
	);
	LUT2 #(
		.INIT('h8)
	) name23409 (
		_w28840_,
		_w28846_,
		_w29236_
	);
	LUT4 #(
		.INIT('h4544)
	) name23410 (
		_w28844_,
		_w28848_,
		_w29235_,
		_w29236_,
		_w29237_
	);
	LUT4 #(
		.INIT('h80b0)
	) name23411 (
		_w28841_,
		_w28842_,
		_w28844_,
		_w28846_,
		_w29238_
	);
	LUT2 #(
		.INIT('h4)
	) name23412 (
		_w29229_,
		_w29238_,
		_w29239_
	);
	LUT3 #(
		.INIT('h01)
	) name23413 (
		_w29237_,
		_w29234_,
		_w29239_,
		_w29240_
	);
	LUT3 #(
		.INIT('h65)
	) name23414 (
		\u0_L7_reg[18]/NET0131 ,
		_w29232_,
		_w29240_,
		_w29241_
	);
	LUT4 #(
		.INIT('hc963)
	) name23415 (
		decrypt_pad,
		\u0_R6_reg[4]/NET0131 ,
		\u0_uk_K_r6_reg[47]/NET0131 ,
		\u0_uk_K_r6_reg[54]/NET0131 ,
		_w29242_
	);
	LUT4 #(
		.INIT('hc963)
	) name23416 (
		decrypt_pad,
		\u0_R6_reg[3]/NET0131 ,
		\u0_uk_K_r6_reg[12]/NET0131 ,
		\u0_uk_K_r6_reg[19]/NET0131 ,
		_w29243_
	);
	LUT4 #(
		.INIT('hc963)
	) name23417 (
		decrypt_pad,
		\u0_R6_reg[5]/NET0131 ,
		\u0_uk_K_r6_reg[18]/NET0131 ,
		\u0_uk_K_r6_reg[25]/NET0131 ,
		_w29244_
	);
	LUT4 #(
		.INIT('hc963)
	) name23418 (
		decrypt_pad,
		\u0_R6_reg[1]/NET0131 ,
		\u0_uk_K_r6_reg[20]/NET0131 ,
		\u0_uk_K_r6_reg[27]/NET0131 ,
		_w29245_
	);
	LUT4 #(
		.INIT('hc963)
	) name23419 (
		decrypt_pad,
		\u0_R6_reg[32]/NET0131 ,
		\u0_uk_K_r6_reg[24]/NET0131 ,
		\u0_uk_K_r6_reg[6]/NET0131 ,
		_w29246_
	);
	LUT4 #(
		.INIT('hc693)
	) name23420 (
		decrypt_pad,
		\u0_R6_reg[2]/NET0131 ,
		\u0_uk_K_r6_reg[10]/NET0131 ,
		\u0_uk_K_r6_reg[3]/NET0131 ,
		_w29247_
	);
	LUT4 #(
		.INIT('hd8dd)
	) name23421 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29248_
	);
	LUT2 #(
		.INIT('h2)
	) name23422 (
		_w29243_,
		_w29248_,
		_w29249_
	);
	LUT4 #(
		.INIT('h2520)
	) name23423 (
		_w29245_,
		_w29243_,
		_w29246_,
		_w29247_,
		_w29250_
	);
	LUT2 #(
		.INIT('h1)
	) name23424 (
		_w29244_,
		_w29245_,
		_w29251_
	);
	LUT4 #(
		.INIT('h0010)
	) name23425 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29252_
	);
	LUT2 #(
		.INIT('h2)
	) name23426 (
		_w29244_,
		_w29246_,
		_w29253_
	);
	LUT2 #(
		.INIT('h2)
	) name23427 (
		_w29243_,
		_w29247_,
		_w29254_
	);
	LUT3 #(
		.INIT('ha2)
	) name23428 (
		_w29245_,
		_w29243_,
		_w29247_,
		_w29255_
	);
	LUT4 #(
		.INIT('h0051)
	) name23429 (
		_w29252_,
		_w29253_,
		_w29255_,
		_w29250_,
		_w29256_
	);
	LUT3 #(
		.INIT('h8a)
	) name23430 (
		_w29242_,
		_w29249_,
		_w29256_,
		_w29257_
	);
	LUT4 #(
		.INIT('h5dbb)
	) name23431 (
		_w29244_,
		_w29245_,
		_w29243_,
		_w29246_,
		_w29258_
	);
	LUT3 #(
		.INIT('h48)
	) name23432 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29259_
	);
	LUT4 #(
		.INIT('h74fc)
	) name23433 (
		_w29243_,
		_w29247_,
		_w29258_,
		_w29259_,
		_w29260_
	);
	LUT2 #(
		.INIT('h9)
	) name23434 (
		_w29246_,
		_w29247_,
		_w29261_
	);
	LUT4 #(
		.INIT('h001d)
	) name23435 (
		_w29244_,
		_w29245_,
		_w29247_,
		_w29242_,
		_w29262_
	);
	LUT4 #(
		.INIT('h7dbb)
	) name23436 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29263_
	);
	LUT4 #(
		.INIT('h4055)
	) name23437 (
		_w29243_,
		_w29261_,
		_w29262_,
		_w29263_,
		_w29264_
	);
	LUT2 #(
		.INIT('h2)
	) name23438 (
		_w29243_,
		_w29246_,
		_w29265_
	);
	LUT3 #(
		.INIT('h20)
	) name23439 (
		_w29243_,
		_w29246_,
		_w29247_,
		_w29266_
	);
	LUT4 #(
		.INIT('h0040)
	) name23440 (
		_w29245_,
		_w29243_,
		_w29246_,
		_w29247_,
		_w29267_
	);
	LUT3 #(
		.INIT('h07)
	) name23441 (
		_w29251_,
		_w29266_,
		_w29267_,
		_w29268_
	);
	LUT4 #(
		.INIT('h3200)
	) name23442 (
		_w29242_,
		_w29264_,
		_w29260_,
		_w29268_,
		_w29269_
	);
	LUT3 #(
		.INIT('h65)
	) name23443 (
		\u0_L6_reg[31]/NET0131 ,
		_w29257_,
		_w29269_,
		_w29270_
	);
	LUT4 #(
		.INIT('hc963)
	) name23444 (
		decrypt_pad,
		\u0_R6_reg[24]/NET0131 ,
		\u0_uk_K_r6_reg[16]/NET0131 ,
		\u0_uk_K_r6_reg[23]/P0001 ,
		_w29271_
	);
	LUT4 #(
		.INIT('hc963)
	) name23445 (
		decrypt_pad,
		\u0_R6_reg[23]/NET0131 ,
		\u0_uk_K_r6_reg[14]/NET0131 ,
		\u0_uk_K_r6_reg[21]/NET0131 ,
		_w29272_
	);
	LUT4 #(
		.INIT('hc963)
	) name23446 (
		decrypt_pad,
		\u0_R6_reg[21]/NET0131 ,
		\u0_uk_K_r6_reg[38]/NET0131 ,
		\u0_uk_K_r6_reg[45]/NET0131 ,
		_w29273_
	);
	LUT4 #(
		.INIT('hc693)
	) name23447 (
		decrypt_pad,
		\u0_R6_reg[20]/NET0131 ,
		\u0_uk_K_r6_reg[2]/NET0131 ,
		\u0_uk_K_r6_reg[50]/NET0131 ,
		_w29274_
	);
	LUT4 #(
		.INIT('hc963)
	) name23448 (
		decrypt_pad,
		\u0_R6_reg[22]/NET0131 ,
		\u0_uk_K_r6_reg[1]/NET0131 ,
		\u0_uk_K_r6_reg[8]/NET0131 ,
		_w29275_
	);
	LUT4 #(
		.INIT('hc963)
	) name23449 (
		decrypt_pad,
		\u0_R6_reg[25]/NET0131 ,
		\u0_uk_K_r6_reg[35]/NET0131 ,
		\u0_uk_K_r6_reg[42]/NET0131 ,
		_w29276_
	);
	LUT4 #(
		.INIT('h0004)
	) name23450 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29277_
	);
	LUT4 #(
		.INIT('h57db)
	) name23451 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29278_
	);
	LUT2 #(
		.INIT('h2)
	) name23452 (
		_w29272_,
		_w29278_,
		_w29279_
	);
	LUT2 #(
		.INIT('h1)
	) name23453 (
		_w29275_,
		_w29272_,
		_w29280_
	);
	LUT4 #(
		.INIT('h0020)
	) name23454 (
		_w29274_,
		_w29275_,
		_w29276_,
		_w29272_,
		_w29281_
	);
	LUT3 #(
		.INIT('h25)
	) name23455 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29282_
	);
	LUT4 #(
		.INIT('h005c)
	) name23456 (
		_w29274_,
		_w29275_,
		_w29276_,
		_w29272_,
		_w29283_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name23457 (
		_w29273_,
		_w29281_,
		_w29282_,
		_w29283_,
		_w29284_
	);
	LUT3 #(
		.INIT('h8a)
	) name23458 (
		_w29271_,
		_w29279_,
		_w29284_,
		_w29285_
	);
	LUT4 #(
		.INIT('h1000)
	) name23459 (
		_w29273_,
		_w29274_,
		_w29276_,
		_w29272_,
		_w29286_
	);
	LUT4 #(
		.INIT('h4000)
	) name23460 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29287_
	);
	LUT2 #(
		.INIT('h2)
	) name23461 (
		_w29274_,
		_w29276_,
		_w29288_
	);
	LUT3 #(
		.INIT('hdc)
	) name23462 (
		_w29273_,
		_w29275_,
		_w29272_,
		_w29289_
	);
	LUT4 #(
		.INIT('h0051)
	) name23463 (
		_w29287_,
		_w29288_,
		_w29289_,
		_w29286_,
		_w29290_
	);
	LUT4 #(
		.INIT('hbcd7)
	) name23464 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29272_,
		_w29291_
	);
	LUT3 #(
		.INIT('h15)
	) name23465 (
		_w29271_,
		_w29290_,
		_w29291_,
		_w29292_
	);
	LUT4 #(
		.INIT('heff7)
	) name23466 (
		_w29273_,
		_w29274_,
		_w29276_,
		_w29272_,
		_w29293_
	);
	LUT2 #(
		.INIT('h1)
	) name23467 (
		_w29275_,
		_w29293_,
		_w29294_
	);
	LUT4 #(
		.INIT('h31f5)
	) name23468 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29295_
	);
	LUT4 #(
		.INIT('hcd00)
	) name23469 (
		_w29274_,
		_w29275_,
		_w29276_,
		_w29272_,
		_w29296_
	);
	LUT3 #(
		.INIT('h01)
	) name23470 (
		_w29273_,
		_w29274_,
		_w29276_,
		_w29297_
	);
	LUT4 #(
		.INIT('h45cf)
	) name23471 (
		_w29280_,
		_w29295_,
		_w29296_,
		_w29297_,
		_w29298_
	);
	LUT2 #(
		.INIT('h4)
	) name23472 (
		_w29294_,
		_w29298_,
		_w29299_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name23473 (
		\u0_L6_reg[11]/NET0131 ,
		_w29292_,
		_w29285_,
		_w29299_,
		_w29300_
	);
	LUT4 #(
		.INIT('hc963)
	) name23474 (
		decrypt_pad,
		\u0_R6_reg[26]/NET0131 ,
		\u0_uk_K_r6_reg[31]/NET0131 ,
		\u0_uk_K_r6_reg[38]/NET0131 ,
		_w29301_
	);
	LUT4 #(
		.INIT('hc963)
	) name23475 (
		decrypt_pad,
		\u0_R6_reg[25]/NET0131 ,
		\u0_uk_K_r6_reg[42]/NET0131 ,
		\u0_uk_K_r6_reg[49]/NET0131 ,
		_w29302_
	);
	LUT4 #(
		.INIT('hc693)
	) name23476 (
		decrypt_pad,
		\u0_R6_reg[24]/NET0131 ,
		\u0_uk_K_r6_reg[14]/NET0131 ,
		\u0_uk_K_r6_reg[7]/NET0131 ,
		_w29303_
	);
	LUT4 #(
		.INIT('hc963)
	) name23477 (
		decrypt_pad,
		\u0_R6_reg[29]/NET0131 ,
		\u0_uk_K_r6_reg[15]/NET0131 ,
		\u0_uk_K_r6_reg[22]/NET0131 ,
		_w29304_
	);
	LUT2 #(
		.INIT('h4)
	) name23478 (
		_w29303_,
		_w29304_,
		_w29305_
	);
	LUT4 #(
		.INIT('h0200)
	) name23479 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29306_
	);
	LUT3 #(
		.INIT('h08)
	) name23480 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29307_
	);
	LUT4 #(
		.INIT('h0008)
	) name23481 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29308_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name23482 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29309_
	);
	LUT3 #(
		.INIT('h40)
	) name23483 (
		_w29301_,
		_w29302_,
		_w29304_,
		_w29310_
	);
	LUT4 #(
		.INIT('hc963)
	) name23484 (
		decrypt_pad,
		\u0_R6_reg[28]/NET0131 ,
		\u0_uk_K_r6_reg[23]/P0001 ,
		\u0_uk_K_r6_reg[30]/P0001 ,
		_w29311_
	);
	LUT4 #(
		.INIT('h9cfc)
	) name23485 (
		_w29301_,
		_w29302_,
		_w29304_,
		_w29311_,
		_w29312_
	);
	LUT4 #(
		.INIT('hc963)
	) name23486 (
		decrypt_pad,
		\u0_R6_reg[27]/NET0131 ,
		\u0_uk_K_r6_reg[36]/NET0131 ,
		\u0_uk_K_r6_reg[43]/NET0131 ,
		_w29313_
	);
	LUT4 #(
		.INIT('h3b00)
	) name23487 (
		_w29303_,
		_w29309_,
		_w29312_,
		_w29313_,
		_w29314_
	);
	LUT4 #(
		.INIT('hee72)
	) name23488 (
		_w29301_,
		_w29302_,
		_w29304_,
		_w29313_,
		_w29315_
	);
	LUT2 #(
		.INIT('h2)
	) name23489 (
		_w29303_,
		_w29315_,
		_w29316_
	);
	LUT4 #(
		.INIT('h0002)
	) name23490 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29317_
	);
	LUT2 #(
		.INIT('h6)
	) name23491 (
		_w29301_,
		_w29303_,
		_w29318_
	);
	LUT3 #(
		.INIT('h8c)
	) name23492 (
		_w29302_,
		_w29304_,
		_w29313_,
		_w29319_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name23493 (
		_w29313_,
		_w29317_,
		_w29318_,
		_w29319_,
		_w29320_
	);
	LUT3 #(
		.INIT('h45)
	) name23494 (
		_w29311_,
		_w29316_,
		_w29320_,
		_w29321_
	);
	LUT4 #(
		.INIT('h1000)
	) name23495 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29322_
	);
	LUT4 #(
		.INIT('he3ff)
	) name23496 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29323_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name23497 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29324_
	);
	LUT4 #(
		.INIT('h02aa)
	) name23498 (
		_w29311_,
		_w29313_,
		_w29323_,
		_w29324_,
		_w29325_
	);
	LUT4 #(
		.INIT('h0084)
	) name23499 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29313_,
		_w29326_
	);
	LUT4 #(
		.INIT('h0100)
	) name23500 (
		_w29301_,
		_w29302_,
		_w29304_,
		_w29313_,
		_w29327_
	);
	LUT2 #(
		.INIT('h1)
	) name23501 (
		_w29326_,
		_w29327_,
		_w29328_
	);
	LUT2 #(
		.INIT('h4)
	) name23502 (
		_w29325_,
		_w29328_,
		_w29329_
	);
	LUT4 #(
		.INIT('h5655)
	) name23503 (
		\u0_L6_reg[22]/NET0131 ,
		_w29314_,
		_w29321_,
		_w29329_,
		_w29330_
	);
	LUT4 #(
		.INIT('hc963)
	) name23504 (
		decrypt_pad,
		\u0_R6_reg[15]/NET0131 ,
		\u0_uk_K_r6_reg[41]/NET0131 ,
		\u0_uk_K_r6_reg[48]/NET0131 ,
		_w29331_
	);
	LUT4 #(
		.INIT('hc963)
	) name23505 (
		decrypt_pad,
		\u0_R6_reg[13]/NET0131 ,
		\u0_uk_K_r6_reg[32]/NET0131 ,
		\u0_uk_K_r6_reg[39]/NET0131 ,
		_w29332_
	);
	LUT4 #(
		.INIT('hc963)
	) name23506 (
		decrypt_pad,
		\u0_R6_reg[12]/NET0131 ,
		\u0_uk_K_r6_reg[13]/NET0131 ,
		\u0_uk_K_r6_reg[20]/NET0131 ,
		_w29333_
	);
	LUT4 #(
		.INIT('hc963)
	) name23507 (
		decrypt_pad,
		\u0_R6_reg[14]/NET0131 ,
		\u0_uk_K_r6_reg[33]/NET0131 ,
		\u0_uk_K_r6_reg[40]/NET0131 ,
		_w29334_
	);
	LUT4 #(
		.INIT('hc693)
	) name23508 (
		decrypt_pad,
		\u0_R6_reg[17]/NET0131 ,
		\u0_uk_K_r6_reg[4]/NET0131 ,
		\u0_uk_K_r6_reg[54]/NET0131 ,
		_w29335_
	);
	LUT3 #(
		.INIT('h01)
	) name23509 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29336_
	);
	LUT4 #(
		.INIT('h0001)
	) name23510 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29337_
	);
	LUT3 #(
		.INIT('h7e)
	) name23511 (
		_w29333_,
		_w29335_,
		_w29332_,
		_w29338_
	);
	LUT3 #(
		.INIT('h0e)
	) name23512 (
		_w29331_,
		_w29337_,
		_w29338_,
		_w29339_
	);
	LUT4 #(
		.INIT('h0200)
	) name23513 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29340_
	);
	LUT4 #(
		.INIT('hc963)
	) name23514 (
		decrypt_pad,
		\u0_R6_reg[16]/NET0131 ,
		\u0_uk_K_r6_reg[17]/NET0131 ,
		\u0_uk_K_r6_reg[24]/NET0131 ,
		_w29341_
	);
	LUT2 #(
		.INIT('h1)
	) name23515 (
		_w29340_,
		_w29341_,
		_w29342_
	);
	LUT4 #(
		.INIT('hf707)
	) name23516 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29343_
	);
	LUT4 #(
		.INIT('h0040)
	) name23517 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29344_
	);
	LUT2 #(
		.INIT('h8)
	) name23518 (
		_w29331_,
		_w29334_,
		_w29345_
	);
	LUT3 #(
		.INIT('h80)
	) name23519 (
		_w29331_,
		_w29334_,
		_w29332_,
		_w29346_
	);
	LUT4 #(
		.INIT('h0800)
	) name23520 (
		_w29331_,
		_w29334_,
		_w29333_,
		_w29332_,
		_w29347_
	);
	LUT4 #(
		.INIT('h0032)
	) name23521 (
		_w29331_,
		_w29344_,
		_w29343_,
		_w29347_,
		_w29348_
	);
	LUT3 #(
		.INIT('h40)
	) name23522 (
		_w29339_,
		_w29342_,
		_w29348_,
		_w29349_
	);
	LUT2 #(
		.INIT('h4)
	) name23523 (
		_w29333_,
		_w29335_,
		_w29350_
	);
	LUT4 #(
		.INIT('h0020)
	) name23524 (
		_w29331_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29351_
	);
	LUT4 #(
		.INIT('h1000)
	) name23525 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29352_
	);
	LUT3 #(
		.INIT('h02)
	) name23526 (
		_w29341_,
		_w29351_,
		_w29352_,
		_w29353_
	);
	LUT2 #(
		.INIT('h2)
	) name23527 (
		_w29334_,
		_w29333_,
		_w29354_
	);
	LUT3 #(
		.INIT('h01)
	) name23528 (
		_w29331_,
		_w29335_,
		_w29332_,
		_w29355_
	);
	LUT2 #(
		.INIT('h2)
	) name23529 (
		_w29333_,
		_w29332_,
		_w29356_
	);
	LUT4 #(
		.INIT('h0110)
	) name23530 (
		_w29331_,
		_w29334_,
		_w29333_,
		_w29332_,
		_w29357_
	);
	LUT3 #(
		.INIT('h07)
	) name23531 (
		_w29354_,
		_w29355_,
		_w29357_,
		_w29358_
	);
	LUT4 #(
		.INIT('h8000)
	) name23532 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29359_
	);
	LUT4 #(
		.INIT('h0800)
	) name23533 (
		_w29331_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29360_
	);
	LUT2 #(
		.INIT('h1)
	) name23534 (
		_w29359_,
		_w29360_,
		_w29361_
	);
	LUT3 #(
		.INIT('h80)
	) name23535 (
		_w29353_,
		_w29358_,
		_w29361_,
		_w29362_
	);
	LUT3 #(
		.INIT('h40)
	) name23536 (
		_w29333_,
		_w29335_,
		_w29332_,
		_w29363_
	);
	LUT4 #(
		.INIT('h0008)
	) name23537 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29364_
	);
	LUT4 #(
		.INIT('h0400)
	) name23538 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29365_
	);
	LUT4 #(
		.INIT('hfbf6)
	) name23539 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29366_
	);
	LUT4 #(
		.INIT('hef45)
	) name23540 (
		_w29331_,
		_w29334_,
		_w29363_,
		_w29366_,
		_w29367_
	);
	LUT4 #(
		.INIT('ha955)
	) name23541 (
		\u0_L6_reg[20]/NET0131 ,
		_w29349_,
		_w29362_,
		_w29367_,
		_w29368_
	);
	LUT4 #(
		.INIT('hc963)
	) name23542 (
		decrypt_pad,
		\u0_R6_reg[31]/P0001 ,
		\u0_uk_K_r6_reg[37]/NET0131 ,
		\u0_uk_K_r6_reg[44]/NET0131 ,
		_w29369_
	);
	LUT4 #(
		.INIT('hc693)
	) name23543 (
		decrypt_pad,
		\u0_R6_reg[30]/NET0131 ,
		\u0_uk_K_r6_reg[1]/NET0131 ,
		\u0_uk_K_r6_reg[49]/NET0131 ,
		_w29370_
	);
	LUT4 #(
		.INIT('hc963)
	) name23544 (
		decrypt_pad,
		\u0_R6_reg[28]/NET0131 ,
		\u0_uk_K_r6_reg[21]/NET0131 ,
		\u0_uk_K_r6_reg[28]/NET0131 ,
		_w29371_
	);
	LUT4 #(
		.INIT('hc693)
	) name23545 (
		decrypt_pad,
		\u0_R6_reg[29]/NET0131 ,
		\u0_uk_K_r6_reg[0]/NET0131 ,
		\u0_uk_K_r6_reg[52]/NET0131 ,
		_w29372_
	);
	LUT4 #(
		.INIT('hc693)
	) name23546 (
		decrypt_pad,
		\u0_R6_reg[1]/NET0131 ,
		\u0_uk_K_r6_reg[16]/NET0131 ,
		\u0_uk_K_r6_reg[9]/NET0131 ,
		_w29373_
	);
	LUT4 #(
		.INIT('h0040)
	) name23547 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29374_
	);
	LUT4 #(
		.INIT('hc963)
	) name23548 (
		decrypt_pad,
		\u0_R6_reg[32]/NET0131 ,
		\u0_uk_K_r6_reg[43]/NET0131 ,
		\u0_uk_K_r6_reg[50]/NET0131 ,
		_w29375_
	);
	LUT2 #(
		.INIT('h4)
	) name23549 (
		_w29370_,
		_w29371_,
		_w29376_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name23550 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29377_
	);
	LUT4 #(
		.INIT('h0200)
	) name23551 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29378_
	);
	LUT4 #(
		.INIT('hf9de)
	) name23552 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29379_
	);
	LUT4 #(
		.INIT('hfd00)
	) name23553 (
		_w29375_,
		_w29374_,
		_w29377_,
		_w29379_,
		_w29380_
	);
	LUT2 #(
		.INIT('h2)
	) name23554 (
		_w29369_,
		_w29380_,
		_w29381_
	);
	LUT4 #(
		.INIT('hfcf7)
	) name23555 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29382_
	);
	LUT2 #(
		.INIT('h4)
	) name23556 (
		_w29382_,
		_w29369_,
		_w29383_
	);
	LUT4 #(
		.INIT('h0fdd)
	) name23557 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29384_
	);
	LUT2 #(
		.INIT('h1)
	) name23558 (
		_w29369_,
		_w29384_,
		_w29385_
	);
	LUT4 #(
		.INIT('h8000)
	) name23559 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29386_
	);
	LUT3 #(
		.INIT('hd0)
	) name23560 (
		_w29372_,
		_w29373_,
		_w29369_,
		_w29387_
	);
	LUT3 #(
		.INIT('h51)
	) name23561 (
		_w29386_,
		_w29376_,
		_w29387_,
		_w29388_
	);
	LUT4 #(
		.INIT('h5455)
	) name23562 (
		_w29375_,
		_w29383_,
		_w29385_,
		_w29388_,
		_w29389_
	);
	LUT4 #(
		.INIT('h2000)
	) name23563 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29390_
	);
	LUT2 #(
		.INIT('h8)
	) name23564 (
		_w29375_,
		_w29390_,
		_w29391_
	);
	LUT4 #(
		.INIT('h0082)
	) name23565 (
		_w29375_,
		_w29370_,
		_w29371_,
		_w29372_,
		_w29392_
	);
	LUT3 #(
		.INIT('h54)
	) name23566 (
		_w29369_,
		_w29392_,
		_w29374_,
		_w29393_
	);
	LUT2 #(
		.INIT('h1)
	) name23567 (
		_w29391_,
		_w29393_,
		_w29394_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name23568 (
		\u0_L6_reg[5]/NET0131 ,
		_w29389_,
		_w29381_,
		_w29394_,
		_w29395_
	);
	LUT4 #(
		.INIT('hc963)
	) name23569 (
		decrypt_pad,
		\u0_R6_reg[8]/NET0131 ,
		\u0_uk_K_r6_reg[48]/NET0131 ,
		\u0_uk_K_r6_reg[55]/P0001 ,
		_w29396_
	);
	LUT4 #(
		.INIT('hc693)
	) name23570 (
		decrypt_pad,
		\u0_R6_reg[6]/NET0131 ,
		\u0_uk_K_r6_reg[13]/NET0131 ,
		\u0_uk_K_r6_reg[6]/NET0131 ,
		_w29397_
	);
	LUT4 #(
		.INIT('hc693)
	) name23571 (
		decrypt_pad,
		\u0_R6_reg[9]/NET0131 ,
		\u0_uk_K_r6_reg[3]/NET0131 ,
		\u0_uk_K_r6_reg[53]/NET0131 ,
		_w29398_
	);
	LUT4 #(
		.INIT('hc963)
	) name23572 (
		decrypt_pad,
		\u0_R6_reg[5]/NET0131 ,
		\u0_uk_K_r6_reg[40]/NET0131 ,
		\u0_uk_K_r6_reg[47]/NET0131 ,
		_w29399_
	);
	LUT4 #(
		.INIT('hc963)
	) name23573 (
		decrypt_pad,
		\u0_R6_reg[7]/NET0131 ,
		\u0_uk_K_r6_reg[25]/NET0131 ,
		\u0_uk_K_r6_reg[32]/NET0131 ,
		_w29400_
	);
	LUT4 #(
		.INIT('h0004)
	) name23574 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29400_,
		_w29401_
	);
	LUT4 #(
		.INIT('hc693)
	) name23575 (
		decrypt_pad,
		\u0_R6_reg[4]/NET0131 ,
		\u0_uk_K_r6_reg[11]/NET0131 ,
		\u0_uk_K_r6_reg[4]/NET0131 ,
		_w29402_
	);
	LUT2 #(
		.INIT('h2)
	) name23576 (
		_w29398_,
		_w29402_,
		_w29403_
	);
	LUT3 #(
		.INIT('h08)
	) name23577 (
		_w29398_,
		_w29399_,
		_w29402_,
		_w29404_
	);
	LUT4 #(
		.INIT('h0080)
	) name23578 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29405_
	);
	LUT2 #(
		.INIT('h1)
	) name23579 (
		_w29401_,
		_w29405_,
		_w29406_
	);
	LUT4 #(
		.INIT('h0800)
	) name23580 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29407_
	);
	LUT4 #(
		.INIT('h0103)
	) name23581 (
		_w29400_,
		_w29401_,
		_w29405_,
		_w29407_,
		_w29408_
	);
	LUT2 #(
		.INIT('h8)
	) name23582 (
		_w29398_,
		_w29402_,
		_w29409_
	);
	LUT4 #(
		.INIT('h1014)
	) name23583 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29410_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name23584 (
		_w29398_,
		_w29399_,
		_w29400_,
		_w29402_,
		_w29411_
	);
	LUT4 #(
		.INIT('h51f3)
	) name23585 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29412_
	);
	LUT3 #(
		.INIT('h51)
	) name23586 (
		_w29410_,
		_w29411_,
		_w29412_,
		_w29413_
	);
	LUT3 #(
		.INIT('h15)
	) name23587 (
		_w29396_,
		_w29408_,
		_w29413_,
		_w29414_
	);
	LUT4 #(
		.INIT('hf7cc)
	) name23588 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29415_
	);
	LUT4 #(
		.INIT('h00c4)
	) name23589 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29416_
	);
	LUT3 #(
		.INIT('h0b)
	) name23590 (
		_w29397_,
		_w29399_,
		_w29400_,
		_w29417_
	);
	LUT4 #(
		.INIT('hf200)
	) name23591 (
		_w29396_,
		_w29415_,
		_w29416_,
		_w29417_,
		_w29418_
	);
	LUT4 #(
		.INIT('h0002)
	) name23592 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29419_
	);
	LUT4 #(
		.INIT('haffd)
	) name23593 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29420_
	);
	LUT2 #(
		.INIT('h2)
	) name23594 (
		_w29400_,
		_w29420_,
		_w29421_
	);
	LUT4 #(
		.INIT('h0100)
	) name23595 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29422_
	);
	LUT4 #(
		.INIT('hc040)
	) name23596 (
		_w29397_,
		_w29399_,
		_w29400_,
		_w29402_,
		_w29423_
	);
	LUT4 #(
		.INIT('h4000)
	) name23597 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29424_
	);
	LUT4 #(
		.INIT('haaa8)
	) name23598 (
		_w29396_,
		_w29422_,
		_w29423_,
		_w29424_,
		_w29425_
	);
	LUT3 #(
		.INIT('h01)
	) name23599 (
		_w29421_,
		_w29425_,
		_w29418_,
		_w29426_
	);
	LUT3 #(
		.INIT('h65)
	) name23600 (
		\u0_L6_reg[2]/NET0131 ,
		_w29414_,
		_w29426_,
		_w29427_
	);
	LUT4 #(
		.INIT('h779a)
	) name23601 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29428_
	);
	LUT4 #(
		.INIT('h0e02)
	) name23602 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29429_
	);
	LUT4 #(
		.INIT('hf17d)
	) name23603 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29430_
	);
	LUT4 #(
		.INIT('h1000)
	) name23604 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29431_
	);
	LUT4 #(
		.INIT('h00e4)
	) name23605 (
		_w29272_,
		_w29430_,
		_w29428_,
		_w29431_,
		_w29432_
	);
	LUT2 #(
		.INIT('h1)
	) name23606 (
		_w29271_,
		_w29432_,
		_w29433_
	);
	LUT4 #(
		.INIT('hdd7d)
	) name23607 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29434_
	);
	LUT2 #(
		.INIT('h2)
	) name23608 (
		_w29272_,
		_w29434_,
		_w29435_
	);
	LUT3 #(
		.INIT('h48)
	) name23609 (
		_w29274_,
		_w29275_,
		_w29276_,
		_w29436_
	);
	LUT4 #(
		.INIT('hab00)
	) name23610 (
		_w29273_,
		_w29275_,
		_w29276_,
		_w29272_,
		_w29437_
	);
	LUT3 #(
		.INIT('h01)
	) name23611 (
		_w29437_,
		_w29429_,
		_w29436_,
		_w29438_
	);
	LUT4 #(
		.INIT('h2000)
	) name23612 (
		_w29273_,
		_w29275_,
		_w29276_,
		_w29272_,
		_w29439_
	);
	LUT2 #(
		.INIT('h1)
	) name23613 (
		_w29277_,
		_w29439_,
		_w29440_
	);
	LUT4 #(
		.INIT('h5700)
	) name23614 (
		_w29271_,
		_w29435_,
		_w29438_,
		_w29440_,
		_w29441_
	);
	LUT3 #(
		.INIT('h9a)
	) name23615 (
		\u0_L6_reg[29]/NET0131 ,
		_w29433_,
		_w29441_,
		_w29442_
	);
	LUT4 #(
		.INIT('hde00)
	) name23616 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29443_
	);
	LUT4 #(
		.INIT('h0205)
	) name23617 (
		_w29244_,
		_w29245_,
		_w29243_,
		_w29246_,
		_w29444_
	);
	LUT4 #(
		.INIT('h9000)
	) name23618 (
		_w29244_,
		_w29245_,
		_w29243_,
		_w29246_,
		_w29445_
	);
	LUT4 #(
		.INIT('hbdff)
	) name23619 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29446_
	);
	LUT4 #(
		.INIT('h0b00)
	) name23620 (
		_w29443_,
		_w29444_,
		_w29445_,
		_w29446_,
		_w29447_
	);
	LUT2 #(
		.INIT('h1)
	) name23621 (
		_w29242_,
		_w29447_,
		_w29448_
	);
	LUT3 #(
		.INIT('hb7)
	) name23622 (
		_w29244_,
		_w29245_,
		_w29247_,
		_w29449_
	);
	LUT2 #(
		.INIT('h2)
	) name23623 (
		_w29265_,
		_w29449_,
		_w29450_
	);
	LUT3 #(
		.INIT('hc8)
	) name23624 (
		_w29245_,
		_w29246_,
		_w29247_,
		_w29451_
	);
	LUT4 #(
		.INIT('h0013)
	) name23625 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29452_
	);
	LUT3 #(
		.INIT('h02)
	) name23626 (
		_w29243_,
		_w29452_,
		_w29451_,
		_w29453_
	);
	LUT4 #(
		.INIT('h0040)
	) name23627 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29454_
	);
	LUT3 #(
		.INIT('h80)
	) name23628 (
		_w29244_,
		_w29245_,
		_w29247_,
		_w29455_
	);
	LUT4 #(
		.INIT('h3001)
	) name23629 (
		_w29245_,
		_w29243_,
		_w29246_,
		_w29247_,
		_w29456_
	);
	LUT3 #(
		.INIT('h01)
	) name23630 (
		_w29455_,
		_w29456_,
		_w29454_,
		_w29457_
	);
	LUT4 #(
		.INIT('h1311)
	) name23631 (
		_w29242_,
		_w29450_,
		_w29453_,
		_w29457_,
		_w29458_
	);
	LUT3 #(
		.INIT('h65)
	) name23632 (
		\u0_L6_reg[17]/NET0131 ,
		_w29448_,
		_w29458_,
		_w29459_
	);
	LUT3 #(
		.INIT('h02)
	) name23633 (
		_w29273_,
		_w29275_,
		_w29276_,
		_w29460_
	);
	LUT4 #(
		.INIT('hfcf4)
	) name23634 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29461_
	);
	LUT2 #(
		.INIT('h1)
	) name23635 (
		_w29272_,
		_w29461_,
		_w29462_
	);
	LUT4 #(
		.INIT('h0002)
	) name23636 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29463_
	);
	LUT3 #(
		.INIT('h80)
	) name23637 (
		_w29273_,
		_w29275_,
		_w29276_,
		_w29464_
	);
	LUT4 #(
		.INIT('h2000)
	) name23638 (
		_w29274_,
		_w29275_,
		_w29276_,
		_w29272_,
		_w29465_
	);
	LUT4 #(
		.INIT('h0002)
	) name23639 (
		_w29271_,
		_w29463_,
		_w29465_,
		_w29464_,
		_w29466_
	);
	LUT2 #(
		.INIT('h4)
	) name23640 (
		_w29462_,
		_w29466_,
		_w29467_
	);
	LUT4 #(
		.INIT('hbc77)
	) name23641 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29468_
	);
	LUT2 #(
		.INIT('h2)
	) name23642 (
		_w29272_,
		_w29468_,
		_w29469_
	);
	LUT4 #(
		.INIT('hefdd)
	) name23643 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29470_
	);
	LUT2 #(
		.INIT('h1)
	) name23644 (
		_w29272_,
		_w29470_,
		_w29471_
	);
	LUT3 #(
		.INIT('h01)
	) name23645 (
		_w29271_,
		_w29277_,
		_w29281_,
		_w29472_
	);
	LUT3 #(
		.INIT('h10)
	) name23646 (
		_w29471_,
		_w29469_,
		_w29472_,
		_w29473_
	);
	LUT4 #(
		.INIT('h70b0)
	) name23647 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29474_
	);
	LUT4 #(
		.INIT('h00cd)
	) name23648 (
		_w29274_,
		_w29275_,
		_w29276_,
		_w29272_,
		_w29475_
	);
	LUT3 #(
		.INIT('hde)
	) name23649 (
		_w29273_,
		_w29274_,
		_w29276_,
		_w29476_
	);
	LUT3 #(
		.INIT('hd6)
	) name23650 (
		_w29273_,
		_w29274_,
		_w29276_,
		_w29477_
	);
	LUT2 #(
		.INIT('h8)
	) name23651 (
		_w29275_,
		_w29272_,
		_w29478_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name23652 (
		_w29474_,
		_w29475_,
		_w29477_,
		_w29478_,
		_w29479_
	);
	LUT4 #(
		.INIT('ha955)
	) name23653 (
		\u0_L6_reg[4]/NET0131 ,
		_w29467_,
		_w29473_,
		_w29479_,
		_w29480_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name23654 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29481_
	);
	LUT2 #(
		.INIT('h2)
	) name23655 (
		_w29313_,
		_w29481_,
		_w29482_
	);
	LUT3 #(
		.INIT('h04)
	) name23656 (
		_w29308_,
		_w29311_,
		_w29322_,
		_w29483_
	);
	LUT2 #(
		.INIT('h9)
	) name23657 (
		_w29303_,
		_w29304_,
		_w29484_
	);
	LUT4 #(
		.INIT('h2022)
	) name23658 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29313_,
		_w29485_
	);
	LUT4 #(
		.INIT('h0400)
	) name23659 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29486_
	);
	LUT3 #(
		.INIT('h0b)
	) name23660 (
		_w29484_,
		_w29485_,
		_w29486_,
		_w29487_
	);
	LUT3 #(
		.INIT('h40)
	) name23661 (
		_w29482_,
		_w29483_,
		_w29487_,
		_w29488_
	);
	LUT3 #(
		.INIT('h08)
	) name23662 (
		_w29301_,
		_w29303_,
		_w29304_,
		_w29489_
	);
	LUT4 #(
		.INIT('h2016)
	) name23663 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29490_
	);
	LUT3 #(
		.INIT('h09)
	) name23664 (
		_w29302_,
		_w29304_,
		_w29313_,
		_w29491_
	);
	LUT3 #(
		.INIT('h47)
	) name23665 (
		_w29301_,
		_w29302_,
		_w29313_,
		_w29492_
	);
	LUT4 #(
		.INIT('h0f07)
	) name23666 (
		_w29301_,
		_w29303_,
		_w29311_,
		_w29313_,
		_w29493_
	);
	LUT4 #(
		.INIT('h0d00)
	) name23667 (
		_w29305_,
		_w29492_,
		_w29491_,
		_w29493_,
		_w29494_
	);
	LUT2 #(
		.INIT('h4)
	) name23668 (
		_w29490_,
		_w29494_,
		_w29495_
	);
	LUT3 #(
		.INIT('ha9)
	) name23669 (
		\u0_L6_reg[12]/NET0131 ,
		_w29488_,
		_w29495_,
		_w29496_
	);
	LUT4 #(
		.INIT('h3b19)
	) name23670 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29497_
	);
	LUT4 #(
		.INIT('h8000)
	) name23671 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29498_
	);
	LUT4 #(
		.INIT('h0e04)
	) name23672 (
		_w29272_,
		_w29476_,
		_w29498_,
		_w29497_,
		_w29499_
	);
	LUT2 #(
		.INIT('h1)
	) name23673 (
		_w29271_,
		_w29499_,
		_w29500_
	);
	LUT4 #(
		.INIT('h2010)
	) name23674 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29501_
	);
	LUT4 #(
		.INIT('he6f7)
	) name23675 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29502_
	);
	LUT2 #(
		.INIT('h2)
	) name23676 (
		_w29272_,
		_w29502_,
		_w29503_
	);
	LUT4 #(
		.INIT('h0100)
	) name23677 (
		_w29273_,
		_w29274_,
		_w29275_,
		_w29276_,
		_w29504_
	);
	LUT3 #(
		.INIT('h04)
	) name23678 (
		_w29273_,
		_w29274_,
		_w29272_,
		_w29505_
	);
	LUT3 #(
		.INIT('h01)
	) name23679 (
		_w29460_,
		_w29504_,
		_w29505_,
		_w29506_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name23680 (
		_w29271_,
		_w29503_,
		_w29501_,
		_w29506_,
		_w29507_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name23681 (
		_w29273_,
		_w29275_,
		_w29293_,
		_w29281_,
		_w29508_
	);
	LUT4 #(
		.INIT('h5655)
	) name23682 (
		\u0_L6_reg[19]/P0001 ,
		_w29507_,
		_w29500_,
		_w29508_,
		_w29509_
	);
	LUT4 #(
		.INIT('hc963)
	) name23683 (
		decrypt_pad,
		\u0_R6_reg[20]/NET0131 ,
		\u0_uk_K_r6_reg[28]/NET0131 ,
		\u0_uk_K_r6_reg[35]/NET0131 ,
		_w29510_
	);
	LUT4 #(
		.INIT('hc693)
	) name23684 (
		decrypt_pad,
		\u0_R6_reg[17]/NET0131 ,
		\u0_uk_K_r6_reg[15]/NET0131 ,
		\u0_uk_K_r6_reg[8]/NET0131 ,
		_w29511_
	);
	LUT4 #(
		.INIT('hc963)
	) name23685 (
		decrypt_pad,
		\u0_R6_reg[16]/NET0131 ,
		\u0_uk_K_r6_reg[45]/NET0131 ,
		\u0_uk_K_r6_reg[52]/NET0131 ,
		_w29512_
	);
	LUT4 #(
		.INIT('hc963)
	) name23686 (
		decrypt_pad,
		\u0_R6_reg[21]/NET0131 ,
		\u0_uk_K_r6_reg[29]/NET0131 ,
		\u0_uk_K_r6_reg[36]/NET0131 ,
		_w29513_
	);
	LUT3 #(
		.INIT('h80)
	) name23687 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29514_
	);
	LUT4 #(
		.INIT('hc963)
	) name23688 (
		decrypt_pad,
		\u0_R6_reg[19]/NET0131 ,
		\u0_uk_K_r6_reg[44]/NET0131 ,
		\u0_uk_K_r6_reg[51]/NET0131 ,
		_w29515_
	);
	LUT4 #(
		.INIT('hc963)
	) name23689 (
		decrypt_pad,
		\u0_R6_reg[18]/NET0131 ,
		\u0_uk_K_r6_reg[2]/NET0131 ,
		\u0_uk_K_r6_reg[9]/NET0131 ,
		_w29516_
	);
	LUT4 #(
		.INIT('h0004)
	) name23690 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29517_
	);
	LUT3 #(
		.INIT('h02)
	) name23691 (
		_w29515_,
		_w29514_,
		_w29517_,
		_w29518_
	);
	LUT4 #(
		.INIT('h2030)
	) name23692 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29519_
	);
	LUT4 #(
		.INIT('h00bf)
	) name23693 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29515_,
		_w29520_
	);
	LUT2 #(
		.INIT('h4)
	) name23694 (
		_w29519_,
		_w29520_,
		_w29521_
	);
	LUT4 #(
		.INIT('hf6dd)
	) name23695 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29522_
	);
	LUT4 #(
		.INIT('h0155)
	) name23696 (
		_w29510_,
		_w29518_,
		_w29521_,
		_w29522_,
		_w29523_
	);
	LUT4 #(
		.INIT('hbfbe)
	) name23697 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29524_
	);
	LUT4 #(
		.INIT('h1200)
	) name23698 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29525_
	);
	LUT2 #(
		.INIT('h1)
	) name23699 (
		_w29515_,
		_w29516_,
		_w29526_
	);
	LUT3 #(
		.INIT('h02)
	) name23700 (
		_w29512_,
		_w29515_,
		_w29516_,
		_w29527_
	);
	LUT4 #(
		.INIT('h0031)
	) name23701 (
		_w29515_,
		_w29525_,
		_w29524_,
		_w29527_,
		_w29528_
	);
	LUT3 #(
		.INIT('h04)
	) name23702 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29529_
	);
	LUT2 #(
		.INIT('h4)
	) name23703 (
		_w29515_,
		_w29516_,
		_w29530_
	);
	LUT4 #(
		.INIT('h1000)
	) name23704 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29531_
	);
	LUT4 #(
		.INIT('he5df)
	) name23705 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29532_
	);
	LUT4 #(
		.INIT('hdf13)
	) name23706 (
		_w29529_,
		_w29515_,
		_w29516_,
		_w29532_,
		_w29533_
	);
	LUT3 #(
		.INIT('hd0)
	) name23707 (
		_w29510_,
		_w29528_,
		_w29533_,
		_w29534_
	);
	LUT3 #(
		.INIT('h65)
	) name23708 (
		\u0_L6_reg[8]/NET0131 ,
		_w29523_,
		_w29534_,
		_w29535_
	);
	LUT4 #(
		.INIT('hf636)
	) name23709 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29536_
	);
	LUT2 #(
		.INIT('h2)
	) name23710 (
		_w29369_,
		_w29536_,
		_w29537_
	);
	LUT4 #(
		.INIT('h0009)
	) name23711 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29538_
	);
	LUT4 #(
		.INIT('h0004)
	) name23712 (
		_w29371_,
		_w29372_,
		_w29373_,
		_w29369_,
		_w29539_
	);
	LUT4 #(
		.INIT('h5155)
	) name23713 (
		_w29375_,
		_w29370_,
		_w29371_,
		_w29372_,
		_w29540_
	);
	LUT2 #(
		.INIT('h4)
	) name23714 (
		_w29539_,
		_w29540_,
		_w29541_
	);
	LUT4 #(
		.INIT('h0020)
	) name23715 (
		_w29370_,
		_w29371_,
		_w29373_,
		_w29369_,
		_w29542_
	);
	LUT3 #(
		.INIT('h73)
	) name23716 (
		_w29372_,
		_w29373_,
		_w29369_,
		_w29543_
	);
	LUT3 #(
		.INIT('h31)
	) name23717 (
		_w29376_,
		_w29542_,
		_w29543_,
		_w29544_
	);
	LUT4 #(
		.INIT('h1000)
	) name23718 (
		_w29538_,
		_w29537_,
		_w29541_,
		_w29544_,
		_w29545_
	);
	LUT4 #(
		.INIT('h0800)
	) name23719 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29546_
	);
	LUT4 #(
		.INIT('h4044)
	) name23720 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29547_
	);
	LUT3 #(
		.INIT('h01)
	) name23721 (
		_w29369_,
		_w29546_,
		_w29547_,
		_w29548_
	);
	LUT4 #(
		.INIT('h3101)
	) name23722 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29549_
	);
	LUT3 #(
		.INIT('h10)
	) name23723 (
		_w29370_,
		_w29372_,
		_w29373_,
		_w29550_
	);
	LUT4 #(
		.INIT('h7f00)
	) name23724 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29369_,
		_w29551_
	);
	LUT3 #(
		.INIT('h10)
	) name23725 (
		_w29549_,
		_w29550_,
		_w29551_,
		_w29552_
	);
	LUT4 #(
		.INIT('h0082)
	) name23726 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29553_
	);
	LUT4 #(
		.INIT('h0100)
	) name23727 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29554_
	);
	LUT3 #(
		.INIT('h02)
	) name23728 (
		_w29375_,
		_w29554_,
		_w29553_,
		_w29555_
	);
	LUT3 #(
		.INIT('he0)
	) name23729 (
		_w29548_,
		_w29552_,
		_w29555_,
		_w29556_
	);
	LUT3 #(
		.INIT('ha9)
	) name23730 (
		\u0_L6_reg[21]/NET0131 ,
		_w29545_,
		_w29556_,
		_w29557_
	);
	LUT3 #(
		.INIT('hd9)
	) name23731 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29558_
	);
	LUT4 #(
		.INIT('he9f9)
	) name23732 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29559_
	);
	LUT2 #(
		.INIT('h1)
	) name23733 (
		_w29243_,
		_w29559_,
		_w29560_
	);
	LUT3 #(
		.INIT('ha2)
	) name23734 (
		_w29243_,
		_w29246_,
		_w29247_,
		_w29561_
	);
	LUT2 #(
		.INIT('h8)
	) name23735 (
		_w29259_,
		_w29561_,
		_w29562_
	);
	LUT4 #(
		.INIT('h0020)
	) name23736 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29563_
	);
	LUT3 #(
		.INIT('h07)
	) name23737 (
		_w29251_,
		_w29266_,
		_w29563_,
		_w29564_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name23738 (
		_w29242_,
		_w29560_,
		_w29562_,
		_w29564_,
		_w29565_
	);
	LUT4 #(
		.INIT('h51ff)
	) name23739 (
		_w29245_,
		_w29243_,
		_w29246_,
		_w29247_,
		_w29566_
	);
	LUT2 #(
		.INIT('h2)
	) name23740 (
		_w29244_,
		_w29566_,
		_w29567_
	);
	LUT4 #(
		.INIT('h0040)
	) name23741 (
		_w29244_,
		_w29245_,
		_w29243_,
		_w29246_,
		_w29568_
	);
	LUT3 #(
		.INIT('h01)
	) name23742 (
		_w29244_,
		_w29245_,
		_w29247_,
		_w29569_
	);
	LUT3 #(
		.INIT('h0e)
	) name23743 (
		_w29244_,
		_w29245_,
		_w29243_,
		_w29570_
	);
	LUT4 #(
		.INIT('h0013)
	) name23744 (
		_w29451_,
		_w29569_,
		_w29570_,
		_w29568_,
		_w29571_
	);
	LUT3 #(
		.INIT('hcb)
	) name23745 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29572_
	);
	LUT4 #(
		.INIT('h7fbd)
	) name23746 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29573_
	);
	LUT4 #(
		.INIT('hfda8)
	) name23747 (
		_w29243_,
		_w29247_,
		_w29572_,
		_w29573_,
		_w29574_
	);
	LUT4 #(
		.INIT('hba00)
	) name23748 (
		_w29242_,
		_w29567_,
		_w29571_,
		_w29574_,
		_w29575_
	);
	LUT3 #(
		.INIT('h9a)
	) name23749 (
		\u0_L6_reg[23]/NET0131 ,
		_w29565_,
		_w29575_,
		_w29576_
	);
	LUT4 #(
		.INIT('hff2e)
	) name23750 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29577_
	);
	LUT3 #(
		.INIT('h02)
	) name23751 (
		_w29397_,
		_w29399_,
		_w29402_,
		_w29578_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name23752 (
		_w29397_,
		_w29399_,
		_w29400_,
		_w29402_,
		_w29579_
	);
	LUT4 #(
		.INIT('h0ef3)
	) name23753 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29580_
	);
	LUT4 #(
		.INIT('h7277)
	) name23754 (
		_w29400_,
		_w29577_,
		_w29578_,
		_w29580_,
		_w29581_
	);
	LUT4 #(
		.INIT('h0802)
	) name23755 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29582_
	);
	LUT4 #(
		.INIT('h2000)
	) name23756 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29583_
	);
	LUT3 #(
		.INIT('h01)
	) name23757 (
		_w29396_,
		_w29583_,
		_w29582_,
		_w29584_
	);
	LUT2 #(
		.INIT('h4)
	) name23758 (
		_w29581_,
		_w29584_,
		_w29585_
	);
	LUT3 #(
		.INIT('h90)
	) name23759 (
		_w29398_,
		_w29399_,
		_w29402_,
		_w29586_
	);
	LUT4 #(
		.INIT('h0020)
	) name23760 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29587_
	);
	LUT3 #(
		.INIT('h02)
	) name23761 (
		_w29400_,
		_w29587_,
		_w29586_,
		_w29588_
	);
	LUT4 #(
		.INIT('hdf2e)
	) name23762 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29589_
	);
	LUT2 #(
		.INIT('h8)
	) name23763 (
		_w29579_,
		_w29589_,
		_w29590_
	);
	LUT2 #(
		.INIT('h8)
	) name23764 (
		_w29400_,
		_w29402_,
		_w29591_
	);
	LUT4 #(
		.INIT('h0dff)
	) name23765 (
		_w29398_,
		_w29399_,
		_w29400_,
		_w29402_,
		_w29592_
	);
	LUT4 #(
		.INIT('h0008)
	) name23766 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29593_
	);
	LUT4 #(
		.INIT('h00a8)
	) name23767 (
		_w29396_,
		_w29397_,
		_w29592_,
		_w29593_,
		_w29594_
	);
	LUT3 #(
		.INIT('he0)
	) name23768 (
		_w29588_,
		_w29590_,
		_w29594_,
		_w29595_
	);
	LUT3 #(
		.INIT('ha9)
	) name23769 (
		\u0_L6_reg[28]/NET0131 ,
		_w29585_,
		_w29595_,
		_w29596_
	);
	LUT4 #(
		.INIT('hc727)
	) name23770 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29597_
	);
	LUT2 #(
		.INIT('h2)
	) name23771 (
		_w29515_,
		_w29597_,
		_w29598_
	);
	LUT3 #(
		.INIT('hde)
	) name23772 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29599_
	);
	LUT2 #(
		.INIT('h2)
	) name23773 (
		_w29526_,
		_w29599_,
		_w29600_
	);
	LUT4 #(
		.INIT('h0440)
	) name23774 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29601_
	);
	LUT4 #(
		.INIT('h0008)
	) name23775 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29602_
	);
	LUT4 #(
		.INIT('h0007)
	) name23776 (
		_w29530_,
		_w29514_,
		_w29602_,
		_w29601_,
		_w29603_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name23777 (
		_w29510_,
		_w29600_,
		_w29598_,
		_w29603_,
		_w29604_
	);
	LUT4 #(
		.INIT('h0080)
	) name23778 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29605_
	);
	LUT4 #(
		.INIT('he56b)
	) name23779 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29606_
	);
	LUT4 #(
		.INIT('h3edc)
	) name23780 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29607_
	);
	LUT4 #(
		.INIT('h4002)
	) name23781 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29608_
	);
	LUT4 #(
		.INIT('h00d8)
	) name23782 (
		_w29515_,
		_w29607_,
		_w29606_,
		_w29608_,
		_w29609_
	);
	LUT4 #(
		.INIT('h0100)
	) name23783 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29610_
	);
	LUT4 #(
		.INIT('heee4)
	) name23784 (
		_w29515_,
		_w29525_,
		_w29602_,
		_w29610_,
		_w29611_
	);
	LUT3 #(
		.INIT('h0e)
	) name23785 (
		_w29510_,
		_w29609_,
		_w29611_,
		_w29612_
	);
	LUT3 #(
		.INIT('h65)
	) name23786 (
		\u0_L6_reg[14]/NET0131 ,
		_w29604_,
		_w29612_,
		_w29613_
	);
	LUT4 #(
		.INIT('h4060)
	) name23787 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29614_
	);
	LUT4 #(
		.INIT('hfc5f)
	) name23788 (
		_w29370_,
		_w29371_,
		_w29373_,
		_w29369_,
		_w29615_
	);
	LUT4 #(
		.INIT('h0032)
	) name23789 (
		_w29372_,
		_w29546_,
		_w29615_,
		_w29614_,
		_w29616_
	);
	LUT2 #(
		.INIT('h2)
	) name23790 (
		_w29375_,
		_w29616_,
		_w29617_
	);
	LUT4 #(
		.INIT('h3c2f)
	) name23791 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29618_
	);
	LUT4 #(
		.INIT('h0004)
	) name23792 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29619_
	);
	LUT4 #(
		.INIT('h5504)
	) name23793 (
		_w29375_,
		_w29369_,
		_w29618_,
		_w29619_,
		_w29620_
	);
	LUT4 #(
		.INIT('he7d6)
	) name23794 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29621_
	);
	LUT2 #(
		.INIT('h1)
	) name23795 (
		_w29369_,
		_w29621_,
		_w29622_
	);
	LUT4 #(
		.INIT('h0004)
	) name23796 (
		_w29375_,
		_w29371_,
		_w29372_,
		_w29369_,
		_w29623_
	);
	LUT3 #(
		.INIT('hb0)
	) name23797 (
		_w29370_,
		_w29372_,
		_w29373_,
		_w29624_
	);
	LUT4 #(
		.INIT('h3100)
	) name23798 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29369_,
		_w29625_
	);
	LUT3 #(
		.INIT('h15)
	) name23799 (
		_w29623_,
		_w29624_,
		_w29625_,
		_w29626_
	);
	LUT3 #(
		.INIT('h10)
	) name23800 (
		_w29620_,
		_w29622_,
		_w29626_,
		_w29627_
	);
	LUT3 #(
		.INIT('h65)
	) name23801 (
		\u0_L6_reg[15]/P0001 ,
		_w29617_,
		_w29627_,
		_w29628_
	);
	LUT4 #(
		.INIT('h9fff)
	) name23802 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29629_
	);
	LUT4 #(
		.INIT('hfec7)
	) name23803 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29630_
	);
	LUT4 #(
		.INIT('h0313)
	) name23804 (
		_w29396_,
		_w29400_,
		_w29629_,
		_w29630_,
		_w29631_
	);
	LUT3 #(
		.INIT('h12)
	) name23805 (
		_w29398_,
		_w29399_,
		_w29402_,
		_w29632_
	);
	LUT4 #(
		.INIT('he0f0)
	) name23806 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29633_
	);
	LUT3 #(
		.INIT('h02)
	) name23807 (
		_w29400_,
		_w29633_,
		_w29632_,
		_w29634_
	);
	LUT3 #(
		.INIT('h54)
	) name23808 (
		_w29397_,
		_w29399_,
		_w29400_,
		_w29635_
	);
	LUT2 #(
		.INIT('h8)
	) name23809 (
		_w29403_,
		_w29635_,
		_w29636_
	);
	LUT3 #(
		.INIT('h8a)
	) name23810 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29637_
	);
	LUT3 #(
		.INIT('h15)
	) name23811 (
		_w29396_,
		_w29591_,
		_w29637_,
		_w29638_
	);
	LUT3 #(
		.INIT('h10)
	) name23812 (
		_w29636_,
		_w29634_,
		_w29638_,
		_w29639_
	);
	LUT3 #(
		.INIT('h02)
	) name23813 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29640_
	);
	LUT3 #(
		.INIT('h08)
	) name23814 (
		_w29397_,
		_w29398_,
		_w29402_,
		_w29641_
	);
	LUT4 #(
		.INIT('hfe00)
	) name23815 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29400_,
		_w29642_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name23816 (
		_w29411_,
		_w29640_,
		_w29641_,
		_w29642_,
		_w29643_
	);
	LUT4 #(
		.INIT('h0010)
	) name23817 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29644_
	);
	LUT3 #(
		.INIT('h08)
	) name23818 (
		_w29396_,
		_w29629_,
		_w29644_,
		_w29645_
	);
	LUT3 #(
		.INIT('h20)
	) name23819 (
		_w29406_,
		_w29643_,
		_w29645_,
		_w29646_
	);
	LUT4 #(
		.INIT('h999a)
	) name23820 (
		\u0_L6_reg[13]/NET0131 ,
		_w29631_,
		_w29639_,
		_w29646_,
		_w29647_
	);
	LUT4 #(
		.INIT('hdfdc)
	) name23821 (
		_w29331_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29648_
	);
	LUT2 #(
		.INIT('h1)
	) name23822 (
		_w29345_,
		_w29648_,
		_w29649_
	);
	LUT3 #(
		.INIT('h8a)
	) name23823 (
		_w29331_,
		_w29334_,
		_w29335_,
		_w29650_
	);
	LUT3 #(
		.INIT('h40)
	) name23824 (
		_w29334_,
		_w29333_,
		_w29332_,
		_w29651_
	);
	LUT4 #(
		.INIT('h1000)
	) name23825 (
		_w29331_,
		_w29334_,
		_w29333_,
		_w29335_,
		_w29652_
	);
	LUT4 #(
		.INIT('h0103)
	) name23826 (
		_w29356_,
		_w29651_,
		_w29652_,
		_w29650_,
		_w29653_
	);
	LUT3 #(
		.INIT('h20)
	) name23827 (
		_w29342_,
		_w29649_,
		_w29653_,
		_w29654_
	);
	LUT4 #(
		.INIT('hfcbf)
	) name23828 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29655_
	);
	LUT2 #(
		.INIT('h2)
	) name23829 (
		_w29331_,
		_w29655_,
		_w29656_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name23830 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29657_
	);
	LUT4 #(
		.INIT('he7f3)
	) name23831 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29658_
	);
	LUT4 #(
		.INIT('hc800)
	) name23832 (
		_w29331_,
		_w29341_,
		_w29658_,
		_w29657_,
		_w29659_
	);
	LUT2 #(
		.INIT('h4)
	) name23833 (
		_w29656_,
		_w29659_,
		_w29660_
	);
	LUT4 #(
		.INIT('he4f5)
	) name23834 (
		_w29331_,
		_w29337_,
		_w29365_,
		_w29657_,
		_w29661_
	);
	LUT2 #(
		.INIT('h1)
	) name23835 (
		_w29347_,
		_w29661_,
		_w29662_
	);
	LUT4 #(
		.INIT('ha955)
	) name23836 (
		\u0_L6_reg[10]/NET0131 ,
		_w29654_,
		_w29660_,
		_w29662_,
		_w29663_
	);
	LUT4 #(
		.INIT('h4104)
	) name23837 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29664_
	);
	LUT4 #(
		.INIT('hffd0)
	) name23838 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29665_
	);
	LUT4 #(
		.INIT('h0504)
	) name23839 (
		_w29331_,
		_w29341_,
		_w29664_,
		_w29665_,
		_w29666_
	);
	LUT3 #(
		.INIT('h02)
	) name23840 (
		_w29331_,
		_w29344_,
		_w29352_,
		_w29667_
	);
	LUT2 #(
		.INIT('h1)
	) name23841 (
		_w29666_,
		_w29667_,
		_w29668_
	);
	LUT4 #(
		.INIT('h5455)
	) name23842 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29669_
	);
	LUT3 #(
		.INIT('h9f)
	) name23843 (
		_w29333_,
		_w29335_,
		_w29332_,
		_w29670_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name23844 (
		_w29331_,
		_w29334_,
		_w29333_,
		_w29335_,
		_w29671_
	);
	LUT3 #(
		.INIT('h15)
	) name23845 (
		_w29669_,
		_w29670_,
		_w29671_,
		_w29672_
	);
	LUT4 #(
		.INIT('h3f2f)
	) name23846 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29673_
	);
	LUT3 #(
		.INIT('h45)
	) name23847 (
		_w29331_,
		_w29334_,
		_w29333_,
		_w29674_
	);
	LUT4 #(
		.INIT('h0002)
	) name23848 (
		_w29331_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29675_
	);
	LUT4 #(
		.INIT('h2022)
	) name23849 (
		_w29341_,
		_w29675_,
		_w29673_,
		_w29674_,
		_w29676_
	);
	LUT3 #(
		.INIT('h04)
	) name23850 (
		_w29334_,
		_w29333_,
		_w29332_,
		_w29677_
	);
	LUT3 #(
		.INIT('h01)
	) name23851 (
		_w29341_,
		_w29352_,
		_w29677_,
		_w29678_
	);
	LUT3 #(
		.INIT('h0b)
	) name23852 (
		_w29350_,
		_w29346_,
		_w29360_,
		_w29679_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name23853 (
		_w29672_,
		_w29676_,
		_w29678_,
		_w29679_,
		_w29680_
	);
	LUT3 #(
		.INIT('h56)
	) name23854 (
		\u0_L6_reg[26]/NET0131 ,
		_w29668_,
		_w29680_,
		_w29681_
	);
	LUT4 #(
		.INIT('h6c6a)
	) name23855 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29682_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name23856 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29683_
	);
	LUT4 #(
		.INIT('h08a0)
	) name23857 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29684_
	);
	LUT4 #(
		.INIT('h00d8)
	) name23858 (
		_w29515_,
		_w29682_,
		_w29683_,
		_w29684_,
		_w29685_
	);
	LUT2 #(
		.INIT('h4)
	) name23859 (
		_w29513_,
		_w29515_,
		_w29686_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name23860 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29687_
	);
	LUT3 #(
		.INIT('hd0)
	) name23861 (
		_w29511_,
		_w29513_,
		_w29515_,
		_w29688_
	);
	LUT4 #(
		.INIT('h00f1)
	) name23862 (
		_w29511_,
		_w29512_,
		_w29515_,
		_w29516_,
		_w29689_
	);
	LUT4 #(
		.INIT('he0ee)
	) name23863 (
		_w29686_,
		_w29687_,
		_w29688_,
		_w29689_,
		_w29690_
	);
	LUT4 #(
		.INIT('hf6ef)
	) name23864 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29691_
	);
	LUT4 #(
		.INIT('h0400)
	) name23865 (
		_w29511_,
		_w29512_,
		_w29515_,
		_w29516_,
		_w29692_
	);
	LUT4 #(
		.INIT('h0031)
	) name23866 (
		_w29515_,
		_w29605_,
		_w29691_,
		_w29692_,
		_w29693_
	);
	LUT4 #(
		.INIT('hd800)
	) name23867 (
		_w29510_,
		_w29685_,
		_w29690_,
		_w29693_,
		_w29694_
	);
	LUT2 #(
		.INIT('h9)
	) name23868 (
		\u0_L6_reg[25]/NET0131 ,
		_w29694_,
		_w29695_
	);
	LUT4 #(
		.INIT('h04c4)
	) name23869 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29696_
	);
	LUT4 #(
		.INIT('hfda8)
	) name23870 (
		_w29331_,
		_w29336_,
		_w29364_,
		_w29696_,
		_w29697_
	);
	LUT4 #(
		.INIT('h6bff)
	) name23871 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29698_
	);
	LUT3 #(
		.INIT('h45)
	) name23872 (
		_w29341_,
		_w29697_,
		_w29698_,
		_w29699_
	);
	LUT4 #(
		.INIT('h8eff)
	) name23873 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29700_
	);
	LUT4 #(
		.INIT('h0800)
	) name23874 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29701_
	);
	LUT4 #(
		.INIT('hf7dd)
	) name23875 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29702_
	);
	LUT4 #(
		.INIT('h04cc)
	) name23876 (
		_w29331_,
		_w29341_,
		_w29700_,
		_w29702_,
		_w29703_
	);
	LUT4 #(
		.INIT('h7ddf)
	) name23877 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29704_
	);
	LUT2 #(
		.INIT('h2)
	) name23878 (
		_w29331_,
		_w29704_,
		_w29705_
	);
	LUT2 #(
		.INIT('h4)
	) name23879 (
		_w29331_,
		_w29701_,
		_w29706_
	);
	LUT4 #(
		.INIT('hff0b)
	) name23880 (
		_w29334_,
		_w29333_,
		_w29335_,
		_w29332_,
		_w29707_
	);
	LUT2 #(
		.INIT('h8)
	) name23881 (
		_w29331_,
		_w29341_,
		_w29708_
	);
	LUT4 #(
		.INIT('h7077)
	) name23882 (
		_w29354_,
		_w29355_,
		_w29707_,
		_w29708_,
		_w29709_
	);
	LUT4 #(
		.INIT('h0100)
	) name23883 (
		_w29705_,
		_w29706_,
		_w29703_,
		_w29709_,
		_w29710_
	);
	LUT3 #(
		.INIT('h65)
	) name23884 (
		\u0_L6_reg[1]/NET0131 ,
		_w29699_,
		_w29710_,
		_w29711_
	);
	LUT4 #(
		.INIT('hd003)
	) name23885 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29712_
	);
	LUT3 #(
		.INIT('h28)
	) name23886 (
		_w29302_,
		_w29303_,
		_w29304_,
		_w29713_
	);
	LUT4 #(
		.INIT('h00d7)
	) name23887 (
		_w29301_,
		_w29303_,
		_w29304_,
		_w29313_,
		_w29714_
	);
	LUT3 #(
		.INIT('h10)
	) name23888 (
		_w29713_,
		_w29712_,
		_w29714_,
		_w29715_
	);
	LUT2 #(
		.INIT('h1)
	) name23889 (
		_w29302_,
		_w29313_,
		_w29716_
	);
	LUT4 #(
		.INIT('hbbfc)
	) name23890 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29717_
	);
	LUT4 #(
		.INIT('h1f13)
	) name23891 (
		_w29302_,
		_w29313_,
		_w29489_,
		_w29717_,
		_w29718_
	);
	LUT3 #(
		.INIT('h8a)
	) name23892 (
		_w29311_,
		_w29715_,
		_w29718_,
		_w29719_
	);
	LUT3 #(
		.INIT('hc4)
	) name23893 (
		_w29301_,
		_w29303_,
		_w29304_,
		_w29720_
	);
	LUT3 #(
		.INIT('h10)
	) name23894 (
		_w29310_,
		_w29716_,
		_w29720_,
		_w29721_
	);
	LUT3 #(
		.INIT('h04)
	) name23895 (
		_w29301_,
		_w29303_,
		_w29304_,
		_w29722_
	);
	LUT3 #(
		.INIT('ha2)
	) name23896 (
		_w29309_,
		_w29491_,
		_w29722_,
		_w29723_
	);
	LUT4 #(
		.INIT('h00a2)
	) name23897 (
		_w29302_,
		_w29303_,
		_w29304_,
		_w29313_,
		_w29724_
	);
	LUT4 #(
		.INIT('h0777)
	) name23898 (
		_w29306_,
		_w29313_,
		_w29318_,
		_w29724_,
		_w29725_
	);
	LUT4 #(
		.INIT('hba00)
	) name23899 (
		_w29311_,
		_w29721_,
		_w29723_,
		_w29725_,
		_w29726_
	);
	LUT3 #(
		.INIT('h65)
	) name23900 (
		\u0_L6_reg[32]/NET0131 ,
		_w29719_,
		_w29726_,
		_w29727_
	);
	LUT4 #(
		.INIT('hce3e)
	) name23901 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29728_
	);
	LUT2 #(
		.INIT('h1)
	) name23902 (
		_w29369_,
		_w29728_,
		_w29729_
	);
	LUT4 #(
		.INIT('h3323)
	) name23903 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29730_
	);
	LUT4 #(
		.INIT('hd500)
	) name23904 (
		_w29371_,
		_w29372_,
		_w29373_,
		_w29369_,
		_w29731_
	);
	LUT4 #(
		.INIT('hdaf7)
	) name23905 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29732_
	);
	LUT3 #(
		.INIT('hb0)
	) name23906 (
		_w29730_,
		_w29731_,
		_w29732_,
		_w29733_
	);
	LUT3 #(
		.INIT('h8a)
	) name23907 (
		_w29375_,
		_w29729_,
		_w29733_,
		_w29734_
	);
	LUT4 #(
		.INIT('hdf00)
	) name23908 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29369_,
		_w29735_
	);
	LUT3 #(
		.INIT('h4b)
	) name23909 (
		_w29370_,
		_w29372_,
		_w29373_,
		_w29736_
	);
	LUT2 #(
		.INIT('h8)
	) name23910 (
		_w29735_,
		_w29736_,
		_w29737_
	);
	LUT4 #(
		.INIT('h0080)
	) name23911 (
		_w29370_,
		_w29371_,
		_w29373_,
		_w29369_,
		_w29738_
	);
	LUT3 #(
		.INIT('h01)
	) name23912 (
		_w29378_,
		_w29539_,
		_w29738_,
		_w29739_
	);
	LUT4 #(
		.INIT('hfb9f)
	) name23913 (
		_w29370_,
		_w29371_,
		_w29372_,
		_w29373_,
		_w29740_
	);
	LUT4 #(
		.INIT('h0200)
	) name23914 (
		_w29370_,
		_w29372_,
		_w29373_,
		_w29369_,
		_w29741_
	);
	LUT3 #(
		.INIT('h0e)
	) name23915 (
		_w29369_,
		_w29740_,
		_w29741_,
		_w29742_
	);
	LUT4 #(
		.INIT('hba00)
	) name23916 (
		_w29375_,
		_w29737_,
		_w29739_,
		_w29742_,
		_w29743_
	);
	LUT3 #(
		.INIT('h65)
	) name23917 (
		\u0_L6_reg[27]/NET0131 ,
		_w29734_,
		_w29743_,
		_w29744_
	);
	LUT4 #(
		.INIT('hc693)
	) name23918 (
		decrypt_pad,
		\u0_R6_reg[8]/NET0131 ,
		\u0_uk_K_r6_reg[12]/NET0131 ,
		\u0_uk_K_r6_reg[5]/NET0131 ,
		_w29745_
	);
	LUT4 #(
		.INIT('hc963)
	) name23919 (
		decrypt_pad,
		\u0_R6_reg[13]/NET0131 ,
		\u0_uk_K_r6_reg[39]/NET0131 ,
		\u0_uk_K_r6_reg[46]/NET0131 ,
		_w29746_
	);
	LUT2 #(
		.INIT('h6)
	) name23920 (
		_w29745_,
		_w29746_,
		_w29747_
	);
	LUT4 #(
		.INIT('hc963)
	) name23921 (
		decrypt_pad,
		\u0_R6_reg[11]/NET0131 ,
		\u0_uk_K_r6_reg[11]/NET0131 ,
		\u0_uk_K_r6_reg[18]/NET0131 ,
		_w29748_
	);
	LUT4 #(
		.INIT('hc963)
	) name23922 (
		decrypt_pad,
		\u0_R6_reg[10]/NET0131 ,
		\u0_uk_K_r6_reg[10]/NET0131 ,
		\u0_uk_K_r6_reg[17]/NET0131 ,
		_w29749_
	);
	LUT4 #(
		.INIT('hc963)
	) name23923 (
		decrypt_pad,
		\u0_R6_reg[9]/NET0131 ,
		\u0_uk_K_r6_reg[34]/NET0131 ,
		\u0_uk_K_r6_reg[41]/NET0131 ,
		_w29750_
	);
	LUT4 #(
		.INIT('h000d)
	) name23924 (
		_w29748_,
		_w29745_,
		_w29749_,
		_w29750_,
		_w29751_
	);
	LUT2 #(
		.INIT('h8)
	) name23925 (
		_w29747_,
		_w29751_,
		_w29752_
	);
	LUT2 #(
		.INIT('h8)
	) name23926 (
		_w29749_,
		_w29750_,
		_w29753_
	);
	LUT4 #(
		.INIT('h2000)
	) name23927 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29754_
	);
	LUT4 #(
		.INIT('hc963)
	) name23928 (
		decrypt_pad,
		\u0_R6_reg[12]/NET0131 ,
		\u0_uk_K_r6_reg[26]/P0001 ,
		\u0_uk_K_r6_reg[33]/NET0131 ,
		_w29755_
	);
	LUT4 #(
		.INIT('h0200)
	) name23929 (
		_w29748_,
		_w29745_,
		_w29749_,
		_w29750_,
		_w29756_
	);
	LUT3 #(
		.INIT('h01)
	) name23930 (
		_w29755_,
		_w29756_,
		_w29754_,
		_w29757_
	);
	LUT4 #(
		.INIT('h4000)
	) name23931 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29758_
	);
	LUT4 #(
		.INIT('h9990)
	) name23932 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29759_
	);
	LUT4 #(
		.INIT('h0990)
	) name23933 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29760_
	);
	LUT3 #(
		.INIT('h0b)
	) name23934 (
		_w29748_,
		_w29758_,
		_w29760_,
		_w29761_
	);
	LUT3 #(
		.INIT('h45)
	) name23935 (
		_w29745_,
		_w29749_,
		_w29750_,
		_w29762_
	);
	LUT3 #(
		.INIT('h41)
	) name23936 (
		_w29748_,
		_w29746_,
		_w29750_,
		_w29763_
	);
	LUT4 #(
		.INIT('h1000)
	) name23937 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29764_
	);
	LUT4 #(
		.INIT('h2022)
	) name23938 (
		_w29755_,
		_w29764_,
		_w29762_,
		_w29763_,
		_w29765_
	);
	LUT4 #(
		.INIT('h00bf)
	) name23939 (
		_w29752_,
		_w29757_,
		_w29761_,
		_w29765_,
		_w29766_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23940 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29767_
	);
	LUT4 #(
		.INIT('h9d33)
	) name23941 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29768_
	);
	LUT3 #(
		.INIT('h08)
	) name23942 (
		_w29746_,
		_w29749_,
		_w29750_,
		_w29769_
	);
	LUT4 #(
		.INIT('h0001)
	) name23943 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29770_
	);
	LUT4 #(
		.INIT('hff3e)
	) name23944 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29771_
	);
	LUT4 #(
		.INIT('h08aa)
	) name23945 (
		_w29748_,
		_w29755_,
		_w29768_,
		_w29771_,
		_w29772_
	);
	LUT3 #(
		.INIT('h56)
	) name23946 (
		\u0_L6_reg[6]/NET0131 ,
		_w29766_,
		_w29772_,
		_w29773_
	);
	LUT3 #(
		.INIT('h02)
	) name23947 (
		_w29515_,
		_w29531_,
		_w29517_,
		_w29774_
	);
	LUT4 #(
		.INIT('h0009)
	) name23948 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29775_
	);
	LUT3 #(
		.INIT('h0e)
	) name23949 (
		_w29526_,
		_w29520_,
		_w29775_,
		_w29776_
	);
	LUT2 #(
		.INIT('h1)
	) name23950 (
		_w29774_,
		_w29776_,
		_w29777_
	);
	LUT4 #(
		.INIT('hf7c7)
	) name23951 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29778_
	);
	LUT2 #(
		.INIT('h2)
	) name23952 (
		_w29515_,
		_w29778_,
		_w29779_
	);
	LUT3 #(
		.INIT('h8c)
	) name23953 (
		_w29511_,
		_w29515_,
		_w29516_,
		_w29780_
	);
	LUT4 #(
		.INIT('h0cbc)
	) name23954 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29781_
	);
	LUT3 #(
		.INIT('h54)
	) name23955 (
		_w29510_,
		_w29780_,
		_w29781_,
		_w29782_
	);
	LUT4 #(
		.INIT('hfd3d)
	) name23956 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29783_
	);
	LUT2 #(
		.INIT('h2)
	) name23957 (
		_w29515_,
		_w29783_,
		_w29784_
	);
	LUT4 #(
		.INIT('h0020)
	) name23958 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29515_,
		_w29785_
	);
	LUT4 #(
		.INIT('h0400)
	) name23959 (
		_w29511_,
		_w29512_,
		_w29513_,
		_w29516_,
		_w29786_
	);
	LUT4 #(
		.INIT('h0002)
	) name23960 (
		_w29510_,
		_w29605_,
		_w29785_,
		_w29786_,
		_w29787_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name23961 (
		_w29779_,
		_w29782_,
		_w29784_,
		_w29787_,
		_w29788_
	);
	LUT3 #(
		.INIT('h56)
	) name23962 (
		\u0_L6_reg[3]/NET0131 ,
		_w29777_,
		_w29788_,
		_w29789_
	);
	LUT2 #(
		.INIT('h4)
	) name23963 (
		_w29311_,
		_w29313_,
		_w29790_
	);
	LUT4 #(
		.INIT('h0880)
	) name23964 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29791_
	);
	LUT4 #(
		.INIT('h877a)
	) name23965 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29792_
	);
	LUT2 #(
		.INIT('h2)
	) name23966 (
		_w29790_,
		_w29792_,
		_w29793_
	);
	LUT4 #(
		.INIT('h7004)
	) name23967 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29794_
	);
	LUT2 #(
		.INIT('h2)
	) name23968 (
		_w29311_,
		_w29313_,
		_w29795_
	);
	LUT2 #(
		.INIT('h9)
	) name23969 (
		_w29311_,
		_w29313_,
		_w29796_
	);
	LUT3 #(
		.INIT('h10)
	) name23970 (
		_w29791_,
		_w29794_,
		_w29796_,
		_w29797_
	);
	LUT4 #(
		.INIT('h2000)
	) name23971 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29798_
	);
	LUT4 #(
		.INIT('hf21e)
	) name23972 (
		_w29301_,
		_w29302_,
		_w29303_,
		_w29304_,
		_w29799_
	);
	LUT4 #(
		.INIT('h0400)
	) name23973 (
		_w29307_,
		_w29795_,
		_w29798_,
		_w29799_,
		_w29800_
	);
	LUT4 #(
		.INIT('h00ab)
	) name23974 (
		_w29317_,
		_w29793_,
		_w29797_,
		_w29800_,
		_w29801_
	);
	LUT2 #(
		.INIT('h6)
	) name23975 (
		\u0_L6_reg[7]/NET0131 ,
		_w29801_,
		_w29802_
	);
	LUT4 #(
		.INIT('h9600)
	) name23976 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29803_
	);
	LUT3 #(
		.INIT('he6)
	) name23977 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29804_
	);
	LUT4 #(
		.INIT('h0031)
	) name23978 (
		_w29254_,
		_w29454_,
		_w29804_,
		_w29803_,
		_w29805_
	);
	LUT4 #(
		.INIT('h2180)
	) name23979 (
		_w29244_,
		_w29245_,
		_w29246_,
		_w29247_,
		_w29806_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name23980 (
		_w29244_,
		_w29245_,
		_w29243_,
		_w29247_,
		_w29807_
	);
	LUT4 #(
		.INIT('h0e06)
	) name23981 (
		_w29244_,
		_w29245_,
		_w29243_,
		_w29246_,
		_w29808_
	);
	LUT4 #(
		.INIT('h3320)
	) name23982 (
		_w29558_,
		_w29806_,
		_w29807_,
		_w29808_,
		_w29809_
	);
	LUT3 #(
		.INIT('h08)
	) name23983 (
		_w29244_,
		_w29245_,
		_w29243_,
		_w29810_
	);
	LUT2 #(
		.INIT('h4)
	) name23984 (
		_w29261_,
		_w29810_,
		_w29811_
	);
	LUT4 #(
		.INIT('h00e4)
	) name23985 (
		_w29242_,
		_w29809_,
		_w29805_,
		_w29811_,
		_w29812_
	);
	LUT2 #(
		.INIT('h9)
	) name23986 (
		\u0_L6_reg[9]/NET0131 ,
		_w29812_,
		_w29813_
	);
	LUT3 #(
		.INIT('h1d)
	) name23987 (
		_w29397_,
		_w29399_,
		_w29400_,
		_w29814_
	);
	LUT3 #(
		.INIT('h0b)
	) name23988 (
		_w29397_,
		_w29399_,
		_w29402_,
		_w29815_
	);
	LUT4 #(
		.INIT('hdefe)
	) name23989 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29402_,
		_w29816_
	);
	LUT4 #(
		.INIT('h3500)
	) name23990 (
		_w29409_,
		_w29815_,
		_w29814_,
		_w29816_,
		_w29817_
	);
	LUT2 #(
		.INIT('h1)
	) name23991 (
		_w29396_,
		_w29817_,
		_w29818_
	);
	LUT4 #(
		.INIT('h4060)
	) name23992 (
		_w29398_,
		_w29399_,
		_w29400_,
		_w29402_,
		_w29819_
	);
	LUT3 #(
		.INIT('ha8)
	) name23993 (
		_w29396_,
		_w29419_,
		_w29819_,
		_w29820_
	);
	LUT3 #(
		.INIT('hb8)
	) name23994 (
		_w29397_,
		_w29398_,
		_w29399_,
		_w29821_
	);
	LUT2 #(
		.INIT('h8)
	) name23995 (
		_w29396_,
		_w29402_,
		_w29822_
	);
	LUT4 #(
		.INIT('h4544)
	) name23996 (
		_w29400_,
		_w29404_,
		_w29821_,
		_w29822_,
		_w29823_
	);
	LUT4 #(
		.INIT('h80b0)
	) name23997 (
		_w29397_,
		_w29398_,
		_w29400_,
		_w29402_,
		_w29824_
	);
	LUT2 #(
		.INIT('h4)
	) name23998 (
		_w29815_,
		_w29824_,
		_w29825_
	);
	LUT3 #(
		.INIT('h01)
	) name23999 (
		_w29823_,
		_w29820_,
		_w29825_,
		_w29826_
	);
	LUT3 #(
		.INIT('h65)
	) name24000 (
		\u0_L6_reg[18]/NET0131 ,
		_w29818_,
		_w29826_,
		_w29827_
	);
	LUT3 #(
		.INIT('h80)
	) name24001 (
		_w29745_,
		_w29746_,
		_w29750_,
		_w29828_
	);
	LUT4 #(
		.INIT('h3dc3)
	) name24002 (
		_w29748_,
		_w29745_,
		_w29746_,
		_w29750_,
		_w29829_
	);
	LUT4 #(
		.INIT('h0104)
	) name24003 (
		_w29748_,
		_w29745_,
		_w29746_,
		_w29749_,
		_w29830_
	);
	LUT4 #(
		.INIT('h0302)
	) name24004 (
		_w29749_,
		_w29758_,
		_w29830_,
		_w29829_,
		_w29831_
	);
	LUT4 #(
		.INIT('h76ba)
	) name24005 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29832_
	);
	LUT4 #(
		.INIT('h2880)
	) name24006 (
		_w29748_,
		_w29745_,
		_w29746_,
		_w29750_,
		_w29833_
	);
	LUT4 #(
		.INIT('h00f2)
	) name24007 (
		_w29748_,
		_w29770_,
		_w29832_,
		_w29833_,
		_w29834_
	);
	LUT4 #(
		.INIT('hdfef)
	) name24008 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29835_
	);
	LUT4 #(
		.INIT('h0040)
	) name24009 (
		_w29748_,
		_w29745_,
		_w29749_,
		_w29750_,
		_w29836_
	);
	LUT3 #(
		.INIT('h0d)
	) name24010 (
		_w29748_,
		_w29835_,
		_w29836_,
		_w29837_
	);
	LUT4 #(
		.INIT('hd800)
	) name24011 (
		_w29755_,
		_w29831_,
		_w29834_,
		_w29837_,
		_w29838_
	);
	LUT2 #(
		.INIT('h9)
	) name24012 (
		\u0_L6_reg[16]/NET0131 ,
		_w29838_,
		_w29839_
	);
	LUT3 #(
		.INIT('h15)
	) name24013 (
		_w29748_,
		_w29745_,
		_w29749_,
		_w29840_
	);
	LUT3 #(
		.INIT('h10)
	) name24014 (
		_w29745_,
		_w29746_,
		_w29750_,
		_w29841_
	);
	LUT4 #(
		.INIT('ha88a)
	) name24015 (
		_w29748_,
		_w29745_,
		_w29746_,
		_w29749_,
		_w29842_
	);
	LUT4 #(
		.INIT('h0002)
	) name24016 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29843_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name24017 (
		_w29840_,
		_w29841_,
		_w29842_,
		_w29843_,
		_w29844_
	);
	LUT2 #(
		.INIT('h2)
	) name24018 (
		_w29755_,
		_w29844_,
		_w29845_
	);
	LUT4 #(
		.INIT('h7c5f)
	) name24019 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29846_
	);
	LUT2 #(
		.INIT('h2)
	) name24020 (
		_w29748_,
		_w29846_,
		_w29847_
	);
	LUT4 #(
		.INIT('h0040)
	) name24021 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29848_
	);
	LUT2 #(
		.INIT('h1)
	) name24022 (
		_w29755_,
		_w29848_,
		_w29849_
	);
	LUT4 #(
		.INIT('h0009)
	) name24023 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29850_
	);
	LUT3 #(
		.INIT('hca)
	) name24024 (
		_w29745_,
		_w29746_,
		_w29750_,
		_w29851_
	);
	LUT3 #(
		.INIT('h13)
	) name24025 (
		_w29840_,
		_w29850_,
		_w29851_,
		_w29852_
	);
	LUT3 #(
		.INIT('h40)
	) name24026 (
		_w29847_,
		_w29849_,
		_w29852_,
		_w29853_
	);
	LUT2 #(
		.INIT('h8)
	) name24027 (
		_w29748_,
		_w29745_,
		_w29854_
	);
	LUT2 #(
		.INIT('h8)
	) name24028 (
		_w29769_,
		_w29854_,
		_w29855_
	);
	LUT2 #(
		.INIT('h4)
	) name24029 (
		_w29748_,
		_w29749_,
		_w29856_
	);
	LUT4 #(
		.INIT('h1000)
	) name24030 (
		_w29748_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29857_
	);
	LUT3 #(
		.INIT('h70)
	) name24031 (
		_w29745_,
		_w29746_,
		_w29755_,
		_w29858_
	);
	LUT3 #(
		.INIT('h13)
	) name24032 (
		_w29753_,
		_w29857_,
		_w29858_,
		_w29859_
	);
	LUT2 #(
		.INIT('h4)
	) name24033 (
		_w29855_,
		_w29859_,
		_w29860_
	);
	LUT4 #(
		.INIT('h56aa)
	) name24034 (
		\u0_L6_reg[30]/NET0131 ,
		_w29845_,
		_w29853_,
		_w29860_,
		_w29861_
	);
	LUT4 #(
		.INIT('hffd6)
	) name24035 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29862_
	);
	LUT3 #(
		.INIT('h40)
	) name24036 (
		_w29748_,
		_w29767_,
		_w29862_,
		_w29863_
	);
	LUT4 #(
		.INIT('hee5f)
	) name24037 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29864_
	);
	LUT2 #(
		.INIT('h8)
	) name24038 (
		_w29842_,
		_w29864_,
		_w29865_
	);
	LUT3 #(
		.INIT('h54)
	) name24039 (
		_w29755_,
		_w29863_,
		_w29865_,
		_w29866_
	);
	LUT2 #(
		.INIT('h2)
	) name24040 (
		_w29748_,
		_w29749_,
		_w29867_
	);
	LUT3 #(
		.INIT('h0b)
	) name24041 (
		_w29745_,
		_w29746_,
		_w29750_,
		_w29868_
	);
	LUT2 #(
		.INIT('h8)
	) name24042 (
		_w29867_,
		_w29868_,
		_w29869_
	);
	LUT3 #(
		.INIT('h70)
	) name24043 (
		_w29747_,
		_w29751_,
		_w29755_,
		_w29870_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name24044 (
		_w29745_,
		_w29746_,
		_w29749_,
		_w29750_,
		_w29871_
	);
	LUT3 #(
		.INIT('hb1)
	) name24045 (
		_w29748_,
		_w29759_,
		_w29871_,
		_w29872_
	);
	LUT3 #(
		.INIT('h40)
	) name24046 (
		_w29869_,
		_w29870_,
		_w29872_,
		_w29873_
	);
	LUT4 #(
		.INIT('h002a)
	) name24047 (
		_w29748_,
		_w29745_,
		_w29746_,
		_w29749_,
		_w29874_
	);
	LUT4 #(
		.INIT('h135f)
	) name24048 (
		_w29828_,
		_w29851_,
		_w29856_,
		_w29874_,
		_w29875_
	);
	LUT4 #(
		.INIT('ha955)
	) name24049 (
		\u0_L6_reg[24]/NET0131 ,
		_w29866_,
		_w29873_,
		_w29875_,
		_w29876_
	);
	LUT4 #(
		.INIT('hc693)
	) name24050 (
		decrypt_pad,
		\u0_R5_reg[28]/NET0131 ,
		\u0_uk_K_r5_reg[44]/NET0131 ,
		\u0_uk_K_r5_reg[9]/NET0131 ,
		_w29877_
	);
	LUT4 #(
		.INIT('hc963)
	) name24051 (
		decrypt_pad,
		\u0_R5_reg[27]/NET0131 ,
		\u0_uk_K_r5_reg[22]/NET0131 ,
		\u0_uk_K_r5_reg[2]/NET0131 ,
		_w29878_
	);
	LUT4 #(
		.INIT('hc693)
	) name24052 (
		decrypt_pad,
		\u0_R5_reg[24]/NET0131 ,
		\u0_uk_K_r5_reg[28]/NET0131 ,
		\u0_uk_K_r5_reg[52]/NET0131 ,
		_w29879_
	);
	LUT4 #(
		.INIT('hc963)
	) name24053 (
		decrypt_pad,
		\u0_R5_reg[26]/NET0131 ,
		\u0_uk_K_r5_reg[44]/NET0131 ,
		\u0_uk_K_r5_reg[52]/NET0131 ,
		_w29880_
	);
	LUT4 #(
		.INIT('hc963)
	) name24054 (
		decrypt_pad,
		\u0_R5_reg[29]/NET0131 ,
		\u0_uk_K_r5_reg[1]/NET0131 ,
		\u0_uk_K_r5_reg[36]/NET0131 ,
		_w29881_
	);
	LUT4 #(
		.INIT('hc963)
	) name24055 (
		decrypt_pad,
		\u0_R5_reg[25]/NET0131 ,
		\u0_uk_K_r5_reg[28]/NET0131 ,
		\u0_uk_K_r5_reg[8]/NET0131 ,
		_w29882_
	);
	LUT4 #(
		.INIT('h0004)
	) name24056 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w29883_
	);
	LUT4 #(
		.INIT('h757b)
	) name24057 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w29884_
	);
	LUT2 #(
		.INIT('h1)
	) name24058 (
		_w29878_,
		_w29884_,
		_w29885_
	);
	LUT2 #(
		.INIT('h1)
	) name24059 (
		_w29880_,
		_w29882_,
		_w29886_
	);
	LUT3 #(
		.INIT('h5d)
	) name24060 (
		_w29879_,
		_w29881_,
		_w29878_,
		_w29887_
	);
	LUT2 #(
		.INIT('h4)
	) name24061 (
		_w29879_,
		_w29881_,
		_w29888_
	);
	LUT4 #(
		.INIT('h0010)
	) name24062 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29878_,
		_w29889_
	);
	LUT2 #(
		.INIT('h6)
	) name24063 (
		_w29879_,
		_w29880_,
		_w29890_
	);
	LUT4 #(
		.INIT('h9000)
	) name24064 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w29891_
	);
	LUT4 #(
		.INIT('h0301)
	) name24065 (
		_w29886_,
		_w29889_,
		_w29891_,
		_w29887_,
		_w29892_
	);
	LUT3 #(
		.INIT('h45)
	) name24066 (
		_w29877_,
		_w29885_,
		_w29892_,
		_w29893_
	);
	LUT4 #(
		.INIT('hafdf)
	) name24067 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w29894_
	);
	LUT2 #(
		.INIT('h1)
	) name24068 (
		_w29878_,
		_w29894_,
		_w29895_
	);
	LUT2 #(
		.INIT('h6)
	) name24069 (
		_w29880_,
		_w29882_,
		_w29896_
	);
	LUT4 #(
		.INIT('ha800)
	) name24070 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29878_,
		_w29897_
	);
	LUT4 #(
		.INIT('h0040)
	) name24071 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w29898_
	);
	LUT4 #(
		.INIT('hffbe)
	) name24072 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w29899_
	);
	LUT3 #(
		.INIT('h70)
	) name24073 (
		_w29896_,
		_w29897_,
		_w29899_,
		_w29900_
	);
	LUT4 #(
		.INIT('hfbb5)
	) name24074 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w29901_
	);
	LUT4 #(
		.INIT('h0100)
	) name24075 (
		_w29880_,
		_w29881_,
		_w29882_,
		_w29878_,
		_w29902_
	);
	LUT4 #(
		.INIT('h0090)
	) name24076 (
		_w29879_,
		_w29880_,
		_w29882_,
		_w29878_,
		_w29903_
	);
	LUT4 #(
		.INIT('h0301)
	) name24077 (
		_w29878_,
		_w29902_,
		_w29903_,
		_w29901_,
		_w29904_
	);
	LUT4 #(
		.INIT('h7500)
	) name24078 (
		_w29877_,
		_w29895_,
		_w29900_,
		_w29904_,
		_w29905_
	);
	LUT3 #(
		.INIT('h65)
	) name24079 (
		\u0_L5_reg[22]/NET0131 ,
		_w29893_,
		_w29905_,
		_w29906_
	);
	LUT4 #(
		.INIT('hc693)
	) name24080 (
		decrypt_pad,
		\u0_R5_reg[4]/NET0131 ,
		\u0_uk_K_r5_reg[11]/NET0131 ,
		\u0_uk_K_r5_reg[33]/NET0131 ,
		_w29907_
	);
	LUT4 #(
		.INIT('hc963)
	) name24081 (
		decrypt_pad,
		\u0_R5_reg[32]/NET0131 ,
		\u0_uk_K_r5_reg[10]/NET0131 ,
		\u0_uk_K_r5_reg[20]/NET0131 ,
		_w29908_
	);
	LUT4 #(
		.INIT('hc693)
	) name24082 (
		decrypt_pad,
		\u0_R5_reg[1]/NET0131 ,
		\u0_uk_K_r5_reg[41]/NET0131 ,
		\u0_uk_K_r5_reg[6]/NET0131 ,
		_w29909_
	);
	LUT4 #(
		.INIT('hc693)
	) name24083 (
		decrypt_pad,
		\u0_R5_reg[2]/NET0131 ,
		\u0_uk_K_r5_reg[24]/NET0131 ,
		\u0_uk_K_r5_reg[46]/NET0131 ,
		_w29910_
	);
	LUT4 #(
		.INIT('hc693)
	) name24084 (
		decrypt_pad,
		\u0_R5_reg[5]/NET0131 ,
		\u0_uk_K_r5_reg[39]/NET0131 ,
		\u0_uk_K_r5_reg[4]/NET0131 ,
		_w29911_
	);
	LUT4 #(
		.INIT('hfe00)
	) name24085 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w29912_
	);
	LUT2 #(
		.INIT('h1)
	) name24086 (
		_w29911_,
		_w29908_,
		_w29913_
	);
	LUT4 #(
		.INIT('hc693)
	) name24087 (
		decrypt_pad,
		\u0_R5_reg[3]/NET0131 ,
		\u0_uk_K_r5_reg[33]/NET0131 ,
		\u0_uk_K_r5_reg[55]/NET0131 ,
		_w29914_
	);
	LUT2 #(
		.INIT('h2)
	) name24088 (
		_w29914_,
		_w29910_,
		_w29915_
	);
	LUT3 #(
		.INIT('ha2)
	) name24089 (
		_w29909_,
		_w29914_,
		_w29910_,
		_w29916_
	);
	LUT3 #(
		.INIT('h01)
	) name24090 (
		_w29913_,
		_w29916_,
		_w29912_,
		_w29917_
	);
	LUT4 #(
		.INIT('hafa3)
	) name24091 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w29918_
	);
	LUT4 #(
		.INIT('h2250)
	) name24092 (
		_w29909_,
		_w29914_,
		_w29910_,
		_w29908_,
		_w29919_
	);
	LUT3 #(
		.INIT('h0d)
	) name24093 (
		_w29914_,
		_w29918_,
		_w29919_,
		_w29920_
	);
	LUT3 #(
		.INIT('h8a)
	) name24094 (
		_w29907_,
		_w29917_,
		_w29920_,
		_w29921_
	);
	LUT4 #(
		.INIT('hfbdc)
	) name24095 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w29922_
	);
	LUT2 #(
		.INIT('h1)
	) name24096 (
		_w29914_,
		_w29922_,
		_w29923_
	);
	LUT2 #(
		.INIT('h8)
	) name24097 (
		_w29914_,
		_w29910_,
		_w29924_
	);
	LUT3 #(
		.INIT('h28)
	) name24098 (
		_w29909_,
		_w29911_,
		_w29908_,
		_w29925_
	);
	LUT4 #(
		.INIT('h2ff5)
	) name24099 (
		_w29909_,
		_w29914_,
		_w29911_,
		_w29908_,
		_w29926_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name24100 (
		_w29914_,
		_w29910_,
		_w29925_,
		_w29926_,
		_w29927_
	);
	LUT3 #(
		.INIT('h45)
	) name24101 (
		_w29907_,
		_w29923_,
		_w29927_,
		_w29928_
	);
	LUT4 #(
		.INIT('h8000)
	) name24102 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w29929_
	);
	LUT4 #(
		.INIT('h0040)
	) name24103 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w29930_
	);
	LUT4 #(
		.INIT('h7dbd)
	) name24104 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w29931_
	);
	LUT2 #(
		.INIT('h1)
	) name24105 (
		_w29914_,
		_w29931_,
		_w29932_
	);
	LUT3 #(
		.INIT('h40)
	) name24106 (
		_w29909_,
		_w29914_,
		_w29910_,
		_w29933_
	);
	LUT4 #(
		.INIT('h0400)
	) name24107 (
		_w29909_,
		_w29914_,
		_w29910_,
		_w29908_,
		_w29934_
	);
	LUT3 #(
		.INIT('h07)
	) name24108 (
		_w29913_,
		_w29933_,
		_w29934_,
		_w29935_
	);
	LUT2 #(
		.INIT('h4)
	) name24109 (
		_w29932_,
		_w29935_,
		_w29936_
	);
	LUT4 #(
		.INIT('h5655)
	) name24110 (
		\u0_L5_reg[31]/NET0131 ,
		_w29928_,
		_w29921_,
		_w29936_,
		_w29937_
	);
	LUT4 #(
		.INIT('hc963)
	) name24111 (
		decrypt_pad,
		\u0_R5_reg[24]/NET0131 ,
		\u0_uk_K_r5_reg[2]/NET0131 ,
		\u0_uk_K_r5_reg[37]/P0001 ,
		_w29938_
	);
	LUT4 #(
		.INIT('hc693)
	) name24112 (
		decrypt_pad,
		\u0_R5_reg[22]/NET0131 ,
		\u0_uk_K_r5_reg[22]/NET0131 ,
		\u0_uk_K_r5_reg[42]/NET0131 ,
		_w29939_
	);
	LUT4 #(
		.INIT('hc693)
	) name24113 (
		decrypt_pad,
		\u0_R5_reg[25]/NET0131 ,
		\u0_uk_K_r5_reg[1]/NET0131 ,
		\u0_uk_K_r5_reg[21]/NET0131 ,
		_w29940_
	);
	LUT4 #(
		.INIT('hc693)
	) name24114 (
		decrypt_pad,
		\u0_R5_reg[20]/NET0131 ,
		\u0_uk_K_r5_reg[16]/NET0131 ,
		\u0_uk_K_r5_reg[36]/NET0131 ,
		_w29941_
	);
	LUT4 #(
		.INIT('hc693)
	) name24115 (
		decrypt_pad,
		\u0_R5_reg[21]/NET0131 ,
		\u0_uk_K_r5_reg[0]/NET0131 ,
		\u0_uk_K_r5_reg[51]/NET0131 ,
		_w29942_
	);
	LUT4 #(
		.INIT('hb080)
	) name24116 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w29943_
	);
	LUT4 #(
		.INIT('hc963)
	) name24117 (
		decrypt_pad,
		\u0_R5_reg[23]/NET0131 ,
		\u0_uk_K_r5_reg[0]/NET0131 ,
		\u0_uk_K_r5_reg[35]/NET0131 ,
		_w29944_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name24118 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w29945_
	);
	LUT3 #(
		.INIT('h01)
	) name24119 (
		_w29944_,
		_w29945_,
		_w29943_,
		_w29946_
	);
	LUT4 #(
		.INIT('h0004)
	) name24120 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w29947_
	);
	LUT4 #(
		.INIT('h47fb)
	) name24121 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w29948_
	);
	LUT4 #(
		.INIT('h0008)
	) name24122 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29944_,
		_w29949_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name24123 (
		_w29942_,
		_w29944_,
		_w29948_,
		_w29949_,
		_w29950_
	);
	LUT3 #(
		.INIT('h8a)
	) name24124 (
		_w29938_,
		_w29946_,
		_w29950_,
		_w29951_
	);
	LUT4 #(
		.INIT('h0060)
	) name24125 (
		_w29941_,
		_w29939_,
		_w29942_,
		_w29944_,
		_w29952_
	);
	LUT2 #(
		.INIT('h8)
	) name24126 (
		_w29939_,
		_w29944_,
		_w29953_
	);
	LUT4 #(
		.INIT('h0800)
	) name24127 (
		_w29941_,
		_w29939_,
		_w29942_,
		_w29944_,
		_w29954_
	);
	LUT4 #(
		.INIT('h0400)
	) name24128 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w29955_
	);
	LUT4 #(
		.INIT('h0004)
	) name24129 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29944_,
		_w29956_
	);
	LUT4 #(
		.INIT('hfcfb)
	) name24130 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29944_,
		_w29957_
	);
	LUT3 #(
		.INIT('h10)
	) name24131 (
		_w29954_,
		_w29955_,
		_w29957_,
		_w29958_
	);
	LUT4 #(
		.INIT('h0200)
	) name24132 (
		_w29940_,
		_w29941_,
		_w29942_,
		_w29944_,
		_w29959_
	);
	LUT4 #(
		.INIT('h0080)
	) name24133 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w29960_
	);
	LUT2 #(
		.INIT('h1)
	) name24134 (
		_w29959_,
		_w29960_,
		_w29961_
	);
	LUT4 #(
		.INIT('h4555)
	) name24135 (
		_w29938_,
		_w29952_,
		_w29958_,
		_w29961_,
		_w29962_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name24136 (
		_w29940_,
		_w29941_,
		_w29942_,
		_w29944_,
		_w29963_
	);
	LUT2 #(
		.INIT('h1)
	) name24137 (
		_w29939_,
		_w29963_,
		_w29964_
	);
	LUT4 #(
		.INIT('h0100)
	) name24138 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w29965_
	);
	LUT4 #(
		.INIT('h7e7f)
	) name24139 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w29966_
	);
	LUT3 #(
		.INIT('h01)
	) name24140 (
		_w29940_,
		_w29941_,
		_w29942_,
		_w29967_
	);
	LUT4 #(
		.INIT('hcacf)
	) name24141 (
		_w29939_,
		_w29966_,
		_w29944_,
		_w29967_,
		_w29968_
	);
	LUT2 #(
		.INIT('h4)
	) name24142 (
		_w29964_,
		_w29968_,
		_w29969_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name24143 (
		\u0_L5_reg[11]/NET0131 ,
		_w29962_,
		_w29951_,
		_w29969_,
		_w29970_
	);
	LUT4 #(
		.INIT('hc963)
	) name24144 (
		decrypt_pad,
		\u0_R5_reg[14]/NET0131 ,
		\u0_uk_K_r5_reg[19]/NET0131 ,
		\u0_uk_K_r5_reg[54]/NET0131 ,
		_w29971_
	);
	LUT4 #(
		.INIT('hc963)
	) name24145 (
		decrypt_pad,
		\u0_R5_reg[13]/NET0131 ,
		\u0_uk_K_r5_reg[18]/NET0131 ,
		\u0_uk_K_r5_reg[53]/NET0131 ,
		_w29972_
	);
	LUT4 #(
		.INIT('hc963)
	) name24146 (
		decrypt_pad,
		\u0_R5_reg[12]/NET0131 ,
		\u0_uk_K_r5_reg[24]/NET0131 ,
		\u0_uk_K_r5_reg[34]/NET0131 ,
		_w29973_
	);
	LUT4 #(
		.INIT('hc693)
	) name24147 (
		decrypt_pad,
		\u0_R5_reg[17]/NET0131 ,
		\u0_uk_K_r5_reg[18]/NET0131 ,
		\u0_uk_K_r5_reg[40]/NET0131 ,
		_w29974_
	);
	LUT4 #(
		.INIT('h8000)
	) name24148 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29975_
	);
	LUT4 #(
		.INIT('hc963)
	) name24149 (
		decrypt_pad,
		\u0_R5_reg[15]/NET0131 ,
		\u0_uk_K_r5_reg[27]/NET0131 ,
		\u0_uk_K_r5_reg[5]/NET0131 ,
		_w29976_
	);
	LUT2 #(
		.INIT('h4)
	) name24150 (
		_w29973_,
		_w29974_,
		_w29977_
	);
	LUT4 #(
		.INIT('h0200)
	) name24151 (
		_w29976_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29978_
	);
	LUT4 #(
		.INIT('h0080)
	) name24152 (
		_w29976_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29979_
	);
	LUT4 #(
		.INIT('h0400)
	) name24153 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29980_
	);
	LUT4 #(
		.INIT('h0001)
	) name24154 (
		_w29978_,
		_w29979_,
		_w29980_,
		_w29975_,
		_w29981_
	);
	LUT4 #(
		.INIT('h0001)
	) name24155 (
		_w29976_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29982_
	);
	LUT4 #(
		.INIT('h0110)
	) name24156 (
		_w29976_,
		_w29971_,
		_w29972_,
		_w29973_,
		_w29983_
	);
	LUT4 #(
		.INIT('hc693)
	) name24157 (
		decrypt_pad,
		\u0_R5_reg[16]/NET0131 ,
		\u0_uk_K_r5_reg[13]/P0001 ,
		\u0_uk_K_r5_reg[3]/NET0131 ,
		_w29984_
	);
	LUT4 #(
		.INIT('h1030)
	) name24158 (
		_w29971_,
		_w29983_,
		_w29984_,
		_w29982_,
		_w29985_
	);
	LUT2 #(
		.INIT('h8)
	) name24159 (
		_w29981_,
		_w29985_,
		_w29986_
	);
	LUT4 #(
		.INIT('haaa8)
	) name24160 (
		_w29976_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29987_
	);
	LUT4 #(
		.INIT('h2aa8)
	) name24161 (
		_w29976_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29988_
	);
	LUT3 #(
		.INIT('h08)
	) name24162 (
		_w29971_,
		_w29973_,
		_w29974_,
		_w29989_
	);
	LUT3 #(
		.INIT('h45)
	) name24163 (
		_w29976_,
		_w29972_,
		_w29974_,
		_w29990_
	);
	LUT3 #(
		.INIT('h45)
	) name24164 (
		_w29988_,
		_w29989_,
		_w29990_,
		_w29991_
	);
	LUT4 #(
		.INIT('h1000)
	) name24165 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29992_
	);
	LUT4 #(
		.INIT('h0001)
	) name24166 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29993_
	);
	LUT3 #(
		.INIT('h01)
	) name24167 (
		_w29984_,
		_w29993_,
		_w29992_,
		_w29994_
	);
	LUT3 #(
		.INIT('h80)
	) name24168 (
		_w29976_,
		_w29971_,
		_w29972_,
		_w29995_
	);
	LUT4 #(
		.INIT('h0080)
	) name24169 (
		_w29976_,
		_w29971_,
		_w29972_,
		_w29973_,
		_w29996_
	);
	LUT3 #(
		.INIT('h02)
	) name24170 (
		_w29972_,
		_w29973_,
		_w29974_,
		_w29997_
	);
	LUT4 #(
		.INIT('h0008)
	) name24171 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w29998_
	);
	LUT2 #(
		.INIT('h1)
	) name24172 (
		_w29996_,
		_w29998_,
		_w29999_
	);
	LUT3 #(
		.INIT('h40)
	) name24173 (
		_w29991_,
		_w29994_,
		_w29999_,
		_w30000_
	);
	LUT4 #(
		.INIT('h0020)
	) name24174 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30001_
	);
	LUT4 #(
		.INIT('heee4)
	) name24175 (
		_w29976_,
		_w29980_,
		_w29993_,
		_w30001_,
		_w30002_
	);
	LUT2 #(
		.INIT('h4)
	) name24176 (
		_w29971_,
		_w29979_,
		_w30003_
	);
	LUT2 #(
		.INIT('h1)
	) name24177 (
		_w30002_,
		_w30003_,
		_w30004_
	);
	LUT4 #(
		.INIT('ha955)
	) name24178 (
		\u0_L5_reg[20]/NET0131 ,
		_w29986_,
		_w30000_,
		_w30004_,
		_w30005_
	);
	LUT4 #(
		.INIT('hc693)
	) name24179 (
		decrypt_pad,
		\u0_R5_reg[28]/NET0131 ,
		\u0_uk_K_r5_reg[42]/NET0131 ,
		\u0_uk_K_r5_reg[7]/NET0131 ,
		_w30006_
	);
	LUT4 #(
		.INIT('hc693)
	) name24180 (
		decrypt_pad,
		\u0_R5_reg[30]/NET0131 ,
		\u0_uk_K_r5_reg[15]/NET0131 ,
		\u0_uk_K_r5_reg[35]/NET0131 ,
		_w30007_
	);
	LUT4 #(
		.INIT('hc693)
	) name24181 (
		decrypt_pad,
		\u0_R5_reg[29]/NET0131 ,
		\u0_uk_K_r5_reg[14]/NET0131 ,
		\u0_uk_K_r5_reg[38]/NET0131 ,
		_w30008_
	);
	LUT4 #(
		.INIT('hc693)
	) name24182 (
		decrypt_pad,
		\u0_R5_reg[1]/NET0131 ,
		\u0_uk_K_r5_reg[30]/NET0131 ,
		\u0_uk_K_r5_reg[50]/NET0131 ,
		_w30009_
	);
	LUT4 #(
		.INIT('hc963)
	) name24183 (
		decrypt_pad,
		\u0_R5_reg[31]/P0001 ,
		\u0_uk_K_r5_reg[23]/NET0131 ,
		\u0_uk_K_r5_reg[31]/NET0131 ,
		_w30010_
	);
	LUT2 #(
		.INIT('h1)
	) name24184 (
		_w30007_,
		_w30010_,
		_w30011_
	);
	LUT4 #(
		.INIT('h7d4c)
	) name24185 (
		_w30008_,
		_w30007_,
		_w30009_,
		_w30010_,
		_w30012_
	);
	LUT2 #(
		.INIT('h2)
	) name24186 (
		_w30006_,
		_w30012_,
		_w30013_
	);
	LUT4 #(
		.INIT('h0020)
	) name24187 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30014_
	);
	LUT4 #(
		.INIT('heedf)
	) name24188 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30015_
	);
	LUT3 #(
		.INIT('h0b)
	) name24189 (
		_w30006_,
		_w30007_,
		_w30009_,
		_w30016_
	);
	LUT3 #(
		.INIT('h0b)
	) name24190 (
		_w30008_,
		_w30009_,
		_w30010_,
		_w30017_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name24191 (
		_w30015_,
		_w30010_,
		_w30016_,
		_w30017_,
		_w30018_
	);
	LUT4 #(
		.INIT('hc963)
	) name24192 (
		decrypt_pad,
		\u0_R5_reg[32]/NET0131 ,
		\u0_uk_K_r5_reg[29]/NET0131 ,
		\u0_uk_K_r5_reg[9]/NET0131 ,
		_w30019_
	);
	LUT3 #(
		.INIT('h0b)
	) name24193 (
		_w30013_,
		_w30018_,
		_w30019_,
		_w30020_
	);
	LUT4 #(
		.INIT('h0008)
	) name24194 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30021_
	);
	LUT4 #(
		.INIT('hf531)
	) name24195 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30022_
	);
	LUT3 #(
		.INIT('h02)
	) name24196 (
		_w30010_,
		_w30022_,
		_w30021_,
		_w30023_
	);
	LUT4 #(
		.INIT('h4000)
	) name24197 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30024_
	);
	LUT4 #(
		.INIT('h0001)
	) name24198 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30010_,
		_w30025_
	);
	LUT2 #(
		.INIT('h1)
	) name24199 (
		_w30024_,
		_w30025_,
		_w30026_
	);
	LUT3 #(
		.INIT('h8a)
	) name24200 (
		_w30019_,
		_w30023_,
		_w30026_,
		_w30027_
	);
	LUT4 #(
		.INIT('h0240)
	) name24201 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30028_
	);
	LUT4 #(
		.INIT('h0001)
	) name24202 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30029_
	);
	LUT4 #(
		.INIT('h1000)
	) name24203 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30030_
	);
	LUT4 #(
		.INIT('hedbe)
	) name24204 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30031_
	);
	LUT2 #(
		.INIT('h2)
	) name24205 (
		_w30010_,
		_w30031_,
		_w30032_
	);
	LUT3 #(
		.INIT('h08)
	) name24206 (
		_w30006_,
		_w30008_,
		_w30009_,
		_w30033_
	);
	LUT3 #(
		.INIT('h20)
	) name24207 (
		_w30006_,
		_w30008_,
		_w30019_,
		_w30034_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24208 (
		_w30007_,
		_w30010_,
		_w30033_,
		_w30034_,
		_w30035_
	);
	LUT2 #(
		.INIT('h4)
	) name24209 (
		_w30032_,
		_w30035_,
		_w30036_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name24210 (
		\u0_L5_reg[5]/NET0131 ,
		_w30020_,
		_w30027_,
		_w30036_,
		_w30037_
	);
	LUT4 #(
		.INIT('h48cc)
	) name24211 (
		_w29909_,
		_w29914_,
		_w29911_,
		_w29908_,
		_w30038_
	);
	LUT3 #(
		.INIT('h41)
	) name24212 (
		_w29909_,
		_w29911_,
		_w29908_,
		_w30039_
	);
	LUT4 #(
		.INIT('h5554)
	) name24213 (
		_w29914_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30040_
	);
	LUT3 #(
		.INIT('h45)
	) name24214 (
		_w30038_,
		_w30039_,
		_w30040_,
		_w30041_
	);
	LUT4 #(
		.INIT('h0800)
	) name24215 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30042_
	);
	LUT3 #(
		.INIT('h01)
	) name24216 (
		_w29907_,
		_w29930_,
		_w30042_,
		_w30043_
	);
	LUT4 #(
		.INIT('h1000)
	) name24217 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30044_
	);
	LUT4 #(
		.INIT('hef11)
	) name24218 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30045_
	);
	LUT2 #(
		.INIT('h2)
	) name24219 (
		_w29914_,
		_w30045_,
		_w30046_
	);
	LUT4 #(
		.INIT('h0200)
	) name24220 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30047_
	);
	LUT4 #(
		.INIT('h3001)
	) name24221 (
		_w29909_,
		_w29914_,
		_w29910_,
		_w29908_,
		_w30048_
	);
	LUT4 #(
		.INIT('h7f00)
	) name24222 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29907_,
		_w30049_
	);
	LUT3 #(
		.INIT('h10)
	) name24223 (
		_w30048_,
		_w30047_,
		_w30049_,
		_w30050_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name24224 (
		_w30041_,
		_w30043_,
		_w30046_,
		_w30050_,
		_w30051_
	);
	LUT3 #(
		.INIT('h08)
	) name24225 (
		_w29909_,
		_w29914_,
		_w29908_,
		_w30052_
	);
	LUT2 #(
		.INIT('h6)
	) name24226 (
		_w29910_,
		_w29911_,
		_w30053_
	);
	LUT2 #(
		.INIT('h8)
	) name24227 (
		_w30052_,
		_w30053_,
		_w30054_
	);
	LUT3 #(
		.INIT('h56)
	) name24228 (
		\u0_L5_reg[17]/NET0131 ,
		_w30051_,
		_w30054_,
		_w30055_
	);
	LUT4 #(
		.INIT('h67ba)
	) name24229 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30056_
	);
	LUT4 #(
		.INIT('hb4f7)
	) name24230 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30057_
	);
	LUT4 #(
		.INIT('h0020)
	) name24231 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30058_
	);
	LUT4 #(
		.INIT('h00e4)
	) name24232 (
		_w29944_,
		_w30057_,
		_w30056_,
		_w30058_,
		_w30059_
	);
	LUT2 #(
		.INIT('h1)
	) name24233 (
		_w29938_,
		_w30059_,
		_w30060_
	);
	LUT4 #(
		.INIT('h6f6e)
	) name24234 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30061_
	);
	LUT2 #(
		.INIT('h1)
	) name24235 (
		_w29944_,
		_w30061_,
		_w30062_
	);
	LUT4 #(
		.INIT('h9cff)
	) name24236 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30063_
	);
	LUT2 #(
		.INIT('h2)
	) name24237 (
		_w29944_,
		_w30063_,
		_w30064_
	);
	LUT4 #(
		.INIT('h0012)
	) name24238 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30065_
	);
	LUT3 #(
		.INIT('h01)
	) name24239 (
		_w29960_,
		_w29956_,
		_w30065_,
		_w30066_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name24240 (
		_w29938_,
		_w30064_,
		_w30062_,
		_w30066_,
		_w30067_
	);
	LUT4 #(
		.INIT('h2000)
	) name24241 (
		_w29940_,
		_w29939_,
		_w29942_,
		_w29944_,
		_w30068_
	);
	LUT2 #(
		.INIT('h1)
	) name24242 (
		_w29947_,
		_w30068_,
		_w30069_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name24243 (
		\u0_L5_reg[29]/NET0131 ,
		_w30067_,
		_w30060_,
		_w30069_,
		_w30070_
	);
	LUT4 #(
		.INIT('hc693)
	) name24244 (
		decrypt_pad,
		\u0_R5_reg[8]/NET0131 ,
		\u0_uk_K_r5_reg[12]/NET0131 ,
		\u0_uk_K_r5_reg[34]/NET0131 ,
		_w30071_
	);
	LUT4 #(
		.INIT('hc963)
	) name24245 (
		decrypt_pad,
		\u0_R5_reg[7]/NET0131 ,
		\u0_uk_K_r5_reg[11]/NET0131 ,
		\u0_uk_K_r5_reg[46]/NET0131 ,
		_w30072_
	);
	LUT4 #(
		.INIT('hc963)
	) name24246 (
		decrypt_pad,
		\u0_R5_reg[5]/NET0131 ,
		\u0_uk_K_r5_reg[26]/NET0131 ,
		\u0_uk_K_r5_reg[4]/NET0131 ,
		_w30073_
	);
	LUT4 #(
		.INIT('hc693)
	) name24247 (
		decrypt_pad,
		\u0_R5_reg[4]/NET0131 ,
		\u0_uk_K_r5_reg[25]/NET0131 ,
		\u0_uk_K_r5_reg[47]/NET0131 ,
		_w30074_
	);
	LUT4 #(
		.INIT('hc693)
	) name24248 (
		decrypt_pad,
		\u0_R5_reg[9]/NET0131 ,
		\u0_uk_K_r5_reg[17]/NET0131 ,
		\u0_uk_K_r5_reg[39]/NET0131 ,
		_w30075_
	);
	LUT4 #(
		.INIT('hc963)
	) name24249 (
		decrypt_pad,
		\u0_R5_reg[6]/NET0131 ,
		\u0_uk_K_r5_reg[17]/NET0131 ,
		\u0_uk_K_r5_reg[27]/NET0131 ,
		_w30076_
	);
	LUT3 #(
		.INIT('h5d)
	) name24250 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30077_
	);
	LUT4 #(
		.INIT('h59fb)
	) name24251 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30078_
	);
	LUT2 #(
		.INIT('h1)
	) name24252 (
		_w30072_,
		_w30078_,
		_w30079_
	);
	LUT4 #(
		.INIT('h0034)
	) name24253 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30080_
	);
	LUT4 #(
		.INIT('h0800)
	) name24254 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30081_
	);
	LUT2 #(
		.INIT('h2)
	) name24255 (
		_w30075_,
		_w30076_,
		_w30082_
	);
	LUT4 #(
		.INIT('h0004)
	) name24256 (
		_w30072_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30083_
	);
	LUT4 #(
		.INIT('h4000)
	) name24257 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30084_
	);
	LUT4 #(
		.INIT('h0007)
	) name24258 (
		_w30072_,
		_w30081_,
		_w30083_,
		_w30084_,
		_w30085_
	);
	LUT4 #(
		.INIT('h5455)
	) name24259 (
		_w30071_,
		_w30079_,
		_w30080_,
		_w30085_,
		_w30086_
	);
	LUT4 #(
		.INIT('h0002)
	) name24260 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30087_
	);
	LUT4 #(
		.INIT('h0001)
	) name24261 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30073_,
		_w30088_
	);
	LUT4 #(
		.INIT('h80a0)
	) name24262 (
		_w30072_,
		_w30074_,
		_w30073_,
		_w30076_,
		_w30089_
	);
	LUT3 #(
		.INIT('h01)
	) name24263 (
		_w30088_,
		_w30089_,
		_w30087_,
		_w30090_
	);
	LUT4 #(
		.INIT('h0080)
	) name24264 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30091_
	);
	LUT4 #(
		.INIT('h4500)
	) name24265 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30076_,
		_w30092_
	);
	LUT3 #(
		.INIT('h13)
	) name24266 (
		_w30077_,
		_w30091_,
		_w30092_,
		_w30093_
	);
	LUT4 #(
		.INIT('h4004)
	) name24267 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30094_
	);
	LUT3 #(
		.INIT('h10)
	) name24268 (
		_w30075_,
		_w30073_,
		_w30076_,
		_w30095_
	);
	LUT4 #(
		.INIT('h0100)
	) name24269 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30096_
	);
	LUT3 #(
		.INIT('h08)
	) name24270 (
		_w30074_,
		_w30073_,
		_w30076_,
		_w30097_
	);
	LUT4 #(
		.INIT('heee4)
	) name24271 (
		_w30072_,
		_w30094_,
		_w30097_,
		_w30096_,
		_w30098_
	);
	LUT4 #(
		.INIT('h00d5)
	) name24272 (
		_w30071_,
		_w30090_,
		_w30093_,
		_w30098_,
		_w30099_
	);
	LUT3 #(
		.INIT('h65)
	) name24273 (
		\u0_L5_reg[2]/NET0131 ,
		_w30086_,
		_w30099_,
		_w30100_
	);
	LUT3 #(
		.INIT('h02)
	) name24274 (
		_w29976_,
		_w29992_,
		_w29997_,
		_w30101_
	);
	LUT4 #(
		.INIT('h00b0)
	) name24275 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30102_
	);
	LUT3 #(
		.INIT('h01)
	) name24276 (
		_w29976_,
		_w29980_,
		_w30102_,
		_w30103_
	);
	LUT4 #(
		.INIT('h7dff)
	) name24277 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30104_
	);
	LUT4 #(
		.INIT('h02aa)
	) name24278 (
		_w29984_,
		_w30101_,
		_w30103_,
		_w30104_,
		_w30105_
	);
	LUT4 #(
		.INIT('h353c)
	) name24279 (
		_w29976_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30106_
	);
	LUT2 #(
		.INIT('h1)
	) name24280 (
		_w29971_,
		_w30106_,
		_w30107_
	);
	LUT4 #(
		.INIT('h1000)
	) name24281 (
		_w29976_,
		_w29971_,
		_w29973_,
		_w29974_,
		_w30108_
	);
	LUT2 #(
		.INIT('h1)
	) name24282 (
		_w29982_,
		_w30108_,
		_w30109_
	);
	LUT3 #(
		.INIT('hdc)
	) name24283 (
		_w29971_,
		_w29972_,
		_w29974_,
		_w30110_
	);
	LUT2 #(
		.INIT('h8)
	) name24284 (
		_w29976_,
		_w29973_,
		_w30111_
	);
	LUT3 #(
		.INIT('h45)
	) name24285 (
		_w29998_,
		_w30110_,
		_w30111_,
		_w30112_
	);
	LUT4 #(
		.INIT('h4555)
	) name24286 (
		_w29984_,
		_w30107_,
		_w30109_,
		_w30112_,
		_w30113_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name24287 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30114_
	);
	LUT2 #(
		.INIT('h1)
	) name24288 (
		_w29976_,
		_w30114_,
		_w30115_
	);
	LUT3 #(
		.INIT('h0b)
	) name24289 (
		_w29971_,
		_w29979_,
		_w29996_,
		_w30116_
	);
	LUT2 #(
		.INIT('h4)
	) name24290 (
		_w30115_,
		_w30116_,
		_w30117_
	);
	LUT4 #(
		.INIT('h5655)
	) name24291 (
		\u0_L5_reg[10]/NET0131 ,
		_w30105_,
		_w30113_,
		_w30117_,
		_w30118_
	);
	LUT4 #(
		.INIT('h0084)
	) name24292 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30119_
	);
	LUT3 #(
		.INIT('h47)
	) name24293 (
		_w29880_,
		_w29882_,
		_w29878_,
		_w30120_
	);
	LUT4 #(
		.INIT('h0051)
	) name24294 (
		_w29877_,
		_w29888_,
		_w30120_,
		_w30119_,
		_w30121_
	);
	LUT4 #(
		.INIT('h0770)
	) name24295 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30122_
	);
	LUT4 #(
		.INIT('h0102)
	) name24296 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30123_
	);
	LUT3 #(
		.INIT('h0e)
	) name24297 (
		_w29878_,
		_w30122_,
		_w30123_,
		_w30124_
	);
	LUT4 #(
		.INIT('h55fe)
	) name24298 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30125_
	);
	LUT2 #(
		.INIT('h2)
	) name24299 (
		_w29878_,
		_w30125_,
		_w30126_
	);
	LUT4 #(
		.INIT('hebd7)
	) name24300 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30127_
	);
	LUT4 #(
		.INIT('ha200)
	) name24301 (
		_w29877_,
		_w29898_,
		_w29878_,
		_w30127_,
		_w30128_
	);
	LUT4 #(
		.INIT('h7077)
	) name24302 (
		_w30121_,
		_w30124_,
		_w30126_,
		_w30128_,
		_w30129_
	);
	LUT2 #(
		.INIT('h6)
	) name24303 (
		\u0_L5_reg[12]/NET0131 ,
		_w30129_,
		_w30130_
	);
	LUT4 #(
		.INIT('hc963)
	) name24304 (
		decrypt_pad,
		\u0_R5_reg[20]/NET0131 ,
		\u0_uk_K_r5_reg[14]/NET0131 ,
		\u0_uk_K_r5_reg[49]/NET0131 ,
		_w30131_
	);
	LUT4 #(
		.INIT('hc693)
	) name24305 (
		decrypt_pad,
		\u0_R5_reg[18]/NET0131 ,
		\u0_uk_K_r5_reg[23]/NET0131 ,
		\u0_uk_K_r5_reg[43]/NET0131 ,
		_w30132_
	);
	LUT4 #(
		.INIT('hc963)
	) name24306 (
		decrypt_pad,
		\u0_R5_reg[19]/NET0131 ,
		\u0_uk_K_r5_reg[30]/NET0131 ,
		\u0_uk_K_r5_reg[38]/NET0131 ,
		_w30133_
	);
	LUT4 #(
		.INIT('hc963)
	) name24307 (
		decrypt_pad,
		\u0_R5_reg[21]/NET0131 ,
		\u0_uk_K_r5_reg[15]/NET0131 ,
		\u0_uk_K_r5_reg[50]/NET0131 ,
		_w30134_
	);
	LUT4 #(
		.INIT('hc693)
	) name24308 (
		decrypt_pad,
		\u0_R5_reg[17]/NET0131 ,
		\u0_uk_K_r5_reg[29]/NET0131 ,
		\u0_uk_K_r5_reg[49]/NET0131 ,
		_w30135_
	);
	LUT4 #(
		.INIT('hc963)
	) name24309 (
		decrypt_pad,
		\u0_R5_reg[16]/NET0131 ,
		\u0_uk_K_r5_reg[31]/NET0131 ,
		\u0_uk_K_r5_reg[7]/NET0131 ,
		_w30136_
	);
	LUT4 #(
		.INIT('h0040)
	) name24310 (
		_w30133_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30137_
	);
	LUT4 #(
		.INIT('hc3be)
	) name24311 (
		_w30133_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30138_
	);
	LUT2 #(
		.INIT('h1)
	) name24312 (
		_w30132_,
		_w30138_,
		_w30139_
	);
	LUT4 #(
		.INIT('h50b0)
	) name24313 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30140_
	);
	LUT4 #(
		.INIT('ha34f)
	) name24314 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30141_
	);
	LUT2 #(
		.INIT('h2)
	) name24315 (
		_w30133_,
		_w30141_,
		_w30142_
	);
	LUT3 #(
		.INIT('h80)
	) name24316 (
		_w30135_,
		_w30134_,
		_w30136_,
		_w30143_
	);
	LUT2 #(
		.INIT('h4)
	) name24317 (
		_w30133_,
		_w30132_,
		_w30144_
	);
	LUT4 #(
		.INIT('h0200)
	) name24318 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30145_
	);
	LUT3 #(
		.INIT('h07)
	) name24319 (
		_w30143_,
		_w30144_,
		_w30145_,
		_w30146_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name24320 (
		_w30131_,
		_w30142_,
		_w30139_,
		_w30146_,
		_w30147_
	);
	LUT4 #(
		.INIT('h4000)
	) name24321 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30148_
	);
	LUT4 #(
		.INIT('h0100)
	) name24322 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30149_
	);
	LUT4 #(
		.INIT('hb6c7)
	) name24323 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30150_
	);
	LUT2 #(
		.INIT('h1)
	) name24324 (
		_w30133_,
		_w30150_,
		_w30151_
	);
	LUT4 #(
		.INIT('h7077)
	) name24325 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30152_
	);
	LUT4 #(
		.INIT('h2004)
	) name24326 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30153_
	);
	LUT4 #(
		.INIT('h0f08)
	) name24327 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30154_
	);
	LUT4 #(
		.INIT('h3331)
	) name24328 (
		_w30133_,
		_w30153_,
		_w30140_,
		_w30154_,
		_w30155_
	);
	LUT4 #(
		.INIT('h0402)
	) name24329 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30156_
	);
	LUT4 #(
		.INIT('h0020)
	) name24330 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30157_
	);
	LUT4 #(
		.INIT('h0028)
	) name24331 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30158_
	);
	LUT3 #(
		.INIT('hd8)
	) name24332 (
		_w30133_,
		_w30156_,
		_w30158_,
		_w30159_
	);
	LUT4 #(
		.INIT('h00ba)
	) name24333 (
		_w30131_,
		_w30151_,
		_w30155_,
		_w30159_,
		_w30160_
	);
	LUT3 #(
		.INIT('h65)
	) name24334 (
		\u0_L5_reg[14]/NET0131 ,
		_w30147_,
		_w30160_,
		_w30161_
	);
	LUT4 #(
		.INIT('h7773)
	) name24335 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30162_
	);
	LUT4 #(
		.INIT('h6673)
	) name24336 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30163_
	);
	LUT4 #(
		.INIT('h0002)
	) name24337 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30164_
	);
	LUT4 #(
		.INIT('h3302)
	) name24338 (
		_w30010_,
		_w30019_,
		_w30163_,
		_w30164_,
		_w30165_
	);
	LUT4 #(
		.INIT('h0040)
	) name24339 (
		_w30008_,
		_w30007_,
		_w30009_,
		_w30010_,
		_w30166_
	);
	LUT4 #(
		.INIT('hf7b7)
	) name24340 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30167_
	);
	LUT4 #(
		.INIT('h0100)
	) name24341 (
		_w30006_,
		_w30008_,
		_w30009_,
		_w30010_,
		_w30168_
	);
	LUT4 #(
		.INIT('h2000)
	) name24342 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30169_
	);
	LUT4 #(
		.INIT('h0100)
	) name24343 (
		_w30168_,
		_w30166_,
		_w30169_,
		_w30167_,
		_w30170_
	);
	LUT3 #(
		.INIT('h02)
	) name24344 (
		_w30006_,
		_w30008_,
		_w30019_,
		_w30171_
	);
	LUT4 #(
		.INIT('hfbbf)
	) name24345 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30172_
	);
	LUT4 #(
		.INIT('h00df)
	) name24346 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30010_,
		_w30173_
	);
	LUT4 #(
		.INIT('h1000)
	) name24347 (
		_w30029_,
		_w30171_,
		_w30173_,
		_w30172_,
		_w30174_
	);
	LUT4 #(
		.INIT('h0100)
	) name24348 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30175_
	);
	LUT3 #(
		.INIT('h02)
	) name24349 (
		_w30010_,
		_w30024_,
		_w30175_,
		_w30176_
	);
	LUT4 #(
		.INIT('hddd0)
	) name24350 (
		_w30019_,
		_w30170_,
		_w30174_,
		_w30176_,
		_w30177_
	);
	LUT3 #(
		.INIT('h65)
	) name24351 (
		\u0_L5_reg[15]/P0001 ,
		_w30165_,
		_w30177_,
		_w30178_
	);
	LUT4 #(
		.INIT('h3ec4)
	) name24352 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30179_
	);
	LUT4 #(
		.INIT('hcfbb)
	) name24353 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30180_
	);
	LUT4 #(
		.INIT('h4840)
	) name24354 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30181_
	);
	LUT4 #(
		.INIT('h00d8)
	) name24355 (
		_w30133_,
		_w30179_,
		_w30180_,
		_w30181_,
		_w30182_
	);
	LUT2 #(
		.INIT('h2)
	) name24356 (
		_w30131_,
		_w30182_,
		_w30183_
	);
	LUT4 #(
		.INIT('hf7ed)
	) name24357 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30184_
	);
	LUT2 #(
		.INIT('h2)
	) name24358 (
		_w30133_,
		_w30184_,
		_w30185_
	);
	LUT3 #(
		.INIT('h15)
	) name24359 (
		_w30133_,
		_w30135_,
		_w30136_,
		_w30186_
	);
	LUT2 #(
		.INIT('h4)
	) name24360 (
		_w30152_,
		_w30186_,
		_w30187_
	);
	LUT4 #(
		.INIT('h0020)
	) name24361 (
		_w30133_,
		_w30132_,
		_w30135_,
		_w30134_,
		_w30188_
	);
	LUT4 #(
		.INIT('h0080)
	) name24362 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30189_
	);
	LUT2 #(
		.INIT('h1)
	) name24363 (
		_w30133_,
		_w30132_,
		_w30190_
	);
	LUT4 #(
		.INIT('h0001)
	) name24364 (
		_w30133_,
		_w30132_,
		_w30135_,
		_w30136_,
		_w30191_
	);
	LUT3 #(
		.INIT('h01)
	) name24365 (
		_w30189_,
		_w30191_,
		_w30188_,
		_w30192_
	);
	LUT4 #(
		.INIT('h0400)
	) name24366 (
		_w30133_,
		_w30132_,
		_w30135_,
		_w30136_,
		_w30193_
	);
	LUT2 #(
		.INIT('h1)
	) name24367 (
		_w30148_,
		_w30193_,
		_w30194_
	);
	LUT4 #(
		.INIT('hba00)
	) name24368 (
		_w30131_,
		_w30187_,
		_w30192_,
		_w30194_,
		_w30195_
	);
	LUT4 #(
		.INIT('h5655)
	) name24369 (
		\u0_L5_reg[25]/NET0131 ,
		_w30183_,
		_w30185_,
		_w30195_,
		_w30196_
	);
	LUT4 #(
		.INIT('h080a)
	) name24370 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30197_
	);
	LUT3 #(
		.INIT('h01)
	) name24371 (
		_w30010_,
		_w30169_,
		_w30197_,
		_w30198_
	);
	LUT4 #(
		.INIT('h8381)
	) name24372 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30199_
	);
	LUT4 #(
		.INIT('hbf00)
	) name24373 (
		_w30006_,
		_w30008_,
		_w30009_,
		_w30010_,
		_w30200_
	);
	LUT2 #(
		.INIT('h4)
	) name24374 (
		_w30199_,
		_w30200_,
		_w30201_
	);
	LUT4 #(
		.INIT('h0090)
	) name24375 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30202_
	);
	LUT3 #(
		.INIT('h02)
	) name24376 (
		_w30019_,
		_w30175_,
		_w30202_,
		_w30203_
	);
	LUT3 #(
		.INIT('he0)
	) name24377 (
		_w30198_,
		_w30201_,
		_w30203_,
		_w30204_
	);
	LUT4 #(
		.INIT('hde56)
	) name24378 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30205_
	);
	LUT2 #(
		.INIT('h2)
	) name24379 (
		_w30010_,
		_w30205_,
		_w30206_
	);
	LUT4 #(
		.INIT('h00bf)
	) name24380 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30019_,
		_w30207_
	);
	LUT2 #(
		.INIT('h4)
	) name24381 (
		_w30014_,
		_w30207_,
		_w30208_
	);
	LUT2 #(
		.INIT('h8)
	) name24382 (
		_w30006_,
		_w30009_,
		_w30209_
	);
	LUT3 #(
		.INIT('hdc)
	) name24383 (
		_w30008_,
		_w30007_,
		_w30010_,
		_w30210_
	);
	LUT2 #(
		.INIT('h2)
	) name24384 (
		_w30209_,
		_w30210_,
		_w30211_
	);
	LUT2 #(
		.INIT('h1)
	) name24385 (
		_w30006_,
		_w30010_,
		_w30212_
	);
	LUT3 #(
		.INIT('h35)
	) name24386 (
		_w30008_,
		_w30007_,
		_w30009_,
		_w30213_
	);
	LUT3 #(
		.INIT('h51)
	) name24387 (
		_w30029_,
		_w30212_,
		_w30213_,
		_w30214_
	);
	LUT4 #(
		.INIT('h1000)
	) name24388 (
		_w30206_,
		_w30211_,
		_w30208_,
		_w30214_,
		_w30215_
	);
	LUT3 #(
		.INIT('ha9)
	) name24389 (
		\u0_L5_reg[21]/NET0131 ,
		_w30204_,
		_w30215_,
		_w30216_
	);
	LUT3 #(
		.INIT('h01)
	) name24390 (
		_w29971_,
		_w29973_,
		_w29974_,
		_w30217_
	);
	LUT3 #(
		.INIT('h02)
	) name24391 (
		_w29976_,
		_w30001_,
		_w30217_,
		_w30218_
	);
	LUT3 #(
		.INIT('h40)
	) name24392 (
		_w29972_,
		_w29973_,
		_w29974_,
		_w30219_
	);
	LUT4 #(
		.INIT('h5545)
	) name24393 (
		_w29976_,
		_w29971_,
		_w29973_,
		_w29974_,
		_w30220_
	);
	LUT2 #(
		.INIT('h4)
	) name24394 (
		_w30219_,
		_w30220_,
		_w30221_
	);
	LUT4 #(
		.INIT('h7bbf)
	) name24395 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30222_
	);
	LUT4 #(
		.INIT('h0155)
	) name24396 (
		_w29984_,
		_w30218_,
		_w30221_,
		_w30222_,
		_w30223_
	);
	LUT4 #(
		.INIT('hb3fb)
	) name24397 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30224_
	);
	LUT4 #(
		.INIT('h0080)
	) name24398 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30225_
	);
	LUT4 #(
		.INIT('hfd7d)
	) name24399 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30226_
	);
	LUT4 #(
		.INIT('h04cc)
	) name24400 (
		_w29976_,
		_w29984_,
		_w30224_,
		_w30226_,
		_w30227_
	);
	LUT4 #(
		.INIT('h7df7)
	) name24401 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30228_
	);
	LUT2 #(
		.INIT('h2)
	) name24402 (
		_w29976_,
		_w30228_,
		_w30229_
	);
	LUT2 #(
		.INIT('h4)
	) name24403 (
		_w29976_,
		_w30225_,
		_w30230_
	);
	LUT4 #(
		.INIT('hccef)
	) name24404 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w30231_
	);
	LUT2 #(
		.INIT('h8)
	) name24405 (
		_w29976_,
		_w29984_,
		_w30232_
	);
	LUT4 #(
		.INIT('h7077)
	) name24406 (
		_w29971_,
		_w29982_,
		_w30231_,
		_w30232_,
		_w30233_
	);
	LUT4 #(
		.INIT('h0100)
	) name24407 (
		_w30229_,
		_w30230_,
		_w30227_,
		_w30233_,
		_w30234_
	);
	LUT3 #(
		.INIT('h65)
	) name24408 (
		\u0_L5_reg[1]/NET0131 ,
		_w30223_,
		_w30234_,
		_w30235_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name24409 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30236_
	);
	LUT2 #(
		.INIT('h2)
	) name24410 (
		_w30072_,
		_w30236_,
		_w30237_
	);
	LUT4 #(
		.INIT('hbfae)
	) name24411 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30238_
	);
	LUT2 #(
		.INIT('h1)
	) name24412 (
		_w30072_,
		_w30238_,
		_w30239_
	);
	LUT2 #(
		.INIT('h8)
	) name24413 (
		_w30072_,
		_w30074_,
		_w30240_
	);
	LUT4 #(
		.INIT('h7737)
	) name24414 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30073_,
		_w30241_
	);
	LUT4 #(
		.INIT('h0400)
	) name24415 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30242_
	);
	LUT3 #(
		.INIT('h0e)
	) name24416 (
		_w30076_,
		_w30241_,
		_w30242_,
		_w30243_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name24417 (
		_w30071_,
		_w30239_,
		_w30237_,
		_w30243_,
		_w30244_
	);
	LUT4 #(
		.INIT('hdaff)
	) name24418 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30245_
	);
	LUT2 #(
		.INIT('h1)
	) name24419 (
		_w30072_,
		_w30245_,
		_w30246_
	);
	LUT3 #(
		.INIT('h02)
	) name24420 (
		_w30074_,
		_w30075_,
		_w30076_,
		_w30247_
	);
	LUT4 #(
		.INIT('h1145)
	) name24421 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30073_,
		_w30248_
	);
	LUT4 #(
		.INIT('h7077)
	) name24422 (
		_w30072_,
		_w30238_,
		_w30247_,
		_w30248_,
		_w30249_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name24423 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30250_
	);
	LUT4 #(
		.INIT('h2322)
	) name24424 (
		_w30071_,
		_w30246_,
		_w30249_,
		_w30250_,
		_w30251_
	);
	LUT3 #(
		.INIT('h65)
	) name24425 (
		\u0_L5_reg[28]/NET0131 ,
		_w30244_,
		_w30251_,
		_w30252_
	);
	LUT4 #(
		.INIT('hb97d)
	) name24426 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30253_
	);
	LUT2 #(
		.INIT('h2)
	) name24427 (
		_w29944_,
		_w30253_,
		_w30254_
	);
	LUT4 #(
		.INIT('heedf)
	) name24428 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30255_
	);
	LUT4 #(
		.INIT('h0302)
	) name24429 (
		_w29944_,
		_w29947_,
		_w29949_,
		_w30255_,
		_w30256_
	);
	LUT3 #(
		.INIT('h45)
	) name24430 (
		_w29938_,
		_w30254_,
		_w30256_,
		_w30257_
	);
	LUT4 #(
		.INIT('h7ebe)
	) name24431 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30258_
	);
	LUT2 #(
		.INIT('h1)
	) name24432 (
		_w29944_,
		_w30258_,
		_w30259_
	);
	LUT4 #(
		.INIT('hf8fc)
	) name24433 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30260_
	);
	LUT2 #(
		.INIT('h1)
	) name24434 (
		_w29944_,
		_w30260_,
		_w30261_
	);
	LUT4 #(
		.INIT('h0800)
	) name24435 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29944_,
		_w30262_
	);
	LUT3 #(
		.INIT('h80)
	) name24436 (
		_w29940_,
		_w29939_,
		_w29942_,
		_w30263_
	);
	LUT3 #(
		.INIT('h01)
	) name24437 (
		_w29965_,
		_w30262_,
		_w30263_,
		_w30264_
	);
	LUT3 #(
		.INIT('h9e)
	) name24438 (
		_w29940_,
		_w29941_,
		_w29942_,
		_w30265_
	);
	LUT2 #(
		.INIT('h2)
	) name24439 (
		_w29953_,
		_w30265_,
		_w30266_
	);
	LUT4 #(
		.INIT('h0075)
	) name24440 (
		_w29938_,
		_w30261_,
		_w30264_,
		_w30266_,
		_w30267_
	);
	LUT4 #(
		.INIT('h5655)
	) name24441 (
		\u0_L5_reg[4]/NET0131 ,
		_w30259_,
		_w30257_,
		_w30267_,
		_w30268_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name24442 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30269_
	);
	LUT4 #(
		.INIT('hcb6d)
	) name24443 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30270_
	);
	LUT2 #(
		.INIT('h1)
	) name24444 (
		_w30072_,
		_w30270_,
		_w30271_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name24445 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30272_
	);
	LUT4 #(
		.INIT('haa82)
	) name24446 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30073_,
		_w30273_
	);
	LUT2 #(
		.INIT('h4)
	) name24447 (
		_w30272_,
		_w30273_,
		_w30274_
	);
	LUT3 #(
		.INIT('hb0)
	) name24448 (
		_w30075_,
		_w30073_,
		_w30076_,
		_w30275_
	);
	LUT2 #(
		.INIT('h8)
	) name24449 (
		_w30240_,
		_w30275_,
		_w30276_
	);
	LUT3 #(
		.INIT('h32)
	) name24450 (
		_w30072_,
		_w30074_,
		_w30073_,
		_w30277_
	);
	LUT3 #(
		.INIT('h15)
	) name24451 (
		_w30071_,
		_w30082_,
		_w30277_,
		_w30278_
	);
	LUT4 #(
		.INIT('h0100)
	) name24452 (
		_w30276_,
		_w30271_,
		_w30274_,
		_w30278_,
		_w30279_
	);
	LUT3 #(
		.INIT('h01)
	) name24453 (
		_w30075_,
		_w30073_,
		_w30076_,
		_w30280_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name24454 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30076_,
		_w30281_
	);
	LUT4 #(
		.INIT('h5515)
	) name24455 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30073_,
		_w30282_
	);
	LUT4 #(
		.INIT('h8acf)
	) name24456 (
		_w30095_,
		_w30280_,
		_w30281_,
		_w30282_,
		_w30283_
	);
	LUT4 #(
		.INIT('h0010)
	) name24457 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30284_
	);
	LUT4 #(
		.INIT('h0002)
	) name24458 (
		_w30071_,
		_w30083_,
		_w30084_,
		_w30284_,
		_w30285_
	);
	LUT3 #(
		.INIT('h20)
	) name24459 (
		_w30269_,
		_w30283_,
		_w30285_,
		_w30286_
	);
	LUT3 #(
		.INIT('h56)
	) name24460 (
		\u0_L5_reg[13]/NET0131 ,
		_w30279_,
		_w30286_,
		_w30287_
	);
	LUT4 #(
		.INIT('hba76)
	) name24461 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30288_
	);
	LUT2 #(
		.INIT('h1)
	) name24462 (
		_w30010_,
		_w30288_,
		_w30289_
	);
	LUT3 #(
		.INIT('hd0)
	) name24463 (
		_w30006_,
		_w30009_,
		_w30010_,
		_w30290_
	);
	LUT4 #(
		.INIT('hbcdf)
	) name24464 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30291_
	);
	LUT3 #(
		.INIT('hb0)
	) name24465 (
		_w30162_,
		_w30290_,
		_w30291_,
		_w30292_
	);
	LUT3 #(
		.INIT('h8a)
	) name24466 (
		_w30019_,
		_w30289_,
		_w30292_,
		_w30293_
	);
	LUT4 #(
		.INIT('hfd00)
	) name24467 (
		_w30008_,
		_w30007_,
		_w30009_,
		_w30010_,
		_w30294_
	);
	LUT4 #(
		.INIT('h0cbf)
	) name24468 (
		_w30006_,
		_w30008_,
		_w30007_,
		_w30009_,
		_w30295_
	);
	LUT2 #(
		.INIT('h8)
	) name24469 (
		_w30294_,
		_w30295_,
		_w30296_
	);
	LUT4 #(
		.INIT('h0080)
	) name24470 (
		_w30006_,
		_w30007_,
		_w30009_,
		_w30010_,
		_w30297_
	);
	LUT4 #(
		.INIT('h0004)
	) name24471 (
		_w30006_,
		_w30008_,
		_w30009_,
		_w30010_,
		_w30298_
	);
	LUT3 #(
		.INIT('h01)
	) name24472 (
		_w30030_,
		_w30298_,
		_w30297_,
		_w30299_
	);
	LUT3 #(
		.INIT('h45)
	) name24473 (
		_w30019_,
		_w30296_,
		_w30299_,
		_w30300_
	);
	LUT2 #(
		.INIT('h4)
	) name24474 (
		_w30010_,
		_w30028_,
		_w30301_
	);
	LUT4 #(
		.INIT('h0400)
	) name24475 (
		_w30008_,
		_w30007_,
		_w30009_,
		_w30010_,
		_w30302_
	);
	LUT3 #(
		.INIT('h07)
	) name24476 (
		_w30011_,
		_w30033_,
		_w30302_,
		_w30303_
	);
	LUT2 #(
		.INIT('h4)
	) name24477 (
		_w30301_,
		_w30303_,
		_w30304_
	);
	LUT4 #(
		.INIT('h5655)
	) name24478 (
		\u0_L5_reg[27]/NET0131 ,
		_w30293_,
		_w30300_,
		_w30304_,
		_w30305_
	);
	LUT3 #(
		.INIT('hb9)
	) name24479 (
		_w29909_,
		_w29911_,
		_w29908_,
		_w30306_
	);
	LUT4 #(
		.INIT('hfba5)
	) name24480 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30307_
	);
	LUT2 #(
		.INIT('h1)
	) name24481 (
		_w29914_,
		_w30307_,
		_w30308_
	);
	LUT3 #(
		.INIT('h8a)
	) name24482 (
		_w29914_,
		_w29910_,
		_w29908_,
		_w30309_
	);
	LUT2 #(
		.INIT('h8)
	) name24483 (
		_w29925_,
		_w30309_,
		_w30310_
	);
	LUT3 #(
		.INIT('h07)
	) name24484 (
		_w29913_,
		_w29933_,
		_w30044_,
		_w30311_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name24485 (
		_w29907_,
		_w30308_,
		_w30310_,
		_w30311_,
		_w30312_
	);
	LUT4 #(
		.INIT('h0080)
	) name24486 (
		_w29914_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30313_
	);
	LUT3 #(
		.INIT('h7e)
	) name24487 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w30314_
	);
	LUT2 #(
		.INIT('h4)
	) name24488 (
		_w30313_,
		_w30314_,
		_w30315_
	);
	LUT4 #(
		.INIT('h0008)
	) name24489 (
		_w29909_,
		_w29914_,
		_w29911_,
		_w29908_,
		_w30316_
	);
	LUT3 #(
		.INIT('h15)
	) name24490 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w30317_
	);
	LUT2 #(
		.INIT('h4)
	) name24491 (
		_w29914_,
		_w29908_,
		_w30318_
	);
	LUT3 #(
		.INIT('h45)
	) name24492 (
		_w30316_,
		_w30317_,
		_w30318_,
		_w30319_
	);
	LUT3 #(
		.INIT('h15)
	) name24493 (
		_w29907_,
		_w30315_,
		_w30319_,
		_w30320_
	);
	LUT4 #(
		.INIT('hfdef)
	) name24494 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30321_
	);
	LUT3 #(
		.INIT('had)
	) name24495 (
		_w29909_,
		_w29911_,
		_w29908_,
		_w30322_
	);
	LUT4 #(
		.INIT('h3120)
	) name24496 (
		_w29914_,
		_w29929_,
		_w30322_,
		_w30321_,
		_w30323_
	);
	LUT2 #(
		.INIT('h1)
	) name24497 (
		_w29924_,
		_w30323_,
		_w30324_
	);
	LUT4 #(
		.INIT('haaa9)
	) name24498 (
		\u0_L5_reg[23]/NET0131 ,
		_w30320_,
		_w30324_,
		_w30312_,
		_w30325_
	);
	LUT4 #(
		.INIT('h0800)
	) name24499 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30326_
	);
	LUT4 #(
		.INIT('h0012)
	) name24500 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30327_
	);
	LUT4 #(
		.INIT('h0080)
	) name24501 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30328_
	);
	LUT4 #(
		.INIT('h00ef)
	) name24502 (
		_w29879_,
		_w29881_,
		_w29882_,
		_w29878_,
		_w30329_
	);
	LUT3 #(
		.INIT('h10)
	) name24503 (
		_w30328_,
		_w30327_,
		_w30329_,
		_w30330_
	);
	LUT4 #(
		.INIT('h3808)
	) name24504 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30331_
	);
	LUT4 #(
		.INIT('hfe00)
	) name24505 (
		_w29879_,
		_w29881_,
		_w29882_,
		_w29878_,
		_w30332_
	);
	LUT2 #(
		.INIT('h4)
	) name24506 (
		_w30331_,
		_w30332_,
		_w30333_
	);
	LUT4 #(
		.INIT('h888a)
	) name24507 (
		_w29877_,
		_w30326_,
		_w30330_,
		_w30333_,
		_w30334_
	);
	LUT4 #(
		.INIT('h0ff2)
	) name24508 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30335_
	);
	LUT2 #(
		.INIT('h1)
	) name24509 (
		_w29878_,
		_w30335_,
		_w30336_
	);
	LUT3 #(
		.INIT('h58)
	) name24510 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w30337_
	);
	LUT4 #(
		.INIT('h3111)
	) name24511 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30338_
	);
	LUT3 #(
		.INIT('h13)
	) name24512 (
		_w29879_,
		_w29882_,
		_w29878_,
		_w30339_
	);
	LUT3 #(
		.INIT('h01)
	) name24513 (
		_w30338_,
		_w30337_,
		_w30339_,
		_w30340_
	);
	LUT2 #(
		.INIT('h2)
	) name24514 (
		_w29877_,
		_w29878_,
		_w30341_
	);
	LUT4 #(
		.INIT('h00d0)
	) name24515 (
		_w29879_,
		_w29881_,
		_w29882_,
		_w29878_,
		_w30342_
	);
	LUT4 #(
		.INIT('h31f5)
	) name24516 (
		_w29898_,
		_w29890_,
		_w30341_,
		_w30342_,
		_w30343_
	);
	LUT4 #(
		.INIT('hab00)
	) name24517 (
		_w29877_,
		_w30336_,
		_w30340_,
		_w30343_,
		_w30344_
	);
	LUT3 #(
		.INIT('h65)
	) name24518 (
		\u0_L5_reg[32]/NET0131 ,
		_w30334_,
		_w30344_,
		_w30345_
	);
	LUT4 #(
		.INIT('h125a)
	) name24519 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30346_
	);
	LUT4 #(
		.INIT('h8404)
	) name24520 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30347_
	);
	LUT2 #(
		.INIT('h4)
	) name24521 (
		_w29877_,
		_w29878_,
		_w30348_
	);
	LUT3 #(
		.INIT('h04)
	) name24522 (
		_w30347_,
		_w30348_,
		_w30346_,
		_w30349_
	);
	LUT4 #(
		.INIT('h69a0)
	) name24523 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30350_
	);
	LUT2 #(
		.INIT('h9)
	) name24524 (
		_w29877_,
		_w29878_,
		_w30351_
	);
	LUT2 #(
		.INIT('h4)
	) name24525 (
		_w30350_,
		_w30351_,
		_w30352_
	);
	LUT3 #(
		.INIT('h60)
	) name24526 (
		_w29879_,
		_w29881_,
		_w29882_,
		_w30353_
	);
	LUT3 #(
		.INIT('h41)
	) name24527 (
		_w29879_,
		_w29880_,
		_w29882_,
		_w30354_
	);
	LUT4 #(
		.INIT('h0888)
	) name24528 (
		_w29879_,
		_w29880_,
		_w29881_,
		_w29882_,
		_w30355_
	);
	LUT4 #(
		.INIT('h0002)
	) name24529 (
		_w30341_,
		_w30355_,
		_w30354_,
		_w30353_,
		_w30356_
	);
	LUT4 #(
		.INIT('h00ab)
	) name24530 (
		_w29883_,
		_w30349_,
		_w30352_,
		_w30356_,
		_w30357_
	);
	LUT2 #(
		.INIT('h6)
	) name24531 (
		\u0_L5_reg[7]/NET0131 ,
		_w30357_,
		_w30358_
	);
	LUT4 #(
		.INIT('hcffe)
	) name24532 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30359_
	);
	LUT3 #(
		.INIT('h10)
	) name24533 (
		_w30133_,
		_w30132_,
		_w30136_,
		_w30360_
	);
	LUT4 #(
		.INIT('h0031)
	) name24534 (
		_w30133_,
		_w30158_,
		_w30359_,
		_w30360_,
		_w30361_
	);
	LUT2 #(
		.INIT('h2)
	) name24535 (
		_w30131_,
		_w30361_,
		_w30362_
	);
	LUT3 #(
		.INIT('h02)
	) name24536 (
		_w30133_,
		_w30149_,
		_w30143_,
		_w30363_
	);
	LUT4 #(
		.INIT('h00d0)
	) name24537 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30364_
	);
	LUT4 #(
		.INIT('h4555)
	) name24538 (
		_w30133_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30365_
	);
	LUT2 #(
		.INIT('h4)
	) name24539 (
		_w30364_,
		_w30365_,
		_w30366_
	);
	LUT4 #(
		.INIT('hf7b9)
	) name24540 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30367_
	);
	LUT4 #(
		.INIT('h0155)
	) name24541 (
		_w30131_,
		_w30363_,
		_w30366_,
		_w30367_,
		_w30368_
	);
	LUT4 #(
		.INIT('hf797)
	) name24542 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30369_
	);
	LUT4 #(
		.INIT('hcf45)
	) name24543 (
		_w30133_,
		_w30134_,
		_w30193_,
		_w30369_,
		_w30370_
	);
	LUT4 #(
		.INIT('h5655)
	) name24544 (
		\u0_L5_reg[8]/NET0131 ,
		_w30368_,
		_w30362_,
		_w30370_,
		_w30371_
	);
	LUT4 #(
		.INIT('hf3dd)
	) name24545 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30372_
	);
	LUT2 #(
		.INIT('h2)
	) name24546 (
		_w29944_,
		_w30372_,
		_w30373_
	);
	LUT3 #(
		.INIT('h02)
	) name24547 (
		_w29941_,
		_w29942_,
		_w29944_,
		_w30374_
	);
	LUT4 #(
		.INIT('hef00)
	) name24548 (
		_w29940_,
		_w29939_,
		_w29942_,
		_w29938_,
		_w30375_
	);
	LUT4 #(
		.INIT('hdfed)
	) name24549 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30376_
	);
	LUT3 #(
		.INIT('h40)
	) name24550 (
		_w30374_,
		_w30375_,
		_w30376_,
		_w30377_
	);
	LUT4 #(
		.INIT('h2e33)
	) name24551 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30378_
	);
	LUT2 #(
		.INIT('h2)
	) name24552 (
		_w29944_,
		_w30378_,
		_w30379_
	);
	LUT4 #(
		.INIT('h0021)
	) name24553 (
		_w29940_,
		_w29941_,
		_w29942_,
		_w29944_,
		_w30380_
	);
	LUT4 #(
		.INIT('h8000)
	) name24554 (
		_w29940_,
		_w29941_,
		_w29939_,
		_w29942_,
		_w30381_
	);
	LUT3 #(
		.INIT('h01)
	) name24555 (
		_w29938_,
		_w30381_,
		_w30380_,
		_w30382_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name24556 (
		_w30373_,
		_w30377_,
		_w30379_,
		_w30382_,
		_w30383_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name24557 (
		_w29939_,
		_w29942_,
		_w29963_,
		_w29949_,
		_w30384_
	);
	LUT3 #(
		.INIT('h65)
	) name24558 (
		\u0_L5_reg[19]/P0001 ,
		_w30383_,
		_w30384_,
		_w30385_
	);
	LUT4 #(
		.INIT('hc693)
	) name24559 (
		decrypt_pad,
		\u0_R5_reg[11]/P0001 ,
		\u0_uk_K_r5_reg[32]/NET0131 ,
		\u0_uk_K_r5_reg[54]/NET0131 ,
		_w30386_
	);
	LUT4 #(
		.INIT('hc963)
	) name24560 (
		decrypt_pad,
		\u0_R5_reg[9]/NET0131 ,
		\u0_uk_K_r5_reg[20]/NET0131 ,
		\u0_uk_K_r5_reg[55]/NET0131 ,
		_w30387_
	);
	LUT4 #(
		.INIT('hc963)
	) name24561 (
		decrypt_pad,
		\u0_R5_reg[13]/NET0131 ,
		\u0_uk_K_r5_reg[25]/NET0131 ,
		\u0_uk_K_r5_reg[3]/NET0131 ,
		_w30388_
	);
	LUT4 #(
		.INIT('hc963)
	) name24562 (
		decrypt_pad,
		\u0_R5_reg[10]/NET0131 ,
		\u0_uk_K_r5_reg[53]/NET0131 ,
		\u0_uk_K_r5_reg[6]/NET0131 ,
		_w30389_
	);
	LUT4 #(
		.INIT('hc693)
	) name24563 (
		decrypt_pad,
		\u0_R5_reg[8]/NET0131 ,
		\u0_uk_K_r5_reg[26]/NET0131 ,
		\u0_uk_K_r5_reg[48]/NET0131 ,
		_w30390_
	);
	LUT4 #(
		.INIT('h9909)
	) name24564 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30391_
	);
	LUT4 #(
		.INIT('hc963)
	) name24565 (
		decrypt_pad,
		\u0_R5_reg[12]/NET0131 ,
		\u0_uk_K_r5_reg[12]/NET0131 ,
		\u0_uk_K_r5_reg[47]/NET0131 ,
		_w30392_
	);
	LUT3 #(
		.INIT('ha8)
	) name24566 (
		_w30392_,
		_w30388_,
		_w30390_,
		_w30393_
	);
	LUT4 #(
		.INIT('h0001)
	) name24567 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30394_
	);
	LUT4 #(
		.INIT('hbfbe)
	) name24568 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30395_
	);
	LUT4 #(
		.INIT('h40cc)
	) name24569 (
		_w30391_,
		_w30386_,
		_w30393_,
		_w30395_,
		_w30396_
	);
	LUT3 #(
		.INIT('h0e)
	) name24570 (
		_w30387_,
		_w30390_,
		_w30386_,
		_w30397_
	);
	LUT4 #(
		.INIT('h0020)
	) name24571 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30398_
	);
	LUT4 #(
		.INIT('haa80)
	) name24572 (
		_w30392_,
		_w30391_,
		_w30397_,
		_w30398_,
		_w30399_
	);
	LUT2 #(
		.INIT('h8)
	) name24573 (
		_w30388_,
		_w30386_,
		_w30400_
	);
	LUT3 #(
		.INIT('h80)
	) name24574 (
		_w30387_,
		_w30388_,
		_w30386_,
		_w30401_
	);
	LUT2 #(
		.INIT('h1)
	) name24575 (
		_w30387_,
		_w30389_,
		_w30402_
	);
	LUT2 #(
		.INIT('h6)
	) name24576 (
		_w30387_,
		_w30389_,
		_w30403_
	);
	LUT2 #(
		.INIT('h9)
	) name24577 (
		_w30388_,
		_w30390_,
		_w30404_
	);
	LUT4 #(
		.INIT('h1248)
	) name24578 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30405_
	);
	LUT2 #(
		.INIT('h4)
	) name24579 (
		_w30401_,
		_w30405_,
		_w30406_
	);
	LUT3 #(
		.INIT('h46)
	) name24580 (
		_w30388_,
		_w30390_,
		_w30386_,
		_w30407_
	);
	LUT3 #(
		.INIT('h54)
	) name24581 (
		_w30392_,
		_w30403_,
		_w30407_,
		_w30408_
	);
	LUT4 #(
		.INIT('h0045)
	) name24582 (
		_w30399_,
		_w30406_,
		_w30408_,
		_w30396_,
		_w30409_
	);
	LUT2 #(
		.INIT('h9)
	) name24583 (
		\u0_L5_reg[6]/NET0131 ,
		_w30409_,
		_w30410_
	);
	LUT3 #(
		.INIT('h29)
	) name24584 (
		_w30388_,
		_w30390_,
		_w30386_,
		_w30411_
	);
	LUT2 #(
		.INIT('h2)
	) name24585 (
		_w30402_,
		_w30411_,
		_w30412_
	);
	LUT3 #(
		.INIT('h0e)
	) name24586 (
		_w30387_,
		_w30389_,
		_w30386_,
		_w30413_
	);
	LUT3 #(
		.INIT('h2a)
	) name24587 (
		_w30392_,
		_w30404_,
		_w30413_,
		_w30414_
	);
	LUT3 #(
		.INIT('hf9)
	) name24588 (
		_w30388_,
		_w30389_,
		_w30390_,
		_w30415_
	);
	LUT3 #(
		.INIT('h40)
	) name24589 (
		_w30387_,
		_w30389_,
		_w30390_,
		_w30416_
	);
	LUT3 #(
		.INIT('h02)
	) name24590 (
		_w30387_,
		_w30388_,
		_w30390_,
		_w30417_
	);
	LUT4 #(
		.INIT('hafc1)
	) name24591 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30418_
	);
	LUT4 #(
		.INIT('h1000)
	) name24592 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30419_
	);
	LUT4 #(
		.INIT('h0501)
	) name24593 (
		_w30392_,
		_w30386_,
		_w30419_,
		_w30418_,
		_w30420_
	);
	LUT3 #(
		.INIT('h0b)
	) name24594 (
		_w30412_,
		_w30414_,
		_w30420_,
		_w30421_
	);
	LUT4 #(
		.INIT('h0108)
	) name24595 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30422_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name24596 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30423_
	);
	LUT4 #(
		.INIT('h00c4)
	) name24597 (
		_w30392_,
		_w30386_,
		_w30423_,
		_w30422_,
		_w30424_
	);
	LUT4 #(
		.INIT('hd93e)
	) name24598 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30425_
	);
	LUT4 #(
		.INIT('h8000)
	) name24599 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30426_
	);
	LUT4 #(
		.INIT('h0032)
	) name24600 (
		_w30392_,
		_w30386_,
		_w30425_,
		_w30426_,
		_w30427_
	);
	LUT2 #(
		.INIT('h1)
	) name24601 (
		_w30424_,
		_w30427_,
		_w30428_
	);
	LUT3 #(
		.INIT('h56)
	) name24602 (
		\u0_L5_reg[24]/NET0131 ,
		_w30421_,
		_w30428_,
		_w30429_
	);
	LUT4 #(
		.INIT('h696b)
	) name24603 (
		_w30387_,
		_w30388_,
		_w30390_,
		_w30386_,
		_w30430_
	);
	LUT4 #(
		.INIT('h0080)
	) name24604 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30431_
	);
	LUT3 #(
		.INIT('h07)
	) name24605 (
		_w30389_,
		_w30390_,
		_w30386_,
		_w30432_
	);
	LUT4 #(
		.INIT('h0014)
	) name24606 (
		_w30388_,
		_w30389_,
		_w30390_,
		_w30386_,
		_w30433_
	);
	LUT4 #(
		.INIT('h0032)
	) name24607 (
		_w30389_,
		_w30431_,
		_w30430_,
		_w30433_,
		_w30434_
	);
	LUT2 #(
		.INIT('h2)
	) name24608 (
		_w30392_,
		_w30434_,
		_w30435_
	);
	LUT4 #(
		.INIT('h4430)
	) name24609 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30436_
	);
	LUT4 #(
		.INIT('h5015)
	) name24610 (
		_w30392_,
		_w30387_,
		_w30388_,
		_w30390_,
		_w30437_
	);
	LUT4 #(
		.INIT('h4544)
	) name24611 (
		_w30386_,
		_w30416_,
		_w30436_,
		_w30437_,
		_w30438_
	);
	LUT4 #(
		.INIT('h6800)
	) name24612 (
		_w30387_,
		_w30388_,
		_w30390_,
		_w30386_,
		_w30439_
	);
	LUT3 #(
		.INIT('h54)
	) name24613 (
		_w30392_,
		_w30394_,
		_w30439_,
		_w30440_
	);
	LUT3 #(
		.INIT('hde)
	) name24614 (
		_w30387_,
		_w30388_,
		_w30390_,
		_w30441_
	);
	LUT2 #(
		.INIT('h8)
	) name24615 (
		_w30389_,
		_w30386_,
		_w30442_
	);
	LUT2 #(
		.INIT('h4)
	) name24616 (
		_w30441_,
		_w30442_,
		_w30443_
	);
	LUT3 #(
		.INIT('h01)
	) name24617 (
		_w30438_,
		_w30440_,
		_w30443_,
		_w30444_
	);
	LUT3 #(
		.INIT('h65)
	) name24618 (
		\u0_L5_reg[16]/NET0131 ,
		_w30435_,
		_w30444_,
		_w30445_
	);
	LUT3 #(
		.INIT('h02)
	) name24619 (
		_w30133_,
		_w30149_,
		_w30157_,
		_w30446_
	);
	LUT4 #(
		.INIT('h0401)
	) name24620 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30447_
	);
	LUT3 #(
		.INIT('h0e)
	) name24621 (
		_w30190_,
		_w30365_,
		_w30447_,
		_w30448_
	);
	LUT2 #(
		.INIT('h1)
	) name24622 (
		_w30446_,
		_w30448_,
		_w30449_
	);
	LUT4 #(
		.INIT('hf3af)
	) name24623 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30450_
	);
	LUT2 #(
		.INIT('h2)
	) name24624 (
		_w30133_,
		_w30450_,
		_w30451_
	);
	LUT4 #(
		.INIT('h4f50)
	) name24625 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30452_
	);
	LUT4 #(
		.INIT('h2022)
	) name24626 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30453_
	);
	LUT4 #(
		.INIT('h0054)
	) name24627 (
		_w30131_,
		_w30133_,
		_w30452_,
		_w30453_,
		_w30454_
	);
	LUT4 #(
		.INIT('ha0f3)
	) name24628 (
		_w30132_,
		_w30135_,
		_w30134_,
		_w30136_,
		_w30455_
	);
	LUT3 #(
		.INIT('h8a)
	) name24629 (
		_w30133_,
		_w30134_,
		_w30136_,
		_w30456_
	);
	LUT2 #(
		.INIT('h4)
	) name24630 (
		_w30455_,
		_w30456_,
		_w30457_
	);
	LUT4 #(
		.INIT('h0002)
	) name24631 (
		_w30131_,
		_w30148_,
		_w30145_,
		_w30137_,
		_w30458_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name24632 (
		_w30451_,
		_w30454_,
		_w30457_,
		_w30458_,
		_w30459_
	);
	LUT3 #(
		.INIT('h56)
	) name24633 (
		\u0_L5_reg[3]/NET0131 ,
		_w30449_,
		_w30459_,
		_w30460_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name24634 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30461_
	);
	LUT4 #(
		.INIT('hdf00)
	) name24635 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30386_,
		_w30462_
	);
	LUT4 #(
		.INIT('hfbbe)
	) name24636 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30463_
	);
	LUT4 #(
		.INIT('h4700)
	) name24637 (
		_w30397_,
		_w30461_,
		_w30462_,
		_w30463_,
		_w30464_
	);
	LUT2 #(
		.INIT('h1)
	) name24638 (
		_w30392_,
		_w30464_,
		_w30465_
	);
	LUT2 #(
		.INIT('h8)
	) name24639 (
		_w30400_,
		_w30416_,
		_w30466_
	);
	LUT4 #(
		.INIT('h0020)
	) name24640 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30386_,
		_w30467_
	);
	LUT2 #(
		.INIT('h1)
	) name24641 (
		_w30392_,
		_w30467_,
		_w30468_
	);
	LUT4 #(
		.INIT('h20a0)
	) name24642 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30469_
	);
	LUT2 #(
		.INIT('h4)
	) name24643 (
		_w30417_,
		_w30432_,
		_w30470_
	);
	LUT4 #(
		.INIT('h0100)
	) name24644 (
		_w30387_,
		_w30388_,
		_w30389_,
		_w30390_,
		_w30471_
	);
	LUT3 #(
		.INIT('h08)
	) name24645 (
		_w30386_,
		_w30415_,
		_w30471_,
		_w30472_
	);
	LUT4 #(
		.INIT('h4445)
	) name24646 (
		_w30468_,
		_w30469_,
		_w30470_,
		_w30472_,
		_w30473_
	);
	LUT4 #(
		.INIT('haaa9)
	) name24647 (
		\u0_L5_reg[30]/NET0131 ,
		_w30466_,
		_w30473_,
		_w30465_,
		_w30474_
	);
	LUT3 #(
		.INIT('h19)
	) name24648 (
		_w29909_,
		_w29911_,
		_w29908_,
		_w30475_
	);
	LUT4 #(
		.INIT('h3212)
	) name24649 (
		_w29909_,
		_w29914_,
		_w29911_,
		_w29908_,
		_w30476_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name24650 (
		_w29909_,
		_w29914_,
		_w29910_,
		_w29911_,
		_w30477_
	);
	LUT4 #(
		.INIT('h9ffb)
	) name24651 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30478_
	);
	LUT4 #(
		.INIT('hec00)
	) name24652 (
		_w30306_,
		_w30476_,
		_w30477_,
		_w30478_,
		_w30479_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name24653 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30480_
	);
	LUT2 #(
		.INIT('h1)
	) name24654 (
		_w29914_,
		_w30480_,
		_w30481_
	);
	LUT4 #(
		.INIT('h8448)
	) name24655 (
		_w29909_,
		_w29910_,
		_w29911_,
		_w29908_,
		_w30482_
	);
	LUT4 #(
		.INIT('h0013)
	) name24656 (
		_w29915_,
		_w30047_,
		_w30475_,
		_w30482_,
		_w30483_
	);
	LUT4 #(
		.INIT('h3120)
	) name24657 (
		_w29907_,
		_w30481_,
		_w30483_,
		_w30479_,
		_w30484_
	);
	LUT2 #(
		.INIT('h9)
	) name24658 (
		\u0_L5_reg[9]/NET0131 ,
		_w30484_,
		_w30485_
	);
	LUT4 #(
		.INIT('h0a20)
	) name24659 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30073_,
		_w30486_
	);
	LUT4 #(
		.INIT('hfd75)
	) name24660 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30487_
	);
	LUT4 #(
		.INIT('h0032)
	) name24661 (
		_w30072_,
		_w30096_,
		_w30487_,
		_w30486_,
		_w30488_
	);
	LUT4 #(
		.INIT('h8000)
	) name24662 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30073_,
		_w30489_
	);
	LUT4 #(
		.INIT('hdffc)
	) name24663 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30490_
	);
	LUT4 #(
		.INIT('h1003)
	) name24664 (
		_w30072_,
		_w30074_,
		_w30073_,
		_w30076_,
		_w30491_
	);
	LUT4 #(
		.INIT('h0100)
	) name24665 (
		_w30081_,
		_w30489_,
		_w30491_,
		_w30490_,
		_w30492_
	);
	LUT4 #(
		.INIT('h1000)
	) name24666 (
		_w30072_,
		_w30074_,
		_w30075_,
		_w30073_,
		_w30493_
	);
	LUT4 #(
		.INIT('h77ef)
	) name24667 (
		_w30074_,
		_w30075_,
		_w30073_,
		_w30076_,
		_w30494_
	);
	LUT3 #(
		.INIT('h31)
	) name24668 (
		_w30072_,
		_w30493_,
		_w30494_,
		_w30495_
	);
	LUT4 #(
		.INIT('hd800)
	) name24669 (
		_w30071_,
		_w30488_,
		_w30492_,
		_w30495_,
		_w30496_
	);
	LUT2 #(
		.INIT('h9)
	) name24670 (
		\u0_L5_reg[18]/NET0131 ,
		_w30496_,
		_w30497_
	);
	LUT4 #(
		.INIT('hc963)
	) name24671 (
		decrypt_pad,
		\u0_R4_reg[4]/NET0131 ,
		\u0_uk_K_r4_reg[19]/NET0131 ,
		\u0_uk_K_r4_reg[25]/NET0131 ,
		_w30498_
	);
	LUT4 #(
		.INIT('hc693)
	) name24672 (
		decrypt_pad,
		\u0_R4_reg[2]/NET0131 ,
		\u0_uk_K_r4_reg[13]/NET0131 ,
		\u0_uk_K_r4_reg[32]/NET0131 ,
		_w30499_
	);
	LUT4 #(
		.INIT('hc963)
	) name24673 (
		decrypt_pad,
		\u0_R4_reg[3]/NET0131 ,
		\u0_uk_K_r4_reg[41]/NET0131 ,
		\u0_uk_K_r4_reg[47]/NET0131 ,
		_w30500_
	);
	LUT4 #(
		.INIT('hc963)
	) name24674 (
		decrypt_pad,
		\u0_R4_reg[1]/NET0131 ,
		\u0_uk_K_r4_reg[17]/NET0131 ,
		\u0_uk_K_r4_reg[55]/NET0131 ,
		_w30501_
	);
	LUT4 #(
		.INIT('hc693)
	) name24675 (
		decrypt_pad,
		\u0_R4_reg[32]/NET0131 ,
		\u0_uk_K_r4_reg[34]/NET0131 ,
		\u0_uk_K_r4_reg[53]/NET0131 ,
		_w30502_
	);
	LUT4 #(
		.INIT('hc963)
	) name24676 (
		decrypt_pad,
		\u0_R4_reg[5]/NET0131 ,
		\u0_uk_K_r4_reg[47]/NET0131 ,
		\u0_uk_K_r4_reg[53]/NET0131 ,
		_w30503_
	);
	LUT4 #(
		.INIT('h73cf)
	) name24677 (
		_w30500_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30504_
	);
	LUT2 #(
		.INIT('h1)
	) name24678 (
		_w30499_,
		_w30504_,
		_w30505_
	);
	LUT2 #(
		.INIT('h4)
	) name24679 (
		_w30502_,
		_w30503_,
		_w30506_
	);
	LUT3 #(
		.INIT('h48)
	) name24680 (
		_w30502_,
		_w30501_,
		_w30503_,
		_w30507_
	);
	LUT4 #(
		.INIT('hefe6)
	) name24681 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30508_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name24682 (
		_w30500_,
		_w30499_,
		_w30507_,
		_w30508_,
		_w30509_
	);
	LUT3 #(
		.INIT('h45)
	) name24683 (
		_w30498_,
		_w30505_,
		_w30509_,
		_w30510_
	);
	LUT4 #(
		.INIT('hafac)
	) name24684 (
		_w30500_,
		_w30499_,
		_w30501_,
		_w30503_,
		_w30511_
	);
	LUT2 #(
		.INIT('h2)
	) name24685 (
		_w30502_,
		_w30511_,
		_w30512_
	);
	LUT2 #(
		.INIT('h2)
	) name24686 (
		_w30500_,
		_w30499_,
		_w30513_
	);
	LUT3 #(
		.INIT('hd0)
	) name24687 (
		_w30500_,
		_w30499_,
		_w30501_,
		_w30514_
	);
	LUT2 #(
		.INIT('h2)
	) name24688 (
		_w30506_,
		_w30514_,
		_w30515_
	);
	LUT3 #(
		.INIT('ha8)
	) name24689 (
		_w30500_,
		_w30499_,
		_w30503_,
		_w30516_
	);
	LUT3 #(
		.INIT('h35)
	) name24690 (
		_w30502_,
		_w30501_,
		_w30503_,
		_w30517_
	);
	LUT3 #(
		.INIT('h02)
	) name24691 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30518_
	);
	LUT3 #(
		.INIT('h07)
	) name24692 (
		_w30516_,
		_w30517_,
		_w30518_,
		_w30519_
	);
	LUT4 #(
		.INIT('hef00)
	) name24693 (
		_w30512_,
		_w30515_,
		_w30519_,
		_w30498_,
		_w30520_
	);
	LUT4 #(
		.INIT('h0200)
	) name24694 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30521_
	);
	LUT4 #(
		.INIT('h7daf)
	) name24695 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30522_
	);
	LUT2 #(
		.INIT('h1)
	) name24696 (
		_w30500_,
		_w30522_,
		_w30523_
	);
	LUT4 #(
		.INIT('h0020)
	) name24697 (
		_w30500_,
		_w30499_,
		_w30502_,
		_w30501_,
		_w30524_
	);
	LUT2 #(
		.INIT('h2)
	) name24698 (
		_w30500_,
		_w30503_,
		_w30525_
	);
	LUT3 #(
		.INIT('h15)
	) name24699 (
		_w30524_,
		_w30518_,
		_w30525_,
		_w30526_
	);
	LUT2 #(
		.INIT('h4)
	) name24700 (
		_w30523_,
		_w30526_,
		_w30527_
	);
	LUT4 #(
		.INIT('h5655)
	) name24701 (
		\u0_L4_reg[31]/NET0131 ,
		_w30520_,
		_w30510_,
		_w30527_,
		_w30528_
	);
	LUT4 #(
		.INIT('hc963)
	) name24702 (
		decrypt_pad,
		\u0_R4_reg[24]/NET0131 ,
		\u0_uk_K_r4_reg[43]/NET0131 ,
		\u0_uk_K_r4_reg[51]/NET0131 ,
		_w30529_
	);
	LUT4 #(
		.INIT('hc963)
	) name24703 (
		decrypt_pad,
		\u0_R4_reg[22]/NET0131 ,
		\u0_uk_K_r4_reg[28]/NET0131 ,
		\u0_uk_K_r4_reg[36]/NET0131 ,
		_w30530_
	);
	LUT4 #(
		.INIT('hc693)
	) name24704 (
		decrypt_pad,
		\u0_R4_reg[21]/NET0131 ,
		\u0_uk_K_r4_reg[14]/NET0131 ,
		\u0_uk_K_r4_reg[37]/NET0131 ,
		_w30531_
	);
	LUT4 #(
		.INIT('hc963)
	) name24705 (
		decrypt_pad,
		\u0_R4_reg[20]/NET0131 ,
		\u0_uk_K_r4_reg[22]/NET0131 ,
		\u0_uk_K_r4_reg[30]/NET0131 ,
		_w30532_
	);
	LUT4 #(
		.INIT('hc693)
	) name24706 (
		decrypt_pad,
		\u0_R4_reg[25]/NET0131 ,
		\u0_uk_K_r4_reg[15]/NET0131 ,
		\u0_uk_K_r4_reg[7]/NET0131 ,
		_w30533_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name24707 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30534_
	);
	LUT3 #(
		.INIT('h40)
	) name24708 (
		_w30532_,
		_w30530_,
		_w30531_,
		_w30535_
	);
	LUT4 #(
		.INIT('hc963)
	) name24709 (
		decrypt_pad,
		\u0_R4_reg[23]/NET0131 ,
		\u0_uk_K_r4_reg[45]/NET0131 ,
		\u0_uk_K_r4_reg[49]/NET0131 ,
		_w30536_
	);
	LUT4 #(
		.INIT('h007f)
	) name24710 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30536_,
		_w30537_
	);
	LUT3 #(
		.INIT('h10)
	) name24711 (
		_w30535_,
		_w30534_,
		_w30537_,
		_w30538_
	);
	LUT4 #(
		.INIT('h0002)
	) name24712 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30539_
	);
	LUT4 #(
		.INIT('h27fd)
	) name24713 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30540_
	);
	LUT2 #(
		.INIT('h1)
	) name24714 (
		_w30530_,
		_w30536_,
		_w30541_
	);
	LUT4 #(
		.INIT('h0008)
	) name24715 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30536_,
		_w30542_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name24716 (
		_w30531_,
		_w30536_,
		_w30540_,
		_w30542_,
		_w30543_
	);
	LUT3 #(
		.INIT('h8a)
	) name24717 (
		_w30529_,
		_w30538_,
		_w30543_,
		_w30544_
	);
	LUT4 #(
		.INIT('h0060)
	) name24718 (
		_w30532_,
		_w30530_,
		_w30531_,
		_w30536_,
		_w30545_
	);
	LUT4 #(
		.INIT('h0200)
	) name24719 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30546_
	);
	LUT2 #(
		.INIT('h8)
	) name24720 (
		_w30530_,
		_w30536_,
		_w30547_
	);
	LUT4 #(
		.INIT('h0800)
	) name24721 (
		_w30532_,
		_w30530_,
		_w30531_,
		_w30536_,
		_w30548_
	);
	LUT4 #(
		.INIT('h0002)
	) name24722 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30536_,
		_w30549_
	);
	LUT4 #(
		.INIT('hfafd)
	) name24723 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30536_,
		_w30550_
	);
	LUT3 #(
		.INIT('h10)
	) name24724 (
		_w30546_,
		_w30548_,
		_w30550_,
		_w30551_
	);
	LUT4 #(
		.INIT('h0400)
	) name24725 (
		_w30532_,
		_w30533_,
		_w30531_,
		_w30536_,
		_w30552_
	);
	LUT4 #(
		.INIT('h0080)
	) name24726 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30553_
	);
	LUT2 #(
		.INIT('h1)
	) name24727 (
		_w30552_,
		_w30553_,
		_w30554_
	);
	LUT4 #(
		.INIT('h4555)
	) name24728 (
		_w30529_,
		_w30545_,
		_w30551_,
		_w30554_,
		_w30555_
	);
	LUT4 #(
		.INIT('hfbdf)
	) name24729 (
		_w30532_,
		_w30533_,
		_w30531_,
		_w30536_,
		_w30556_
	);
	LUT2 #(
		.INIT('h1)
	) name24730 (
		_w30530_,
		_w30556_,
		_w30557_
	);
	LUT4 #(
		.INIT('h0100)
	) name24731 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30558_
	);
	LUT4 #(
		.INIT('h7e7f)
	) name24732 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30559_
	);
	LUT3 #(
		.INIT('h01)
	) name24733 (
		_w30532_,
		_w30533_,
		_w30531_,
		_w30560_
	);
	LUT4 #(
		.INIT('hcacf)
	) name24734 (
		_w30530_,
		_w30559_,
		_w30536_,
		_w30560_,
		_w30561_
	);
	LUT2 #(
		.INIT('h4)
	) name24735 (
		_w30557_,
		_w30561_,
		_w30562_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name24736 (
		\u0_L4_reg[11]/NET0131 ,
		_w30555_,
		_w30544_,
		_w30562_,
		_w30563_
	);
	LUT4 #(
		.INIT('hc963)
	) name24737 (
		decrypt_pad,
		\u0_R4_reg[24]/NET0131 ,
		\u0_uk_K_r4_reg[38]/NET0131 ,
		\u0_uk_K_r4_reg[42]/NET0131 ,
		_w30564_
	);
	LUT4 #(
		.INIT('hc963)
	) name24738 (
		decrypt_pad,
		\u0_R4_reg[25]/NET0131 ,
		\u0_uk_K_r4_reg[14]/NET0131 ,
		\u0_uk_K_r4_reg[22]/NET0131 ,
		_w30565_
	);
	LUT4 #(
		.INIT('hc963)
	) name24739 (
		decrypt_pad,
		\u0_R4_reg[26]/NET0131 ,
		\u0_uk_K_r4_reg[30]/NET0131 ,
		\u0_uk_K_r4_reg[7]/NET0131 ,
		_w30566_
	);
	LUT4 #(
		.INIT('hc963)
	) name24740 (
		decrypt_pad,
		\u0_R4_reg[29]/NET0131 ,
		\u0_uk_K_r4_reg[42]/NET0131 ,
		\u0_uk_K_r4_reg[50]/NET0131 ,
		_w30567_
	);
	LUT4 #(
		.INIT('h0201)
	) name24741 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30568_
	);
	LUT4 #(
		.INIT('hc693)
	) name24742 (
		decrypt_pad,
		\u0_R4_reg[28]/NET0131 ,
		\u0_uk_K_r4_reg[31]/P0001 ,
		\u0_uk_K_r4_reg[50]/NET0131 ,
		_w30569_
	);
	LUT2 #(
		.INIT('h4)
	) name24743 (
		_w30568_,
		_w30569_,
		_w30570_
	);
	LUT3 #(
		.INIT('h72)
	) name24744 (
		_w30566_,
		_w30565_,
		_w30567_,
		_w30571_
	);
	LUT4 #(
		.INIT('hc693)
	) name24745 (
		decrypt_pad,
		\u0_R4_reg[27]/NET0131 ,
		\u0_uk_K_r4_reg[16]/NET0131 ,
		\u0_uk_K_r4_reg[8]/NET0131 ,
		_w30572_
	);
	LUT4 #(
		.INIT('hc800)
	) name24746 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30572_,
		_w30573_
	);
	LUT2 #(
		.INIT('h6)
	) name24747 (
		_w30564_,
		_w30565_,
		_w30574_
	);
	LUT4 #(
		.INIT('h0700)
	) name24748 (
		_w30566_,
		_w30564_,
		_w30572_,
		_w30567_,
		_w30575_
	);
	LUT4 #(
		.INIT('h0777)
	) name24749 (
		_w30571_,
		_w30573_,
		_w30574_,
		_w30575_,
		_w30576_
	);
	LUT2 #(
		.INIT('h8)
	) name24750 (
		_w30570_,
		_w30576_,
		_w30577_
	);
	LUT3 #(
		.INIT('h35)
	) name24751 (
		_w30566_,
		_w30564_,
		_w30572_,
		_w30578_
	);
	LUT4 #(
		.INIT('h0407)
	) name24752 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30579_
	);
	LUT2 #(
		.INIT('h4)
	) name24753 (
		_w30578_,
		_w30579_,
		_w30580_
	);
	LUT2 #(
		.INIT('h6)
	) name24754 (
		_w30566_,
		_w30564_,
		_w30581_
	);
	LUT3 #(
		.INIT('hb0)
	) name24755 (
		_w30565_,
		_w30572_,
		_w30567_,
		_w30582_
	);
	LUT2 #(
		.INIT('h4)
	) name24756 (
		_w30581_,
		_w30582_,
		_w30583_
	);
	LUT2 #(
		.INIT('h2)
	) name24757 (
		_w30564_,
		_w30572_,
		_w30584_
	);
	LUT3 #(
		.INIT('h45)
	) name24758 (
		_w30569_,
		_w30571_,
		_w30584_,
		_w30585_
	);
	LUT3 #(
		.INIT('h10)
	) name24759 (
		_w30580_,
		_w30583_,
		_w30585_,
		_w30586_
	);
	LUT4 #(
		.INIT('h006f)
	) name24760 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30572_,
		_w30587_
	);
	LUT4 #(
		.INIT('h0200)
	) name24761 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30588_
	);
	LUT4 #(
		.INIT('hfddf)
	) name24762 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30589_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name24763 (
		_w30564_,
		_w30565_,
		_w30572_,
		_w30567_,
		_w30590_
	);
	LUT4 #(
		.INIT('h0010)
	) name24764 (
		_w30566_,
		_w30565_,
		_w30572_,
		_w30567_,
		_w30591_
	);
	LUT4 #(
		.INIT('h00ea)
	) name24765 (
		_w30587_,
		_w30589_,
		_w30590_,
		_w30591_,
		_w30592_
	);
	LUT4 #(
		.INIT('ha955)
	) name24766 (
		\u0_L4_reg[22]/NET0131 ,
		_w30577_,
		_w30586_,
		_w30592_,
		_w30593_
	);
	LUT4 #(
		.INIT('h0400)
	) name24767 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30594_
	);
	LUT4 #(
		.INIT('hc9cd)
	) name24768 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30595_
	);
	LUT2 #(
		.INIT('h2)
	) name24769 (
		_w30500_,
		_w30595_,
		_w30596_
	);
	LUT4 #(
		.INIT('h4041)
	) name24770 (
		_w30500_,
		_w30499_,
		_w30502_,
		_w30501_,
		_w30597_
	);
	LUT4 #(
		.INIT('h0040)
	) name24771 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30598_
	);
	LUT3 #(
		.INIT('h80)
	) name24772 (
		_w30499_,
		_w30501_,
		_w30503_,
		_w30599_
	);
	LUT4 #(
		.INIT('h0002)
	) name24773 (
		_w30498_,
		_w30598_,
		_w30597_,
		_w30599_,
		_w30600_
	);
	LUT2 #(
		.INIT('h4)
	) name24774 (
		_w30596_,
		_w30600_,
		_w30601_
	);
	LUT4 #(
		.INIT('h0c13)
	) name24775 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30602_
	);
	LUT2 #(
		.INIT('h1)
	) name24776 (
		_w30500_,
		_w30602_,
		_w30603_
	);
	LUT4 #(
		.INIT('h0020)
	) name24777 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30604_
	);
	LUT3 #(
		.INIT('h82)
	) name24778 (
		_w30502_,
		_w30501_,
		_w30503_,
		_w30605_
	);
	LUT4 #(
		.INIT('h1000)
	) name24779 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30606_
	);
	LUT4 #(
		.INIT('h0002)
	) name24780 (
		_w30500_,
		_w30606_,
		_w30605_,
		_w30604_,
		_w30607_
	);
	LUT2 #(
		.INIT('h8)
	) name24781 (
		_w30499_,
		_w30502_,
		_w30608_
	);
	LUT4 #(
		.INIT('h0080)
	) name24782 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30609_
	);
	LUT3 #(
		.INIT('h01)
	) name24783 (
		_w30498_,
		_w30521_,
		_w30609_,
		_w30610_
	);
	LUT3 #(
		.INIT('he0)
	) name24784 (
		_w30603_,
		_w30607_,
		_w30610_,
		_w30611_
	);
	LUT3 #(
		.INIT('ha9)
	) name24785 (
		\u0_L4_reg[17]/NET0131 ,
		_w30601_,
		_w30611_,
		_w30612_
	);
	LUT4 #(
		.INIT('hc963)
	) name24786 (
		decrypt_pad,
		\u0_R4_reg[8]/NET0131 ,
		\u0_uk_K_r4_reg[20]/NET0131 ,
		\u0_uk_K_r4_reg[26]/NET0131 ,
		_w30613_
	);
	LUT4 #(
		.INIT('hc693)
	) name24787 (
		decrypt_pad,
		\u0_R4_reg[7]/NET0131 ,
		\u0_uk_K_r4_reg[3]/NET0131 ,
		\u0_uk_K_r4_reg[54]/NET0131 ,
		_w30614_
	);
	LUT4 #(
		.INIT('hc963)
	) name24788 (
		decrypt_pad,
		\u0_R4_reg[5]/NET0131 ,
		\u0_uk_K_r4_reg[12]/NET0131 ,
		\u0_uk_K_r4_reg[18]/NET0131 ,
		_w30615_
	);
	LUT4 #(
		.INIT('hc963)
	) name24789 (
		decrypt_pad,
		\u0_R4_reg[4]/NET0131 ,
		\u0_uk_K_r4_reg[33]/NET0131 ,
		\u0_uk_K_r4_reg[39]/NET0131 ,
		_w30616_
	);
	LUT4 #(
		.INIT('hc963)
	) name24790 (
		decrypt_pad,
		\u0_R4_reg[9]/NET0131 ,
		\u0_uk_K_r4_reg[25]/NET0131 ,
		\u0_uk_K_r4_reg[6]/NET0131 ,
		_w30617_
	);
	LUT3 #(
		.INIT('h04)
	) name24791 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30618_
	);
	LUT4 #(
		.INIT('hc963)
	) name24792 (
		decrypt_pad,
		\u0_R4_reg[6]/NET0131 ,
		\u0_uk_K_r4_reg[3]/NET0131 ,
		\u0_uk_K_r4_reg[41]/NET0131 ,
		_w30619_
	);
	LUT4 #(
		.INIT('h59fb)
	) name24793 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30620_
	);
	LUT2 #(
		.INIT('h1)
	) name24794 (
		_w30614_,
		_w30620_,
		_w30621_
	);
	LUT4 #(
		.INIT('h0034)
	) name24795 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30622_
	);
	LUT4 #(
		.INIT('h0800)
	) name24796 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30623_
	);
	LUT2 #(
		.INIT('h2)
	) name24797 (
		_w30617_,
		_w30619_,
		_w30624_
	);
	LUT4 #(
		.INIT('h0004)
	) name24798 (
		_w30614_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30625_
	);
	LUT4 #(
		.INIT('h4000)
	) name24799 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30626_
	);
	LUT4 #(
		.INIT('h0007)
	) name24800 (
		_w30614_,
		_w30623_,
		_w30625_,
		_w30626_,
		_w30627_
	);
	LUT4 #(
		.INIT('h5455)
	) name24801 (
		_w30613_,
		_w30621_,
		_w30622_,
		_w30627_,
		_w30628_
	);
	LUT4 #(
		.INIT('he6ee)
	) name24802 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30629_
	);
	LUT4 #(
		.INIT('h4044)
	) name24803 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30630_
	);
	LUT3 #(
		.INIT('h51)
	) name24804 (
		_w30614_,
		_w30615_,
		_w30619_,
		_w30631_
	);
	LUT4 #(
		.INIT('hf200)
	) name24805 (
		_w30613_,
		_w30629_,
		_w30630_,
		_w30631_,
		_w30632_
	);
	LUT3 #(
		.INIT('h10)
	) name24806 (
		_w30617_,
		_w30615_,
		_w30619_,
		_w30633_
	);
	LUT4 #(
		.INIT('h0100)
	) name24807 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30634_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name24808 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30635_
	);
	LUT2 #(
		.INIT('h2)
	) name24809 (
		_w30614_,
		_w30635_,
		_w30636_
	);
	LUT4 #(
		.INIT('h0002)
	) name24810 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30637_
	);
	LUT4 #(
		.INIT('h0080)
	) name24811 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30638_
	);
	LUT4 #(
		.INIT('h80a0)
	) name24812 (
		_w30614_,
		_w30616_,
		_w30615_,
		_w30619_,
		_w30639_
	);
	LUT4 #(
		.INIT('haaa8)
	) name24813 (
		_w30613_,
		_w30637_,
		_w30638_,
		_w30639_,
		_w30640_
	);
	LUT3 #(
		.INIT('h01)
	) name24814 (
		_w30636_,
		_w30640_,
		_w30632_,
		_w30641_
	);
	LUT3 #(
		.INIT('h65)
	) name24815 (
		\u0_L4_reg[2]/NET0131 ,
		_w30628_,
		_w30641_,
		_w30642_
	);
	LUT4 #(
		.INIT('hd97b)
	) name24816 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30643_
	);
	LUT2 #(
		.INIT('h2)
	) name24817 (
		_w30536_,
		_w30643_,
		_w30644_
	);
	LUT4 #(
		.INIT('h0040)
	) name24818 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30645_
	);
	LUT4 #(
		.INIT('heebf)
	) name24819 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30646_
	);
	LUT4 #(
		.INIT('h0302)
	) name24820 (
		_w30536_,
		_w30539_,
		_w30542_,
		_w30646_,
		_w30647_
	);
	LUT3 #(
		.INIT('h45)
	) name24821 (
		_w30529_,
		_w30644_,
		_w30647_,
		_w30648_
	);
	LUT3 #(
		.INIT('h8a)
	) name24822 (
		_w30532_,
		_w30533_,
		_w30531_,
		_w30649_
	);
	LUT2 #(
		.INIT('h2)
	) name24823 (
		_w30541_,
		_w30649_,
		_w30650_
	);
	LUT3 #(
		.INIT('h80)
	) name24824 (
		_w30533_,
		_w30530_,
		_w30531_,
		_w30651_
	);
	LUT4 #(
		.INIT('h0800)
	) name24825 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30536_,
		_w30652_
	);
	LUT3 #(
		.INIT('h01)
	) name24826 (
		_w30558_,
		_w30651_,
		_w30652_,
		_w30653_
	);
	LUT3 #(
		.INIT('h9e)
	) name24827 (
		_w30532_,
		_w30533_,
		_w30531_,
		_w30654_
	);
	LUT4 #(
		.INIT('h70d0)
	) name24828 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30655_
	);
	LUT4 #(
		.INIT('h00f1)
	) name24829 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30536_,
		_w30656_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name24830 (
		_w30547_,
		_w30654_,
		_w30655_,
		_w30656_,
		_w30657_
	);
	LUT4 #(
		.INIT('h7500)
	) name24831 (
		_w30529_,
		_w30650_,
		_w30653_,
		_w30657_,
		_w30658_
	);
	LUT3 #(
		.INIT('h65)
	) name24832 (
		\u0_L4_reg[4]/NET0131 ,
		_w30648_,
		_w30658_,
		_w30659_
	);
	LUT4 #(
		.INIT('hc693)
	) name24833 (
		decrypt_pad,
		\u0_R4_reg[31]/P0001 ,
		\u0_uk_K_r4_reg[45]/NET0131 ,
		\u0_uk_K_r4_reg[9]/NET0131 ,
		_w30660_
	);
	LUT4 #(
		.INIT('hc693)
	) name24834 (
		decrypt_pad,
		\u0_R4_reg[29]/NET0131 ,
		\u0_uk_K_r4_reg[28]/NET0131 ,
		\u0_uk_K_r4_reg[51]/NET0131 ,
		_w30661_
	);
	LUT4 #(
		.INIT('hc963)
	) name24835 (
		decrypt_pad,
		\u0_R4_reg[30]/NET0131 ,
		\u0_uk_K_r4_reg[21]/NET0131 ,
		\u0_uk_K_r4_reg[29]/NET0131 ,
		_w30662_
	);
	LUT4 #(
		.INIT('hc963)
	) name24836 (
		decrypt_pad,
		\u0_R4_reg[1]/NET0131 ,
		\u0_uk_K_r4_reg[36]/NET0131 ,
		\u0_uk_K_r4_reg[44]/NET0131 ,
		_w30663_
	);
	LUT4 #(
		.INIT('hc693)
	) name24837 (
		decrypt_pad,
		\u0_R4_reg[28]/NET0131 ,
		\u0_uk_K_r4_reg[1]/NET0131 ,
		\u0_uk_K_r4_reg[52]/NET0131 ,
		_w30664_
	);
	LUT4 #(
		.INIT('h0200)
	) name24838 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30665_
	);
	LUT4 #(
		.INIT('hc963)
	) name24839 (
		decrypt_pad,
		\u0_R4_reg[32]/NET0131 ,
		\u0_uk_K_r4_reg[15]/NET0131 ,
		\u0_uk_K_r4_reg[23]/P0001 ,
		_w30666_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name24840 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30667_
	);
	LUT4 #(
		.INIT('h0040)
	) name24841 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30668_
	);
	LUT4 #(
		.INIT('h0020)
	) name24842 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30669_
	);
	LUT3 #(
		.INIT('h01)
	) name24843 (
		_w30661_,
		_w30662_,
		_w30664_,
		_w30670_
	);
	LUT4 #(
		.INIT('h0001)
	) name24844 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30671_
	);
	LUT4 #(
		.INIT('hfb9e)
	) name24845 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30672_
	);
	LUT4 #(
		.INIT('hfd00)
	) name24846 (
		_w30666_,
		_w30667_,
		_w30665_,
		_w30672_,
		_w30673_
	);
	LUT2 #(
		.INIT('h2)
	) name24847 (
		_w30660_,
		_w30673_,
		_w30674_
	);
	LUT4 #(
		.INIT('haaa2)
	) name24848 (
		_w30660_,
		_w30661_,
		_w30663_,
		_w30662_,
		_w30675_
	);
	LUT4 #(
		.INIT('h00a2)
	) name24849 (
		_w30660_,
		_w30661_,
		_w30663_,
		_w30662_,
		_w30676_
	);
	LUT4 #(
		.INIT('h8f00)
	) name24850 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30677_
	);
	LUT2 #(
		.INIT('h4)
	) name24851 (
		_w30676_,
		_w30677_,
		_w30678_
	);
	LUT3 #(
		.INIT('h04)
	) name24852 (
		_w30663_,
		_w30662_,
		_w30664_,
		_w30679_
	);
	LUT3 #(
		.INIT('h15)
	) name24853 (
		_w30660_,
		_w30661_,
		_w30663_,
		_w30680_
	);
	LUT3 #(
		.INIT('h10)
	) name24854 (
		_w30665_,
		_w30679_,
		_w30680_,
		_w30681_
	);
	LUT4 #(
		.INIT('h1000)
	) name24855 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30682_
	);
	LUT4 #(
		.INIT('haa8a)
	) name24856 (
		_w30660_,
		_w30661_,
		_w30663_,
		_w30664_,
		_w30683_
	);
	LUT2 #(
		.INIT('h4)
	) name24857 (
		_w30682_,
		_w30683_,
		_w30684_
	);
	LUT4 #(
		.INIT('h0054)
	) name24858 (
		_w30666_,
		_w30681_,
		_w30684_,
		_w30678_,
		_w30685_
	);
	LUT4 #(
		.INIT('hadfa)
	) name24859 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30686_
	);
	LUT4 #(
		.INIT('h0080)
	) name24860 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30687_
	);
	LUT4 #(
		.INIT('h00c8)
	) name24861 (
		_w30660_,
		_w30666_,
		_w30686_,
		_w30687_,
		_w30688_
	);
	LUT4 #(
		.INIT('h999a)
	) name24862 (
		\u0_L4_reg[5]/NET0131 ,
		_w30674_,
		_w30685_,
		_w30688_,
		_w30689_
	);
	LUT4 #(
		.INIT('h67dc)
	) name24863 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30690_
	);
	LUT2 #(
		.INIT('h2)
	) name24864 (
		_w30536_,
		_w30690_,
		_w30691_
	);
	LUT4 #(
		.INIT('h2500)
	) name24865 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30692_
	);
	LUT4 #(
		.INIT('h0203)
	) name24866 (
		_w30536_,
		_w30542_,
		_w30645_,
		_w30692_,
		_w30693_
	);
	LUT3 #(
		.INIT('h45)
	) name24867 (
		_w30529_,
		_w30691_,
		_w30693_,
		_w30694_
	);
	LUT4 #(
		.INIT('h6f6e)
	) name24868 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30695_
	);
	LUT2 #(
		.INIT('h1)
	) name24869 (
		_w30536_,
		_w30695_,
		_w30696_
	);
	LUT4 #(
		.INIT('h9aff)
	) name24870 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30697_
	);
	LUT2 #(
		.INIT('h2)
	) name24871 (
		_w30536_,
		_w30697_,
		_w30698_
	);
	LUT4 #(
		.INIT('hffeb)
	) name24872 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30699_
	);
	LUT3 #(
		.INIT('h10)
	) name24873 (
		_w30553_,
		_w30549_,
		_w30699_,
		_w30700_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name24874 (
		_w30529_,
		_w30698_,
		_w30696_,
		_w30700_,
		_w30701_
	);
	LUT4 #(
		.INIT('h2000)
	) name24875 (
		_w30533_,
		_w30530_,
		_w30531_,
		_w30536_,
		_w30702_
	);
	LUT2 #(
		.INIT('h1)
	) name24876 (
		_w30539_,
		_w30702_,
		_w30703_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name24877 (
		\u0_L4_reg[29]/NET0131 ,
		_w30701_,
		_w30694_,
		_w30703_,
		_w30704_
	);
	LUT4 #(
		.INIT('hc693)
	) name24878 (
		decrypt_pad,
		\u0_R4_reg[13]/NET0131 ,
		\u0_uk_K_r4_reg[10]/NET0131 ,
		\u0_uk_K_r4_reg[4]/NET0131 ,
		_w30705_
	);
	LUT4 #(
		.INIT('hc963)
	) name24879 (
		decrypt_pad,
		\u0_R4_reg[15]/NET0131 ,
		\u0_uk_K_r4_reg[13]/NET0131 ,
		\u0_uk_K_r4_reg[19]/NET0131 ,
		_w30706_
	);
	LUT4 #(
		.INIT('hc693)
	) name24880 (
		decrypt_pad,
		\u0_R4_reg[14]/NET0131 ,
		\u0_uk_K_r4_reg[11]/NET0131 ,
		\u0_uk_K_r4_reg[5]/NET0131 ,
		_w30707_
	);
	LUT3 #(
		.INIT('h80)
	) name24881 (
		_w30705_,
		_w30706_,
		_w30707_,
		_w30708_
	);
	LUT4 #(
		.INIT('hc963)
	) name24882 (
		decrypt_pad,
		\u0_R4_reg[12]/NET0131 ,
		\u0_uk_K_r4_reg[10]/NET0131 ,
		\u0_uk_K_r4_reg[48]/NET0131 ,
		_w30709_
	);
	LUT4 #(
		.INIT('h0080)
	) name24883 (
		_w30705_,
		_w30706_,
		_w30707_,
		_w30709_,
		_w30710_
	);
	LUT4 #(
		.INIT('hc963)
	) name24884 (
		decrypt_pad,
		\u0_R4_reg[17]/NET0131 ,
		\u0_uk_K_r4_reg[26]/NET0131 ,
		\u0_uk_K_r4_reg[32]/NET0131 ,
		_w30711_
	);
	LUT4 #(
		.INIT('h8000)
	) name24885 (
		_w30705_,
		_w30706_,
		_w30709_,
		_w30711_,
		_w30712_
	);
	LUT4 #(
		.INIT('hc693)
	) name24886 (
		decrypt_pad,
		\u0_R4_reg[16]/NET0131 ,
		\u0_uk_K_r4_reg[27]/P0001 ,
		\u0_uk_K_r4_reg[46]/NET0131 ,
		_w30713_
	);
	LUT2 #(
		.INIT('h4)
	) name24887 (
		_w30705_,
		_w30706_,
		_w30714_
	);
	LUT4 #(
		.INIT('h0004)
	) name24888 (
		_w30705_,
		_w30706_,
		_w30709_,
		_w30711_,
		_w30715_
	);
	LUT2 #(
		.INIT('h4)
	) name24889 (
		_w30707_,
		_w30709_,
		_w30716_
	);
	LUT4 #(
		.INIT('h1000)
	) name24890 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30717_
	);
	LUT4 #(
		.INIT('h0001)
	) name24891 (
		_w30712_,
		_w30715_,
		_w30713_,
		_w30717_,
		_w30718_
	);
	LUT4 #(
		.INIT('hfff6)
	) name24892 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30719_
	);
	LUT4 #(
		.INIT('haa3f)
	) name24893 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30720_
	);
	LUT3 #(
		.INIT('hc8)
	) name24894 (
		_w30706_,
		_w30719_,
		_w30720_,
		_w30721_
	);
	LUT3 #(
		.INIT('h40)
	) name24895 (
		_w30710_,
		_w30718_,
		_w30721_,
		_w30722_
	);
	LUT4 #(
		.INIT('h0400)
	) name24896 (
		_w30705_,
		_w30706_,
		_w30709_,
		_w30711_,
		_w30723_
	);
	LUT4 #(
		.INIT('h0102)
	) name24897 (
		_w30705_,
		_w30706_,
		_w30707_,
		_w30709_,
		_w30724_
	);
	LUT4 #(
		.INIT('h8000)
	) name24898 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30725_
	);
	LUT4 #(
		.INIT('h0002)
	) name24899 (
		_w30713_,
		_w30724_,
		_w30725_,
		_w30723_,
		_w30726_
	);
	LUT4 #(
		.INIT('h0001)
	) name24900 (
		_w30705_,
		_w30706_,
		_w30709_,
		_w30711_,
		_w30727_
	);
	LUT4 #(
		.INIT('h0080)
	) name24901 (
		_w30705_,
		_w30706_,
		_w30709_,
		_w30711_,
		_w30728_
	);
	LUT2 #(
		.INIT('h4)
	) name24902 (
		_w30709_,
		_w30711_,
		_w30729_
	);
	LUT3 #(
		.INIT('h20)
	) name24903 (
		_w30705_,
		_w30709_,
		_w30711_,
		_w30730_
	);
	LUT4 #(
		.INIT('h0200)
	) name24904 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30731_
	);
	LUT2 #(
		.INIT('h1)
	) name24905 (
		_w30728_,
		_w30731_,
		_w30732_
	);
	LUT4 #(
		.INIT('h0207)
	) name24906 (
		_w30707_,
		_w30727_,
		_w30728_,
		_w30730_,
		_w30733_
	);
	LUT2 #(
		.INIT('h8)
	) name24907 (
		_w30726_,
		_w30733_,
		_w30734_
	);
	LUT3 #(
		.INIT('h01)
	) name24908 (
		_w30707_,
		_w30709_,
		_w30711_,
		_w30735_
	);
	LUT3 #(
		.INIT('hf6)
	) name24909 (
		_w30707_,
		_w30709_,
		_w30711_,
		_w30736_
	);
	LUT2 #(
		.INIT('h2)
	) name24910 (
		_w30714_,
		_w30736_,
		_w30737_
	);
	LUT4 #(
		.INIT('hcecf)
	) name24911 (
		_w30706_,
		_w30707_,
		_w30728_,
		_w30730_,
		_w30738_
	);
	LUT2 #(
		.INIT('h4)
	) name24912 (
		_w30737_,
		_w30738_,
		_w30739_
	);
	LUT4 #(
		.INIT('ha955)
	) name24913 (
		\u0_L4_reg[20]/NET0131 ,
		_w30722_,
		_w30734_,
		_w30739_,
		_w30740_
	);
	LUT4 #(
		.INIT('hebed)
	) name24914 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30741_
	);
	LUT2 #(
		.INIT('h1)
	) name24915 (
		_w30614_,
		_w30741_,
		_w30742_
	);
	LUT4 #(
		.INIT('haaa2)
	) name24916 (
		_w30614_,
		_w30616_,
		_w30617_,
		_w30615_,
		_w30743_
	);
	LUT4 #(
		.INIT('h0b2b)
	) name24917 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30744_
	);
	LUT2 #(
		.INIT('h8)
	) name24918 (
		_w30743_,
		_w30744_,
		_w30745_
	);
	LUT2 #(
		.INIT('h8)
	) name24919 (
		_w30614_,
		_w30616_,
		_w30746_
	);
	LUT3 #(
		.INIT('hb0)
	) name24920 (
		_w30617_,
		_w30615_,
		_w30619_,
		_w30747_
	);
	LUT3 #(
		.INIT('h32)
	) name24921 (
		_w30614_,
		_w30616_,
		_w30615_,
		_w30748_
	);
	LUT4 #(
		.INIT('h153f)
	) name24922 (
		_w30624_,
		_w30746_,
		_w30747_,
		_w30748_,
		_w30749_
	);
	LUT4 #(
		.INIT('h5455)
	) name24923 (
		_w30613_,
		_w30742_,
		_w30745_,
		_w30749_,
		_w30750_
	);
	LUT4 #(
		.INIT('h2000)
	) name24924 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30751_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name24925 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30752_
	);
	LUT2 #(
		.INIT('h1)
	) name24926 (
		_w30614_,
		_w30752_,
		_w30753_
	);
	LUT4 #(
		.INIT('h5515)
	) name24927 (
		_w30614_,
		_w30616_,
		_w30617_,
		_w30615_,
		_w30754_
	);
	LUT3 #(
		.INIT('h40)
	) name24928 (
		_w30616_,
		_w30617_,
		_w30619_,
		_w30755_
	);
	LUT4 #(
		.INIT('haaa8)
	) name24929 (
		_w30614_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30756_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name24930 (
		_w30633_,
		_w30754_,
		_w30755_,
		_w30756_,
		_w30757_
	);
	LUT4 #(
		.INIT('h0010)
	) name24931 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30758_
	);
	LUT4 #(
		.INIT('h0010)
	) name24932 (
		_w30625_,
		_w30626_,
		_w30752_,
		_w30758_,
		_w30759_
	);
	LUT4 #(
		.INIT('h1311)
	) name24933 (
		_w30613_,
		_w30753_,
		_w30757_,
		_w30759_,
		_w30760_
	);
	LUT3 #(
		.INIT('h9a)
	) name24934 (
		\u0_L4_reg[13]/NET0131 ,
		_w30750_,
		_w30760_,
		_w30761_
	);
	LUT3 #(
		.INIT('h20)
	) name24935 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30762_
	);
	LUT4 #(
		.INIT('h1000)
	) name24936 (
		_w30706_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30763_
	);
	LUT3 #(
		.INIT('h01)
	) name24937 (
		_w30727_,
		_w30762_,
		_w30763_,
		_w30764_
	);
	LUT2 #(
		.INIT('h4)
	) name24938 (
		_w30707_,
		_w30711_,
		_w30765_
	);
	LUT3 #(
		.INIT('h40)
	) name24939 (
		_w30705_,
		_w30706_,
		_w30709_,
		_w30766_
	);
	LUT4 #(
		.INIT('h0200)
	) name24940 (
		_w30706_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30767_
	);
	LUT3 #(
		.INIT('h0b)
	) name24941 (
		_w30765_,
		_w30766_,
		_w30767_,
		_w30768_
	);
	LUT4 #(
		.INIT('h1555)
	) name24942 (
		_w30713_,
		_w30719_,
		_w30764_,
		_w30768_,
		_w30769_
	);
	LUT4 #(
		.INIT('heff5)
	) name24943 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30770_
	);
	LUT2 #(
		.INIT('h2)
	) name24944 (
		_w30706_,
		_w30770_,
		_w30771_
	);
	LUT3 #(
		.INIT('hd0)
	) name24945 (
		_w30705_,
		_w30707_,
		_w30711_,
		_w30772_
	);
	LUT3 #(
		.INIT('h54)
	) name24946 (
		_w30706_,
		_w30709_,
		_w30711_,
		_w30773_
	);
	LUT4 #(
		.INIT('h8400)
	) name24947 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30774_
	);
	LUT4 #(
		.INIT('h00ef)
	) name24948 (
		_w30772_,
		_w30762_,
		_w30773_,
		_w30774_,
		_w30775_
	);
	LUT3 #(
		.INIT('h8a)
	) name24949 (
		_w30713_,
		_w30771_,
		_w30775_,
		_w30776_
	);
	LUT4 #(
		.INIT('h7bfe)
	) name24950 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30777_
	);
	LUT2 #(
		.INIT('h1)
	) name24951 (
		_w30706_,
		_w30777_,
		_w30778_
	);
	LUT3 #(
		.INIT('h23)
	) name24952 (
		_w30707_,
		_w30710_,
		_w30728_,
		_w30779_
	);
	LUT2 #(
		.INIT('h4)
	) name24953 (
		_w30778_,
		_w30779_,
		_w30780_
	);
	LUT4 #(
		.INIT('h5655)
	) name24954 (
		\u0_L4_reg[10]/NET0131 ,
		_w30776_,
		_w30769_,
		_w30780_,
		_w30781_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name24955 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30782_
	);
	LUT2 #(
		.INIT('h2)
	) name24956 (
		_w30572_,
		_w30782_,
		_w30783_
	);
	LUT4 #(
		.INIT('h1428)
	) name24957 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30784_
	);
	LUT4 #(
		.INIT('h00b0)
	) name24958 (
		_w30572_,
		_w30588_,
		_w30569_,
		_w30784_,
		_w30785_
	);
	LUT4 #(
		.INIT('h2816)
	) name24959 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30786_
	);
	LUT3 #(
		.INIT('h21)
	) name24960 (
		_w30565_,
		_w30572_,
		_w30567_,
		_w30787_
	);
	LUT3 #(
		.INIT('h08)
	) name24961 (
		_w30566_,
		_w30564_,
		_w30572_,
		_w30788_
	);
	LUT4 #(
		.INIT('h1000)
	) name24962 (
		_w30564_,
		_w30565_,
		_w30572_,
		_w30567_,
		_w30789_
	);
	LUT4 #(
		.INIT('h0001)
	) name24963 (
		_w30569_,
		_w30789_,
		_w30787_,
		_w30788_,
		_w30790_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name24964 (
		_w30783_,
		_w30785_,
		_w30786_,
		_w30790_,
		_w30791_
	);
	LUT2 #(
		.INIT('h6)
	) name24965 (
		\u0_L4_reg[12]/NET0131 ,
		_w30791_,
		_w30792_
	);
	LUT4 #(
		.INIT('h373f)
	) name24966 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30793_
	);
	LUT2 #(
		.INIT('h1)
	) name24967 (
		_w30500_,
		_w30793_,
		_w30794_
	);
	LUT4 #(
		.INIT('h0020)
	) name24968 (
		_w30500_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30795_
	);
	LUT4 #(
		.INIT('h00fe)
	) name24969 (
		_w30499_,
		_w30501_,
		_w30503_,
		_w30498_,
		_w30796_
	);
	LUT4 #(
		.INIT('h0800)
	) name24970 (
		_w30500_,
		_w30499_,
		_w30502_,
		_w30503_,
		_w30797_
	);
	LUT4 #(
		.INIT('h0100)
	) name24971 (
		_w30599_,
		_w30797_,
		_w30795_,
		_w30796_,
		_w30798_
	);
	LUT2 #(
		.INIT('h8)
	) name24972 (
		_w30516_,
		_w30507_,
		_w30799_
	);
	LUT4 #(
		.INIT('h004c)
	) name24973 (
		_w30518_,
		_w30498_,
		_w30525_,
		_w30594_,
		_w30800_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name24974 (
		_w30794_,
		_w30798_,
		_w30799_,
		_w30800_,
		_w30801_
	);
	LUT4 #(
		.INIT('hfcc7)
	) name24975 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30802_
	);
	LUT4 #(
		.INIT('h0140)
	) name24976 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w30803_
	);
	LUT4 #(
		.INIT('h5504)
	) name24977 (
		_w30500_,
		_w30498_,
		_w30802_,
		_w30803_,
		_w30804_
	);
	LUT3 #(
		.INIT('h40)
	) name24978 (
		_w30500_,
		_w30501_,
		_w30503_,
		_w30805_
	);
	LUT3 #(
		.INIT('hd9)
	) name24979 (
		_w30502_,
		_w30501_,
		_w30503_,
		_w30806_
	);
	LUT4 #(
		.INIT('h3f15)
	) name24980 (
		_w30513_,
		_w30608_,
		_w30805_,
		_w30806_,
		_w30807_
	);
	LUT2 #(
		.INIT('h4)
	) name24981 (
		_w30804_,
		_w30807_,
		_w30808_
	);
	LUT3 #(
		.INIT('h9a)
	) name24982 (
		\u0_L4_reg[23]/NET0131 ,
		_w30801_,
		_w30808_,
		_w30809_
	);
	LUT4 #(
		.INIT('h55b9)
	) name24983 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30810_
	);
	LUT4 #(
		.INIT('h0100)
	) name24984 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30811_
	);
	LUT4 #(
		.INIT('h3302)
	) name24985 (
		_w30660_,
		_w30666_,
		_w30810_,
		_w30811_,
		_w30812_
	);
	LUT4 #(
		.INIT('h0008)
	) name24986 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30813_
	);
	LUT4 #(
		.INIT('h4050)
	) name24987 (
		_w30661_,
		_w30662_,
		_w30664_,
		_w30666_,
		_w30814_
	);
	LUT4 #(
		.INIT('h0001)
	) name24988 (
		_w30669_,
		_w30671_,
		_w30814_,
		_w30813_,
		_w30815_
	);
	LUT2 #(
		.INIT('h1)
	) name24989 (
		_w30660_,
		_w30815_,
		_w30816_
	);
	LUT4 #(
		.INIT('h0004)
	) name24990 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30817_
	);
	LUT4 #(
		.INIT('hff7b)
	) name24991 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30818_
	);
	LUT2 #(
		.INIT('h2)
	) name24992 (
		_w30660_,
		_w30818_,
		_w30819_
	);
	LUT4 #(
		.INIT('h0002)
	) name24993 (
		_w30660_,
		_w30661_,
		_w30663_,
		_w30664_,
		_w30820_
	);
	LUT2 #(
		.INIT('h1)
	) name24994 (
		_w30669_,
		_w30820_,
		_w30821_
	);
	LUT4 #(
		.INIT('h4000)
	) name24995 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30822_
	);
	LUT3 #(
		.INIT('h20)
	) name24996 (
		_w30661_,
		_w30662_,
		_w30664_,
		_w30823_
	);
	LUT2 #(
		.INIT('h4)
	) name24997 (
		_w30660_,
		_w30663_,
		_w30824_
	);
	LUT4 #(
		.INIT('h1000)
	) name24998 (
		_w30660_,
		_w30661_,
		_w30663_,
		_w30662_,
		_w30825_
	);
	LUT3 #(
		.INIT('h01)
	) name24999 (
		_w30823_,
		_w30825_,
		_w30822_,
		_w30826_
	);
	LUT4 #(
		.INIT('h3111)
	) name25000 (
		_w30666_,
		_w30819_,
		_w30821_,
		_w30826_,
		_w30827_
	);
	LUT4 #(
		.INIT('h5655)
	) name25001 (
		\u0_L4_reg[15]/P0001 ,
		_w30812_,
		_w30816_,
		_w30827_,
		_w30828_
	);
	LUT4 #(
		.INIT('hbfae)
	) name25002 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30829_
	);
	LUT2 #(
		.INIT('h8)
	) name25003 (
		_w30614_,
		_w30829_,
		_w30830_
	);
	LUT3 #(
		.INIT('h10)
	) name25004 (
		_w30616_,
		_w30615_,
		_w30619_,
		_w30831_
	);
	LUT4 #(
		.INIT('h5b59)
	) name25005 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30832_
	);
	LUT4 #(
		.INIT('h0100)
	) name25006 (
		_w30614_,
		_w30751_,
		_w30831_,
		_w30832_,
		_w30833_
	);
	LUT4 #(
		.INIT('h0900)
	) name25007 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30834_
	);
	LUT3 #(
		.INIT('h01)
	) name25008 (
		_w30613_,
		_w30751_,
		_w30834_,
		_w30835_
	);
	LUT3 #(
		.INIT('he0)
	) name25009 (
		_w30830_,
		_w30833_,
		_w30835_,
		_w30836_
	);
	LUT4 #(
		.INIT('h0010)
	) name25010 (
		_w30614_,
		_w30751_,
		_w30829_,
		_w30831_,
		_w30837_
	);
	LUT4 #(
		.INIT('h1000)
	) name25011 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w30838_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name25012 (
		_w30614_,
		_w30616_,
		_w30617_,
		_w30615_,
		_w30839_
	);
	LUT2 #(
		.INIT('h4)
	) name25013 (
		_w30838_,
		_w30839_,
		_w30840_
	);
	LUT4 #(
		.INIT('h7737)
	) name25014 (
		_w30614_,
		_w30616_,
		_w30617_,
		_w30615_,
		_w30841_
	);
	LUT4 #(
		.INIT('h2a08)
	) name25015 (
		_w30613_,
		_w30619_,
		_w30618_,
		_w30841_,
		_w30842_
	);
	LUT3 #(
		.INIT('he0)
	) name25016 (
		_w30837_,
		_w30840_,
		_w30842_,
		_w30843_
	);
	LUT3 #(
		.INIT('ha9)
	) name25017 (
		\u0_L4_reg[28]/NET0131 ,
		_w30836_,
		_w30843_,
		_w30844_
	);
	LUT4 #(
		.INIT('hc963)
	) name25018 (
		decrypt_pad,
		\u0_R4_reg[21]/NET0131 ,
		\u0_uk_K_r4_reg[1]/NET0131 ,
		\u0_uk_K_r4_reg[9]/NET0131 ,
		_w30845_
	);
	LUT4 #(
		.INIT('hc693)
	) name25019 (
		decrypt_pad,
		\u0_R4_reg[16]/NET0131 ,
		\u0_uk_K_r4_reg[21]/NET0131 ,
		\u0_uk_K_r4_reg[44]/NET0131 ,
		_w30846_
	);
	LUT4 #(
		.INIT('hc963)
	) name25020 (
		decrypt_pad,
		\u0_R4_reg[17]/NET0131 ,
		\u0_uk_K_r4_reg[35]/NET0131 ,
		\u0_uk_K_r4_reg[43]/NET0131 ,
		_w30847_
	);
	LUT4 #(
		.INIT('hc963)
	) name25021 (
		decrypt_pad,
		\u0_R4_reg[18]/NET0131 ,
		\u0_uk_K_r4_reg[29]/NET0131 ,
		\u0_uk_K_r4_reg[37]/NET0131 ,
		_w30848_
	);
	LUT4 #(
		.INIT('h0400)
	) name25022 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30849_
	);
	LUT4 #(
		.INIT('hc963)
	) name25023 (
		decrypt_pad,
		\u0_R4_reg[19]/NET0131 ,
		\u0_uk_K_r4_reg[16]/NET0131 ,
		\u0_uk_K_r4_reg[52]/NET0131 ,
		_w30850_
	);
	LUT4 #(
		.INIT('h0200)
	) name25024 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30851_
	);
	LUT2 #(
		.INIT('h2)
	) name25025 (
		_w30847_,
		_w30848_,
		_w30852_
	);
	LUT4 #(
		.INIT('hafdf)
	) name25026 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30853_
	);
	LUT4 #(
		.INIT('he2ee)
	) name25027 (
		_w30849_,
		_w30850_,
		_w30851_,
		_w30853_,
		_w30854_
	);
	LUT4 #(
		.INIT('h0001)
	) name25028 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30855_
	);
	LUT4 #(
		.INIT('hf7f6)
	) name25029 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30856_
	);
	LUT4 #(
		.INIT('h1200)
	) name25030 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30857_
	);
	LUT4 #(
		.INIT('hc963)
	) name25031 (
		decrypt_pad,
		\u0_R4_reg[20]/NET0131 ,
		\u0_uk_K_r4_reg[0]/P0001 ,
		\u0_uk_K_r4_reg[8]/NET0131 ,
		_w30858_
	);
	LUT4 #(
		.INIT('hfd00)
	) name25032 (
		_w30846_,
		_w30848_,
		_w30850_,
		_w30858_,
		_w30859_
	);
	LUT4 #(
		.INIT('h0d00)
	) name25033 (
		_w30850_,
		_w30856_,
		_w30857_,
		_w30859_,
		_w30860_
	);
	LUT4 #(
		.INIT('h0004)
	) name25034 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30861_
	);
	LUT4 #(
		.INIT('h7f00)
	) name25035 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30850_,
		_w30862_
	);
	LUT4 #(
		.INIT('h2022)
	) name25036 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30863_
	);
	LUT4 #(
		.INIT('h00f7)
	) name25037 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30850_,
		_w30864_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name25038 (
		_w30861_,
		_w30862_,
		_w30863_,
		_w30864_,
		_w30865_
	);
	LUT4 #(
		.INIT('h0100)
	) name25039 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30866_
	);
	LUT4 #(
		.INIT('hbeff)
	) name25040 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30867_
	);
	LUT4 #(
		.INIT('h00fb)
	) name25041 (
		_w30846_,
		_w30847_,
		_w30848_,
		_w30858_,
		_w30868_
	);
	LUT2 #(
		.INIT('h8)
	) name25042 (
		_w30867_,
		_w30868_,
		_w30869_
	);
	LUT4 #(
		.INIT('h4544)
	) name25043 (
		_w30854_,
		_w30860_,
		_w30865_,
		_w30869_,
		_w30870_
	);
	LUT2 #(
		.INIT('h9)
	) name25044 (
		\u0_L4_reg[8]/NET0131 ,
		_w30870_,
		_w30871_
	);
	LUT4 #(
		.INIT('h5030)
	) name25045 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30872_
	);
	LUT4 #(
		.INIT('h0040)
	) name25046 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30873_
	);
	LUT4 #(
		.INIT('hfad8)
	) name25047 (
		_w30706_,
		_w30735_,
		_w30872_,
		_w30873_,
		_w30874_
	);
	LUT4 #(
		.INIT('h7ddf)
	) name25048 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30875_
	);
	LUT3 #(
		.INIT('h45)
	) name25049 (
		_w30713_,
		_w30874_,
		_w30875_,
		_w30876_
	);
	LUT3 #(
		.INIT('h10)
	) name25050 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30877_
	);
	LUT4 #(
		.INIT('haaef)
	) name25051 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30878_
	);
	LUT4 #(
		.INIT('h7bf7)
	) name25052 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30879_
	);
	LUT4 #(
		.INIT('h08aa)
	) name25053 (
		_w30706_,
		_w30713_,
		_w30878_,
		_w30879_,
		_w30880_
	);
	LUT4 #(
		.INIT('h0080)
	) name25054 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30881_
	);
	LUT4 #(
		.INIT('hd5fd)
	) name25055 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30882_
	);
	LUT4 #(
		.INIT('h5054)
	) name25056 (
		_w30706_,
		_w30713_,
		_w30881_,
		_w30882_,
		_w30883_
	);
	LUT4 #(
		.INIT('hfb7b)
	) name25057 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30884_
	);
	LUT4 #(
		.INIT('h5f13)
	) name25058 (
		_w30707_,
		_w30713_,
		_w30727_,
		_w30884_,
		_w30885_
	);
	LUT3 #(
		.INIT('h10)
	) name25059 (
		_w30883_,
		_w30880_,
		_w30885_,
		_w30886_
	);
	LUT3 #(
		.INIT('h65)
	) name25060 (
		\u0_L4_reg[1]/NET0131 ,
		_w30876_,
		_w30886_,
		_w30887_
	);
	LUT4 #(
		.INIT('h7fde)
	) name25061 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30888_
	);
	LUT2 #(
		.INIT('h1)
	) name25062 (
		_w30850_,
		_w30888_,
		_w30889_
	);
	LUT3 #(
		.INIT('h08)
	) name25063 (
		_w30847_,
		_w30848_,
		_w30850_,
		_w30890_
	);
	LUT4 #(
		.INIT('h4440)
	) name25064 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30891_
	);
	LUT2 #(
		.INIT('h4)
	) name25065 (
		_w30890_,
		_w30891_,
		_w30892_
	);
	LUT2 #(
		.INIT('h2)
	) name25066 (
		_w30847_,
		_w30850_,
		_w30893_
	);
	LUT3 #(
		.INIT('h08)
	) name25067 (
		_w30845_,
		_w30846_,
		_w30848_,
		_w30894_
	);
	LUT3 #(
		.INIT('h20)
	) name25068 (
		_w30845_,
		_w30846_,
		_w30850_,
		_w30895_
	);
	LUT4 #(
		.INIT('h8acf)
	) name25069 (
		_w30852_,
		_w30893_,
		_w30894_,
		_w30895_,
		_w30896_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name25070 (
		_w30858_,
		_w30889_,
		_w30892_,
		_w30896_,
		_w30897_
	);
	LUT4 #(
		.INIT('h0810)
	) name25071 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30898_
	);
	LUT4 #(
		.INIT('h0080)
	) name25072 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30899_
	);
	LUT4 #(
		.INIT('h00fd)
	) name25073 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30850_,
		_w30900_
	);
	LUT4 #(
		.INIT('haffb)
	) name25074 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30901_
	);
	LUT3 #(
		.INIT('h40)
	) name25075 (
		_w30899_,
		_w30900_,
		_w30901_,
		_w30902_
	);
	LUT4 #(
		.INIT('hfb00)
	) name25076 (
		_w30846_,
		_w30847_,
		_w30848_,
		_w30850_,
		_w30903_
	);
	LUT4 #(
		.INIT('h76fe)
	) name25077 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30904_
	);
	LUT2 #(
		.INIT('h8)
	) name25078 (
		_w30903_,
		_w30904_,
		_w30905_
	);
	LUT4 #(
		.INIT('h4445)
	) name25079 (
		_w30858_,
		_w30898_,
		_w30902_,
		_w30905_,
		_w30906_
	);
	LUT4 #(
		.INIT('h0040)
	) name25080 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30907_
	);
	LUT4 #(
		.INIT('heee4)
	) name25081 (
		_w30850_,
		_w30857_,
		_w30866_,
		_w30907_,
		_w30908_
	);
	LUT4 #(
		.INIT('h5556)
	) name25082 (
		\u0_L4_reg[14]/NET0131 ,
		_w30906_,
		_w30897_,
		_w30908_,
		_w30909_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name25083 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30910_
	);
	LUT2 #(
		.INIT('h2)
	) name25084 (
		_w30536_,
		_w30910_,
		_w30911_
	);
	LUT4 #(
		.INIT('hef00)
	) name25085 (
		_w30533_,
		_w30530_,
		_w30531_,
		_w30529_,
		_w30912_
	);
	LUT4 #(
		.INIT('h4000)
	) name25086 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30913_
	);
	LUT3 #(
		.INIT('h02)
	) name25087 (
		_w30532_,
		_w30531_,
		_w30536_,
		_w30914_
	);
	LUT4 #(
		.INIT('h0200)
	) name25088 (
		_w30699_,
		_w30913_,
		_w30914_,
		_w30912_,
		_w30915_
	);
	LUT3 #(
		.INIT('h45)
	) name25089 (
		_w30532_,
		_w30533_,
		_w30531_,
		_w30916_
	);
	LUT4 #(
		.INIT('hdf00)
	) name25090 (
		_w30532_,
		_w30530_,
		_w30531_,
		_w30536_,
		_w30917_
	);
	LUT2 #(
		.INIT('h4)
	) name25091 (
		_w30916_,
		_w30917_,
		_w30918_
	);
	LUT4 #(
		.INIT('h0041)
	) name25092 (
		_w30532_,
		_w30533_,
		_w30531_,
		_w30536_,
		_w30919_
	);
	LUT4 #(
		.INIT('h8000)
	) name25093 (
		_w30532_,
		_w30533_,
		_w30530_,
		_w30531_,
		_w30920_
	);
	LUT3 #(
		.INIT('h01)
	) name25094 (
		_w30529_,
		_w30919_,
		_w30920_,
		_w30921_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name25095 (
		_w30911_,
		_w30915_,
		_w30918_,
		_w30921_,
		_w30922_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name25096 (
		_w30530_,
		_w30531_,
		_w30556_,
		_w30542_,
		_w30923_
	);
	LUT3 #(
		.INIT('h65)
	) name25097 (
		\u0_L4_reg[19]/NET0131 ,
		_w30922_,
		_w30923_,
		_w30924_
	);
	LUT4 #(
		.INIT('h6c78)
	) name25098 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30925_
	);
	LUT4 #(
		.INIT('hf7c7)
	) name25099 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30926_
	);
	LUT4 #(
		.INIT('hbf5f)
	) name25100 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30927_
	);
	LUT4 #(
		.INIT('hd800)
	) name25101 (
		_w30850_,
		_w30925_,
		_w30926_,
		_w30927_,
		_w30928_
	);
	LUT2 #(
		.INIT('h2)
	) name25102 (
		_w30858_,
		_w30928_,
		_w30929_
	);
	LUT4 #(
		.INIT('hbefd)
	) name25103 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w30930_
	);
	LUT2 #(
		.INIT('h2)
	) name25104 (
		_w30850_,
		_w30930_,
		_w30931_
	);
	LUT3 #(
		.INIT('h0b)
	) name25105 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30932_
	);
	LUT3 #(
		.INIT('h8c)
	) name25106 (
		_w30846_,
		_w30847_,
		_w30848_,
		_w30933_
	);
	LUT2 #(
		.INIT('h4)
	) name25107 (
		_w30845_,
		_w30850_,
		_w30934_
	);
	LUT3 #(
		.INIT('h01)
	) name25108 (
		_w30933_,
		_w30932_,
		_w30934_,
		_w30935_
	);
	LUT3 #(
		.INIT('hb0)
	) name25109 (
		_w30845_,
		_w30847_,
		_w30850_,
		_w30936_
	);
	LUT4 #(
		.INIT('h0f01)
	) name25110 (
		_w30846_,
		_w30847_,
		_w30848_,
		_w30850_,
		_w30937_
	);
	LUT2 #(
		.INIT('h4)
	) name25111 (
		_w30936_,
		_w30937_,
		_w30938_
	);
	LUT4 #(
		.INIT('h0020)
	) name25112 (
		_w30846_,
		_w30847_,
		_w30848_,
		_w30850_,
		_w30939_
	);
	LUT2 #(
		.INIT('h1)
	) name25113 (
		_w30899_,
		_w30939_,
		_w30940_
	);
	LUT4 #(
		.INIT('hab00)
	) name25114 (
		_w30858_,
		_w30935_,
		_w30938_,
		_w30940_,
		_w30941_
	);
	LUT4 #(
		.INIT('h5655)
	) name25115 (
		\u0_L4_reg[25]/NET0131 ,
		_w30929_,
		_w30931_,
		_w30941_,
		_w30942_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name25116 (
		_w30705_,
		_w30706_,
		_w30709_,
		_w30711_,
		_w30943_
	);
	LUT3 #(
		.INIT('h31)
	) name25117 (
		_w30707_,
		_w30715_,
		_w30943_,
		_w30944_
	);
	LUT4 #(
		.INIT('h0eff)
	) name25118 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30945_
	);
	LUT3 #(
		.INIT('h45)
	) name25119 (
		_w30706_,
		_w30707_,
		_w30709_,
		_w30946_
	);
	LUT4 #(
		.INIT('h0082)
	) name25120 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30947_
	);
	LUT3 #(
		.INIT('h0b)
	) name25121 (
		_w30945_,
		_w30946_,
		_w30947_,
		_w30948_
	);
	LUT3 #(
		.INIT('h2a)
	) name25122 (
		_w30713_,
		_w30944_,
		_w30948_,
		_w30949_
	);
	LUT3 #(
		.INIT('h0d)
	) name25123 (
		_w30708_,
		_w30729_,
		_w30877_,
		_w30950_
	);
	LUT3 #(
		.INIT('h15)
	) name25124 (
		_w30713_,
		_w30732_,
		_w30950_,
		_w30951_
	);
	LUT4 #(
		.INIT('hfbaa)
	) name25125 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30952_
	);
	LUT4 #(
		.INIT('h2002)
	) name25126 (
		_w30705_,
		_w30707_,
		_w30709_,
		_w30711_,
		_w30953_
	);
	LUT4 #(
		.INIT('h5501)
	) name25127 (
		_w30706_,
		_w30713_,
		_w30952_,
		_w30953_,
		_w30954_
	);
	LUT3 #(
		.INIT('hbe)
	) name25128 (
		_w30705_,
		_w30706_,
		_w30711_,
		_w30955_
	);
	LUT4 #(
		.INIT('h5f13)
	) name25129 (
		_w30705_,
		_w30716_,
		_w30767_,
		_w30955_,
		_w30956_
	);
	LUT2 #(
		.INIT('h4)
	) name25130 (
		_w30954_,
		_w30956_,
		_w30957_
	);
	LUT4 #(
		.INIT('h5655)
	) name25131 (
		\u0_L4_reg[26]/NET0131 ,
		_w30949_,
		_w30951_,
		_w30957_,
		_w30958_
	);
	LUT4 #(
		.INIT('haa2a)
	) name25132 (
		_w30660_,
		_w30661_,
		_w30663_,
		_w30664_,
		_w30959_
	);
	LUT4 #(
		.INIT('h5bfb)
	) name25133 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30960_
	);
	LUT4 #(
		.INIT('h5455)
	) name25134 (
		_w30660_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30961_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name25135 (
		_w30822_,
		_w30959_,
		_w30960_,
		_w30961_,
		_w30962_
	);
	LUT4 #(
		.INIT('h2010)
	) name25136 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30963_
	);
	LUT3 #(
		.INIT('h02)
	) name25137 (
		_w30666_,
		_w30817_,
		_w30963_,
		_w30964_
	);
	LUT4 #(
		.INIT('h1001)
	) name25138 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30965_
	);
	LUT4 #(
		.INIT('h0004)
	) name25139 (
		_w30660_,
		_w30661_,
		_w30663_,
		_w30664_,
		_w30966_
	);
	LUT3 #(
		.INIT('h01)
	) name25140 (
		_w30666_,
		_w30965_,
		_w30966_,
		_w30967_
	);
	LUT4 #(
		.INIT('h8dff)
	) name25141 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30968_
	);
	LUT4 #(
		.INIT('hf31f)
	) name25142 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30969_
	);
	LUT4 #(
		.INIT('hf520)
	) name25143 (
		_w30660_,
		_w30661_,
		_w30968_,
		_w30969_,
		_w30970_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name25144 (
		_w30962_,
		_w30964_,
		_w30967_,
		_w30970_,
		_w30971_
	);
	LUT4 #(
		.INIT('h0002)
	) name25145 (
		_w30660_,
		_w30661_,
		_w30662_,
		_w30664_,
		_w30972_
	);
	LUT3 #(
		.INIT('h07)
	) name25146 (
		_w30823_,
		_w30824_,
		_w30972_,
		_w30973_
	);
	LUT3 #(
		.INIT('h65)
	) name25147 (
		\u0_L4_reg[21]/NET0131 ,
		_w30971_,
		_w30973_,
		_w30974_
	);
	LUT4 #(
		.INIT('h8802)
	) name25148 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30975_
	);
	LUT3 #(
		.INIT('hd7)
	) name25149 (
		_w30661_,
		_w30663_,
		_w30664_,
		_w30976_
	);
	LUT4 #(
		.INIT('he4f5)
	) name25150 (
		_w30660_,
		_w30670_,
		_w30975_,
		_w30976_,
		_w30977_
	);
	LUT4 #(
		.INIT('heb7b)
	) name25151 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30978_
	);
	LUT3 #(
		.INIT('h8a)
	) name25152 (
		_w30666_,
		_w30977_,
		_w30978_,
		_w30979_
	);
	LUT4 #(
		.INIT('hc4e4)
	) name25153 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30980_
	);
	LUT2 #(
		.INIT('h2)
	) name25154 (
		_w30675_,
		_w30980_,
		_w30981_
	);
	LUT4 #(
		.INIT('h4000)
	) name25155 (
		_w30660_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30982_
	);
	LUT3 #(
		.INIT('h01)
	) name25156 (
		_w30668_,
		_w30966_,
		_w30982_,
		_w30983_
	);
	LUT4 #(
		.INIT('hf9df)
	) name25157 (
		_w30661_,
		_w30663_,
		_w30662_,
		_w30664_,
		_w30984_
	);
	LUT4 #(
		.INIT('h0200)
	) name25158 (
		_w30660_,
		_w30661_,
		_w30663_,
		_w30662_,
		_w30985_
	);
	LUT3 #(
		.INIT('h0e)
	) name25159 (
		_w30660_,
		_w30984_,
		_w30985_,
		_w30986_
	);
	LUT4 #(
		.INIT('hba00)
	) name25160 (
		_w30666_,
		_w30981_,
		_w30983_,
		_w30986_,
		_w30987_
	);
	LUT3 #(
		.INIT('h65)
	) name25161 (
		\u0_L4_reg[27]/NET0131 ,
		_w30979_,
		_w30987_,
		_w30988_
	);
	LUT4 #(
		.INIT('h0002)
	) name25162 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30989_
	);
	LUT2 #(
		.INIT('h2)
	) name25163 (
		_w30572_,
		_w30569_,
		_w30990_
	);
	LUT4 #(
		.INIT('h936e)
	) name25164 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30991_
	);
	LUT2 #(
		.INIT('h2)
	) name25165 (
		_w30990_,
		_w30991_,
		_w30992_
	);
	LUT4 #(
		.INIT('h4410)
	) name25166 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30993_
	);
	LUT4 #(
		.INIT('h0800)
	) name25167 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30994_
	);
	LUT4 #(
		.INIT('hd77f)
	) name25168 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30995_
	);
	LUT2 #(
		.INIT('h4)
	) name25169 (
		_w30572_,
		_w30569_,
		_w30996_
	);
	LUT2 #(
		.INIT('h9)
	) name25170 (
		_w30572_,
		_w30569_,
		_w30997_
	);
	LUT3 #(
		.INIT('h20)
	) name25171 (
		_w30995_,
		_w30993_,
		_w30997_,
		_w30998_
	);
	LUT4 #(
		.INIT('h31e9)
	) name25172 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w30999_
	);
	LUT3 #(
		.INIT('h08)
	) name25173 (
		_w30995_,
		_w30996_,
		_w30999_,
		_w31000_
	);
	LUT4 #(
		.INIT('h00ab)
	) name25174 (
		_w30989_,
		_w30992_,
		_w30998_,
		_w31000_,
		_w31001_
	);
	LUT2 #(
		.INIT('h6)
	) name25175 (
		\u0_L4_reg[7]/NET0131 ,
		_w31001_,
		_w31002_
	);
	LUT4 #(
		.INIT('hf7bf)
	) name25176 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w31003_
	);
	LUT3 #(
		.INIT('h10)
	) name25177 (
		_w30850_,
		_w30855_,
		_w31003_,
		_w31004_
	);
	LUT3 #(
		.INIT('h02)
	) name25178 (
		_w30850_,
		_w30851_,
		_w30861_,
		_w31005_
	);
	LUT2 #(
		.INIT('h1)
	) name25179 (
		_w31004_,
		_w31005_,
		_w31006_
	);
	LUT4 #(
		.INIT('hbf9d)
	) name25180 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w31007_
	);
	LUT2 #(
		.INIT('h2)
	) name25181 (
		_w30850_,
		_w31007_,
		_w31008_
	);
	LUT3 #(
		.INIT('hb0)
	) name25182 (
		_w30847_,
		_w30848_,
		_w30850_,
		_w31009_
	);
	LUT4 #(
		.INIT('h44e6)
	) name25183 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w31010_
	);
	LUT3 #(
		.INIT('h54)
	) name25184 (
		_w30858_,
		_w31009_,
		_w31010_,
		_w31011_
	);
	LUT4 #(
		.INIT('hef67)
	) name25185 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30848_,
		_w31012_
	);
	LUT2 #(
		.INIT('h2)
	) name25186 (
		_w30850_,
		_w31012_,
		_w31013_
	);
	LUT4 #(
		.INIT('h0020)
	) name25187 (
		_w30845_,
		_w30846_,
		_w30847_,
		_w30850_,
		_w31014_
	);
	LUT4 #(
		.INIT('h0004)
	) name25188 (
		_w30849_,
		_w30858_,
		_w30899_,
		_w31014_,
		_w31015_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name25189 (
		_w31008_,
		_w31011_,
		_w31013_,
		_w31015_,
		_w31016_
	);
	LUT3 #(
		.INIT('h56)
	) name25190 (
		\u0_L4_reg[3]/NET0131 ,
		_w31006_,
		_w31016_,
		_w31017_
	);
	LUT4 #(
		.INIT('hc963)
	) name25191 (
		decrypt_pad,
		\u0_R4_reg[13]/NET0131 ,
		\u0_uk_K_r4_reg[11]/NET0131 ,
		\u0_uk_K_r4_reg[17]/NET0131 ,
		_w31018_
	);
	LUT4 #(
		.INIT('hc693)
	) name25192 (
		decrypt_pad,
		\u0_R4_reg[9]/NET0131 ,
		\u0_uk_K_r4_reg[12]/NET0131 ,
		\u0_uk_K_r4_reg[6]/NET0131 ,
		_w31019_
	);
	LUT2 #(
		.INIT('h9)
	) name25193 (
		_w31018_,
		_w31019_,
		_w31020_
	);
	LUT4 #(
		.INIT('hc963)
	) name25194 (
		decrypt_pad,
		\u0_R4_reg[11]/NET0131 ,
		\u0_uk_K_r4_reg[40]/NET0131 ,
		\u0_uk_K_r4_reg[46]/NET0131 ,
		_w31021_
	);
	LUT4 #(
		.INIT('hc963)
	) name25195 (
		decrypt_pad,
		\u0_R4_reg[8]/NET0131 ,
		\u0_uk_K_r4_reg[34]/NET0131 ,
		\u0_uk_K_r4_reg[40]/NET0131 ,
		_w31022_
	);
	LUT4 #(
		.INIT('hc693)
	) name25196 (
		decrypt_pad,
		\u0_R4_reg[10]/NET0131 ,
		\u0_uk_K_r4_reg[20]/NET0131 ,
		\u0_uk_K_r4_reg[39]/NET0131 ,
		_w31023_
	);
	LUT4 #(
		.INIT('h00ae)
	) name25197 (
		_w31022_,
		_w31019_,
		_w31023_,
		_w31021_,
		_w31024_
	);
	LUT4 #(
		.INIT('h1000)
	) name25198 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31025_
	);
	LUT4 #(
		.INIT('hc693)
	) name25199 (
		decrypt_pad,
		\u0_R4_reg[12]/NET0131 ,
		\u0_uk_K_r4_reg[4]/NET0131 ,
		\u0_uk_K_r4_reg[55]/NET0131 ,
		_w31026_
	);
	LUT4 #(
		.INIT('h1500)
	) name25200 (
		_w31025_,
		_w31020_,
		_w31024_,
		_w31026_,
		_w31027_
	);
	LUT2 #(
		.INIT('h6)
	) name25201 (
		_w31022_,
		_w31018_,
		_w31028_
	);
	LUT4 #(
		.INIT('h9990)
	) name25202 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31029_
	);
	LUT4 #(
		.INIT('h0990)
	) name25203 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31030_
	);
	LUT2 #(
		.INIT('h4)
	) name25204 (
		_w31022_,
		_w31018_,
		_w31031_
	);
	LUT3 #(
		.INIT('h08)
	) name25205 (
		_w31019_,
		_w31023_,
		_w31021_,
		_w31032_
	);
	LUT4 #(
		.INIT('h0400)
	) name25206 (
		_w31022_,
		_w31019_,
		_w31023_,
		_w31021_,
		_w31033_
	);
	LUT4 #(
		.INIT('h0015)
	) name25207 (
		_w31026_,
		_w31031_,
		_w31032_,
		_w31033_,
		_w31034_
	);
	LUT4 #(
		.INIT('h2000)
	) name25208 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31035_
	);
	LUT4 #(
		.INIT('h0203)
	) name25209 (
		_w31022_,
		_w31019_,
		_w31023_,
		_w31021_,
		_w31036_
	);
	LUT3 #(
		.INIT('h13)
	) name25210 (
		_w31028_,
		_w31035_,
		_w31036_,
		_w31037_
	);
	LUT4 #(
		.INIT('h4555)
	) name25211 (
		_w31027_,
		_w31030_,
		_w31034_,
		_w31037_,
		_w31038_
	);
	LUT4 #(
		.INIT('h93d3)
	) name25212 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31039_
	);
	LUT4 #(
		.INIT('h0001)
	) name25213 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31040_
	);
	LUT4 #(
		.INIT('hf3fe)
	) name25214 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31041_
	);
	LUT4 #(
		.INIT('h08aa)
	) name25215 (
		_w31021_,
		_w31026_,
		_w31039_,
		_w31041_,
		_w31042_
	);
	LUT3 #(
		.INIT('h56)
	) name25216 (
		\u0_L4_reg[6]/NET0131 ,
		_w31038_,
		_w31042_,
		_w31043_
	);
	LUT4 #(
		.INIT('h0080)
	) name25217 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w31044_
	);
	LUT4 #(
		.INIT('h0104)
	) name25218 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w31045_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name25219 (
		_w30564_,
		_w30565_,
		_w30572_,
		_w30567_,
		_w31046_
	);
	LUT3 #(
		.INIT('h10)
	) name25220 (
		_w30994_,
		_w31045_,
		_w31046_,
		_w31047_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name25221 (
		_w30564_,
		_w30565_,
		_w30572_,
		_w30567_,
		_w31048_
	);
	LUT4 #(
		.INIT('haf77)
	) name25222 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w31049_
	);
	LUT2 #(
		.INIT('h8)
	) name25223 (
		_w31048_,
		_w31049_,
		_w31050_
	);
	LUT4 #(
		.INIT('h888a)
	) name25224 (
		_w30569_,
		_w31044_,
		_w31047_,
		_w31050_,
		_w31051_
	);
	LUT3 #(
		.INIT('h04)
	) name25225 (
		_w30566_,
		_w30564_,
		_w30567_,
		_w31052_
	);
	LUT4 #(
		.INIT('hf3bb)
	) name25226 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w31053_
	);
	LUT2 #(
		.INIT('h2)
	) name25227 (
		_w30572_,
		_w31053_,
		_w31054_
	);
	LUT4 #(
		.INIT('h7d9f)
	) name25228 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w31055_
	);
	LUT3 #(
		.INIT('hd0)
	) name25229 (
		_w30787_,
		_w31052_,
		_w31055_,
		_w31056_
	);
	LUT4 #(
		.INIT('h8fcf)
	) name25230 (
		_w30566_,
		_w30564_,
		_w30565_,
		_w30567_,
		_w31057_
	);
	LUT3 #(
		.INIT('h0e)
	) name25231 (
		_w30566_,
		_w30564_,
		_w30572_,
		_w31058_
	);
	LUT4 #(
		.INIT('h7077)
	) name25232 (
		_w30566_,
		_w30789_,
		_w31057_,
		_w31058_,
		_w31059_
	);
	LUT4 #(
		.INIT('hba00)
	) name25233 (
		_w30569_,
		_w31054_,
		_w31056_,
		_w31059_,
		_w31060_
	);
	LUT3 #(
		.INIT('h65)
	) name25234 (
		\u0_L4_reg[32]/NET0131 ,
		_w31051_,
		_w31060_,
		_w31061_
	);
	LUT3 #(
		.INIT('h43)
	) name25235 (
		_w30502_,
		_w30501_,
		_w30503_,
		_w31062_
	);
	LUT4 #(
		.INIT('h1005)
	) name25236 (
		_w30500_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w31063_
	);
	LUT2 #(
		.INIT('h1)
	) name25237 (
		_w30498_,
		_w31063_,
		_w31064_
	);
	LUT3 #(
		.INIT('h40)
	) name25238 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w31065_
	);
	LUT4 #(
		.INIT('h4802)
	) name25239 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w31066_
	);
	LUT3 #(
		.INIT('h28)
	) name25240 (
		_w30500_,
		_w30501_,
		_w30503_,
		_w31067_
	);
	LUT3 #(
		.INIT('h23)
	) name25241 (
		_w31065_,
		_w31066_,
		_w31067_,
		_w31068_
	);
	LUT4 #(
		.INIT('h8228)
	) name25242 (
		_w30499_,
		_w30502_,
		_w30501_,
		_w30503_,
		_w31069_
	);
	LUT4 #(
		.INIT('h040c)
	) name25243 (
		_w30513_,
		_w30498_,
		_w30598_,
		_w31062_,
		_w31070_
	);
	LUT4 #(
		.INIT('h7077)
	) name25244 (
		_w31064_,
		_w31068_,
		_w31069_,
		_w31070_,
		_w31071_
	);
	LUT2 #(
		.INIT('h6)
	) name25245 (
		_w30499_,
		_w30502_,
		_w31072_
	);
	LUT2 #(
		.INIT('h8)
	) name25246 (
		_w30805_,
		_w31072_,
		_w31073_
	);
	LUT3 #(
		.INIT('h56)
	) name25247 (
		\u0_L4_reg[9]/NET0131 ,
		_w31071_,
		_w31073_,
		_w31074_
	);
	LUT4 #(
		.INIT('h45cf)
	) name25248 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31075_
	);
	LUT4 #(
		.INIT('hbf00)
	) name25249 (
		_w31018_,
		_w31019_,
		_w31023_,
		_w31021_,
		_w31076_
	);
	LUT3 #(
		.INIT('h0e)
	) name25250 (
		_w31022_,
		_w31019_,
		_w31021_,
		_w31077_
	);
	LUT4 #(
		.INIT('hfbf6)
	) name25251 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31078_
	);
	LUT4 #(
		.INIT('h2700)
	) name25252 (
		_w31075_,
		_w31077_,
		_w31076_,
		_w31078_,
		_w31079_
	);
	LUT2 #(
		.INIT('h1)
	) name25253 (
		_w31026_,
		_w31079_,
		_w31080_
	);
	LUT3 #(
		.INIT('heb)
	) name25254 (
		_w31022_,
		_w31018_,
		_w31023_,
		_w31081_
	);
	LUT4 #(
		.INIT('h0002)
	) name25255 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31082_
	);
	LUT3 #(
		.INIT('h08)
	) name25256 (
		_w31021_,
		_w31081_,
		_w31082_,
		_w31083_
	);
	LUT3 #(
		.INIT('h10)
	) name25257 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31084_
	);
	LUT3 #(
		.INIT('h07)
	) name25258 (
		_w31022_,
		_w31023_,
		_w31021_,
		_w31085_
	);
	LUT3 #(
		.INIT('h8a)
	) name25259 (
		_w31026_,
		_w31084_,
		_w31085_,
		_w31086_
	);
	LUT3 #(
		.INIT('h20)
	) name25260 (
		_w31022_,
		_w31019_,
		_w31023_,
		_w31087_
	);
	LUT2 #(
		.INIT('h8)
	) name25261 (
		_w31018_,
		_w31021_,
		_w31088_
	);
	LUT3 #(
		.INIT('h0e)
	) name25262 (
		_w31018_,
		_w31021_,
		_w31026_,
		_w31089_
	);
	LUT4 #(
		.INIT('h7000)
	) name25263 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31090_
	);
	LUT4 #(
		.INIT('h7077)
	) name25264 (
		_w31087_,
		_w31088_,
		_w31089_,
		_w31090_,
		_w31091_
	);
	LUT3 #(
		.INIT('hb0)
	) name25265 (
		_w31083_,
		_w31086_,
		_w31091_,
		_w31092_
	);
	LUT3 #(
		.INIT('h9a)
	) name25266 (
		\u0_L4_reg[30]/NET0131 ,
		_w31080_,
		_w31092_,
		_w31093_
	);
	LUT4 #(
		.INIT('h6979)
	) name25267 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31021_,
		_w31094_
	);
	LUT4 #(
		.INIT('h4000)
	) name25268 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31095_
	);
	LUT4 #(
		.INIT('h0012)
	) name25269 (
		_w31022_,
		_w31018_,
		_w31023_,
		_w31021_,
		_w31096_
	);
	LUT4 #(
		.INIT('h0032)
	) name25270 (
		_w31023_,
		_w31095_,
		_w31094_,
		_w31096_,
		_w31097_
	);
	LUT4 #(
		.INIT('h7b6a)
	) name25271 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31098_
	);
	LUT4 #(
		.INIT('h6800)
	) name25272 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31021_,
		_w31099_
	);
	LUT4 #(
		.INIT('h0032)
	) name25273 (
		_w31021_,
		_w31040_,
		_w31098_,
		_w31099_,
		_w31100_
	);
	LUT4 #(
		.INIT('hdeff)
	) name25274 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31101_
	);
	LUT4 #(
		.INIT('h0020)
	) name25275 (
		_w31022_,
		_w31019_,
		_w31023_,
		_w31021_,
		_w31102_
	);
	LUT3 #(
		.INIT('h0d)
	) name25276 (
		_w31021_,
		_w31101_,
		_w31102_,
		_w31103_
	);
	LUT4 #(
		.INIT('hd800)
	) name25277 (
		_w31026_,
		_w31097_,
		_w31100_,
		_w31103_,
		_w31104_
	);
	LUT2 #(
		.INIT('h9)
	) name25278 (
		\u0_L4_reg[16]/NET0131 ,
		_w31104_,
		_w31105_
	);
	LUT4 #(
		.INIT('h1003)
	) name25279 (
		_w30614_,
		_w30616_,
		_w30615_,
		_w30619_,
		_w31106_
	);
	LUT4 #(
		.INIT('hf7fc)
	) name25280 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w31107_
	);
	LUT4 #(
		.INIT('h8000)
	) name25281 (
		_w30614_,
		_w30616_,
		_w30617_,
		_w30615_,
		_w31108_
	);
	LUT4 #(
		.INIT('h0100)
	) name25282 (
		_w30613_,
		_w30751_,
		_w31108_,
		_w31107_,
		_w31109_
	);
	LUT4 #(
		.INIT('hfd75)
	) name25283 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w31110_
	);
	LUT2 #(
		.INIT('h1)
	) name25284 (
		_w30614_,
		_w31110_,
		_w31111_
	);
	LUT4 #(
		.INIT('h0a20)
	) name25285 (
		_w30614_,
		_w30616_,
		_w30617_,
		_w30615_,
		_w31112_
	);
	LUT3 #(
		.INIT('h02)
	) name25286 (
		_w30613_,
		_w30634_,
		_w31112_,
		_w31113_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name25287 (
		_w31106_,
		_w31109_,
		_w31111_,
		_w31113_,
		_w31114_
	);
	LUT4 #(
		.INIT('h77ef)
	) name25288 (
		_w30616_,
		_w30617_,
		_w30615_,
		_w30619_,
		_w31115_
	);
	LUT4 #(
		.INIT('h1000)
	) name25289 (
		_w30614_,
		_w30616_,
		_w30617_,
		_w30615_,
		_w31116_
	);
	LUT3 #(
		.INIT('h0d)
	) name25290 (
		_w30614_,
		_w31115_,
		_w31116_,
		_w31117_
	);
	LUT3 #(
		.INIT('h65)
	) name25291 (
		\u0_L4_reg[18]/NET0131 ,
		_w31114_,
		_w31117_,
		_w31118_
	);
	LUT4 #(
		.INIT('h0200)
	) name25292 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31119_
	);
	LUT4 #(
		.INIT('he4ab)
	) name25293 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31120_
	);
	LUT4 #(
		.INIT('h3032)
	) name25294 (
		_w31021_,
		_w31026_,
		_w31119_,
		_w31120_,
		_w31121_
	);
	LUT2 #(
		.INIT('h4)
	) name25295 (
		_w31021_,
		_w31029_,
		_w31122_
	);
	LUT4 #(
		.INIT('h1bff)
	) name25296 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31123_
	);
	LUT2 #(
		.INIT('h2)
	) name25297 (
		_w31021_,
		_w31123_,
		_w31124_
	);
	LUT2 #(
		.INIT('h4)
	) name25298 (
		_w31023_,
		_w31021_,
		_w31125_
	);
	LUT3 #(
		.INIT('h0b)
	) name25299 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31126_
	);
	LUT4 #(
		.INIT('h0777)
	) name25300 (
		_w31028_,
		_w31036_,
		_w31125_,
		_w31126_,
		_w31127_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name25301 (
		_w31026_,
		_w31124_,
		_w31122_,
		_w31127_,
		_w31128_
	);
	LUT4 #(
		.INIT('h9bd6)
	) name25302 (
		_w31022_,
		_w31018_,
		_w31019_,
		_w31023_,
		_w31129_
	);
	LUT2 #(
		.INIT('h1)
	) name25303 (
		_w31021_,
		_w31026_,
		_w31130_
	);
	LUT2 #(
		.INIT('h4)
	) name25304 (
		_w31129_,
		_w31130_,
		_w31131_
	);
	LUT4 #(
		.INIT('h0900)
	) name25305 (
		_w31018_,
		_w31019_,
		_w31023_,
		_w31021_,
		_w31132_
	);
	LUT4 #(
		.INIT('h197f)
	) name25306 (
		_w31022_,
		_w31018_,
		_w31032_,
		_w31132_,
		_w31133_
	);
	LUT2 #(
		.INIT('h4)
	) name25307 (
		_w31131_,
		_w31133_,
		_w31134_
	);
	LUT4 #(
		.INIT('h5655)
	) name25308 (
		\u0_L4_reg[24]/NET0131 ,
		_w31128_,
		_w31121_,
		_w31134_,
		_w31135_
	);
	LUT4 #(
		.INIT('hc963)
	) name25309 (
		decrypt_pad,
		\u0_R3_reg[28]/NET0131 ,
		\u0_uk_K_r3_reg[36]/NET0131 ,
		\u0_uk_K_r3_reg[45]/P0001 ,
		_w31136_
	);
	LUT4 #(
		.INIT('hc693)
	) name25310 (
		decrypt_pad,
		\u0_R3_reg[27]/NET0131 ,
		\u0_uk_K_r3_reg[30]/NET0131 ,
		\u0_uk_K_r3_reg[49]/NET0131 ,
		_w31137_
	);
	LUT4 #(
		.INIT('hc963)
	) name25311 (
		decrypt_pad,
		\u0_R3_reg[26]/NET0131 ,
		\u0_uk_K_r3_reg[16]/NET0131 ,
		\u0_uk_K_r3_reg[21]/NET0131 ,
		_w31138_
	);
	LUT4 #(
		.INIT('hc693)
	) name25312 (
		decrypt_pad,
		\u0_R3_reg[24]/NET0131 ,
		\u0_uk_K_r3_reg[1]/NET0131 ,
		\u0_uk_K_r3_reg[51]/NET0131 ,
		_w31139_
	);
	LUT4 #(
		.INIT('hc963)
	) name25313 (
		decrypt_pad,
		\u0_R3_reg[29]/NET0131 ,
		\u0_uk_K_r3_reg[28]/NET0131 ,
		\u0_uk_K_r3_reg[9]/NET0131 ,
		_w31140_
	);
	LUT2 #(
		.INIT('h4)
	) name25314 (
		_w31139_,
		_w31140_,
		_w31141_
	);
	LUT4 #(
		.INIT('hc963)
	) name25315 (
		decrypt_pad,
		\u0_R3_reg[25]/NET0131 ,
		\u0_uk_K_r3_reg[0]/NET0131 ,
		\u0_uk_K_r3_reg[36]/NET0131 ,
		_w31142_
	);
	LUT4 #(
		.INIT('h5f67)
	) name25316 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31143_
	);
	LUT2 #(
		.INIT('h1)
	) name25317 (
		_w31137_,
		_w31143_,
		_w31144_
	);
	LUT4 #(
		.INIT('hbdad)
	) name25318 (
		_w31139_,
		_w31142_,
		_w31140_,
		_w31137_,
		_w31145_
	);
	LUT4 #(
		.INIT('h8000)
	) name25319 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31146_
	);
	LUT4 #(
		.INIT('h0200)
	) name25320 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31137_,
		_w31147_
	);
	LUT4 #(
		.INIT('h0032)
	) name25321 (
		_w31138_,
		_w31146_,
		_w31145_,
		_w31147_,
		_w31148_
	);
	LUT3 #(
		.INIT('h45)
	) name25322 (
		_w31136_,
		_w31144_,
		_w31148_,
		_w31149_
	);
	LUT2 #(
		.INIT('h6)
	) name25323 (
		_w31142_,
		_w31138_,
		_w31150_
	);
	LUT4 #(
		.INIT('ha800)
	) name25324 (
		_w31139_,
		_w31138_,
		_w31140_,
		_w31137_,
		_w31151_
	);
	LUT2 #(
		.INIT('h8)
	) name25325 (
		_w31150_,
		_w31151_,
		_w31152_
	);
	LUT4 #(
		.INIT('h1001)
	) name25326 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31153_
	);
	LUT2 #(
		.INIT('h9)
	) name25327 (
		_w31139_,
		_w31142_,
		_w31154_
	);
	LUT4 #(
		.INIT('h0070)
	) name25328 (
		_w31139_,
		_w31138_,
		_w31140_,
		_w31137_,
		_w31155_
	);
	LUT3 #(
		.INIT('h45)
	) name25329 (
		_w31153_,
		_w31154_,
		_w31155_,
		_w31156_
	);
	LUT4 #(
		.INIT('h1000)
	) name25330 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31157_
	);
	LUT4 #(
		.INIT('hef9d)
	) name25331 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31158_
	);
	LUT4 #(
		.INIT('h0100)
	) name25332 (
		_w31142_,
		_w31138_,
		_w31140_,
		_w31137_,
		_w31159_
	);
	LUT4 #(
		.INIT('h0084)
	) name25333 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31137_,
		_w31160_
	);
	LUT4 #(
		.INIT('h0031)
	) name25334 (
		_w31137_,
		_w31159_,
		_w31158_,
		_w31160_,
		_w31161_
	);
	LUT4 #(
		.INIT('h7500)
	) name25335 (
		_w31136_,
		_w31152_,
		_w31156_,
		_w31161_,
		_w31162_
	);
	LUT3 #(
		.INIT('h65)
	) name25336 (
		\u0_L3_reg[22]/NET0131 ,
		_w31149_,
		_w31162_,
		_w31163_
	);
	LUT4 #(
		.INIT('hc693)
	) name25337 (
		decrypt_pad,
		\u0_R3_reg[4]/NET0131 ,
		\u0_uk_K_r3_reg[39]/NET0131 ,
		\u0_uk_K_r3_reg[5]/NET0131 ,
		_w31164_
	);
	LUT4 #(
		.INIT('hc963)
	) name25338 (
		decrypt_pad,
		\u0_R3_reg[3]/NET0131 ,
		\u0_uk_K_r3_reg[27]/NET0131 ,
		\u0_uk_K_r3_reg[4]/NET0131 ,
		_w31165_
	);
	LUT4 #(
		.INIT('hc963)
	) name25339 (
		decrypt_pad,
		\u0_R3_reg[32]/NET0131 ,
		\u0_uk_K_r3_reg[39]/NET0131 ,
		\u0_uk_K_r3_reg[48]/NET0131 ,
		_w31166_
	);
	LUT4 #(
		.INIT('hc693)
	) name25340 (
		decrypt_pad,
		\u0_R3_reg[1]/NET0131 ,
		\u0_uk_K_r3_reg[12]/NET0131 ,
		\u0_uk_K_r3_reg[3]/NET0131 ,
		_w31167_
	);
	LUT4 #(
		.INIT('hc693)
	) name25341 (
		decrypt_pad,
		\u0_R3_reg[5]/NET0131 ,
		\u0_uk_K_r3_reg[10]/NET0131 ,
		\u0_uk_K_r3_reg[33]/NET0131 ,
		_w31168_
	);
	LUT4 #(
		.INIT('hc963)
	) name25342 (
		decrypt_pad,
		\u0_R3_reg[2]/NET0131 ,
		\u0_uk_K_r3_reg[18]/NET0131 ,
		\u0_uk_K_r3_reg[27]/NET0131 ,
		_w31169_
	);
	LUT4 #(
		.INIT('h2000)
	) name25343 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31170_
	);
	LUT4 #(
		.INIT('h9fff)
	) name25344 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31171_
	);
	LUT2 #(
		.INIT('h2)
	) name25345 (
		_w31165_,
		_w31171_,
		_w31172_
	);
	LUT4 #(
		.INIT('h0010)
	) name25346 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31173_
	);
	LUT2 #(
		.INIT('h8)
	) name25347 (
		_w31166_,
		_w31168_,
		_w31174_
	);
	LUT2 #(
		.INIT('h4)
	) name25348 (
		_w31169_,
		_w31165_,
		_w31175_
	);
	LUT3 #(
		.INIT('hce)
	) name25349 (
		_w31167_,
		_w31169_,
		_w31165_,
		_w31176_
	);
	LUT3 #(
		.INIT('h51)
	) name25350 (
		_w31173_,
		_w31174_,
		_w31176_,
		_w31177_
	);
	LUT3 #(
		.INIT('h45)
	) name25351 (
		_w31164_,
		_w31172_,
		_w31177_,
		_w31178_
	);
	LUT2 #(
		.INIT('h1)
	) name25352 (
		_w31166_,
		_w31168_,
		_w31179_
	);
	LUT3 #(
		.INIT('h01)
	) name25353 (
		_w31168_,
		_w31167_,
		_w31169_,
		_w31180_
	);
	LUT4 #(
		.INIT('h1511)
	) name25354 (
		_w31166_,
		_w31167_,
		_w31169_,
		_w31165_,
		_w31181_
	);
	LUT3 #(
		.INIT('h54)
	) name25355 (
		_w31179_,
		_w31180_,
		_w31181_,
		_w31182_
	);
	LUT3 #(
		.INIT('h10)
	) name25356 (
		_w31166_,
		_w31168_,
		_w31169_,
		_w31183_
	);
	LUT4 #(
		.INIT('he2f3)
	) name25357 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31184_
	);
	LUT4 #(
		.INIT('h1098)
	) name25358 (
		_w31166_,
		_w31167_,
		_w31169_,
		_w31165_,
		_w31185_
	);
	LUT3 #(
		.INIT('h0d)
	) name25359 (
		_w31165_,
		_w31184_,
		_w31185_,
		_w31186_
	);
	LUT3 #(
		.INIT('hb0)
	) name25360 (
		_w31182_,
		_w31186_,
		_w31164_,
		_w31187_
	);
	LUT4 #(
		.INIT('h0400)
	) name25361 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31188_
	);
	LUT4 #(
		.INIT('h7bcf)
	) name25362 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31189_
	);
	LUT2 #(
		.INIT('h1)
	) name25363 (
		_w31165_,
		_w31189_,
		_w31190_
	);
	LUT3 #(
		.INIT('hd0)
	) name25364 (
		_w31166_,
		_w31167_,
		_w31169_,
		_w31191_
	);
	LUT3 #(
		.INIT('h0d)
	) name25365 (
		_w31166_,
		_w31169_,
		_w31165_,
		_w31192_
	);
	LUT3 #(
		.INIT('h0d)
	) name25366 (
		_w31168_,
		_w31167_,
		_w31164_,
		_w31193_
	);
	LUT3 #(
		.INIT('h20)
	) name25367 (
		_w31192_,
		_w31191_,
		_w31193_,
		_w31194_
	);
	LUT4 #(
		.INIT('h0200)
	) name25368 (
		_w31166_,
		_w31167_,
		_w31169_,
		_w31165_,
		_w31195_
	);
	LUT2 #(
		.INIT('h4)
	) name25369 (
		_w31166_,
		_w31165_,
		_w31196_
	);
	LUT3 #(
		.INIT('h10)
	) name25370 (
		_w31168_,
		_w31167_,
		_w31169_,
		_w31197_
	);
	LUT3 #(
		.INIT('h15)
	) name25371 (
		_w31195_,
		_w31196_,
		_w31197_,
		_w31198_
	);
	LUT3 #(
		.INIT('h10)
	) name25372 (
		_w31194_,
		_w31190_,
		_w31198_,
		_w31199_
	);
	LUT4 #(
		.INIT('h5655)
	) name25373 (
		\u0_L3_reg[31]/NET0131 ,
		_w31187_,
		_w31178_,
		_w31199_,
		_w31200_
	);
	LUT4 #(
		.INIT('hc963)
	) name25374 (
		decrypt_pad,
		\u0_R3_reg[15]/NET0131 ,
		\u0_uk_K_r3_reg[24]/NET0131 ,
		\u0_uk_K_r3_reg[33]/NET0131 ,
		_w31201_
	);
	LUT4 #(
		.INIT('hc693)
	) name25375 (
		decrypt_pad,
		\u0_R3_reg[13]/NET0131 ,
		\u0_uk_K_r3_reg[24]/NET0131 ,
		\u0_uk_K_r3_reg[47]/NET0131 ,
		_w31202_
	);
	LUT4 #(
		.INIT('hc963)
	) name25376 (
		decrypt_pad,
		\u0_R3_reg[12]/NET0131 ,
		\u0_uk_K_r3_reg[53]/NET0131 ,
		\u0_uk_K_r3_reg[5]/NET0131 ,
		_w31203_
	);
	LUT4 #(
		.INIT('hc693)
	) name25377 (
		decrypt_pad,
		\u0_R3_reg[14]/NET0131 ,
		\u0_uk_K_r3_reg[25]/NET0131 ,
		\u0_uk_K_r3_reg[48]/NET0131 ,
		_w31204_
	);
	LUT4 #(
		.INIT('hc963)
	) name25378 (
		decrypt_pad,
		\u0_R3_reg[17]/NET0131 ,
		\u0_uk_K_r3_reg[12]/NET0131 ,
		\u0_uk_K_r3_reg[46]/NET0131 ,
		_w31205_
	);
	LUT4 #(
		.INIT('h0200)
	) name25379 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31206_
	);
	LUT2 #(
		.INIT('h1)
	) name25380 (
		_w31201_,
		_w31206_,
		_w31207_
	);
	LUT4 #(
		.INIT('h0001)
	) name25381 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31208_
	);
	LUT4 #(
		.INIT('h0040)
	) name25382 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31209_
	);
	LUT4 #(
		.INIT('h0008)
	) name25383 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31210_
	);
	LUT4 #(
		.INIT('h0002)
	) name25384 (
		_w31201_,
		_w31209_,
		_w31210_,
		_w31208_,
		_w31211_
	);
	LUT2 #(
		.INIT('h1)
	) name25385 (
		_w31207_,
		_w31211_,
		_w31212_
	);
	LUT4 #(
		.INIT('h0200)
	) name25386 (
		_w31201_,
		_w31202_,
		_w31203_,
		_w31205_,
		_w31213_
	);
	LUT4 #(
		.INIT('hc963)
	) name25387 (
		decrypt_pad,
		\u0_R3_reg[16]/NET0131 ,
		\u0_uk_K_r3_reg[32]/NET0131 ,
		\u0_uk_K_r3_reg[41]/NET0131 ,
		_w31214_
	);
	LUT4 #(
		.INIT('h0080)
	) name25388 (
		_w31201_,
		_w31202_,
		_w31203_,
		_w31205_,
		_w31215_
	);
	LUT2 #(
		.INIT('h4)
	) name25389 (
		_w31202_,
		_w31203_,
		_w31216_
	);
	LUT4 #(
		.INIT('h0014)
	) name25390 (
		_w31201_,
		_w31202_,
		_w31203_,
		_w31204_,
		_w31217_
	);
	LUT4 #(
		.INIT('h0004)
	) name25391 (
		_w31213_,
		_w31214_,
		_w31215_,
		_w31217_,
		_w31218_
	);
	LUT4 #(
		.INIT('h7dff)
	) name25392 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31219_
	);
	LUT4 #(
		.INIT('h0001)
	) name25393 (
		_w31201_,
		_w31202_,
		_w31203_,
		_w31205_,
		_w31220_
	);
	LUT3 #(
		.INIT('h4c)
	) name25394 (
		_w31204_,
		_w31219_,
		_w31220_,
		_w31221_
	);
	LUT4 #(
		.INIT('h2aa8)
	) name25395 (
		_w31201_,
		_w31202_,
		_w31203_,
		_w31205_,
		_w31222_
	);
	LUT3 #(
		.INIT('h08)
	) name25396 (
		_w31203_,
		_w31204_,
		_w31205_,
		_w31223_
	);
	LUT3 #(
		.INIT('h45)
	) name25397 (
		_w31201_,
		_w31202_,
		_w31205_,
		_w31224_
	);
	LUT3 #(
		.INIT('h45)
	) name25398 (
		_w31222_,
		_w31223_,
		_w31224_,
		_w31225_
	);
	LUT4 #(
		.INIT('hffde)
	) name25399 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31226_
	);
	LUT2 #(
		.INIT('h8)
	) name25400 (
		_w31201_,
		_w31204_,
		_w31227_
	);
	LUT4 #(
		.INIT('h0800)
	) name25401 (
		_w31201_,
		_w31202_,
		_w31203_,
		_w31204_,
		_w31228_
	);
	LUT4 #(
		.INIT('h0400)
	) name25402 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31229_
	);
	LUT4 #(
		.INIT('h0004)
	) name25403 (
		_w31214_,
		_w31226_,
		_w31229_,
		_w31228_,
		_w31230_
	);
	LUT4 #(
		.INIT('h7077)
	) name25404 (
		_w31218_,
		_w31221_,
		_w31225_,
		_w31230_,
		_w31231_
	);
	LUT3 #(
		.INIT('h56)
	) name25405 (
		\u0_L3_reg[20]/NET0131 ,
		_w31212_,
		_w31231_,
		_w31232_
	);
	LUT4 #(
		.INIT('hc963)
	) name25406 (
		decrypt_pad,
		\u0_R3_reg[32]/NET0131 ,
		\u0_uk_K_r3_reg[1]/NET0131 ,
		\u0_uk_K_r3_reg[37]/NET0131 ,
		_w31233_
	);
	LUT4 #(
		.INIT('hc693)
	) name25407 (
		decrypt_pad,
		\u0_R3_reg[28]/NET0131 ,
		\u0_uk_K_r3_reg[15]/NET0131 ,
		\u0_uk_K_r3_reg[38]/NET0131 ,
		_w31234_
	);
	LUT4 #(
		.INIT('hc963)
	) name25408 (
		decrypt_pad,
		\u0_R3_reg[1]/NET0131 ,
		\u0_uk_K_r3_reg[22]/NET0131 ,
		\u0_uk_K_r3_reg[31]/NET0131 ,
		_w31235_
	);
	LUT4 #(
		.INIT('hc693)
	) name25409 (
		decrypt_pad,
		\u0_R3_reg[30]/NET0131 ,
		\u0_uk_K_r3_reg[43]/NET0131 ,
		\u0_uk_K_r3_reg[7]/NET0131 ,
		_w31236_
	);
	LUT4 #(
		.INIT('hc963)
	) name25410 (
		decrypt_pad,
		\u0_R3_reg[29]/NET0131 ,
		\u0_uk_K_r3_reg[37]/NET0131 ,
		\u0_uk_K_r3_reg[42]/NET0131 ,
		_w31237_
	);
	LUT4 #(
		.INIT('hc693)
	) name25411 (
		decrypt_pad,
		\u0_R3_reg[31]/P0001 ,
		\u0_uk_K_r3_reg[0]/NET0131 ,
		\u0_uk_K_r3_reg[50]/NET0131 ,
		_w31238_
	);
	LUT2 #(
		.INIT('h1)
	) name25412 (
		_w31236_,
		_w31238_,
		_w31239_
	);
	LUT4 #(
		.INIT('h72ba)
	) name25413 (
		_w31236_,
		_w31237_,
		_w31238_,
		_w31235_,
		_w31240_
	);
	LUT2 #(
		.INIT('h2)
	) name25414 (
		_w31234_,
		_w31240_,
		_w31241_
	);
	LUT4 #(
		.INIT('h0008)
	) name25415 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31242_
	);
	LUT4 #(
		.INIT('he0f0)
	) name25416 (
		_w31234_,
		_w31237_,
		_w31238_,
		_w31235_,
		_w31243_
	);
	LUT3 #(
		.INIT('h04)
	) name25417 (
		_w31234_,
		_w31236_,
		_w31235_,
		_w31244_
	);
	LUT3 #(
		.INIT('h13)
	) name25418 (
		_w31237_,
		_w31238_,
		_w31235_,
		_w31245_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name25419 (
		_w31242_,
		_w31243_,
		_w31244_,
		_w31245_,
		_w31246_
	);
	LUT3 #(
		.INIT('h54)
	) name25420 (
		_w31233_,
		_w31241_,
		_w31246_,
		_w31247_
	);
	LUT4 #(
		.INIT('h0009)
	) name25421 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31238_,
		_w31248_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name25422 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31249_
	);
	LUT4 #(
		.INIT('h4000)
	) name25423 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31250_
	);
	LUT3 #(
		.INIT('h20)
	) name25424 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31251_
	);
	LUT4 #(
		.INIT('h0020)
	) name25425 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31252_
	);
	LUT4 #(
		.INIT('h00f2)
	) name25426 (
		_w31238_,
		_w31249_,
		_w31250_,
		_w31252_,
		_w31253_
	);
	LUT4 #(
		.INIT('h0040)
	) name25427 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31254_
	);
	LUT3 #(
		.INIT('h10)
	) name25428 (
		_w31236_,
		_w31237_,
		_w31235_,
		_w31255_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name25429 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31256_
	);
	LUT4 #(
		.INIT('h0400)
	) name25430 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31257_
	);
	LUT4 #(
		.INIT('hf9be)
	) name25431 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31258_
	);
	LUT2 #(
		.INIT('h1)
	) name25432 (
		_w31238_,
		_w31235_,
		_w31259_
	);
	LUT4 #(
		.INIT('hef45)
	) name25433 (
		_w31238_,
		_w31235_,
		_w31251_,
		_w31258_,
		_w31260_
	);
	LUT4 #(
		.INIT('h1f00)
	) name25434 (
		_w31248_,
		_w31253_,
		_w31233_,
		_w31260_,
		_w31261_
	);
	LUT3 #(
		.INIT('h9a)
	) name25435 (
		\u0_L3_reg[5]/NET0131 ,
		_w31247_,
		_w31261_,
		_w31262_
	);
	LUT4 #(
		.INIT('hc963)
	) name25436 (
		decrypt_pad,
		\u0_R3_reg[24]/NET0131 ,
		\u0_uk_K_r3_reg[29]/NET0131 ,
		\u0_uk_K_r3_reg[38]/NET0131 ,
		_w31263_
	);
	LUT4 #(
		.INIT('hc963)
	) name25437 (
		decrypt_pad,
		\u0_R3_reg[22]/NET0131 ,
		\u0_uk_K_r3_reg[14]/NET0131 ,
		\u0_uk_K_r3_reg[50]/NET0131 ,
		_w31264_
	);
	LUT4 #(
		.INIT('hc693)
	) name25438 (
		decrypt_pad,
		\u0_R3_reg[20]/NET0131 ,
		\u0_uk_K_r3_reg[44]/NET0131 ,
		\u0_uk_K_r3_reg[8]/NET0131 ,
		_w31265_
	);
	LUT4 #(
		.INIT('hc963)
	) name25439 (
		decrypt_pad,
		\u0_R3_reg[21]/NET0131 ,
		\u0_uk_K_r3_reg[23]/NET0131 ,
		\u0_uk_K_r3_reg[28]/NET0131 ,
		_w31266_
	);
	LUT4 #(
		.INIT('hc693)
	) name25440 (
		decrypt_pad,
		\u0_R3_reg[25]/NET0131 ,
		\u0_uk_K_r3_reg[29]/NET0131 ,
		\u0_uk_K_r3_reg[52]/NET0131 ,
		_w31267_
	);
	LUT4 #(
		.INIT('ha820)
	) name25441 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31268_
	);
	LUT4 #(
		.INIT('hc963)
	) name25442 (
		decrypt_pad,
		\u0_R3_reg[23]/NET0131 ,
		\u0_uk_K_r3_reg[31]/NET0131 ,
		\u0_uk_K_r3_reg[8]/NET0131 ,
		_w31269_
	);
	LUT4 #(
		.INIT('h4555)
	) name25443 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31270_
	);
	LUT3 #(
		.INIT('h01)
	) name25444 (
		_w31269_,
		_w31270_,
		_w31268_,
		_w31271_
	);
	LUT4 #(
		.INIT('h0040)
	) name25445 (
		_w31264_,
		_w31265_,
		_w31267_,
		_w31269_,
		_w31272_
	);
	LUT2 #(
		.INIT('h2)
	) name25446 (
		_w31266_,
		_w31267_,
		_w31273_
	);
	LUT4 #(
		.INIT('hf700)
	) name25447 (
		_w31265_,
		_w31266_,
		_w31267_,
		_w31269_,
		_w31274_
	);
	LUT4 #(
		.INIT('he0e4)
	) name25448 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31275_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name25449 (
		_w31266_,
		_w31272_,
		_w31274_,
		_w31275_,
		_w31276_
	);
	LUT3 #(
		.INIT('h8a)
	) name25450 (
		_w31263_,
		_w31271_,
		_w31276_,
		_w31277_
	);
	LUT4 #(
		.INIT('heeae)
	) name25451 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31278_
	);
	LUT4 #(
		.INIT('he0ee)
	) name25452 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31279_
	);
	LUT3 #(
		.INIT('h8a)
	) name25453 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31280_
	);
	LUT4 #(
		.INIT('h002e)
	) name25454 (
		_w31279_,
		_w31269_,
		_w31278_,
		_w31280_,
		_w31281_
	);
	LUT3 #(
		.INIT('h07)
	) name25455 (
		_w31265_,
		_w31267_,
		_w31269_,
		_w31282_
	);
	LUT4 #(
		.INIT('h0a08)
	) name25456 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31283_
	);
	LUT2 #(
		.INIT('h4)
	) name25457 (
		_w31282_,
		_w31283_,
		_w31284_
	);
	LUT3 #(
		.INIT('h54)
	) name25458 (
		_w31263_,
		_w31281_,
		_w31284_,
		_w31285_
	);
	LUT4 #(
		.INIT('h1000)
	) name25459 (
		_w31265_,
		_w31266_,
		_w31267_,
		_w31269_,
		_w31286_
	);
	LUT4 #(
		.INIT('heff7)
	) name25460 (
		_w31265_,
		_w31266_,
		_w31267_,
		_w31269_,
		_w31287_
	);
	LUT2 #(
		.INIT('h1)
	) name25461 (
		_w31264_,
		_w31287_,
		_w31288_
	);
	LUT4 #(
		.INIT('h0001)
	) name25462 (
		_w31264_,
		_w31265_,
		_w31267_,
		_w31269_,
		_w31289_
	);
	LUT4 #(
		.INIT('h0010)
	) name25463 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31290_
	);
	LUT4 #(
		.INIT('h77ef)
	) name25464 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31291_
	);
	LUT4 #(
		.INIT('haf23)
	) name25465 (
		_w31266_,
		_w31269_,
		_w31289_,
		_w31291_,
		_w31292_
	);
	LUT2 #(
		.INIT('h4)
	) name25466 (
		_w31288_,
		_w31292_,
		_w31293_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name25467 (
		\u0_L3_reg[11]/NET0131 ,
		_w31285_,
		_w31277_,
		_w31293_,
		_w31294_
	);
	LUT4 #(
		.INIT('h0100)
	) name25468 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31238_,
		_w31295_
	);
	LUT2 #(
		.INIT('h1)
	) name25469 (
		_w31233_,
		_w31295_,
		_w31296_
	);
	LUT4 #(
		.INIT('hd080)
	) name25470 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31297_
	);
	LUT4 #(
		.INIT('hfe00)
	) name25471 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31238_,
		_w31298_
	);
	LUT3 #(
		.INIT('h10)
	) name25472 (
		_w31255_,
		_w31297_,
		_w31298_,
		_w31299_
	);
	LUT4 #(
		.INIT('h0800)
	) name25473 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31300_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name25474 (
		_w31234_,
		_w31236_,
		_w31238_,
		_w31235_,
		_w31301_
	);
	LUT2 #(
		.INIT('h4)
	) name25475 (
		_w31300_,
		_w31301_,
		_w31302_
	);
	LUT4 #(
		.INIT('hfe7b)
	) name25476 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31303_
	);
	LUT4 #(
		.INIT('h0155)
	) name25477 (
		_w31296_,
		_w31299_,
		_w31302_,
		_w31303_,
		_w31304_
	);
	LUT3 #(
		.INIT('h80)
	) name25478 (
		_w31234_,
		_w31237_,
		_w31235_,
		_w31305_
	);
	LUT2 #(
		.INIT('h8)
	) name25479 (
		_w31239_,
		_w31305_,
		_w31306_
	);
	LUT2 #(
		.INIT('h4)
	) name25480 (
		_w31237_,
		_w31238_,
		_w31307_
	);
	LUT4 #(
		.INIT('h4440)
	) name25481 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31308_
	);
	LUT4 #(
		.INIT('h0004)
	) name25482 (
		_w31234_,
		_w31237_,
		_w31238_,
		_w31235_,
		_w31309_
	);
	LUT3 #(
		.INIT('h20)
	) name25483 (
		_w31234_,
		_w31236_,
		_w31235_,
		_w31310_
	);
	LUT4 #(
		.INIT('h5554)
	) name25484 (
		_w31307_,
		_w31309_,
		_w31308_,
		_w31310_,
		_w31311_
	);
	LUT4 #(
		.INIT('hf757)
	) name25485 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31312_
	);
	LUT4 #(
		.INIT('hfff6)
	) name25486 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31313_
	);
	LUT3 #(
		.INIT('hd0)
	) name25487 (
		_w31238_,
		_w31312_,
		_w31313_,
		_w31314_
	);
	LUT4 #(
		.INIT('h2322)
	) name25488 (
		_w31233_,
		_w31306_,
		_w31311_,
		_w31314_,
		_w31315_
	);
	LUT3 #(
		.INIT('h65)
	) name25489 (
		\u0_L3_reg[21]/NET0131 ,
		_w31304_,
		_w31315_,
		_w31316_
	);
	LUT4 #(
		.INIT('hc693)
	) name25490 (
		decrypt_pad,
		\u0_R3_reg[20]/NET0131 ,
		\u0_uk_K_r3_reg[22]/NET0131 ,
		\u0_uk_K_r3_reg[45]/P0001 ,
		_w31317_
	);
	LUT4 #(
		.INIT('hc963)
	) name25491 (
		decrypt_pad,
		\u0_R3_reg[19]/NET0131 ,
		\u0_uk_K_r3_reg[2]/NET0131 ,
		\u0_uk_K_r3_reg[7]/NET0131 ,
		_w31318_
	);
	LUT4 #(
		.INIT('hc963)
	) name25492 (
		decrypt_pad,
		\u0_R3_reg[17]/NET0131 ,
		\u0_uk_K_r3_reg[21]/NET0131 ,
		\u0_uk_K_r3_reg[2]/NET0131 ,
		_w31319_
	);
	LUT4 #(
		.INIT('hc963)
	) name25493 (
		decrypt_pad,
		\u0_R3_reg[16]/NET0131 ,
		\u0_uk_K_r3_reg[30]/NET0131 ,
		\u0_uk_K_r3_reg[35]/NET0131 ,
		_w31320_
	);
	LUT4 #(
		.INIT('hc693)
	) name25494 (
		decrypt_pad,
		\u0_R3_reg[21]/NET0131 ,
		\u0_uk_K_r3_reg[23]/NET0131 ,
		\u0_uk_K_r3_reg[42]/NET0131 ,
		_w31321_
	);
	LUT4 #(
		.INIT('hc963)
	) name25495 (
		decrypt_pad,
		\u0_R3_reg[18]/NET0131 ,
		\u0_uk_K_r3_reg[15]/NET0131 ,
		\u0_uk_K_r3_reg[51]/NET0131 ,
		_w31322_
	);
	LUT4 #(
		.INIT('hc25f)
	) name25496 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31323_
	);
	LUT2 #(
		.INIT('h2)
	) name25497 (
		_w31318_,
		_w31323_,
		_w31324_
	);
	LUT3 #(
		.INIT('hde)
	) name25498 (
		_w31319_,
		_w31320_,
		_w31321_,
		_w31325_
	);
	LUT2 #(
		.INIT('h1)
	) name25499 (
		_w31322_,
		_w31318_,
		_w31326_
	);
	LUT2 #(
		.INIT('h4)
	) name25500 (
		_w31325_,
		_w31326_,
		_w31327_
	);
	LUT2 #(
		.INIT('h8)
	) name25501 (
		_w31320_,
		_w31321_,
		_w31328_
	);
	LUT3 #(
		.INIT('he6)
	) name25502 (
		_w31319_,
		_w31322_,
		_w31318_,
		_w31329_
	);
	LUT4 #(
		.INIT('h0020)
	) name25503 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31330_
	);
	LUT4 #(
		.INIT('h0040)
	) name25504 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31331_
	);
	LUT4 #(
		.INIT('hff9f)
	) name25505 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31332_
	);
	LUT3 #(
		.INIT('hd0)
	) name25506 (
		_w31328_,
		_w31329_,
		_w31332_,
		_w31333_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name25507 (
		_w31317_,
		_w31324_,
		_w31327_,
		_w31333_,
		_w31334_
	);
	LUT4 #(
		.INIT('h0010)
	) name25508 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31335_
	);
	LUT3 #(
		.INIT('h08)
	) name25509 (
		_w31319_,
		_w31322_,
		_w31321_,
		_w31336_
	);
	LUT4 #(
		.INIT('hda67)
	) name25510 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31337_
	);
	LUT4 #(
		.INIT('h3df8)
	) name25511 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31338_
	);
	LUT3 #(
		.INIT('h40)
	) name25512 (
		_w31319_,
		_w31320_,
		_w31321_,
		_w31339_
	);
	LUT4 #(
		.INIT('h4000)
	) name25513 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31340_
	);
	LUT4 #(
		.INIT('hbffd)
	) name25514 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31341_
	);
	LUT4 #(
		.INIT('he400)
	) name25515 (
		_w31318_,
		_w31337_,
		_w31338_,
		_w31341_,
		_w31342_
	);
	LUT4 #(
		.INIT('hffdb)
	) name25516 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31343_
	);
	LUT4 #(
		.INIT('h0400)
	) name25517 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31344_
	);
	LUT4 #(
		.INIT('hfbf7)
	) name25518 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31345_
	);
	LUT3 #(
		.INIT('hd8)
	) name25519 (
		_w31318_,
		_w31343_,
		_w31345_,
		_w31346_
	);
	LUT3 #(
		.INIT('he0)
	) name25520 (
		_w31317_,
		_w31342_,
		_w31346_,
		_w31347_
	);
	LUT3 #(
		.INIT('h65)
	) name25521 (
		\u0_L3_reg[14]/NET0131 ,
		_w31334_,
		_w31347_,
		_w31348_
	);
	LUT4 #(
		.INIT('hc693)
	) name25522 (
		decrypt_pad,
		\u0_R3_reg[8]/NET0131 ,
		\u0_uk_K_r3_reg[40]/NET0131 ,
		\u0_uk_K_r3_reg[6]/NET0131 ,
		_w31349_
	);
	LUT4 #(
		.INIT('hc963)
	) name25523 (
		decrypt_pad,
		\u0_R3_reg[6]/NET0131 ,
		\u0_uk_K_r3_reg[46]/NET0131 ,
		\u0_uk_K_r3_reg[55]/NET0131 ,
		_w31350_
	);
	LUT4 #(
		.INIT('hc963)
	) name25524 (
		decrypt_pad,
		\u0_R3_reg[9]/NET0131 ,
		\u0_uk_K_r3_reg[11]/NET0131 ,
		\u0_uk_K_r3_reg[20]/NET0131 ,
		_w31351_
	);
	LUT4 #(
		.INIT('hc693)
	) name25525 (
		decrypt_pad,
		\u0_R3_reg[5]/NET0131 ,
		\u0_uk_K_r3_reg[32]/NET0131 ,
		\u0_uk_K_r3_reg[55]/NET0131 ,
		_w31352_
	);
	LUT4 #(
		.INIT('hc693)
	) name25526 (
		decrypt_pad,
		\u0_R3_reg[7]/NET0131 ,
		\u0_uk_K_r3_reg[17]/NET0131 ,
		\u0_uk_K_r3_reg[40]/NET0131 ,
		_w31353_
	);
	LUT4 #(
		.INIT('h0004)
	) name25527 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31353_,
		_w31354_
	);
	LUT4 #(
		.INIT('hc963)
	) name25528 (
		decrypt_pad,
		\u0_R3_reg[4]/NET0131 ,
		\u0_uk_K_r3_reg[19]/NET0131 ,
		\u0_uk_K_r3_reg[53]/NET0131 ,
		_w31355_
	);
	LUT2 #(
		.INIT('h2)
	) name25529 (
		_w31351_,
		_w31355_,
		_w31356_
	);
	LUT3 #(
		.INIT('h08)
	) name25530 (
		_w31351_,
		_w31352_,
		_w31355_,
		_w31357_
	);
	LUT4 #(
		.INIT('h0080)
	) name25531 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31358_
	);
	LUT2 #(
		.INIT('h1)
	) name25532 (
		_w31354_,
		_w31358_,
		_w31359_
	);
	LUT4 #(
		.INIT('h0800)
	) name25533 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31360_
	);
	LUT4 #(
		.INIT('h0103)
	) name25534 (
		_w31353_,
		_w31354_,
		_w31358_,
		_w31360_,
		_w31361_
	);
	LUT2 #(
		.INIT('h8)
	) name25535 (
		_w31351_,
		_w31355_,
		_w31362_
	);
	LUT4 #(
		.INIT('h1014)
	) name25536 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31363_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name25537 (
		_w31351_,
		_w31352_,
		_w31353_,
		_w31355_,
		_w31364_
	);
	LUT4 #(
		.INIT('h51f3)
	) name25538 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31365_
	);
	LUT3 #(
		.INIT('h51)
	) name25539 (
		_w31363_,
		_w31364_,
		_w31365_,
		_w31366_
	);
	LUT3 #(
		.INIT('h15)
	) name25540 (
		_w31349_,
		_w31361_,
		_w31366_,
		_w31367_
	);
	LUT4 #(
		.INIT('hf7cc)
	) name25541 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31368_
	);
	LUT4 #(
		.INIT('h00c4)
	) name25542 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31369_
	);
	LUT3 #(
		.INIT('h0b)
	) name25543 (
		_w31350_,
		_w31352_,
		_w31353_,
		_w31370_
	);
	LUT4 #(
		.INIT('hf200)
	) name25544 (
		_w31349_,
		_w31368_,
		_w31369_,
		_w31370_,
		_w31371_
	);
	LUT4 #(
		.INIT('h0002)
	) name25545 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31372_
	);
	LUT4 #(
		.INIT('haffd)
	) name25546 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31373_
	);
	LUT2 #(
		.INIT('h2)
	) name25547 (
		_w31353_,
		_w31373_,
		_w31374_
	);
	LUT4 #(
		.INIT('h0100)
	) name25548 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31375_
	);
	LUT4 #(
		.INIT('hc040)
	) name25549 (
		_w31350_,
		_w31352_,
		_w31353_,
		_w31355_,
		_w31376_
	);
	LUT4 #(
		.INIT('h4000)
	) name25550 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31377_
	);
	LUT4 #(
		.INIT('haaa8)
	) name25551 (
		_w31349_,
		_w31375_,
		_w31376_,
		_w31377_,
		_w31378_
	);
	LUT3 #(
		.INIT('h01)
	) name25552 (
		_w31374_,
		_w31378_,
		_w31371_,
		_w31379_
	);
	LUT3 #(
		.INIT('h65)
	) name25553 (
		\u0_L3_reg[2]/NET0131 ,
		_w31367_,
		_w31379_,
		_w31380_
	);
	LUT4 #(
		.INIT('h0200)
	) name25554 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31381_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name25555 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31382_
	);
	LUT2 #(
		.INIT('h1)
	) name25556 (
		_w31269_,
		_w31382_,
		_w31383_
	);
	LUT4 #(
		.INIT('he63f)
	) name25557 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31384_
	);
	LUT4 #(
		.INIT('h0004)
	) name25558 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31385_
	);
	LUT4 #(
		.INIT('h0031)
	) name25559 (
		_w31269_,
		_w31272_,
		_w31384_,
		_w31385_,
		_w31386_
	);
	LUT3 #(
		.INIT('h45)
	) name25560 (
		_w31263_,
		_w31383_,
		_w31386_,
		_w31387_
	);
	LUT2 #(
		.INIT('h1)
	) name25561 (
		_w31269_,
		_w31278_,
		_w31388_
	);
	LUT3 #(
		.INIT('h80)
	) name25562 (
		_w31264_,
		_w31266_,
		_w31267_,
		_w31389_
	);
	LUT4 #(
		.INIT('h4000)
	) name25563 (
		_w31264_,
		_w31265_,
		_w31267_,
		_w31269_,
		_w31390_
	);
	LUT3 #(
		.INIT('h01)
	) name25564 (
		_w31290_,
		_w31390_,
		_w31389_,
		_w31391_
	);
	LUT4 #(
		.INIT('h007d)
	) name25565 (
		_w31265_,
		_w31266_,
		_w31267_,
		_w31269_,
		_w31392_
	);
	LUT4 #(
		.INIT('hb600)
	) name25566 (
		_w31265_,
		_w31266_,
		_w31267_,
		_w31269_,
		_w31393_
	);
	LUT4 #(
		.INIT('h3331)
	) name25567 (
		_w31264_,
		_w31289_,
		_w31393_,
		_w31392_,
		_w31394_
	);
	LUT4 #(
		.INIT('h7500)
	) name25568 (
		_w31263_,
		_w31388_,
		_w31391_,
		_w31394_,
		_w31395_
	);
	LUT3 #(
		.INIT('h65)
	) name25569 (
		\u0_L3_reg[4]/NET0131 ,
		_w31387_,
		_w31395_,
		_w31396_
	);
	LUT4 #(
		.INIT('hefaa)
	) name25570 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31397_
	);
	LUT2 #(
		.INIT('h1)
	) name25571 (
		_w31201_,
		_w31397_,
		_w31398_
	);
	LUT3 #(
		.INIT('h8a)
	) name25572 (
		_w31202_,
		_w31203_,
		_w31205_,
		_w31399_
	);
	LUT4 #(
		.INIT('hf9fb)
	) name25573 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31400_
	);
	LUT4 #(
		.INIT('h1500)
	) name25574 (
		_w31215_,
		_w31227_,
		_w31399_,
		_w31400_,
		_w31401_
	);
	LUT3 #(
		.INIT('h45)
	) name25575 (
		_w31214_,
		_w31398_,
		_w31401_,
		_w31402_
	);
	LUT4 #(
		.INIT('hcfee)
	) name25576 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31403_
	);
	LUT3 #(
		.INIT('h01)
	) name25577 (
		_w31203_,
		_w31204_,
		_w31205_,
		_w31404_
	);
	LUT4 #(
		.INIT('h0002)
	) name25578 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31405_
	);
	LUT3 #(
		.INIT('h0d)
	) name25579 (
		_w31201_,
		_w31403_,
		_w31405_,
		_w31406_
	);
	LUT4 #(
		.INIT('h2080)
	) name25580 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31407_
	);
	LUT4 #(
		.INIT('h32ff)
	) name25581 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31408_
	);
	LUT3 #(
		.INIT('h51)
	) name25582 (
		_w31201_,
		_w31203_,
		_w31204_,
		_w31409_
	);
	LUT3 #(
		.INIT('h45)
	) name25583 (
		_w31407_,
		_w31408_,
		_w31409_,
		_w31410_
	);
	LUT4 #(
		.INIT('h1541)
	) name25584 (
		_w31201_,
		_w31202_,
		_w31203_,
		_w31205_,
		_w31411_
	);
	LUT4 #(
		.INIT('h82aa)
	) name25585 (
		_w31201_,
		_w31202_,
		_w31203_,
		_w31205_,
		_w31412_
	);
	LUT3 #(
		.INIT('h01)
	) name25586 (
		_w31204_,
		_w31412_,
		_w31411_,
		_w31413_
	);
	LUT4 #(
		.INIT('h00d5)
	) name25587 (
		_w31214_,
		_w31406_,
		_w31410_,
		_w31413_,
		_w31414_
	);
	LUT3 #(
		.INIT('h65)
	) name25588 (
		\u0_L3_reg[26]/NET0131 ,
		_w31402_,
		_w31414_,
		_w31415_
	);
	LUT4 #(
		.INIT('h0002)
	) name25589 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31416_
	);
	LUT4 #(
		.INIT('h5a4f)
	) name25590 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31417_
	);
	LUT4 #(
		.INIT('h3032)
	) name25591 (
		_w31238_,
		_w31233_,
		_w31416_,
		_w31417_,
		_w31418_
	);
	LUT4 #(
		.INIT('hdf9f)
	) name25592 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31419_
	);
	LUT4 #(
		.INIT('h0200)
	) name25593 (
		_w31236_,
		_w31237_,
		_w31238_,
		_w31235_,
		_w31420_
	);
	LUT4 #(
		.INIT('h0010)
	) name25594 (
		_w31234_,
		_w31237_,
		_w31238_,
		_w31235_,
		_w31421_
	);
	LUT4 #(
		.INIT('h0100)
	) name25595 (
		_w31300_,
		_w31420_,
		_w31421_,
		_w31419_,
		_w31422_
	);
	LUT4 #(
		.INIT('hbeff)
	) name25596 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31423_
	);
	LUT2 #(
		.INIT('h2)
	) name25597 (
		_w31238_,
		_w31423_,
		_w31424_
	);
	LUT4 #(
		.INIT('h1001)
	) name25598 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31425_
	);
	LUT4 #(
		.INIT('h080a)
	) name25599 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31233_,
		_w31426_
	);
	LUT4 #(
		.INIT('h5554)
	) name25600 (
		_w31238_,
		_w31254_,
		_w31426_,
		_w31425_,
		_w31427_
	);
	LUT4 #(
		.INIT('h0031)
	) name25601 (
		_w31233_,
		_w31424_,
		_w31422_,
		_w31427_,
		_w31428_
	);
	LUT3 #(
		.INIT('h65)
	) name25602 (
		\u0_L3_reg[15]/P0001 ,
		_w31418_,
		_w31428_,
		_w31429_
	);
	LUT4 #(
		.INIT('h440c)
	) name25603 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31430_
	);
	LUT4 #(
		.INIT('hfda8)
	) name25604 (
		_w31201_,
		_w31209_,
		_w31404_,
		_w31430_,
		_w31431_
	);
	LUT4 #(
		.INIT('h7df7)
	) name25605 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31432_
	);
	LUT3 #(
		.INIT('h45)
	) name25606 (
		_w31214_,
		_w31431_,
		_w31432_,
		_w31433_
	);
	LUT4 #(
		.INIT('hd5fd)
	) name25607 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31434_
	);
	LUT4 #(
		.INIT('h0080)
	) name25608 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31435_
	);
	LUT4 #(
		.INIT('hef6f)
	) name25609 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31436_
	);
	LUT4 #(
		.INIT('h04cc)
	) name25610 (
		_w31201_,
		_w31214_,
		_w31434_,
		_w31436_,
		_w31437_
	);
	LUT4 #(
		.INIT('h6fff)
	) name25611 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31438_
	);
	LUT4 #(
		.INIT('h6fdf)
	) name25612 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31439_
	);
	LUT2 #(
		.INIT('h2)
	) name25613 (
		_w31201_,
		_w31439_,
		_w31440_
	);
	LUT2 #(
		.INIT('h4)
	) name25614 (
		_w31201_,
		_w31435_,
		_w31441_
	);
	LUT4 #(
		.INIT('haafb)
	) name25615 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31442_
	);
	LUT2 #(
		.INIT('h8)
	) name25616 (
		_w31201_,
		_w31214_,
		_w31443_
	);
	LUT4 #(
		.INIT('h7077)
	) name25617 (
		_w31204_,
		_w31220_,
		_w31442_,
		_w31443_,
		_w31444_
	);
	LUT4 #(
		.INIT('h0100)
	) name25618 (
		_w31440_,
		_w31441_,
		_w31437_,
		_w31444_,
		_w31445_
	);
	LUT3 #(
		.INIT('h65)
	) name25619 (
		\u0_L3_reg[1]/NET0131 ,
		_w31433_,
		_w31445_,
		_w31446_
	);
	LUT4 #(
		.INIT('hff2e)
	) name25620 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31447_
	);
	LUT3 #(
		.INIT('h02)
	) name25621 (
		_w31350_,
		_w31352_,
		_w31355_,
		_w31448_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name25622 (
		_w31350_,
		_w31352_,
		_w31353_,
		_w31355_,
		_w31449_
	);
	LUT4 #(
		.INIT('h0ef3)
	) name25623 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31450_
	);
	LUT4 #(
		.INIT('h7277)
	) name25624 (
		_w31353_,
		_w31447_,
		_w31448_,
		_w31450_,
		_w31451_
	);
	LUT4 #(
		.INIT('h0802)
	) name25625 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31452_
	);
	LUT4 #(
		.INIT('h2000)
	) name25626 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31453_
	);
	LUT3 #(
		.INIT('h01)
	) name25627 (
		_w31349_,
		_w31453_,
		_w31452_,
		_w31454_
	);
	LUT2 #(
		.INIT('h4)
	) name25628 (
		_w31451_,
		_w31454_,
		_w31455_
	);
	LUT3 #(
		.INIT('h90)
	) name25629 (
		_w31351_,
		_w31352_,
		_w31355_,
		_w31456_
	);
	LUT4 #(
		.INIT('h0020)
	) name25630 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31457_
	);
	LUT3 #(
		.INIT('h02)
	) name25631 (
		_w31353_,
		_w31457_,
		_w31456_,
		_w31458_
	);
	LUT4 #(
		.INIT('hdf2e)
	) name25632 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31459_
	);
	LUT2 #(
		.INIT('h8)
	) name25633 (
		_w31449_,
		_w31459_,
		_w31460_
	);
	LUT2 #(
		.INIT('h8)
	) name25634 (
		_w31353_,
		_w31355_,
		_w31461_
	);
	LUT4 #(
		.INIT('h0dff)
	) name25635 (
		_w31351_,
		_w31352_,
		_w31353_,
		_w31355_,
		_w31462_
	);
	LUT4 #(
		.INIT('h0008)
	) name25636 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31463_
	);
	LUT4 #(
		.INIT('h00a8)
	) name25637 (
		_w31349_,
		_w31350_,
		_w31462_,
		_w31463_,
		_w31464_
	);
	LUT3 #(
		.INIT('he0)
	) name25638 (
		_w31458_,
		_w31460_,
		_w31464_,
		_w31465_
	);
	LUT3 #(
		.INIT('ha9)
	) name25639 (
		\u0_L3_reg[28]/NET0131 ,
		_w31455_,
		_w31465_,
		_w31466_
	);
	LUT4 #(
		.INIT('h0400)
	) name25640 (
		_w31201_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31467_
	);
	LUT3 #(
		.INIT('h08)
	) name25641 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31468_
	);
	LUT3 #(
		.INIT('h01)
	) name25642 (
		_w31220_,
		_w31467_,
		_w31468_,
		_w31469_
	);
	LUT4 #(
		.INIT('h0200)
	) name25643 (
		_w31201_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31470_
	);
	LUT3 #(
		.INIT('h8a)
	) name25644 (
		_w31201_,
		_w31204_,
		_w31205_,
		_w31471_
	);
	LUT3 #(
		.INIT('h13)
	) name25645 (
		_w31216_,
		_w31470_,
		_w31471_,
		_w31472_
	);
	LUT4 #(
		.INIT('h1555)
	) name25646 (
		_w31214_,
		_w31226_,
		_w31469_,
		_w31472_,
		_w31473_
	);
	LUT4 #(
		.INIT('hfd3b)
	) name25647 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31474_
	);
	LUT4 #(
		.INIT('hfbdd)
	) name25648 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31475_
	);
	LUT4 #(
		.INIT('hc480)
	) name25649 (
		_w31201_,
		_w31438_,
		_w31475_,
		_w31474_,
		_w31476_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name25650 (
		_w31202_,
		_w31203_,
		_w31204_,
		_w31205_,
		_w31477_
	);
	LUT4 #(
		.INIT('h0702)
	) name25651 (
		_w31201_,
		_w31210_,
		_w31228_,
		_w31477_,
		_w31478_
	);
	LUT3 #(
		.INIT('hd0)
	) name25652 (
		_w31214_,
		_w31476_,
		_w31478_,
		_w31479_
	);
	LUT3 #(
		.INIT('h65)
	) name25653 (
		\u0_L3_reg[10]/NET0131 ,
		_w31473_,
		_w31479_,
		_w31480_
	);
	LUT4 #(
		.INIT('h5410)
	) name25654 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31481_
	);
	LUT4 #(
		.INIT('hab6f)
	) name25655 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31482_
	);
	LUT2 #(
		.INIT('h1)
	) name25656 (
		_w31269_,
		_w31482_,
		_w31483_
	);
	LUT4 #(
		.INIT('h3fd2)
	) name25657 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31484_
	);
	LUT4 #(
		.INIT('h0501)
	) name25658 (
		_w31263_,
		_w31269_,
		_w31381_,
		_w31484_,
		_w31485_
	);
	LUT3 #(
		.INIT('h28)
	) name25659 (
		_w31264_,
		_w31265_,
		_w31267_,
		_w31486_
	);
	LUT4 #(
		.INIT('hcd00)
	) name25660 (
		_w31264_,
		_w31266_,
		_w31267_,
		_w31269_,
		_w31487_
	);
	LUT3 #(
		.INIT('h01)
	) name25661 (
		_w31481_,
		_w31487_,
		_w31486_,
		_w31488_
	);
	LUT4 #(
		.INIT('hcf6f)
	) name25662 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31489_
	);
	LUT3 #(
		.INIT('ha2)
	) name25663 (
		_w31263_,
		_w31269_,
		_w31489_,
		_w31490_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name25664 (
		_w31483_,
		_w31485_,
		_w31488_,
		_w31490_,
		_w31491_
	);
	LUT4 #(
		.INIT('h4000)
	) name25665 (
		_w31264_,
		_w31266_,
		_w31267_,
		_w31269_,
		_w31492_
	);
	LUT2 #(
		.INIT('h1)
	) name25666 (
		_w31385_,
		_w31492_,
		_w31493_
	);
	LUT3 #(
		.INIT('h9a)
	) name25667 (
		\u0_L3_reg[29]/NET0131 ,
		_w31491_,
		_w31493_,
		_w31494_
	);
	LUT3 #(
		.INIT('h82)
	) name25668 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31495_
	);
	LUT3 #(
		.INIT('h69)
	) name25669 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31496_
	);
	LUT3 #(
		.INIT('h8a)
	) name25670 (
		_w31166_,
		_w31168_,
		_w31169_,
		_w31497_
	);
	LUT4 #(
		.INIT('h7500)
	) name25671 (
		_w31166_,
		_w31168_,
		_w31169_,
		_w31164_,
		_w31498_
	);
	LUT4 #(
		.INIT('h0020)
	) name25672 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31499_
	);
	LUT4 #(
		.INIT('h7fdb)
	) name25673 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31500_
	);
	LUT4 #(
		.INIT('h1055)
	) name25674 (
		_w31165_,
		_w31496_,
		_w31498_,
		_w31500_,
		_w31501_
	);
	LUT4 #(
		.INIT('h007e)
	) name25675 (
		_w31168_,
		_w31167_,
		_w31169_,
		_w31164_,
		_w31502_
	);
	LUT3 #(
		.INIT('h13)
	) name25676 (
		_w31168_,
		_w31167_,
		_w31169_,
		_w31503_
	);
	LUT3 #(
		.INIT('h1b)
	) name25677 (
		_w31168_,
		_w31167_,
		_w31169_,
		_w31504_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name25678 (
		_w31166_,
		_w31165_,
		_w31503_,
		_w31504_,
		_w31505_
	);
	LUT2 #(
		.INIT('h8)
	) name25679 (
		_w31167_,
		_w31165_,
		_w31506_
	);
	LUT3 #(
		.INIT('h10)
	) name25680 (
		_w31183_,
		_w31497_,
		_w31506_,
		_w31507_
	);
	LUT4 #(
		.INIT('h0008)
	) name25681 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31508_
	);
	LUT4 #(
		.INIT('h002a)
	) name25682 (
		_w31164_,
		_w31196_,
		_w31197_,
		_w31508_,
		_w31509_
	);
	LUT4 #(
		.INIT('h7077)
	) name25683 (
		_w31502_,
		_w31505_,
		_w31507_,
		_w31509_,
		_w31510_
	);
	LUT4 #(
		.INIT('haaa9)
	) name25684 (
		\u0_L3_reg[23]/NET0131 ,
		_w31195_,
		_w31510_,
		_w31501_,
		_w31511_
	);
	LUT4 #(
		.INIT('h0001)
	) name25685 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31512_
	);
	LUT4 #(
		.INIT('haffe)
	) name25686 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31513_
	);
	LUT4 #(
		.INIT('haa8a)
	) name25687 (
		_w31317_,
		_w31322_,
		_w31320_,
		_w31318_,
		_w31514_
	);
	LUT4 #(
		.INIT('hc400)
	) name25688 (
		_w31318_,
		_w31345_,
		_w31513_,
		_w31514_,
		_w31515_
	);
	LUT4 #(
		.INIT('h5fef)
	) name25689 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31516_
	);
	LUT4 #(
		.INIT('h5551)
	) name25690 (
		_w31317_,
		_w31319_,
		_w31322_,
		_w31320_,
		_w31517_
	);
	LUT3 #(
		.INIT('hd0)
	) name25691 (
		_w31318_,
		_w31516_,
		_w31517_,
		_w31518_
	);
	LUT4 #(
		.INIT('ha4ff)
	) name25692 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31519_
	);
	LUT4 #(
		.INIT('hff7b)
	) name25693 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31520_
	);
	LUT3 #(
		.INIT('he0)
	) name25694 (
		_w31318_,
		_w31519_,
		_w31520_,
		_w31521_
	);
	LUT3 #(
		.INIT('h15)
	) name25695 (
		_w31515_,
		_w31518_,
		_w31521_,
		_w31522_
	);
	LUT2 #(
		.INIT('h1)
	) name25696 (
		_w31318_,
		_w31331_,
		_w31523_
	);
	LUT4 #(
		.INIT('h0200)
	) name25697 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31524_
	);
	LUT4 #(
		.INIT('h0002)
	) name25698 (
		_w31318_,
		_w31336_,
		_w31344_,
		_w31524_,
		_w31525_
	);
	LUT2 #(
		.INIT('h1)
	) name25699 (
		_w31523_,
		_w31525_,
		_w31526_
	);
	LUT3 #(
		.INIT('h56)
	) name25700 (
		\u0_L3_reg[8]/NET0131 ,
		_w31522_,
		_w31526_,
		_w31527_
	);
	LUT4 #(
		.INIT('h2146)
	) name25701 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31528_
	);
	LUT3 #(
		.INIT('h01)
	) name25702 (
		_w31139_,
		_w31142_,
		_w31140_,
		_w31529_
	);
	LUT4 #(
		.INIT('hf35f)
	) name25703 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31530_
	);
	LUT4 #(
		.INIT('he4ee)
	) name25704 (
		_w31137_,
		_w31528_,
		_w31529_,
		_w31530_,
		_w31531_
	);
	LUT4 #(
		.INIT('h0080)
	) name25705 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31532_
	);
	LUT3 #(
		.INIT('ha8)
	) name25706 (
		_w31136_,
		_w31531_,
		_w31532_,
		_w31533_
	);
	LUT3 #(
		.INIT('h02)
	) name25707 (
		_w31139_,
		_w31138_,
		_w31140_,
		_w31534_
	);
	LUT4 #(
		.INIT('hddf5)
	) name25708 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31535_
	);
	LUT2 #(
		.INIT('h2)
	) name25709 (
		_w31137_,
		_w31535_,
		_w31536_
	);
	LUT3 #(
		.INIT('h09)
	) name25710 (
		_w31142_,
		_w31140_,
		_w31137_,
		_w31537_
	);
	LUT4 #(
		.INIT('h6fb7)
	) name25711 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31538_
	);
	LUT3 #(
		.INIT('hb0)
	) name25712 (
		_w31534_,
		_w31537_,
		_w31538_,
		_w31539_
	);
	LUT4 #(
		.INIT('hb3bb)
	) name25713 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31540_
	);
	LUT3 #(
		.INIT('h0e)
	) name25714 (
		_w31139_,
		_w31138_,
		_w31137_,
		_w31541_
	);
	LUT4 #(
		.INIT('h7077)
	) name25715 (
		_w31137_,
		_w31157_,
		_w31540_,
		_w31541_,
		_w31542_
	);
	LUT4 #(
		.INIT('hba00)
	) name25716 (
		_w31136_,
		_w31536_,
		_w31539_,
		_w31542_,
		_w31543_
	);
	LUT3 #(
		.INIT('h65)
	) name25717 (
		\u0_L3_reg[32]/NET0131 ,
		_w31533_,
		_w31543_,
		_w31544_
	);
	LUT4 #(
		.INIT('hbf00)
	) name25718 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31269_,
		_w31545_
	);
	LUT3 #(
		.INIT('ha8)
	) name25719 (
		_w31265_,
		_w31389_,
		_w31545_,
		_w31546_
	);
	LUT4 #(
		.INIT('h0041)
	) name25720 (
		_w31265_,
		_w31266_,
		_w31267_,
		_w31269_,
		_w31547_
	);
	LUT3 #(
		.INIT('h07)
	) name25721 (
		_w31273_,
		_w31545_,
		_w31547_,
		_w31548_
	);
	LUT3 #(
		.INIT('h45)
	) name25722 (
		_w31263_,
		_w31546_,
		_w31548_,
		_w31549_
	);
	LUT4 #(
		.INIT('h400c)
	) name25723 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31269_,
		_w31550_
	);
	LUT4 #(
		.INIT('h2002)
	) name25724 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31551_
	);
	LUT4 #(
		.INIT('h0150)
	) name25725 (
		_w31264_,
		_w31265_,
		_w31266_,
		_w31267_,
		_w31552_
	);
	LUT4 #(
		.INIT('h0001)
	) name25726 (
		_w31286_,
		_w31551_,
		_w31550_,
		_w31552_,
		_w31553_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name25727 (
		_w31264_,
		_w31266_,
		_w31287_,
		_w31272_,
		_w31554_
	);
	LUT3 #(
		.INIT('hd0)
	) name25728 (
		_w31263_,
		_w31553_,
		_w31554_,
		_w31555_
	);
	LUT3 #(
		.INIT('h65)
	) name25729 (
		\u0_L3_reg[19]/P0001 ,
		_w31549_,
		_w31555_,
		_w31556_
	);
	LUT4 #(
		.INIT('h0010)
	) name25730 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31557_
	);
	LUT4 #(
		.INIT('h70f0)
	) name25731 (
		_w31234_,
		_w31237_,
		_w31238_,
		_w31235_,
		_w31558_
	);
	LUT3 #(
		.INIT('h48)
	) name25732 (
		_w31234_,
		_w31237_,
		_w31235_,
		_w31559_
	);
	LUT4 #(
		.INIT('h00fe)
	) name25733 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31238_,
		_w31560_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name25734 (
		_w31557_,
		_w31558_,
		_w31559_,
		_w31560_,
		_w31561_
	);
	LUT4 #(
		.INIT('hbcf7)
	) name25735 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31562_
	);
	LUT3 #(
		.INIT('h8a)
	) name25736 (
		_w31233_,
		_w31561_,
		_w31562_,
		_w31563_
	);
	LUT4 #(
		.INIT('hcf40)
	) name25737 (
		_w31234_,
		_w31236_,
		_w31237_,
		_w31235_,
		_w31564_
	);
	LUT4 #(
		.INIT('hf0b0)
	) name25738 (
		_w31236_,
		_w31237_,
		_w31238_,
		_w31235_,
		_w31565_
	);
	LUT2 #(
		.INIT('h4)
	) name25739 (
		_w31564_,
		_w31565_,
		_w31566_
	);
	LUT4 #(
		.INIT('h0800)
	) name25740 (
		_w31234_,
		_w31236_,
		_w31238_,
		_w31235_,
		_w31567_
	);
	LUT3 #(
		.INIT('h01)
	) name25741 (
		_w31257_,
		_w31309_,
		_w31567_,
		_w31568_
	);
	LUT3 #(
		.INIT('h45)
	) name25742 (
		_w31233_,
		_w31566_,
		_w31568_,
		_w31569_
	);
	LUT2 #(
		.INIT('h1)
	) name25743 (
		_w31238_,
		_w31256_,
		_w31570_
	);
	LUT4 #(
		.INIT('h0020)
	) name25744 (
		_w31236_,
		_w31237_,
		_w31238_,
		_w31235_,
		_w31571_
	);
	LUT3 #(
		.INIT('h07)
	) name25745 (
		_w31251_,
		_w31259_,
		_w31571_,
		_w31572_
	);
	LUT2 #(
		.INIT('h4)
	) name25746 (
		_w31570_,
		_w31572_,
		_w31573_
	);
	LUT4 #(
		.INIT('h5655)
	) name25747 (
		\u0_L3_reg[27]/NET0131 ,
		_w31563_,
		_w31569_,
		_w31573_,
		_w31574_
	);
	LUT4 #(
		.INIT('hc963)
	) name25748 (
		decrypt_pad,
		\u0_R3_reg[11]/NET0131 ,
		\u0_uk_K_r3_reg[26]/NET0131 ,
		\u0_uk_K_r3_reg[3]/NET0131 ,
		_w31575_
	);
	LUT4 #(
		.INIT('hc693)
	) name25749 (
		decrypt_pad,
		\u0_R3_reg[12]/NET0131 ,
		\u0_uk_K_r3_reg[18]/NET0131 ,
		\u0_uk_K_r3_reg[41]/NET0131 ,
		_w31576_
	);
	LUT4 #(
		.INIT('hc963)
	) name25750 (
		decrypt_pad,
		\u0_R3_reg[13]/NET0131 ,
		\u0_uk_K_r3_reg[54]/NET0131 ,
		\u0_uk_K_r3_reg[6]/NET0131 ,
		_w31577_
	);
	LUT4 #(
		.INIT('hc963)
	) name25751 (
		decrypt_pad,
		\u0_R3_reg[9]/NET0131 ,
		\u0_uk_K_r3_reg[17]/NET0131 ,
		\u0_uk_K_r3_reg[26]/NET0131 ,
		_w31578_
	);
	LUT4 #(
		.INIT('hc963)
	) name25752 (
		decrypt_pad,
		\u0_R3_reg[10]/NET0131 ,
		\u0_uk_K_r3_reg[25]/NET0131 ,
		\u0_uk_K_r3_reg[34]/NET0131 ,
		_w31579_
	);
	LUT4 #(
		.INIT('hc963)
	) name25753 (
		decrypt_pad,
		\u0_R3_reg[8]/NET0131 ,
		\u0_uk_K_r3_reg[20]/NET0131 ,
		\u0_uk_K_r3_reg[54]/NET0131 ,
		_w31580_
	);
	LUT2 #(
		.INIT('h2)
	) name25754 (
		_w31577_,
		_w31580_,
		_w31581_
	);
	LUT4 #(
		.INIT('h95b5)
	) name25755 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31582_
	);
	LUT4 #(
		.INIT('h0001)
	) name25756 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31583_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name25757 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31584_
	);
	LUT4 #(
		.INIT('h08cc)
	) name25758 (
		_w31576_,
		_w31575_,
		_w31582_,
		_w31584_,
		_w31585_
	);
	LUT2 #(
		.INIT('h1)
	) name25759 (
		_w31578_,
		_w31579_,
		_w31586_
	);
	LUT2 #(
		.INIT('h6)
	) name25760 (
		_w31578_,
		_w31579_,
		_w31587_
	);
	LUT2 #(
		.INIT('h1)
	) name25761 (
		_w31577_,
		_w31580_,
		_w31588_
	);
	LUT2 #(
		.INIT('h8)
	) name25762 (
		_w31577_,
		_w31580_,
		_w31589_
	);
	LUT2 #(
		.INIT('h6)
	) name25763 (
		_w31577_,
		_w31580_,
		_w31590_
	);
	LUT3 #(
		.INIT('h46)
	) name25764 (
		_w31577_,
		_w31580_,
		_w31575_,
		_w31591_
	);
	LUT2 #(
		.INIT('h1)
	) name25765 (
		_w31587_,
		_w31591_,
		_w31592_
	);
	LUT4 #(
		.INIT('h383c)
	) name25766 (
		_w31580_,
		_w31578_,
		_w31579_,
		_w31575_,
		_w31593_
	);
	LUT3 #(
		.INIT('h15)
	) name25767 (
		_w31576_,
		_w31590_,
		_w31593_,
		_w31594_
	);
	LUT3 #(
		.INIT('h80)
	) name25768 (
		_w31578_,
		_w31579_,
		_w31576_,
		_w31595_
	);
	LUT3 #(
		.INIT('h51)
	) name25769 (
		_w31580_,
		_w31578_,
		_w31579_,
		_w31596_
	);
	LUT4 #(
		.INIT('h0090)
	) name25770 (
		_w31577_,
		_w31578_,
		_w31576_,
		_w31575_,
		_w31597_
	);
	LUT4 #(
		.INIT('h7077)
	) name25771 (
		_w31588_,
		_w31595_,
		_w31596_,
		_w31597_,
		_w31598_
	);
	LUT4 #(
		.INIT('h4500)
	) name25772 (
		_w31585_,
		_w31592_,
		_w31594_,
		_w31598_,
		_w31599_
	);
	LUT2 #(
		.INIT('h9)
	) name25773 (
		\u0_L3_reg[6]/NET0131 ,
		_w31599_,
		_w31600_
	);
	LUT4 #(
		.INIT('hba16)
	) name25774 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31601_
	);
	LUT2 #(
		.INIT('h1)
	) name25775 (
		_w31137_,
		_w31601_,
		_w31602_
	);
	LUT4 #(
		.INIT('h6080)
	) name25776 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31603_
	);
	LUT4 #(
		.INIT('h0a04)
	) name25777 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31604_
	);
	LUT4 #(
		.INIT('h020a)
	) name25778 (
		_w31136_,
		_w31137_,
		_w31603_,
		_w31604_,
		_w31605_
	);
	LUT4 #(
		.INIT('h4080)
	) name25779 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31606_
	);
	LUT4 #(
		.INIT('h2a05)
	) name25780 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31607_
	);
	LUT4 #(
		.INIT('h5551)
	) name25781 (
		_w31136_,
		_w31137_,
		_w31607_,
		_w31606_,
		_w31608_
	);
	LUT3 #(
		.INIT('h0b)
	) name25782 (
		_w31602_,
		_w31605_,
		_w31608_,
		_w31609_
	);
	LUT2 #(
		.INIT('h4)
	) name25783 (
		_w31137_,
		_w31603_,
		_w31610_
	);
	LUT2 #(
		.INIT('h2)
	) name25784 (
		_w31136_,
		_w31137_,
		_w31611_
	);
	LUT4 #(
		.INIT('h0010)
	) name25785 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w31612_
	);
	LUT4 #(
		.INIT('h0f04)
	) name25786 (
		_w31137_,
		_w31604_,
		_w31611_,
		_w31612_,
		_w31613_
	);
	LUT2 #(
		.INIT('h1)
	) name25787 (
		_w31610_,
		_w31613_,
		_w31614_
	);
	LUT3 #(
		.INIT('h65)
	) name25788 (
		\u0_L3_reg[7]/NET0131 ,
		_w31609_,
		_w31614_,
		_w31615_
	);
	LUT4 #(
		.INIT('h9fff)
	) name25789 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31616_
	);
	LUT4 #(
		.INIT('hfec7)
	) name25790 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31617_
	);
	LUT4 #(
		.INIT('h0313)
	) name25791 (
		_w31349_,
		_w31353_,
		_w31616_,
		_w31617_,
		_w31618_
	);
	LUT3 #(
		.INIT('h12)
	) name25792 (
		_w31351_,
		_w31352_,
		_w31355_,
		_w31619_
	);
	LUT4 #(
		.INIT('he0f0)
	) name25793 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31620_
	);
	LUT3 #(
		.INIT('h02)
	) name25794 (
		_w31353_,
		_w31620_,
		_w31619_,
		_w31621_
	);
	LUT3 #(
		.INIT('h54)
	) name25795 (
		_w31350_,
		_w31352_,
		_w31353_,
		_w31622_
	);
	LUT2 #(
		.INIT('h8)
	) name25796 (
		_w31356_,
		_w31622_,
		_w31623_
	);
	LUT3 #(
		.INIT('h8a)
	) name25797 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31624_
	);
	LUT3 #(
		.INIT('h15)
	) name25798 (
		_w31349_,
		_w31461_,
		_w31624_,
		_w31625_
	);
	LUT3 #(
		.INIT('h10)
	) name25799 (
		_w31623_,
		_w31621_,
		_w31625_,
		_w31626_
	);
	LUT3 #(
		.INIT('h02)
	) name25800 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31627_
	);
	LUT3 #(
		.INIT('h08)
	) name25801 (
		_w31350_,
		_w31351_,
		_w31355_,
		_w31628_
	);
	LUT4 #(
		.INIT('hfe00)
	) name25802 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31353_,
		_w31629_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name25803 (
		_w31364_,
		_w31627_,
		_w31628_,
		_w31629_,
		_w31630_
	);
	LUT4 #(
		.INIT('h0010)
	) name25804 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31631_
	);
	LUT3 #(
		.INIT('h08)
	) name25805 (
		_w31349_,
		_w31616_,
		_w31631_,
		_w31632_
	);
	LUT3 #(
		.INIT('h20)
	) name25806 (
		_w31359_,
		_w31630_,
		_w31632_,
		_w31633_
	);
	LUT4 #(
		.INIT('h999a)
	) name25807 (
		\u0_L3_reg[13]/NET0131 ,
		_w31618_,
		_w31626_,
		_w31633_,
		_w31634_
	);
	LUT4 #(
		.INIT('h300a)
	) name25808 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31635_
	);
	LUT3 #(
		.INIT('h02)
	) name25809 (
		_w31317_,
		_w31331_,
		_w31635_,
		_w31636_
	);
	LUT4 #(
		.INIT('h4404)
	) name25810 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31637_
	);
	LUT4 #(
		.INIT('hfc5f)
	) name25811 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31638_
	);
	LUT3 #(
		.INIT('h10)
	) name25812 (
		_w31317_,
		_w31637_,
		_w31638_,
		_w31639_
	);
	LUT3 #(
		.INIT('h02)
	) name25813 (
		_w31318_,
		_w31335_,
		_w31344_,
		_w31640_
	);
	LUT3 #(
		.INIT('he0)
	) name25814 (
		_w31636_,
		_w31639_,
		_w31640_,
		_w31641_
	);
	LUT4 #(
		.INIT('h23f0)
	) name25815 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31642_
	);
	LUT3 #(
		.INIT('h10)
	) name25816 (
		_w31317_,
		_w31637_,
		_w31642_,
		_w31643_
	);
	LUT4 #(
		.INIT('hd5ff)
	) name25817 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w31644_
	);
	LUT3 #(
		.INIT('h20)
	) name25818 (
		_w31317_,
		_w31331_,
		_w31644_,
		_w31645_
	);
	LUT4 #(
		.INIT('h0001)
	) name25819 (
		_w31318_,
		_w31340_,
		_w31330_,
		_w31512_,
		_w31646_
	);
	LUT3 #(
		.INIT('he0)
	) name25820 (
		_w31643_,
		_w31645_,
		_w31646_,
		_w31647_
	);
	LUT3 #(
		.INIT('ha9)
	) name25821 (
		\u0_L3_reg[3]/NET0131 ,
		_w31641_,
		_w31647_,
		_w31648_
	);
	LUT3 #(
		.INIT('h20)
	) name25822 (
		_w31580_,
		_w31578_,
		_w31579_,
		_w31649_
	);
	LUT4 #(
		.INIT('h0400)
	) name25823 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31650_
	);
	LUT3 #(
		.INIT('hed)
	) name25824 (
		_w31577_,
		_w31580_,
		_w31579_,
		_w31651_
	);
	LUT3 #(
		.INIT('h10)
	) name25825 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31652_
	);
	LUT4 #(
		.INIT('he2cd)
	) name25826 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31653_
	);
	LUT4 #(
		.INIT('h5054)
	) name25827 (
		_w31576_,
		_w31575_,
		_w31650_,
		_w31653_,
		_w31654_
	);
	LUT2 #(
		.INIT('h8)
	) name25828 (
		_w31586_,
		_w31591_,
		_w31655_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name25829 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31656_
	);
	LUT3 #(
		.INIT('he0)
	) name25830 (
		_w31578_,
		_w31579_,
		_w31575_,
		_w31657_
	);
	LUT4 #(
		.INIT('h0302)
	) name25831 (
		_w31575_,
		_w31581_,
		_w31657_,
		_w31656_,
		_w31658_
	);
	LUT3 #(
		.INIT('ha8)
	) name25832 (
		_w31576_,
		_w31655_,
		_w31658_,
		_w31659_
	);
	LUT4 #(
		.INIT('h1dff)
	) name25833 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31660_
	);
	LUT4 #(
		.INIT('h0024)
	) name25834 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31661_
	);
	LUT4 #(
		.INIT('hcc08)
	) name25835 (
		_w31576_,
		_w31575_,
		_w31660_,
		_w31661_,
		_w31662_
	);
	LUT3 #(
		.INIT('h80)
	) name25836 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31663_
	);
	LUT2 #(
		.INIT('h2)
	) name25837 (
		_w31579_,
		_w31575_,
		_w31664_
	);
	LUT4 #(
		.INIT('h0009)
	) name25838 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31665_
	);
	LUT4 #(
		.INIT('h9db6)
	) name25839 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31666_
	);
	LUT2 #(
		.INIT('h1)
	) name25840 (
		_w31576_,
		_w31575_,
		_w31667_
	);
	LUT4 #(
		.INIT('h7077)
	) name25841 (
		_w31663_,
		_w31664_,
		_w31666_,
		_w31667_,
		_w31668_
	);
	LUT2 #(
		.INIT('h4)
	) name25842 (
		_w31662_,
		_w31668_,
		_w31669_
	);
	LUT4 #(
		.INIT('h5655)
	) name25843 (
		\u0_L3_reg[24]/NET0131 ,
		_w31654_,
		_w31659_,
		_w31669_,
		_w31670_
	);
	LUT4 #(
		.INIT('h0004)
	) name25844 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31671_
	);
	LUT3 #(
		.INIT('h08)
	) name25845 (
		_w31575_,
		_w31651_,
		_w31671_,
		_w31672_
	);
	LUT3 #(
		.INIT('h07)
	) name25846 (
		_w31580_,
		_w31579_,
		_w31575_,
		_w31673_
	);
	LUT2 #(
		.INIT('h4)
	) name25847 (
		_w31652_,
		_w31673_,
		_w31674_
	);
	LUT3 #(
		.INIT('ha8)
	) name25848 (
		_w31576_,
		_w31672_,
		_w31674_,
		_w31675_
	);
	LUT4 #(
		.INIT('h20ac)
	) name25849 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31676_
	);
	LUT4 #(
		.INIT('h8c00)
	) name25850 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31677_
	);
	LUT3 #(
		.INIT('h04)
	) name25851 (
		_w31577_,
		_w31578_,
		_w31579_,
		_w31678_
	);
	LUT4 #(
		.INIT('heee4)
	) name25852 (
		_w31575_,
		_w31676_,
		_w31678_,
		_w31677_,
		_w31679_
	);
	LUT4 #(
		.INIT('h0200)
	) name25853 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31680_
	);
	LUT3 #(
		.INIT('h01)
	) name25854 (
		_w31576_,
		_w31665_,
		_w31680_,
		_w31681_
	);
	LUT2 #(
		.INIT('h4)
	) name25855 (
		_w31679_,
		_w31681_,
		_w31682_
	);
	LUT2 #(
		.INIT('h8)
	) name25856 (
		_w31579_,
		_w31575_,
		_w31683_
	);
	LUT3 #(
		.INIT('h08)
	) name25857 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31684_
	);
	LUT2 #(
		.INIT('h8)
	) name25858 (
		_w31683_,
		_w31684_,
		_w31685_
	);
	LUT4 #(
		.INIT('h0040)
	) name25859 (
		_w31577_,
		_w31578_,
		_w31579_,
		_w31575_,
		_w31686_
	);
	LUT3 #(
		.INIT('h0d)
	) name25860 (
		_w31595_,
		_w31589_,
		_w31686_,
		_w31687_
	);
	LUT2 #(
		.INIT('h4)
	) name25861 (
		_w31685_,
		_w31687_,
		_w31688_
	);
	LUT4 #(
		.INIT('h56aa)
	) name25862 (
		\u0_L3_reg[30]/NET0131 ,
		_w31675_,
		_w31682_,
		_w31688_,
		_w31689_
	);
	LUT4 #(
		.INIT('h9600)
	) name25863 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31690_
	);
	LUT3 #(
		.INIT('h43)
	) name25864 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31691_
	);
	LUT4 #(
		.INIT('h0013)
	) name25865 (
		_w31175_,
		_w31499_,
		_w31691_,
		_w31690_,
		_w31692_
	);
	LUT4 #(
		.INIT('h0043)
	) name25866 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31165_,
		_w31693_
	);
	LUT3 #(
		.INIT('h08)
	) name25867 (
		_w31166_,
		_w31167_,
		_w31169_,
		_w31694_
	);
	LUT3 #(
		.INIT('h60)
	) name25868 (
		_w31168_,
		_w31167_,
		_w31165_,
		_w31695_
	);
	LUT4 #(
		.INIT('hf67f)
	) name25869 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31696_
	);
	LUT4 #(
		.INIT('h0b00)
	) name25870 (
		_w31694_,
		_w31695_,
		_w31693_,
		_w31696_,
		_w31697_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name25871 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w31698_
	);
	LUT2 #(
		.INIT('h1)
	) name25872 (
		_w31165_,
		_w31698_,
		_w31699_
	);
	LUT4 #(
		.INIT('h0e04)
	) name25873 (
		_w31164_,
		_w31697_,
		_w31699_,
		_w31692_,
		_w31700_
	);
	LUT2 #(
		.INIT('h9)
	) name25874 (
		\u0_L3_reg[9]/NET0131 ,
		_w31700_,
		_w31701_
	);
	LUT4 #(
		.INIT('h7d6c)
	) name25875 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31702_
	);
	LUT4 #(
		.INIT('h6800)
	) name25876 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31575_,
		_w31703_
	);
	LUT4 #(
		.INIT('h0032)
	) name25877 (
		_w31575_,
		_w31583_,
		_w31702_,
		_w31703_,
		_w31704_
	);
	LUT2 #(
		.INIT('h1)
	) name25878 (
		_w31576_,
		_w31704_,
		_w31705_
	);
	LUT4 #(
		.INIT('h6979)
	) name25879 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31575_,
		_w31706_
	);
	LUT4 #(
		.INIT('h2000)
	) name25880 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31579_,
		_w31707_
	);
	LUT4 #(
		.INIT('hcc04)
	) name25881 (
		_w31579_,
		_w31576_,
		_w31706_,
		_w31707_,
		_w31708_
	);
	LUT4 #(
		.INIT('h1400)
	) name25882 (
		_w31577_,
		_w31580_,
		_w31579_,
		_w31576_,
		_w31709_
	);
	LUT3 #(
		.INIT('h54)
	) name25883 (
		_w31575_,
		_w31649_,
		_w31709_,
		_w31710_
	);
	LUT3 #(
		.INIT('hbe)
	) name25884 (
		_w31577_,
		_w31580_,
		_w31578_,
		_w31711_
	);
	LUT2 #(
		.INIT('h2)
	) name25885 (
		_w31683_,
		_w31711_,
		_w31712_
	);
	LUT3 #(
		.INIT('h01)
	) name25886 (
		_w31708_,
		_w31710_,
		_w31712_,
		_w31713_
	);
	LUT3 #(
		.INIT('h65)
	) name25887 (
		\u0_L3_reg[16]/NET0131 ,
		_w31705_,
		_w31713_,
		_w31714_
	);
	LUT3 #(
		.INIT('h1d)
	) name25888 (
		_w31350_,
		_w31352_,
		_w31353_,
		_w31715_
	);
	LUT3 #(
		.INIT('h0b)
	) name25889 (
		_w31350_,
		_w31352_,
		_w31355_,
		_w31716_
	);
	LUT4 #(
		.INIT('hdefe)
	) name25890 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31355_,
		_w31717_
	);
	LUT4 #(
		.INIT('h3500)
	) name25891 (
		_w31362_,
		_w31716_,
		_w31715_,
		_w31717_,
		_w31718_
	);
	LUT2 #(
		.INIT('h1)
	) name25892 (
		_w31349_,
		_w31718_,
		_w31719_
	);
	LUT4 #(
		.INIT('h4060)
	) name25893 (
		_w31351_,
		_w31352_,
		_w31353_,
		_w31355_,
		_w31720_
	);
	LUT3 #(
		.INIT('ha8)
	) name25894 (
		_w31349_,
		_w31372_,
		_w31720_,
		_w31721_
	);
	LUT3 #(
		.INIT('hb8)
	) name25895 (
		_w31350_,
		_w31351_,
		_w31352_,
		_w31722_
	);
	LUT2 #(
		.INIT('h8)
	) name25896 (
		_w31349_,
		_w31355_,
		_w31723_
	);
	LUT4 #(
		.INIT('h4544)
	) name25897 (
		_w31353_,
		_w31357_,
		_w31722_,
		_w31723_,
		_w31724_
	);
	LUT4 #(
		.INIT('h80b0)
	) name25898 (
		_w31350_,
		_w31351_,
		_w31353_,
		_w31355_,
		_w31725_
	);
	LUT2 #(
		.INIT('h4)
	) name25899 (
		_w31716_,
		_w31725_,
		_w31726_
	);
	LUT3 #(
		.INIT('h01)
	) name25900 (
		_w31724_,
		_w31721_,
		_w31726_,
		_w31727_
	);
	LUT3 #(
		.INIT('h65)
	) name25901 (
		\u0_L3_reg[18]/NET0131 ,
		_w31719_,
		_w31727_,
		_w31728_
	);
	LUT4 #(
		.INIT('hc963)
	) name25902 (
		decrypt_pad,
		\u0_R2_reg[4]/NET0131 ,
		\u0_uk_K_r2_reg[48]/NET0131 ,
		\u0_uk_K_r2_reg[53]/P0001 ,
		_w31729_
	);
	LUT4 #(
		.INIT('hc963)
	) name25903 (
		decrypt_pad,
		\u0_R2_reg[3]/NET0131 ,
		\u0_uk_K_r2_reg[13]/NET0131 ,
		\u0_uk_K_r2_reg[18]/NET0131 ,
		_w31730_
	);
	LUT4 #(
		.INIT('hc693)
	) name25904 (
		decrypt_pad,
		\u0_R2_reg[1]/NET0131 ,
		\u0_uk_K_r2_reg[26]/NET0131 ,
		\u0_uk_K_r2_reg[46]/NET0131 ,
		_w31731_
	);
	LUT4 #(
		.INIT('hc963)
	) name25905 (
		decrypt_pad,
		\u0_R2_reg[5]/NET0131 ,
		\u0_uk_K_r2_reg[19]/NET0131 ,
		\u0_uk_K_r2_reg[24]/NET0131 ,
		_w31732_
	);
	LUT4 #(
		.INIT('hc693)
	) name25906 (
		decrypt_pad,
		\u0_R2_reg[2]/NET0131 ,
		\u0_uk_K_r2_reg[41]/NET0131 ,
		\u0_uk_K_r2_reg[4]/NET0131 ,
		_w31733_
	);
	LUT4 #(
		.INIT('hc963)
	) name25907 (
		decrypt_pad,
		\u0_R2_reg[32]/NET0131 ,
		\u0_uk_K_r2_reg[25]/NET0131 ,
		\u0_uk_K_r2_reg[5]/NET0131 ,
		_w31734_
	);
	LUT4 #(
		.INIT('hccf5)
	) name25908 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31735_
	);
	LUT2 #(
		.INIT('h2)
	) name25909 (
		_w31730_,
		_w31735_,
		_w31736_
	);
	LUT2 #(
		.INIT('h4)
	) name25910 (
		_w31733_,
		_w31734_,
		_w31737_
	);
	LUT4 #(
		.INIT('h0212)
	) name25911 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31738_
	);
	LUT3 #(
		.INIT('h40)
	) name25912 (
		_w31730_,
		_w31731_,
		_w31734_,
		_w31739_
	);
	LUT2 #(
		.INIT('h4)
	) name25913 (
		_w31734_,
		_w31732_,
		_w31740_
	);
	LUT2 #(
		.INIT('h4)
	) name25914 (
		_w31733_,
		_w31730_,
		_w31741_
	);
	LUT3 #(
		.INIT('hb0)
	) name25915 (
		_w31733_,
		_w31730_,
		_w31731_,
		_w31742_
	);
	LUT4 #(
		.INIT('h0051)
	) name25916 (
		_w31739_,
		_w31740_,
		_w31742_,
		_w31738_,
		_w31743_
	);
	LUT3 #(
		.INIT('h8a)
	) name25917 (
		_w31729_,
		_w31736_,
		_w31743_,
		_w31744_
	);
	LUT4 #(
		.INIT('h0880)
	) name25918 (
		_w31730_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31745_
	);
	LUT2 #(
		.INIT('h8)
	) name25919 (
		_w31733_,
		_w31745_,
		_w31746_
	);
	LUT4 #(
		.INIT('h1013)
	) name25920 (
		_w31733_,
		_w31730_,
		_w31731_,
		_w31732_,
		_w31747_
	);
	LUT4 #(
		.INIT('h4ff3)
	) name25921 (
		_w31730_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31748_
	);
	LUT4 #(
		.INIT('h6f2a)
	) name25922 (
		_w31733_,
		_w31734_,
		_w31747_,
		_w31748_,
		_w31749_
	);
	LUT3 #(
		.INIT('h45)
	) name25923 (
		_w31729_,
		_w31746_,
		_w31749_,
		_w31750_
	);
	LUT4 #(
		.INIT('h7dbb)
	) name25924 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31751_
	);
	LUT2 #(
		.INIT('h1)
	) name25925 (
		_w31730_,
		_w31751_,
		_w31752_
	);
	LUT4 #(
		.INIT('h0400)
	) name25926 (
		_w31733_,
		_w31730_,
		_w31731_,
		_w31734_,
		_w31753_
	);
	LUT2 #(
		.INIT('h1)
	) name25927 (
		_w31731_,
		_w31732_,
		_w31754_
	);
	LUT3 #(
		.INIT('h08)
	) name25928 (
		_w31733_,
		_w31730_,
		_w31734_,
		_w31755_
	);
	LUT3 #(
		.INIT('h15)
	) name25929 (
		_w31753_,
		_w31754_,
		_w31755_,
		_w31756_
	);
	LUT2 #(
		.INIT('h4)
	) name25930 (
		_w31752_,
		_w31756_,
		_w31757_
	);
	LUT4 #(
		.INIT('h5655)
	) name25931 (
		\u0_L2_reg[31]/NET0131 ,
		_w31750_,
		_w31744_,
		_w31757_,
		_w31758_
	);
	LUT4 #(
		.INIT('hc963)
	) name25932 (
		decrypt_pad,
		\u0_R2_reg[24]/NET0131 ,
		\u0_uk_K_r2_reg[15]/NET0131 ,
		\u0_uk_K_r2_reg[52]/NET0131 ,
		_w31759_
	);
	LUT4 #(
		.INIT('hc693)
	) name25933 (
		decrypt_pad,
		\u0_R2_reg[23]/NET0131 ,
		\u0_uk_K_r2_reg[22]/NET0131 ,
		\u0_uk_K_r2_reg[44]/NET0131 ,
		_w31760_
	);
	LUT4 #(
		.INIT('hc963)
	) name25934 (
		decrypt_pad,
		\u0_R2_reg[22]/NET0131 ,
		\u0_uk_K_r2_reg[0]/NET0131 ,
		\u0_uk_K_r2_reg[9]/NET0131 ,
		_w31761_
	);
	LUT4 #(
		.INIT('hc693)
	) name25935 (
		decrypt_pad,
		\u0_R2_reg[21]/NET0131 ,
		\u0_uk_K_r2_reg[42]/NET0131 ,
		\u0_uk_K_r2_reg[9]/NET0131 ,
		_w31762_
	);
	LUT4 #(
		.INIT('hc693)
	) name25936 (
		decrypt_pad,
		\u0_R2_reg[20]/NET0131 ,
		\u0_uk_K_r2_reg[31]/NET0131 ,
		\u0_uk_K_r2_reg[49]/NET0131 ,
		_w31763_
	);
	LUT4 #(
		.INIT('hc963)
	) name25937 (
		decrypt_pad,
		\u0_R2_reg[25]/NET0131 ,
		\u0_uk_K_r2_reg[38]/NET0131 ,
		\u0_uk_K_r2_reg[43]/NET0131 ,
		_w31764_
	);
	LUT4 #(
		.INIT('h0010)
	) name25938 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31765_
	);
	LUT3 #(
		.INIT('h08)
	) name25939 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31766_
	);
	LUT4 #(
		.INIT('h57e7)
	) name25940 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31767_
	);
	LUT2 #(
		.INIT('h2)
	) name25941 (
		_w31760_,
		_w31767_,
		_w31768_
	);
	LUT4 #(
		.INIT('h0040)
	) name25942 (
		_w31761_,
		_w31763_,
		_w31764_,
		_w31760_,
		_w31769_
	);
	LUT2 #(
		.INIT('h4)
	) name25943 (
		_w31762_,
		_w31769_,
		_w31770_
	);
	LUT3 #(
		.INIT('h13)
	) name25944 (
		_w31762_,
		_w31761_,
		_w31764_,
		_w31771_
	);
	LUT3 #(
		.INIT('h07)
	) name25945 (
		_w31763_,
		_w31764_,
		_w31760_,
		_w31772_
	);
	LUT3 #(
		.INIT('h10)
	) name25946 (
		_w31766_,
		_w31771_,
		_w31772_,
		_w31773_
	);
	LUT4 #(
		.INIT('haaa8)
	) name25947 (
		_w31759_,
		_w31768_,
		_w31770_,
		_w31773_,
		_w31774_
	);
	LUT3 #(
		.INIT('h20)
	) name25948 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31775_
	);
	LUT4 #(
		.INIT('h0028)
	) name25949 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31760_,
		_w31776_
	);
	LUT4 #(
		.INIT('h0020)
	) name25950 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31777_
	);
	LUT4 #(
		.INIT('h4000)
	) name25951 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31760_,
		_w31778_
	);
	LUT4 #(
		.INIT('heefb)
	) name25952 (
		_w31761_,
		_w31763_,
		_w31764_,
		_w31760_,
		_w31779_
	);
	LUT3 #(
		.INIT('h10)
	) name25953 (
		_w31777_,
		_w31778_,
		_w31779_,
		_w31780_
	);
	LUT4 #(
		.INIT('h4000)
	) name25954 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31781_
	);
	LUT4 #(
		.INIT('h1000)
	) name25955 (
		_w31762_,
		_w31763_,
		_w31764_,
		_w31760_,
		_w31782_
	);
	LUT2 #(
		.INIT('h1)
	) name25956 (
		_w31781_,
		_w31782_,
		_w31783_
	);
	LUT4 #(
		.INIT('h4555)
	) name25957 (
		_w31759_,
		_w31776_,
		_w31780_,
		_w31783_,
		_w31784_
	);
	LUT4 #(
		.INIT('heff7)
	) name25958 (
		_w31762_,
		_w31763_,
		_w31764_,
		_w31760_,
		_w31785_
	);
	LUT2 #(
		.INIT('h1)
	) name25959 (
		_w31761_,
		_w31785_,
		_w31786_
	);
	LUT3 #(
		.INIT('h01)
	) name25960 (
		_w31762_,
		_w31763_,
		_w31764_,
		_w31787_
	);
	LUT4 #(
		.INIT('h0002)
	) name25961 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31788_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name25962 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31789_
	);
	LUT4 #(
		.INIT('hef23)
	) name25963 (
		_w31761_,
		_w31760_,
		_w31787_,
		_w31789_,
		_w31790_
	);
	LUT2 #(
		.INIT('h4)
	) name25964 (
		_w31786_,
		_w31790_,
		_w31791_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name25965 (
		\u0_L2_reg[11]/NET0131 ,
		_w31784_,
		_w31774_,
		_w31791_,
		_w31792_
	);
	LUT4 #(
		.INIT('hc963)
	) name25966 (
		decrypt_pad,
		\u0_R2_reg[26]/NET0131 ,
		\u0_uk_K_r2_reg[2]/NET0131 ,
		\u0_uk_K_r2_reg[35]/NET0131 ,
		_w31793_
	);
	LUT4 #(
		.INIT('hc963)
	) name25967 (
		decrypt_pad,
		\u0_R2_reg[25]/NET0131 ,
		\u0_uk_K_r2_reg[45]/NET0131 ,
		\u0_uk_K_r2_reg[50]/NET0131 ,
		_w31794_
	);
	LUT4 #(
		.INIT('hc693)
	) name25968 (
		decrypt_pad,
		\u0_R2_reg[24]/NET0131 ,
		\u0_uk_K_r2_reg[15]/NET0131 ,
		\u0_uk_K_r2_reg[37]/NET0131 ,
		_w31795_
	);
	LUT4 #(
		.INIT('hc963)
	) name25969 (
		decrypt_pad,
		\u0_R2_reg[29]/NET0131 ,
		\u0_uk_K_r2_reg[14]/NET0131 ,
		\u0_uk_K_r2_reg[23]/NET0131 ,
		_w31796_
	);
	LUT2 #(
		.INIT('h4)
	) name25970 (
		_w31795_,
		_w31796_,
		_w31797_
	);
	LUT4 #(
		.INIT('h0200)
	) name25971 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w31798_
	);
	LUT4 #(
		.INIT('h0008)
	) name25972 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w31799_
	);
	LUT4 #(
		.INIT('hfdf7)
	) name25973 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w31800_
	);
	LUT4 #(
		.INIT('hc693)
	) name25974 (
		decrypt_pad,
		\u0_R2_reg[28]/NET0131 ,
		\u0_uk_K_r2_reg[0]/NET0131 ,
		\u0_uk_K_r2_reg[22]/NET0131 ,
		_w31801_
	);
	LUT4 #(
		.INIT('h9cfc)
	) name25975 (
		_w31793_,
		_w31794_,
		_w31796_,
		_w31801_,
		_w31802_
	);
	LUT4 #(
		.INIT('hc963)
	) name25976 (
		decrypt_pad,
		\u0_R2_reg[27]/NET0131 ,
		\u0_uk_K_r2_reg[35]/NET0131 ,
		\u0_uk_K_r2_reg[44]/NET0131 ,
		_w31803_
	);
	LUT4 #(
		.INIT('h3b00)
	) name25977 (
		_w31795_,
		_w31800_,
		_w31802_,
		_w31803_,
		_w31804_
	);
	LUT4 #(
		.INIT('hee72)
	) name25978 (
		_w31793_,
		_w31794_,
		_w31796_,
		_w31803_,
		_w31805_
	);
	LUT2 #(
		.INIT('h2)
	) name25979 (
		_w31795_,
		_w31805_,
		_w31806_
	);
	LUT4 #(
		.INIT('h0002)
	) name25980 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w31807_
	);
	LUT2 #(
		.INIT('h6)
	) name25981 (
		_w31793_,
		_w31795_,
		_w31808_
	);
	LUT3 #(
		.INIT('h8c)
	) name25982 (
		_w31794_,
		_w31796_,
		_w31803_,
		_w31809_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name25983 (
		_w31803_,
		_w31807_,
		_w31808_,
		_w31809_,
		_w31810_
	);
	LUT3 #(
		.INIT('h45)
	) name25984 (
		_w31801_,
		_w31806_,
		_w31810_,
		_w31811_
	);
	LUT4 #(
		.INIT('h1000)
	) name25985 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w31812_
	);
	LUT4 #(
		.INIT('he3ff)
	) name25986 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w31813_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name25987 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w31814_
	);
	LUT4 #(
		.INIT('h02aa)
	) name25988 (
		_w31801_,
		_w31803_,
		_w31813_,
		_w31814_,
		_w31815_
	);
	LUT4 #(
		.INIT('h0084)
	) name25989 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31803_,
		_w31816_
	);
	LUT4 #(
		.INIT('h0100)
	) name25990 (
		_w31793_,
		_w31794_,
		_w31796_,
		_w31803_,
		_w31817_
	);
	LUT2 #(
		.INIT('h1)
	) name25991 (
		_w31816_,
		_w31817_,
		_w31818_
	);
	LUT2 #(
		.INIT('h4)
	) name25992 (
		_w31815_,
		_w31818_,
		_w31819_
	);
	LUT4 #(
		.INIT('h5655)
	) name25993 (
		\u0_L2_reg[22]/NET0131 ,
		_w31804_,
		_w31811_,
		_w31819_,
		_w31820_
	);
	LUT4 #(
		.INIT('hc963)
	) name25994 (
		decrypt_pad,
		\u0_R2_reg[8]/NET0131 ,
		\u0_uk_K_r2_reg[17]/NET0131 ,
		\u0_uk_K_r2_reg[54]/NET0131 ,
		_w31821_
	);
	LUT4 #(
		.INIT('hc693)
	) name25995 (
		decrypt_pad,
		\u0_R2_reg[4]/NET0131 ,
		\u0_uk_K_r2_reg[10]/NET0131 ,
		\u0_uk_K_r2_reg[5]/NET0131 ,
		_w31822_
	);
	LUT4 #(
		.INIT('hc693)
	) name25996 (
		decrypt_pad,
		\u0_R2_reg[9]/NET0131 ,
		\u0_uk_K_r2_reg[34]/NET0131 ,
		\u0_uk_K_r2_reg[54]/NET0131 ,
		_w31823_
	);
	LUT4 #(
		.INIT('hc963)
	) name25997 (
		decrypt_pad,
		\u0_R2_reg[5]/NET0131 ,
		\u0_uk_K_r2_reg[41]/NET0131 ,
		\u0_uk_K_r2_reg[46]/NET0131 ,
		_w31824_
	);
	LUT4 #(
		.INIT('hc693)
	) name25998 (
		decrypt_pad,
		\u0_R2_reg[6]/NET0131 ,
		\u0_uk_K_r2_reg[12]/NET0131 ,
		\u0_uk_K_r2_reg[32]/NET0131 ,
		_w31825_
	);
	LUT4 #(
		.INIT('h59fb)
	) name25999 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31826_
	);
	LUT4 #(
		.INIT('hc963)
	) name26000 (
		decrypt_pad,
		\u0_R2_reg[7]/NET0131 ,
		\u0_uk_K_r2_reg[26]/NET0131 ,
		\u0_uk_K_r2_reg[6]/NET0131 ,
		_w31827_
	);
	LUT2 #(
		.INIT('h1)
	) name26001 (
		_w31826_,
		_w31827_,
		_w31828_
	);
	LUT4 #(
		.INIT('hbf00)
	) name26002 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31829_
	);
	LUT2 #(
		.INIT('h1)
	) name26003 (
		_w31824_,
		_w31827_,
		_w31830_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name26004 (
		_w31823_,
		_w31824_,
		_w31825_,
		_w31827_,
		_w31831_
	);
	LUT2 #(
		.INIT('h1)
	) name26005 (
		_w31829_,
		_w31831_,
		_w31832_
	);
	LUT4 #(
		.INIT('h0034)
	) name26006 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31833_
	);
	LUT2 #(
		.INIT('h8)
	) name26007 (
		_w31822_,
		_w31823_,
		_w31834_
	);
	LUT4 #(
		.INIT('h0800)
	) name26008 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31835_
	);
	LUT3 #(
		.INIT('h15)
	) name26009 (
		_w31833_,
		_w31827_,
		_w31835_,
		_w31836_
	);
	LUT4 #(
		.INIT('h5455)
	) name26010 (
		_w31821_,
		_w31828_,
		_w31832_,
		_w31836_,
		_w31837_
	);
	LUT4 #(
		.INIT('he6ee)
	) name26011 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31838_
	);
	LUT4 #(
		.INIT('h4044)
	) name26012 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31839_
	);
	LUT3 #(
		.INIT('h0d)
	) name26013 (
		_w31824_,
		_w31825_,
		_w31827_,
		_w31840_
	);
	LUT4 #(
		.INIT('hf200)
	) name26014 (
		_w31821_,
		_w31838_,
		_w31839_,
		_w31840_,
		_w31841_
	);
	LUT4 #(
		.INIT('hfe5f)
	) name26015 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31842_
	);
	LUT2 #(
		.INIT('h2)
	) name26016 (
		_w31827_,
		_w31842_,
		_w31843_
	);
	LUT4 #(
		.INIT('h0080)
	) name26017 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31844_
	);
	LUT4 #(
		.INIT('h0002)
	) name26018 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31845_
	);
	LUT4 #(
		.INIT('h8c00)
	) name26019 (
		_w31822_,
		_w31824_,
		_w31825_,
		_w31827_,
		_w31846_
	);
	LUT4 #(
		.INIT('haaa8)
	) name26020 (
		_w31821_,
		_w31845_,
		_w31846_,
		_w31844_,
		_w31847_
	);
	LUT3 #(
		.INIT('h01)
	) name26021 (
		_w31843_,
		_w31847_,
		_w31841_,
		_w31848_
	);
	LUT3 #(
		.INIT('h65)
	) name26022 (
		\u0_L2_reg[2]/NET0131 ,
		_w31837_,
		_w31848_,
		_w31849_
	);
	LUT4 #(
		.INIT('h8aa8)
	) name26023 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31850_
	);
	LUT4 #(
		.INIT('h1005)
	) name26024 (
		_w31730_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31851_
	);
	LUT4 #(
		.INIT('h8020)
	) name26025 (
		_w31730_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31852_
	);
	LUT4 #(
		.INIT('hfd7f)
	) name26026 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31853_
	);
	LUT4 #(
		.INIT('h0b00)
	) name26027 (
		_w31850_,
		_w31851_,
		_w31852_,
		_w31853_,
		_w31854_
	);
	LUT2 #(
		.INIT('h1)
	) name26028 (
		_w31729_,
		_w31854_,
		_w31855_
	);
	LUT2 #(
		.INIT('h1)
	) name26029 (
		_w31733_,
		_w31731_,
		_w31856_
	);
	LUT4 #(
		.INIT('h1000)
	) name26030 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31857_
	);
	LUT4 #(
		.INIT('he1f1)
	) name26031 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31858_
	);
	LUT2 #(
		.INIT('h2)
	) name26032 (
		_w31730_,
		_w31858_,
		_w31859_
	);
	LUT4 #(
		.INIT('h0040)
	) name26033 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w31860_
	);
	LUT4 #(
		.INIT('h2201)
	) name26034 (
		_w31733_,
		_w31730_,
		_w31731_,
		_w31734_,
		_w31861_
	);
	LUT3 #(
		.INIT('h80)
	) name26035 (
		_w31733_,
		_w31731_,
		_w31732_,
		_w31862_
	);
	LUT3 #(
		.INIT('h01)
	) name26036 (
		_w31861_,
		_w31860_,
		_w31862_,
		_w31863_
	);
	LUT3 #(
		.INIT('hb7)
	) name26037 (
		_w31733_,
		_w31731_,
		_w31732_,
		_w31864_
	);
	LUT2 #(
		.INIT('h2)
	) name26038 (
		_w31730_,
		_w31734_,
		_w31865_
	);
	LUT2 #(
		.INIT('h4)
	) name26039 (
		_w31864_,
		_w31865_,
		_w31866_
	);
	LUT4 #(
		.INIT('h0075)
	) name26040 (
		_w31729_,
		_w31859_,
		_w31863_,
		_w31866_,
		_w31867_
	);
	LUT3 #(
		.INIT('h65)
	) name26041 (
		\u0_L2_reg[17]/NET0131 ,
		_w31855_,
		_w31867_,
		_w31868_
	);
	LUT4 #(
		.INIT('h5fa6)
	) name26042 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31869_
	);
	LUT4 #(
		.INIT('h3202)
	) name26043 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31870_
	);
	LUT4 #(
		.INIT('hcd7d)
	) name26044 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31871_
	);
	LUT4 #(
		.INIT('h0400)
	) name26045 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31872_
	);
	LUT4 #(
		.INIT('h00e4)
	) name26046 (
		_w31760_,
		_w31871_,
		_w31869_,
		_w31872_,
		_w31873_
	);
	LUT2 #(
		.INIT('h1)
	) name26047 (
		_w31759_,
		_w31873_,
		_w31874_
	);
	LUT4 #(
		.INIT('hf57d)
	) name26048 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31875_
	);
	LUT2 #(
		.INIT('h2)
	) name26049 (
		_w31760_,
		_w31875_,
		_w31876_
	);
	LUT4 #(
		.INIT('hab00)
	) name26050 (
		_w31762_,
		_w31761_,
		_w31764_,
		_w31760_,
		_w31877_
	);
	LUT3 #(
		.INIT('h28)
	) name26051 (
		_w31761_,
		_w31763_,
		_w31764_,
		_w31878_
	);
	LUT3 #(
		.INIT('h01)
	) name26052 (
		_w31877_,
		_w31878_,
		_w31870_,
		_w31879_
	);
	LUT4 #(
		.INIT('h2000)
	) name26053 (
		_w31762_,
		_w31761_,
		_w31764_,
		_w31760_,
		_w31880_
	);
	LUT2 #(
		.INIT('h1)
	) name26054 (
		_w31765_,
		_w31880_,
		_w31881_
	);
	LUT4 #(
		.INIT('h5700)
	) name26055 (
		_w31759_,
		_w31876_,
		_w31879_,
		_w31881_,
		_w31882_
	);
	LUT3 #(
		.INIT('h9a)
	) name26056 (
		\u0_L2_reg[29]/NET0131 ,
		_w31874_,
		_w31882_,
		_w31883_
	);
	LUT4 #(
		.INIT('hfbf5)
	) name26057 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31884_
	);
	LUT2 #(
		.INIT('h1)
	) name26058 (
		_w31760_,
		_w31884_,
		_w31885_
	);
	LUT4 #(
		.INIT('hbc5f)
	) name26059 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31886_
	);
	LUT4 #(
		.INIT('h0301)
	) name26060 (
		_w31760_,
		_w31765_,
		_w31769_,
		_w31886_,
		_w31887_
	);
	LUT3 #(
		.INIT('h45)
	) name26061 (
		_w31759_,
		_w31885_,
		_w31887_,
		_w31888_
	);
	LUT3 #(
		.INIT('h02)
	) name26062 (
		_w31762_,
		_w31761_,
		_w31764_,
		_w31889_
	);
	LUT4 #(
		.INIT('hfcdc)
	) name26063 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31890_
	);
	LUT2 #(
		.INIT('h1)
	) name26064 (
		_w31760_,
		_w31890_,
		_w31891_
	);
	LUT4 #(
		.INIT('h4000)
	) name26065 (
		_w31761_,
		_w31763_,
		_w31764_,
		_w31760_,
		_w31892_
	);
	LUT3 #(
		.INIT('h80)
	) name26066 (
		_w31762_,
		_w31761_,
		_w31764_,
		_w31893_
	);
	LUT3 #(
		.INIT('h01)
	) name26067 (
		_w31788_,
		_w31892_,
		_w31893_,
		_w31894_
	);
	LUT4 #(
		.INIT('h7fbc)
	) name26068 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w31895_
	);
	LUT3 #(
		.INIT('hd6)
	) name26069 (
		_w31762_,
		_w31763_,
		_w31764_,
		_w31896_
	);
	LUT4 #(
		.INIT('hfc74)
	) name26070 (
		_w31761_,
		_w31760_,
		_w31895_,
		_w31896_,
		_w31897_
	);
	LUT4 #(
		.INIT('h7500)
	) name26071 (
		_w31759_,
		_w31891_,
		_w31894_,
		_w31897_,
		_w31898_
	);
	LUT3 #(
		.INIT('h65)
	) name26072 (
		\u0_L2_reg[4]/NET0131 ,
		_w31888_,
		_w31898_,
		_w31899_
	);
	LUT4 #(
		.INIT('hc693)
	) name26073 (
		decrypt_pad,
		\u0_R2_reg[31]/NET0131 ,
		\u0_uk_K_r2_reg[14]/NET0131 ,
		\u0_uk_K_r2_reg[36]/NET0131 ,
		_w31900_
	);
	LUT4 #(
		.INIT('hc693)
	) name26074 (
		decrypt_pad,
		\u0_R2_reg[28]/NET0131 ,
		\u0_uk_K_r2_reg[29]/NET0131 ,
		\u0_uk_K_r2_reg[51]/NET0131 ,
		_w31901_
	);
	LUT4 #(
		.INIT('hc693)
	) name26075 (
		decrypt_pad,
		\u0_R2_reg[30]/NET0131 ,
		\u0_uk_K_r2_reg[2]/NET0131 ,
		\u0_uk_K_r2_reg[52]/NET0131 ,
		_w31902_
	);
	LUT2 #(
		.INIT('h2)
	) name26076 (
		_w31901_,
		_w31902_,
		_w31903_
	);
	LUT4 #(
		.INIT('hc693)
	) name26077 (
		decrypt_pad,
		\u0_R2_reg[1]/NET0131 ,
		\u0_uk_K_r2_reg[45]/NET0131 ,
		\u0_uk_K_r2_reg[8]/NET0131 ,
		_w31904_
	);
	LUT4 #(
		.INIT('hc693)
	) name26078 (
		decrypt_pad,
		\u0_R2_reg[29]/NET0131 ,
		\u0_uk_K_r2_reg[1]/NET0131 ,
		\u0_uk_K_r2_reg[23]/NET0131 ,
		_w31905_
	);
	LUT2 #(
		.INIT('h4)
	) name26079 (
		_w31904_,
		_w31905_,
		_w31906_
	);
	LUT4 #(
		.INIT('hc963)
	) name26080 (
		decrypt_pad,
		\u0_R2_reg[32]/NET0131 ,
		\u0_uk_K_r2_reg[42]/NET0131 ,
		\u0_uk_K_r2_reg[51]/NET0131 ,
		_w31907_
	);
	LUT4 #(
		.INIT('h0020)
	) name26081 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31908_
	);
	LUT4 #(
		.INIT('h1000)
	) name26082 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31909_
	);
	LUT2 #(
		.INIT('h1)
	) name26083 (
		_w31905_,
		_w31902_,
		_w31910_
	);
	LUT4 #(
		.INIT('heff7)
	) name26084 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31911_
	);
	LUT4 #(
		.INIT('h0400)
	) name26085 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31912_
	);
	LUT3 #(
		.INIT('h01)
	) name26086 (
		_w31901_,
		_w31905_,
		_w31902_,
		_w31913_
	);
	LUT4 #(
		.INIT('h0001)
	) name26087 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31914_
	);
	LUT4 #(
		.INIT('hebf6)
	) name26088 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31915_
	);
	LUT4 #(
		.INIT('hd700)
	) name26089 (
		_w31907_,
		_w31903_,
		_w31906_,
		_w31915_,
		_w31916_
	);
	LUT2 #(
		.INIT('h2)
	) name26090 (
		_w31900_,
		_w31916_,
		_w31917_
	);
	LUT4 #(
		.INIT('h0200)
	) name26091 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31918_
	);
	LUT4 #(
		.INIT('haa8a)
	) name26092 (
		_w31900_,
		_w31901_,
		_w31904_,
		_w31905_,
		_w31919_
	);
	LUT3 #(
		.INIT('h10)
	) name26093 (
		_w31901_,
		_w31904_,
		_w31902_,
		_w31920_
	);
	LUT3 #(
		.INIT('h15)
	) name26094 (
		_w31900_,
		_w31904_,
		_w31905_,
		_w31921_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name26095 (
		_w31918_,
		_w31919_,
		_w31920_,
		_w31921_,
		_w31922_
	);
	LUT4 #(
		.INIT('h8000)
	) name26096 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31923_
	);
	LUT3 #(
		.INIT('h04)
	) name26097 (
		_w31900_,
		_w31901_,
		_w31902_,
		_w31924_
	);
	LUT3 #(
		.INIT('h01)
	) name26098 (
		_w31908_,
		_w31924_,
		_w31923_,
		_w31925_
	);
	LUT3 #(
		.INIT('h45)
	) name26099 (
		_w31907_,
		_w31922_,
		_w31925_,
		_w31926_
	);
	LUT2 #(
		.INIT('h4)
	) name26100 (
		_w31900_,
		_w31908_,
		_w31927_
	);
	LUT4 #(
		.INIT('h4000)
	) name26101 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31928_
	);
	LUT4 #(
		.INIT('hb5fa)
	) name26102 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w31929_
	);
	LUT4 #(
		.INIT('h00a2)
	) name26103 (
		_w31907_,
		_w31900_,
		_w31928_,
		_w31929_,
		_w31930_
	);
	LUT2 #(
		.INIT('h1)
	) name26104 (
		_w31927_,
		_w31930_,
		_w31931_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name26105 (
		\u0_L2_reg[5]/NET0131 ,
		_w31926_,
		_w31917_,
		_w31931_,
		_w31932_
	);
	LUT4 #(
		.INIT('hc963)
	) name26106 (
		decrypt_pad,
		\u0_R2_reg[16]/NET0131 ,
		\u0_uk_K_r2_reg[18]/NET0131 ,
		\u0_uk_K_r2_reg[55]/NET0131 ,
		_w31933_
	);
	LUT4 #(
		.INIT('hc693)
	) name26107 (
		decrypt_pad,
		\u0_R2_reg[12]/NET0131 ,
		\u0_uk_K_r2_reg[19]/NET0131 ,
		\u0_uk_K_r2_reg[39]/NET0131 ,
		_w31934_
	);
	LUT4 #(
		.INIT('hc963)
	) name26108 (
		decrypt_pad,
		\u0_R2_reg[15]/NET0131 ,
		\u0_uk_K_r2_reg[10]/NET0131 ,
		\u0_uk_K_r2_reg[47]/NET0131 ,
		_w31935_
	);
	LUT4 #(
		.INIT('hc693)
	) name26109 (
		decrypt_pad,
		\u0_R2_reg[13]/NET0131 ,
		\u0_uk_K_r2_reg[13]/NET0131 ,
		\u0_uk_K_r2_reg[33]/NET0131 ,
		_w31936_
	);
	LUT4 #(
		.INIT('hc963)
	) name26110 (
		decrypt_pad,
		\u0_R2_reg[14]/NET0131 ,
		\u0_uk_K_r2_reg[34]/NET0131 ,
		\u0_uk_K_r2_reg[39]/NET0131 ,
		_w31937_
	);
	LUT3 #(
		.INIT('h80)
	) name26111 (
		_w31935_,
		_w31936_,
		_w31937_,
		_w31938_
	);
	LUT4 #(
		.INIT('h0800)
	) name26112 (
		_w31935_,
		_w31936_,
		_w31934_,
		_w31937_,
		_w31939_
	);
	LUT4 #(
		.INIT('hc693)
	) name26113 (
		decrypt_pad,
		\u0_R2_reg[17]/NET0131 ,
		\u0_uk_K_r2_reg[3]/NET0131 ,
		\u0_uk_K_r2_reg[55]/NET0131 ,
		_w31940_
	);
	LUT4 #(
		.INIT('h0002)
	) name26114 (
		_w31935_,
		_w31936_,
		_w31934_,
		_w31940_,
		_w31941_
	);
	LUT2 #(
		.INIT('h8)
	) name26115 (
		_w31934_,
		_w31940_,
		_w31942_
	);
	LUT3 #(
		.INIT('h74)
	) name26116 (
		_w31935_,
		_w31936_,
		_w31937_,
		_w31943_
	);
	LUT4 #(
		.INIT('h0031)
	) name26117 (
		_w31942_,
		_w31941_,
		_w31943_,
		_w31939_,
		_w31944_
	);
	LUT4 #(
		.INIT('h0200)
	) name26118 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31945_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name26119 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31946_
	);
	LUT4 #(
		.INIT('ha3af)
	) name26120 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31947_
	);
	LUT3 #(
		.INIT('hc8)
	) name26121 (
		_w31935_,
		_w31946_,
		_w31947_,
		_w31948_
	);
	LUT3 #(
		.INIT('h15)
	) name26122 (
		_w31933_,
		_w31944_,
		_w31948_,
		_w31949_
	);
	LUT3 #(
		.INIT('h04)
	) name26123 (
		_w31936_,
		_w31934_,
		_w31937_,
		_w31950_
	);
	LUT3 #(
		.INIT('hf9)
	) name26124 (
		_w31936_,
		_w31934_,
		_w31937_,
		_w31951_
	);
	LUT4 #(
		.INIT('h0100)
	) name26125 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31952_
	);
	LUT4 #(
		.INIT('hfe99)
	) name26126 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31953_
	);
	LUT2 #(
		.INIT('h1)
	) name26127 (
		_w31935_,
		_w31953_,
		_w31954_
	);
	LUT4 #(
		.INIT('h0080)
	) name26128 (
		_w31935_,
		_w31936_,
		_w31934_,
		_w31940_,
		_w31955_
	);
	LUT4 #(
		.INIT('h0020)
	) name26129 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31956_
	);
	LUT2 #(
		.INIT('h1)
	) name26130 (
		_w31955_,
		_w31956_,
		_w31957_
	);
	LUT4 #(
		.INIT('h8000)
	) name26131 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31958_
	);
	LUT2 #(
		.INIT('h4)
	) name26132 (
		_w31934_,
		_w31940_,
		_w31959_
	);
	LUT4 #(
		.INIT('h0200)
	) name26133 (
		_w31935_,
		_w31936_,
		_w31934_,
		_w31940_,
		_w31960_
	);
	LUT4 #(
		.INIT('h0001)
	) name26134 (
		_w31955_,
		_w31956_,
		_w31958_,
		_w31960_,
		_w31961_
	);
	LUT3 #(
		.INIT('h8a)
	) name26135 (
		_w31933_,
		_w31954_,
		_w31961_,
		_w31962_
	);
	LUT4 #(
		.INIT('h0400)
	) name26136 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31963_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name26137 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31964_
	);
	LUT2 #(
		.INIT('h2)
	) name26138 (
		_w31935_,
		_w31964_,
		_w31965_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name26139 (
		_w31935_,
		_w31955_,
		_w31937_,
		_w31956_,
		_w31966_
	);
	LUT2 #(
		.INIT('h4)
	) name26140 (
		_w31965_,
		_w31966_,
		_w31967_
	);
	LUT4 #(
		.INIT('h5655)
	) name26141 (
		\u0_L2_reg[20]/NET0131 ,
		_w31962_,
		_w31949_,
		_w31967_,
		_w31968_
	);
	LUT2 #(
		.INIT('h1)
	) name26142 (
		_w31822_,
		_w31825_,
		_w31969_
	);
	LUT4 #(
		.INIT('h6d7d)
	) name26143 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31970_
	);
	LUT2 #(
		.INIT('h2)
	) name26144 (
		_w31827_,
		_w31970_,
		_w31971_
	);
	LUT4 #(
		.INIT('hbfae)
	) name26145 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31972_
	);
	LUT2 #(
		.INIT('h1)
	) name26146 (
		_w31827_,
		_w31972_,
		_w31973_
	);
	LUT2 #(
		.INIT('h8)
	) name26147 (
		_w31822_,
		_w31827_,
		_w31974_
	);
	LUT4 #(
		.INIT('h55f7)
	) name26148 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31827_,
		_w31975_
	);
	LUT4 #(
		.INIT('h0400)
	) name26149 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31976_
	);
	LUT3 #(
		.INIT('h0e)
	) name26150 (
		_w31825_,
		_w31975_,
		_w31976_,
		_w31977_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name26151 (
		_w31821_,
		_w31971_,
		_w31973_,
		_w31977_,
		_w31978_
	);
	LUT4 #(
		.INIT('hdaff)
	) name26152 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31979_
	);
	LUT2 #(
		.INIT('h1)
	) name26153 (
		_w31827_,
		_w31979_,
		_w31980_
	);
	LUT4 #(
		.INIT('h5b59)
	) name26154 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31981_
	);
	LUT4 #(
		.INIT('hd6ff)
	) name26155 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w31982_
	);
	LUT4 #(
		.INIT('he400)
	) name26156 (
		_w31827_,
		_w31981_,
		_w31972_,
		_w31982_,
		_w31983_
	);
	LUT3 #(
		.INIT('h32)
	) name26157 (
		_w31821_,
		_w31980_,
		_w31983_,
		_w31984_
	);
	LUT3 #(
		.INIT('h65)
	) name26158 (
		\u0_L2_reg[28]/NET0131 ,
		_w31978_,
		_w31984_,
		_w31985_
	);
	LUT4 #(
		.INIT('h0800)
	) name26159 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31986_
	);
	LUT3 #(
		.INIT('h01)
	) name26160 (
		_w31935_,
		_w31952_,
		_w31986_,
		_w31987_
	);
	LUT4 #(
		.INIT('hafab)
	) name26161 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31988_
	);
	LUT2 #(
		.INIT('h2)
	) name26162 (
		_w31933_,
		_w31988_,
		_w31989_
	);
	LUT4 #(
		.INIT('h6fff)
	) name26163 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31990_
	);
	LUT3 #(
		.INIT('h20)
	) name26164 (
		_w31935_,
		_w31945_,
		_w31990_,
		_w31991_
	);
	LUT3 #(
		.INIT('h45)
	) name26165 (
		_w31987_,
		_w31989_,
		_w31991_,
		_w31992_
	);
	LUT4 #(
		.INIT('hdf55)
	) name26166 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w31993_
	);
	LUT3 #(
		.INIT('h51)
	) name26167 (
		_w31935_,
		_w31934_,
		_w31940_,
		_w31994_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name26168 (
		_w31933_,
		_w31936_,
		_w31934_,
		_w31937_,
		_w31995_
	);
	LUT4 #(
		.INIT('h4500)
	) name26169 (
		_w31986_,
		_w31993_,
		_w31994_,
		_w31995_,
		_w31996_
	);
	LUT3 #(
		.INIT('h01)
	) name26170 (
		_w31934_,
		_w31940_,
		_w31937_,
		_w31997_
	);
	LUT3 #(
		.INIT('h02)
	) name26171 (
		_w31935_,
		_w31963_,
		_w31997_,
		_w31998_
	);
	LUT3 #(
		.INIT('h40)
	) name26172 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31999_
	);
	LUT4 #(
		.INIT('h5551)
	) name26173 (
		_w31935_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32000_
	);
	LUT2 #(
		.INIT('h4)
	) name26174 (
		_w31999_,
		_w32000_,
		_w32001_
	);
	LUT4 #(
		.INIT('h8008)
	) name26175 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32002_
	);
	LUT3 #(
		.INIT('h01)
	) name26176 (
		_w31933_,
		_w31956_,
		_w32002_,
		_w32003_
	);
	LUT4 #(
		.INIT('h0155)
	) name26177 (
		_w31996_,
		_w31998_,
		_w32001_,
		_w32003_,
		_w32004_
	);
	LUT3 #(
		.INIT('h56)
	) name26178 (
		\u0_L2_reg[1]/NET0131 ,
		_w31992_,
		_w32004_,
		_w32005_
	);
	LUT4 #(
		.INIT('hf3db)
	) name26179 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32006_
	);
	LUT4 #(
		.INIT('hfdbd)
	) name26180 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32007_
	);
	LUT4 #(
		.INIT('hc480)
	) name26181 (
		_w31935_,
		_w31990_,
		_w32007_,
		_w32006_,
		_w32008_
	);
	LUT2 #(
		.INIT('h2)
	) name26182 (
		_w31933_,
		_w32008_,
		_w32009_
	);
	LUT4 #(
		.INIT('hdd31)
	) name26183 (
		_w31935_,
		_w31936_,
		_w31940_,
		_w31937_,
		_w32010_
	);
	LUT2 #(
		.INIT('h2)
	) name26184 (
		_w31934_,
		_w32010_,
		_w32011_
	);
	LUT4 #(
		.INIT('h0060)
	) name26185 (
		_w31935_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32012_
	);
	LUT4 #(
		.INIT('h0001)
	) name26186 (
		_w31935_,
		_w31936_,
		_w31934_,
		_w31940_,
		_w32013_
	);
	LUT3 #(
		.INIT('h02)
	) name26187 (
		_w31946_,
		_w32013_,
		_w32012_,
		_w32014_
	);
	LUT3 #(
		.INIT('h45)
	) name26188 (
		_w31933_,
		_w32011_,
		_w32014_,
		_w32015_
	);
	LUT4 #(
		.INIT('h6ffe)
	) name26189 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32016_
	);
	LUT2 #(
		.INIT('h1)
	) name26190 (
		_w31935_,
		_w32016_,
		_w32017_
	);
	LUT3 #(
		.INIT('h0d)
	) name26191 (
		_w31955_,
		_w31937_,
		_w31939_,
		_w32018_
	);
	LUT2 #(
		.INIT('h4)
	) name26192 (
		_w32017_,
		_w32018_,
		_w32019_
	);
	LUT4 #(
		.INIT('h5655)
	) name26193 (
		\u0_L2_reg[10]/NET0131 ,
		_w32015_,
		_w32009_,
		_w32019_,
		_w32020_
	);
	LUT4 #(
		.INIT('hc963)
	) name26194 (
		decrypt_pad,
		\u0_R2_reg[20]/NET0131 ,
		\u0_uk_K_r2_reg[31]/NET0131 ,
		\u0_uk_K_r2_reg[36]/NET0131 ,
		_w32021_
	);
	LUT4 #(
		.INIT('hc693)
	) name26195 (
		decrypt_pad,
		\u0_R2_reg[19]/NET0131 ,
		\u0_uk_K_r2_reg[21]/NET0131 ,
		\u0_uk_K_r2_reg[43]/NET0131 ,
		_w32022_
	);
	LUT4 #(
		.INIT('hc963)
	) name26196 (
		decrypt_pad,
		\u0_R2_reg[16]/NET0131 ,
		\u0_uk_K_r2_reg[16]/NET0131 ,
		\u0_uk_K_r2_reg[49]/NET0131 ,
		_w32023_
	);
	LUT4 #(
		.INIT('hc693)
	) name26197 (
		decrypt_pad,
		\u0_R2_reg[17]/NET0131 ,
		\u0_uk_K_r2_reg[16]/NET0131 ,
		\u0_uk_K_r2_reg[7]/NET0131 ,
		_w32024_
	);
	LUT4 #(
		.INIT('hc963)
	) name26198 (
		decrypt_pad,
		\u0_R2_reg[21]/NET0131 ,
		\u0_uk_K_r2_reg[28]/NET0131 ,
		\u0_uk_K_r2_reg[37]/NET0131 ,
		_w32025_
	);
	LUT4 #(
		.INIT('hc963)
	) name26199 (
		decrypt_pad,
		\u0_R2_reg[18]/NET0131 ,
		\u0_uk_K_r2_reg[1]/NET0131 ,
		\u0_uk_K_r2_reg[38]/NET0131 ,
		_w32026_
	);
	LUT3 #(
		.INIT('h04)
	) name26200 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32027_
	);
	LUT3 #(
		.INIT('h70)
	) name26201 (
		_w32026_,
		_w32023_,
		_w32025_,
		_w32028_
	);
	LUT4 #(
		.INIT('ha43f)
	) name26202 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32029_
	);
	LUT2 #(
		.INIT('h2)
	) name26203 (
		_w32022_,
		_w32029_,
		_w32030_
	);
	LUT2 #(
		.INIT('h1)
	) name26204 (
		_w32022_,
		_w32026_,
		_w32031_
	);
	LUT3 #(
		.INIT('hde)
	) name26205 (
		_w32024_,
		_w32023_,
		_w32025_,
		_w32032_
	);
	LUT2 #(
		.INIT('h2)
	) name26206 (
		_w32031_,
		_w32032_,
		_w32033_
	);
	LUT4 #(
		.INIT('h0020)
	) name26207 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32034_
	);
	LUT4 #(
		.INIT('h0040)
	) name26208 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32035_
	);
	LUT2 #(
		.INIT('h4)
	) name26209 (
		_w32022_,
		_w32024_,
		_w32036_
	);
	LUT3 #(
		.INIT('h8c)
	) name26210 (
		_w32022_,
		_w32026_,
		_w32024_,
		_w32037_
	);
	LUT4 #(
		.INIT('hb000)
	) name26211 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32038_
	);
	LUT4 #(
		.INIT('h0045)
	) name26212 (
		_w32035_,
		_w32037_,
		_w32038_,
		_w32034_,
		_w32039_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name26213 (
		_w32021_,
		_w32033_,
		_w32030_,
		_w32039_,
		_w32040_
	);
	LUT4 #(
		.INIT('h0010)
	) name26214 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32041_
	);
	LUT4 #(
		.INIT('hbc67)
	) name26215 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32042_
	);
	LUT4 #(
		.INIT('h5bf8)
	) name26216 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32043_
	);
	LUT4 #(
		.INIT('h2004)
	) name26217 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32044_
	);
	LUT4 #(
		.INIT('h00d8)
	) name26218 (
		_w32022_,
		_w32043_,
		_w32042_,
		_w32044_,
		_w32045_
	);
	LUT4 #(
		.INIT('h0208)
	) name26219 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32046_
	);
	LUT4 #(
		.INIT('hffbd)
	) name26220 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32047_
	);
	LUT3 #(
		.INIT('hb1)
	) name26221 (
		_w32022_,
		_w32046_,
		_w32047_,
		_w32048_
	);
	LUT3 #(
		.INIT('he0)
	) name26222 (
		_w32045_,
		_w32021_,
		_w32048_,
		_w32049_
	);
	LUT3 #(
		.INIT('h65)
	) name26223 (
		\u0_L2_reg[14]/NET0131 ,
		_w32040_,
		_w32049_,
		_w32050_
	);
	LUT4 #(
		.INIT('hbbfc)
	) name26224 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w32051_
	);
	LUT2 #(
		.INIT('h2)
	) name26225 (
		_w31827_,
		_w32051_,
		_w32052_
	);
	LUT3 #(
		.INIT('h47)
	) name26226 (
		_w31822_,
		_w31823_,
		_w31825_,
		_w32053_
	);
	LUT4 #(
		.INIT('h0010)
	) name26227 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w32054_
	);
	LUT4 #(
		.INIT('h0a02)
	) name26228 (
		_w31821_,
		_w31830_,
		_w32054_,
		_w32053_,
		_w32055_
	);
	LUT3 #(
		.INIT('h10)
	) name26229 (
		_w31832_,
		_w32052_,
		_w32055_,
		_w32056_
	);
	LUT3 #(
		.INIT('ha8)
	) name26230 (
		_w31823_,
		_w31824_,
		_w31827_,
		_w32057_
	);
	LUT2 #(
		.INIT('h8)
	) name26231 (
		_w31969_,
		_w32057_,
		_w32058_
	);
	LUT3 #(
		.INIT('hb0)
	) name26232 (
		_w31823_,
		_w31824_,
		_w31825_,
		_w32059_
	);
	LUT3 #(
		.INIT('h15)
	) name26233 (
		_w31821_,
		_w31974_,
		_w32059_,
		_w32060_
	);
	LUT3 #(
		.INIT('h10)
	) name26234 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w32061_
	);
	LUT4 #(
		.INIT('h0001)
	) name26235 (
		_w31827_,
		_w31845_,
		_w31976_,
		_w32061_,
		_w32062_
	);
	LUT3 #(
		.INIT('h40)
	) name26236 (
		_w32058_,
		_w32060_,
		_w32062_,
		_w32063_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name26237 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w32064_
	);
	LUT4 #(
		.INIT('h0929)
	) name26238 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w32065_
	);
	LUT2 #(
		.INIT('h2)
	) name26239 (
		_w31827_,
		_w32065_,
		_w32066_
	);
	LUT3 #(
		.INIT('h40)
	) name26240 (
		_w32058_,
		_w32060_,
		_w32066_,
		_w32067_
	);
	LUT4 #(
		.INIT('h001f)
	) name26241 (
		_w32056_,
		_w32063_,
		_w32064_,
		_w32067_,
		_w32068_
	);
	LUT2 #(
		.INIT('h9)
	) name26242 (
		\u0_L2_reg[13]/NET0131 ,
		_w32068_,
		_w32069_
	);
	LUT4 #(
		.INIT('h5b4b)
	) name26243 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32070_
	);
	LUT4 #(
		.INIT('h0002)
	) name26244 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32071_
	);
	LUT4 #(
		.INIT('h5504)
	) name26245 (
		_w31907_,
		_w31900_,
		_w32070_,
		_w32071_,
		_w32072_
	);
	LUT4 #(
		.INIT('h0004)
	) name26246 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32073_
	);
	LUT3 #(
		.INIT('h02)
	) name26247 (
		_w31900_,
		_w31928_,
		_w32073_,
		_w32074_
	);
	LUT4 #(
		.INIT('h0040)
	) name26248 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32075_
	);
	LUT4 #(
		.INIT('h0c04)
	) name26249 (
		_w31907_,
		_w31901_,
		_w31905_,
		_w31902_,
		_w32076_
	);
	LUT4 #(
		.INIT('h0001)
	) name26250 (
		_w31900_,
		_w31909_,
		_w32075_,
		_w32076_,
		_w32077_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name26251 (
		_w31900_,
		_w31901_,
		_w31904_,
		_w31902_,
		_w32078_
	);
	LUT3 #(
		.INIT('h0e)
	) name26252 (
		_w31900_,
		_w31904_,
		_w31905_,
		_w32079_
	);
	LUT4 #(
		.INIT('h0800)
	) name26253 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32080_
	);
	LUT4 #(
		.INIT('he75f)
	) name26254 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32081_
	);
	LUT4 #(
		.INIT('h20aa)
	) name26255 (
		_w31907_,
		_w32078_,
		_w32079_,
		_w32081_,
		_w32082_
	);
	LUT4 #(
		.INIT('h00dc)
	) name26256 (
		_w31914_,
		_w32074_,
		_w32077_,
		_w32082_,
		_w32083_
	);
	LUT3 #(
		.INIT('h65)
	) name26257 (
		\u0_L2_reg[15]/P0001 ,
		_w32072_,
		_w32083_,
		_w32084_
	);
	LUT4 #(
		.INIT('h5551)
	) name26258 (
		_w31900_,
		_w31901_,
		_w31904_,
		_w31902_,
		_w32085_
	);
	LUT4 #(
		.INIT('he040)
	) name26259 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32086_
	);
	LUT4 #(
		.INIT('haaa2)
	) name26260 (
		_w31900_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32087_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name26261 (
		_w32080_,
		_w32085_,
		_w32086_,
		_w32087_,
		_w32088_
	);
	LUT4 #(
		.INIT('h2100)
	) name26262 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32089_
	);
	LUT3 #(
		.INIT('h02)
	) name26263 (
		_w31907_,
		_w32073_,
		_w32089_,
		_w32090_
	);
	LUT2 #(
		.INIT('h4)
	) name26264 (
		_w32088_,
		_w32090_,
		_w32091_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name26265 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32092_
	);
	LUT4 #(
		.INIT('h0040)
	) name26266 (
		_w31900_,
		_w31901_,
		_w31904_,
		_w31902_,
		_w32093_
	);
	LUT4 #(
		.INIT('h0888)
	) name26267 (
		_w31900_,
		_w31901_,
		_w31904_,
		_w31905_,
		_w32094_
	);
	LUT4 #(
		.INIT('h2300)
	) name26268 (
		_w31910_,
		_w32093_,
		_w32094_,
		_w32092_,
		_w32095_
	);
	LUT4 #(
		.INIT('hccef)
	) name26269 (
		_w31900_,
		_w31901_,
		_w31904_,
		_w31905_,
		_w32096_
	);
	LUT2 #(
		.INIT('h2)
	) name26270 (
		_w31902_,
		_w32096_,
		_w32097_
	);
	LUT4 #(
		.INIT('h0080)
	) name26271 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32098_
	);
	LUT4 #(
		.INIT('h0100)
	) name26272 (
		_w31900_,
		_w31901_,
		_w31904_,
		_w31905_,
		_w32099_
	);
	LUT3 #(
		.INIT('h01)
	) name26273 (
		_w31907_,
		_w32099_,
		_w32098_,
		_w32100_
	);
	LUT3 #(
		.INIT('h40)
	) name26274 (
		_w32097_,
		_w32100_,
		_w32095_,
		_w32101_
	);
	LUT4 #(
		.INIT('h0002)
	) name26275 (
		_w31900_,
		_w31901_,
		_w31905_,
		_w31902_,
		_w32102_
	);
	LUT3 #(
		.INIT('h0b)
	) name26276 (
		_w31900_,
		_w32098_,
		_w32102_,
		_w32103_
	);
	LUT4 #(
		.INIT('ha955)
	) name26277 (
		\u0_L2_reg[21]/NET0131 ,
		_w32091_,
		_w32101_,
		_w32103_,
		_w32104_
	);
	LUT3 #(
		.INIT('had)
	) name26278 (
		_w31731_,
		_w31734_,
		_w31732_,
		_w32105_
	);
	LUT4 #(
		.INIT('hfcd3)
	) name26279 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w32106_
	);
	LUT2 #(
		.INIT('h1)
	) name26280 (
		_w31730_,
		_w32106_,
		_w32107_
	);
	LUT2 #(
		.INIT('h4)
	) name26281 (
		_w31737_,
		_w31745_,
		_w32108_
	);
	LUT3 #(
		.INIT('h07)
	) name26282 (
		_w31754_,
		_w31755_,
		_w31857_,
		_w32109_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name26283 (
		_w31729_,
		_w32107_,
		_w32108_,
		_w32109_,
		_w32110_
	);
	LUT4 #(
		.INIT('h5f57)
	) name26284 (
		_w31733_,
		_w31730_,
		_w31731_,
		_w31734_,
		_w32111_
	);
	LUT2 #(
		.INIT('h2)
	) name26285 (
		_w31732_,
		_w32111_,
		_w32112_
	);
	LUT4 #(
		.INIT('h5040)
	) name26286 (
		_w31730_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w32113_
	);
	LUT3 #(
		.INIT('h01)
	) name26287 (
		_w31733_,
		_w31731_,
		_w31732_,
		_w32114_
	);
	LUT4 #(
		.INIT('h0008)
	) name26288 (
		_w31730_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w32115_
	);
	LUT4 #(
		.INIT('h0203)
	) name26289 (
		_w31856_,
		_w32114_,
		_w32115_,
		_w32113_,
		_w32116_
	);
	LUT3 #(
		.INIT('hb9)
	) name26290 (
		_w31731_,
		_w31734_,
		_w31732_,
		_w32117_
	);
	LUT4 #(
		.INIT('h7ebf)
	) name26291 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w32118_
	);
	LUT4 #(
		.INIT('hfbc8)
	) name26292 (
		_w31733_,
		_w31730_,
		_w32117_,
		_w32118_,
		_w32119_
	);
	LUT4 #(
		.INIT('hba00)
	) name26293 (
		_w31729_,
		_w32112_,
		_w32116_,
		_w32119_,
		_w32120_
	);
	LUT3 #(
		.INIT('h9a)
	) name26294 (
		\u0_L2_reg[23]/NET0131 ,
		_w32110_,
		_w32120_,
		_w32121_
	);
	LUT4 #(
		.INIT('hce00)
	) name26295 (
		_w31762_,
		_w31763_,
		_w31764_,
		_w31760_,
		_w32122_
	);
	LUT4 #(
		.INIT('h0021)
	) name26296 (
		_w31762_,
		_w31763_,
		_w31764_,
		_w31760_,
		_w32123_
	);
	LUT4 #(
		.INIT('h8000)
	) name26297 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w32124_
	);
	LUT4 #(
		.INIT('h0203)
	) name26298 (
		_w31775_,
		_w32123_,
		_w32124_,
		_w32122_,
		_w32125_
	);
	LUT2 #(
		.INIT('h1)
	) name26299 (
		_w31759_,
		_w32125_,
		_w32126_
	);
	LUT4 #(
		.INIT('h0104)
	) name26300 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w32127_
	);
	LUT3 #(
		.INIT('h04)
	) name26301 (
		_w31762_,
		_w31763_,
		_w31760_,
		_w32128_
	);
	LUT3 #(
		.INIT('h01)
	) name26302 (
		_w31782_,
		_w31889_,
		_w32128_,
		_w32129_
	);
	LUT4 #(
		.INIT('h2000)
	) name26303 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31760_,
		_w32130_
	);
	LUT4 #(
		.INIT('h0800)
	) name26304 (
		_w31762_,
		_w31761_,
		_w31763_,
		_w31764_,
		_w32131_
	);
	LUT2 #(
		.INIT('h1)
	) name26305 (
		_w32130_,
		_w32131_,
		_w32132_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name26306 (
		_w31759_,
		_w32127_,
		_w32129_,
		_w32132_,
		_w32133_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name26307 (
		_w31762_,
		_w31761_,
		_w31785_,
		_w31769_,
		_w32134_
	);
	LUT4 #(
		.INIT('h5655)
	) name26308 (
		\u0_L2_reg[19]/P0001 ,
		_w32133_,
		_w32126_,
		_w32134_,
		_w32135_
	);
	LUT4 #(
		.INIT('h4555)
	) name26309 (
		_w32022_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32136_
	);
	LUT4 #(
		.INIT('h001b)
	) name26310 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32137_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name26311 (
		_w32022_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32138_
	);
	LUT4 #(
		.INIT('h28a8)
	) name26312 (
		_w32022_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32139_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name26313 (
		_w32027_,
		_w32136_,
		_w32137_,
		_w32139_,
		_w32140_
	);
	LUT4 #(
		.INIT('hbb7f)
	) name26314 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32141_
	);
	LUT3 #(
		.INIT('h8a)
	) name26315 (
		_w32021_,
		_w32140_,
		_w32141_,
		_w32142_
	);
	LUT3 #(
		.INIT('ha2)
	) name26316 (
		_w32022_,
		_w32024_,
		_w32025_,
		_w32143_
	);
	LUT4 #(
		.INIT('h2223)
	) name26317 (
		_w32022_,
		_w32026_,
		_w32024_,
		_w32023_,
		_w32144_
	);
	LUT2 #(
		.INIT('h4)
	) name26318 (
		_w32143_,
		_w32144_,
		_w32145_
	);
	LUT4 #(
		.INIT('h0800)
	) name26319 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32146_
	);
	LUT4 #(
		.INIT('hf7c7)
	) name26320 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32147_
	);
	LUT3 #(
		.INIT('h32)
	) name26321 (
		_w32022_,
		_w32146_,
		_w32147_,
		_w32148_
	);
	LUT4 #(
		.INIT('hff7d)
	) name26322 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32149_
	);
	LUT4 #(
		.INIT('hfe7d)
	) name26323 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32150_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name26324 (
		_w32022_,
		_w32026_,
		_w32024_,
		_w32025_,
		_w32151_
	);
	LUT4 #(
		.INIT('hf531)
	) name26325 (
		_w32022_,
		_w32023_,
		_w32150_,
		_w32151_,
		_w32152_
	);
	LUT4 #(
		.INIT('hba00)
	) name26326 (
		_w32021_,
		_w32145_,
		_w32148_,
		_w32152_,
		_w32153_
	);
	LUT3 #(
		.INIT('h65)
	) name26327 (
		\u0_L2_reg[25]/NET0131 ,
		_w32142_,
		_w32153_,
		_w32154_
	);
	LUT4 #(
		.INIT('h0002)
	) name26328 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32155_
	);
	LUT3 #(
		.INIT('h01)
	) name26329 (
		_w31941_,
		_w31986_,
		_w32155_,
		_w32156_
	);
	LUT4 #(
		.INIT('h3fef)
	) name26330 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32157_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name26331 (
		_w31935_,
		_w31936_,
		_w31934_,
		_w31940_,
		_w32158_
	);
	LUT4 #(
		.INIT('hfa32)
	) name26332 (
		_w31935_,
		_w31937_,
		_w32157_,
		_w32158_,
		_w32159_
	);
	LUT3 #(
		.INIT('h2a)
	) name26333 (
		_w31933_,
		_w32156_,
		_w32159_,
		_w32160_
	);
	LUT4 #(
		.INIT('heafa)
	) name26334 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32161_
	);
	LUT4 #(
		.INIT('h0086)
	) name26335 (
		_w31936_,
		_w31934_,
		_w31940_,
		_w31937_,
		_w32162_
	);
	LUT4 #(
		.INIT('h3301)
	) name26336 (
		_w31933_,
		_w31935_,
		_w32161_,
		_w32162_,
		_w32163_
	);
	LUT3 #(
		.INIT('h45)
	) name26337 (
		_w31950_,
		_w31959_,
		_w31938_,
		_w32164_
	);
	LUT2 #(
		.INIT('h8)
	) name26338 (
		_w31935_,
		_w31940_,
		_w32165_
	);
	LUT2 #(
		.INIT('h4)
	) name26339 (
		_w31951_,
		_w32165_,
		_w32166_
	);
	LUT4 #(
		.INIT('h00ea)
	) name26340 (
		_w31933_,
		_w31957_,
		_w32164_,
		_w32166_,
		_w32167_
	);
	LUT4 #(
		.INIT('h5655)
	) name26341 (
		\u0_L2_reg[26]/NET0131 ,
		_w32160_,
		_w32163_,
		_w32167_,
		_w32168_
	);
	LUT4 #(
		.INIT('h0200)
	) name26342 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32169_
	);
	LUT4 #(
		.INIT('hfb77)
	) name26343 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32170_
	);
	LUT4 #(
		.INIT('he4ee)
	) name26344 (
		_w32022_,
		_w32034_,
		_w32169_,
		_w32170_,
		_w32171_
	);
	LUT4 #(
		.INIT('hcffe)
	) name26345 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32172_
	);
	LUT4 #(
		.INIT('hef00)
	) name26346 (
		_w32022_,
		_w32026_,
		_w32023_,
		_w32021_,
		_w32173_
	);
	LUT4 #(
		.INIT('h3100)
	) name26347 (
		_w32022_,
		_w32046_,
		_w32172_,
		_w32173_,
		_w32174_
	);
	LUT4 #(
		.INIT('h0d00)
	) name26348 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32175_
	);
	LUT4 #(
		.INIT('haf23)
	) name26349 (
		_w32041_,
		_w32136_,
		_w32138_,
		_w32175_,
		_w32176_
	);
	LUT4 #(
		.INIT('h00fb)
	) name26350 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32021_,
		_w32177_
	);
	LUT2 #(
		.INIT('h8)
	) name26351 (
		_w32149_,
		_w32177_,
		_w32178_
	);
	LUT4 #(
		.INIT('h4544)
	) name26352 (
		_w32171_,
		_w32174_,
		_w32176_,
		_w32178_,
		_w32179_
	);
	LUT2 #(
		.INIT('h9)
	) name26353 (
		\u0_L2_reg[8]/NET0131 ,
		_w32179_,
		_w32180_
	);
	LUT4 #(
		.INIT('h3f3e)
	) name26354 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32181_
	);
	LUT2 #(
		.INIT('h2)
	) name26355 (
		_w31803_,
		_w32181_,
		_w32182_
	);
	LUT3 #(
		.INIT('h04)
	) name26356 (
		_w31799_,
		_w31801_,
		_w31812_,
		_w32183_
	);
	LUT4 #(
		.INIT('h0400)
	) name26357 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32184_
	);
	LUT2 #(
		.INIT('h6)
	) name26358 (
		_w31795_,
		_w31796_,
		_w32185_
	);
	LUT4 #(
		.INIT('h2022)
	) name26359 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31803_,
		_w32186_
	);
	LUT3 #(
		.INIT('h15)
	) name26360 (
		_w32184_,
		_w32185_,
		_w32186_,
		_w32187_
	);
	LUT3 #(
		.INIT('h40)
	) name26361 (
		_w32182_,
		_w32183_,
		_w32187_,
		_w32188_
	);
	LUT3 #(
		.INIT('h47)
	) name26362 (
		_w31793_,
		_w31794_,
		_w31803_,
		_w32189_
	);
	LUT4 #(
		.INIT('h0006)
	) name26363 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32190_
	);
	LUT4 #(
		.INIT('h0301)
	) name26364 (
		_w31797_,
		_w31801_,
		_w32190_,
		_w32189_,
		_w32191_
	);
	LUT2 #(
		.INIT('h6)
	) name26365 (
		_w31794_,
		_w31796_,
		_w32192_
	);
	LUT4 #(
		.INIT('h134c)
	) name26366 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32193_
	);
	LUT3 #(
		.INIT('h04)
	) name26367 (
		_w31793_,
		_w31795_,
		_w31796_,
		_w32194_
	);
	LUT4 #(
		.INIT('h2010)
	) name26368 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32195_
	);
	LUT3 #(
		.INIT('h0e)
	) name26369 (
		_w31803_,
		_w32193_,
		_w32195_,
		_w32196_
	);
	LUT2 #(
		.INIT('h8)
	) name26370 (
		_w32191_,
		_w32196_,
		_w32197_
	);
	LUT3 #(
		.INIT('ha9)
	) name26371 (
		\u0_L2_reg[12]/NET0131 ,
		_w32188_,
		_w32197_,
		_w32198_
	);
	LUT4 #(
		.INIT('hc693)
	) name26372 (
		decrypt_pad,
		\u0_R2_reg[13]/NET0131 ,
		\u0_uk_K_r2_reg[20]/NET0131 ,
		\u0_uk_K_r2_reg[40]/NET0131 ,
		_w32199_
	);
	LUT4 #(
		.INIT('hc963)
	) name26373 (
		decrypt_pad,
		\u0_R2_reg[10]/NET0131 ,
		\u0_uk_K_r2_reg[11]/NET0131 ,
		\u0_uk_K_r2_reg[48]/NET0131 ,
		_w32200_
	);
	LUT4 #(
		.INIT('hc693)
	) name26374 (
		decrypt_pad,
		\u0_R2_reg[8]/NET0131 ,
		\u0_uk_K_r2_reg[11]/NET0131 ,
		\u0_uk_K_r2_reg[6]/NET0131 ,
		_w32201_
	);
	LUT4 #(
		.INIT('hc963)
	) name26375 (
		decrypt_pad,
		\u0_R2_reg[9]/NET0131 ,
		\u0_uk_K_r2_reg[3]/NET0131 ,
		\u0_uk_K_r2_reg[40]/NET0131 ,
		_w32202_
	);
	LUT4 #(
		.INIT('h0010)
	) name26376 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32203_
	);
	LUT2 #(
		.INIT('h2)
	) name26377 (
		_w32199_,
		_w32201_,
		_w32204_
	);
	LUT4 #(
		.INIT('hc963)
	) name26378 (
		decrypt_pad,
		\u0_R2_reg[11]/NET0131 ,
		\u0_uk_K_r2_reg[12]/NET0131 ,
		\u0_uk_K_r2_reg[17]/NET0131 ,
		_w32205_
	);
	LUT3 #(
		.INIT('h01)
	) name26379 (
		_w32200_,
		_w32202_,
		_w32205_,
		_w32206_
	);
	LUT3 #(
		.INIT('h15)
	) name26380 (
		_w32203_,
		_w32204_,
		_w32206_,
		_w32207_
	);
	LUT4 #(
		.INIT('h4000)
	) name26381 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32208_
	);
	LUT4 #(
		.INIT('hc963)
	) name26382 (
		decrypt_pad,
		\u0_R2_reg[12]/NET0131 ,
		\u0_uk_K_r2_reg[27]/P0001 ,
		\u0_uk_K_r2_reg[32]/NET0131 ,
		_w32209_
	);
	LUT2 #(
		.INIT('h1)
	) name26383 (
		_w32208_,
		_w32209_,
		_w32210_
	);
	LUT2 #(
		.INIT('h4)
	) name26384 (
		_w32200_,
		_w32205_,
		_w32211_
	);
	LUT2 #(
		.INIT('h2)
	) name26385 (
		_w32200_,
		_w32205_,
		_w32212_
	);
	LUT3 #(
		.INIT('hc7)
	) name26386 (
		_w32199_,
		_w32200_,
		_w32205_,
		_w32213_
	);
	LUT2 #(
		.INIT('h4)
	) name26387 (
		_w32201_,
		_w32202_,
		_w32214_
	);
	LUT2 #(
		.INIT('h8)
	) name26388 (
		_w32199_,
		_w32201_,
		_w32215_
	);
	LUT4 #(
		.INIT('ha584)
	) name26389 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32216_
	);
	LUT4 #(
		.INIT('h2184)
	) name26390 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32217_
	);
	LUT3 #(
		.INIT('h0b)
	) name26391 (
		_w32213_,
		_w32214_,
		_w32217_,
		_w32218_
	);
	LUT4 #(
		.INIT('ha251)
	) name26392 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32219_
	);
	LUT3 #(
		.INIT('h0e)
	) name26393 (
		_w32201_,
		_w32202_,
		_w32205_,
		_w32220_
	);
	LUT4 #(
		.INIT('h0400)
	) name26394 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32221_
	);
	LUT4 #(
		.INIT('h0222)
	) name26395 (
		_w32209_,
		_w32221_,
		_w32219_,
		_w32220_,
		_w32222_
	);
	LUT4 #(
		.INIT('h007f)
	) name26396 (
		_w32207_,
		_w32210_,
		_w32218_,
		_w32222_,
		_w32223_
	);
	LUT3 #(
		.INIT('he0)
	) name26397 (
		_w32199_,
		_w32201_,
		_w32209_,
		_w32224_
	);
	LUT4 #(
		.INIT('h0001)
	) name26398 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32225_
	);
	LUT4 #(
		.INIT('hff76)
	) name26399 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32226_
	);
	LUT4 #(
		.INIT('h20aa)
	) name26400 (
		_w32205_,
		_w32219_,
		_w32224_,
		_w32226_,
		_w32227_
	);
	LUT3 #(
		.INIT('h56)
	) name26401 (
		\u0_L2_reg[6]/NET0131 ,
		_w32223_,
		_w32227_,
		_w32228_
	);
	LUT4 #(
		.INIT('h8090)
	) name26402 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32229_
	);
	LUT3 #(
		.INIT('h60)
	) name26403 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w32230_
	);
	LUT4 #(
		.INIT('hf5e4)
	) name26404 (
		_w31900_,
		_w31913_,
		_w32229_,
		_w32230_,
		_w32231_
	);
	LUT4 #(
		.INIT('hbdf3)
	) name26405 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32232_
	);
	LUT3 #(
		.INIT('h8a)
	) name26406 (
		_w31907_,
		_w32231_,
		_w32232_,
		_w32233_
	);
	LUT4 #(
		.INIT('hdc0c)
	) name26407 (
		_w31901_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32234_
	);
	LUT4 #(
		.INIT('haa8a)
	) name26408 (
		_w31900_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32235_
	);
	LUT4 #(
		.INIT('h4544)
	) name26409 (
		_w31907_,
		_w31912_,
		_w32234_,
		_w32235_,
		_w32236_
	);
	LUT2 #(
		.INIT('h1)
	) name26410 (
		_w31900_,
		_w31911_,
		_w32237_
	);
	LUT4 #(
		.INIT('h4000)
	) name26411 (
		_w31900_,
		_w31901_,
		_w31904_,
		_w31902_,
		_w32238_
	);
	LUT3 #(
		.INIT('h54)
	) name26412 (
		_w31907_,
		_w32099_,
		_w32238_,
		_w32239_
	);
	LUT4 #(
		.INIT('h0200)
	) name26413 (
		_w31900_,
		_w31904_,
		_w31905_,
		_w31902_,
		_w32240_
	);
	LUT3 #(
		.INIT('h0b)
	) name26414 (
		_w31900_,
		_w31908_,
		_w32240_,
		_w32241_
	);
	LUT4 #(
		.INIT('h0100)
	) name26415 (
		_w32236_,
		_w32237_,
		_w32239_,
		_w32241_,
		_w32242_
	);
	LUT3 #(
		.INIT('h65)
	) name26416 (
		\u0_L2_reg[27]/NET0131 ,
		_w32233_,
		_w32242_,
		_w32243_
	);
	LUT4 #(
		.INIT('haff3)
	) name26417 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32244_
	);
	LUT2 #(
		.INIT('h2)
	) name26418 (
		_w32022_,
		_w32244_,
		_w32245_
	);
	LUT3 #(
		.INIT('h07)
	) name26419 (
		_w32028_,
		_w32036_,
		_w32034_,
		_w32246_
	);
	LUT3 #(
		.INIT('h8a)
	) name26420 (
		_w32021_,
		_w32245_,
		_w32246_,
		_w32247_
	);
	LUT4 #(
		.INIT('h45f0)
	) name26421 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32248_
	);
	LUT2 #(
		.INIT('h1)
	) name26422 (
		_w32021_,
		_w32248_,
		_w32249_
	);
	LUT4 #(
		.INIT('hffbe)
	) name26423 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32250_
	);
	LUT3 #(
		.INIT('he0)
	) name26424 (
		_w32031_,
		_w32136_,
		_w32250_,
		_w32251_
	);
	LUT4 #(
		.INIT('hd83d)
	) name26425 (
		_w32026_,
		_w32024_,
		_w32023_,
		_w32025_,
		_w32252_
	);
	LUT2 #(
		.INIT('h1)
	) name26426 (
		_w32021_,
		_w32252_,
		_w32253_
	);
	LUT3 #(
		.INIT('h02)
	) name26427 (
		_w32022_,
		_w32041_,
		_w32169_,
		_w32254_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name26428 (
		_w32249_,
		_w32251_,
		_w32253_,
		_w32254_,
		_w32255_
	);
	LUT3 #(
		.INIT('h56)
	) name26429 (
		\u0_L2_reg[3]/NET0131 ,
		_w32247_,
		_w32255_,
		_w32256_
	);
	LUT4 #(
		.INIT('h8228)
	) name26430 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w32257_
	);
	LUT3 #(
		.INIT('hda)
	) name26431 (
		_w31731_,
		_w31734_,
		_w31732_,
		_w32258_
	);
	LUT4 #(
		.INIT('h0031)
	) name26432 (
		_w31741_,
		_w31860_,
		_w32258_,
		_w32257_,
		_w32259_
	);
	LUT4 #(
		.INIT('h1555)
	) name26433 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w32260_
	);
	LUT4 #(
		.INIT('h6002)
	) name26434 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w32261_
	);
	LUT4 #(
		.INIT('h5144)
	) name26435 (
		_w31730_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w32262_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name26436 (
		_w31733_,
		_w31730_,
		_w31731_,
		_w31732_,
		_w32263_
	);
	LUT4 #(
		.INIT('h3230)
	) name26437 (
		_w32105_,
		_w32261_,
		_w32262_,
		_w32263_,
		_w32264_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name26438 (
		_w31733_,
		_w31731_,
		_w31734_,
		_w31732_,
		_w32265_
	);
	LUT3 #(
		.INIT('h01)
	) name26439 (
		_w31730_,
		_w32260_,
		_w32265_,
		_w32266_
	);
	LUT4 #(
		.INIT('h00e4)
	) name26440 (
		_w31729_,
		_w32264_,
		_w32259_,
		_w32266_,
		_w32267_
	);
	LUT2 #(
		.INIT('h9)
	) name26441 (
		\u0_L2_reg[9]/NET0131 ,
		_w32267_,
		_w32268_
	);
	LUT3 #(
		.INIT('h41)
	) name26442 (
		_w31793_,
		_w31795_,
		_w31796_,
		_w32269_
	);
	LUT4 #(
		.INIT('h5004)
	) name26443 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32270_
	);
	LUT2 #(
		.INIT('h2)
	) name26444 (
		_w31803_,
		_w32270_,
		_w32271_
	);
	LUT3 #(
		.INIT('h09)
	) name26445 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w32272_
	);
	LUT3 #(
		.INIT('h28)
	) name26446 (
		_w31794_,
		_w31795_,
		_w31796_,
		_w32273_
	);
	LUT4 #(
		.INIT('h00f7)
	) name26447 (
		_w31793_,
		_w31795_,
		_w31796_,
		_w31803_,
		_w32274_
	);
	LUT3 #(
		.INIT('h10)
	) name26448 (
		_w32273_,
		_w32272_,
		_w32274_,
		_w32275_
	);
	LUT3 #(
		.INIT('h40)
	) name26449 (
		_w31794_,
		_w31795_,
		_w31796_,
		_w32276_
	);
	LUT4 #(
		.INIT('h2880)
	) name26450 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32277_
	);
	LUT2 #(
		.INIT('h2)
	) name26451 (
		_w31801_,
		_w32277_,
		_w32278_
	);
	LUT4 #(
		.INIT('h0880)
	) name26452 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32279_
	);
	LUT4 #(
		.INIT('hbf00)
	) name26453 (
		_w31794_,
		_w31795_,
		_w31796_,
		_w31803_,
		_w32280_
	);
	LUT4 #(
		.INIT('h5545)
	) name26454 (
		_w31801_,
		_w32269_,
		_w32280_,
		_w32279_,
		_w32281_
	);
	LUT4 #(
		.INIT('h001f)
	) name26455 (
		_w32271_,
		_w32275_,
		_w32278_,
		_w32281_,
		_w32282_
	);
	LUT2 #(
		.INIT('h4)
	) name26456 (
		_w31803_,
		_w32277_,
		_w32283_
	);
	LUT2 #(
		.INIT('h2)
	) name26457 (
		_w31801_,
		_w31803_,
		_w32284_
	);
	LUT4 #(
		.INIT('h00dc)
	) name26458 (
		_w31803_,
		_w31807_,
		_w32270_,
		_w32284_,
		_w32285_
	);
	LUT2 #(
		.INIT('h1)
	) name26459 (
		_w32283_,
		_w32285_,
		_w32286_
	);
	LUT3 #(
		.INIT('h65)
	) name26460 (
		\u0_L2_reg[7]/NET0131 ,
		_w32282_,
		_w32286_,
		_w32287_
	);
	LUT4 #(
		.INIT('h2110)
	) name26461 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32288_
	);
	LUT4 #(
		.INIT('h00fd)
	) name26462 (
		_w31794_,
		_w31795_,
		_w31796_,
		_w31803_,
		_w32289_
	);
	LUT4 #(
		.INIT('hbf00)
	) name26463 (
		_w31793_,
		_w31794_,
		_w31796_,
		_w31803_,
		_w32290_
	);
	LUT4 #(
		.INIT('hff5c)
	) name26464 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32291_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name26465 (
		_w32288_,
		_w32289_,
		_w32290_,
		_w32291_,
		_w32292_
	);
	LUT4 #(
		.INIT('h0080)
	) name26466 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32293_
	);
	LUT3 #(
		.INIT('ha8)
	) name26467 (
		_w31801_,
		_w32292_,
		_w32293_,
		_w32294_
	);
	LUT4 #(
		.INIT('haba1)
	) name26468 (
		_w31803_,
		_w32192_,
		_w32194_,
		_w32276_,
		_w32295_
	);
	LUT4 #(
		.INIT('h7db7)
	) name26469 (
		_w31793_,
		_w31794_,
		_w31795_,
		_w31796_,
		_w32296_
	);
	LUT4 #(
		.INIT('h00a2)
	) name26470 (
		_w31794_,
		_w31795_,
		_w31796_,
		_w31803_,
		_w32297_
	);
	LUT4 #(
		.INIT('h0777)
	) name26471 (
		_w31798_,
		_w31803_,
		_w31808_,
		_w32297_,
		_w32298_
	);
	LUT4 #(
		.INIT('hba00)
	) name26472 (
		_w31801_,
		_w32295_,
		_w32296_,
		_w32298_,
		_w32299_
	);
	LUT3 #(
		.INIT('h65)
	) name26473 (
		\u0_L2_reg[32]/NET0131 ,
		_w32294_,
		_w32299_,
		_w32300_
	);
	LUT4 #(
		.INIT('h0021)
	) name26474 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32301_
	);
	LUT3 #(
		.INIT('h08)
	) name26475 (
		_w32200_,
		_w32201_,
		_w32202_,
		_w32302_
	);
	LUT4 #(
		.INIT('ha7b7)
	) name26476 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32303_
	);
	LUT3 #(
		.INIT('h10)
	) name26477 (
		_w32205_,
		_w32301_,
		_w32303_,
		_w32304_
	);
	LUT3 #(
		.INIT('hf9)
	) name26478 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32305_
	);
	LUT3 #(
		.INIT('h10)
	) name26479 (
		_w32199_,
		_w32201_,
		_w32202_,
		_w32306_
	);
	LUT4 #(
		.INIT('hf700)
	) name26480 (
		_w32200_,
		_w32201_,
		_w32202_,
		_w32205_,
		_w32307_
	);
	LUT3 #(
		.INIT('h20)
	) name26481 (
		_w32305_,
		_w32306_,
		_w32307_,
		_w32308_
	);
	LUT3 #(
		.INIT('h54)
	) name26482 (
		_w32209_,
		_w32304_,
		_w32308_,
		_w32309_
	);
	LUT3 #(
		.INIT('h0d)
	) name26483 (
		_w32199_,
		_w32201_,
		_w32202_,
		_w32310_
	);
	LUT3 #(
		.INIT('h4c)
	) name26484 (
		_w32211_,
		_w32209_,
		_w32310_,
		_w32311_
	);
	LUT4 #(
		.INIT('h37f7)
	) name26485 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32312_
	);
	LUT3 #(
		.INIT('hb1)
	) name26486 (
		_w32205_,
		_w32216_,
		_w32312_,
		_w32313_
	);
	LUT3 #(
		.INIT('h80)
	) name26487 (
		_w32207_,
		_w32311_,
		_w32313_,
		_w32314_
	);
	LUT3 #(
		.INIT('h80)
	) name26488 (
		_w32199_,
		_w32201_,
		_w32202_,
		_w32315_
	);
	LUT3 #(
		.INIT('hac)
	) name26489 (
		_w32199_,
		_w32201_,
		_w32202_,
		_w32316_
	);
	LUT4 #(
		.INIT('h1300)
	) name26490 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32205_,
		_w32317_
	);
	LUT4 #(
		.INIT('h0777)
	) name26491 (
		_w32212_,
		_w32315_,
		_w32316_,
		_w32317_,
		_w32318_
	);
	LUT4 #(
		.INIT('ha955)
	) name26492 (
		\u0_L2_reg[24]/NET0131 ,
		_w32309_,
		_w32314_,
		_w32318_,
		_w32319_
	);
	LUT4 #(
		.INIT('h6979)
	) name26493 (
		_w32199_,
		_w32201_,
		_w32202_,
		_w32205_,
		_w32320_
	);
	LUT2 #(
		.INIT('h1)
	) name26494 (
		_w32200_,
		_w32320_,
		_w32321_
	);
	LUT4 #(
		.INIT('h0014)
	) name26495 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32205_,
		_w32322_
	);
	LUT4 #(
		.INIT('h0800)
	) name26496 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32323_
	);
	LUT3 #(
		.INIT('h02)
	) name26497 (
		_w32209_,
		_w32323_,
		_w32322_,
		_w32324_
	);
	LUT4 #(
		.INIT('h5ef4)
	) name26498 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32325_
	);
	LUT2 #(
		.INIT('h1)
	) name26499 (
		_w32205_,
		_w32325_,
		_w32326_
	);
	LUT4 #(
		.INIT('h6800)
	) name26500 (
		_w32199_,
		_w32201_,
		_w32202_,
		_w32205_,
		_w32327_
	);
	LUT3 #(
		.INIT('h01)
	) name26501 (
		_w32209_,
		_w32225_,
		_w32327_,
		_w32328_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name26502 (
		_w32321_,
		_w32324_,
		_w32326_,
		_w32328_,
		_w32329_
	);
	LUT4 #(
		.INIT('h0008)
	) name26503 (
		_w32200_,
		_w32201_,
		_w32202_,
		_w32205_,
		_w32330_
	);
	LUT4 #(
		.INIT('hbffb)
	) name26504 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32331_
	);
	LUT3 #(
		.INIT('h31)
	) name26505 (
		_w32205_,
		_w32330_,
		_w32331_,
		_w32332_
	);
	LUT3 #(
		.INIT('h65)
	) name26506 (
		\u0_L2_reg[16]/NET0131 ,
		_w32329_,
		_w32332_,
		_w32333_
	);
	LUT3 #(
		.INIT('h07)
	) name26507 (
		_w32200_,
		_w32201_,
		_w32205_,
		_w32334_
	);
	LUT2 #(
		.INIT('h4)
	) name26508 (
		_w32306_,
		_w32334_,
		_w32335_
	);
	LUT3 #(
		.INIT('h40)
	) name26509 (
		_w32203_,
		_w32205_,
		_w32305_,
		_w32336_
	);
	LUT3 #(
		.INIT('ha8)
	) name26510 (
		_w32209_,
		_w32335_,
		_w32336_,
		_w32337_
	);
	LUT4 #(
		.INIT('h6e3f)
	) name26511 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32338_
	);
	LUT2 #(
		.INIT('h2)
	) name26512 (
		_w32205_,
		_w32338_,
		_w32339_
	);
	LUT2 #(
		.INIT('h8)
	) name26513 (
		_w32316_,
		_w32334_,
		_w32340_
	);
	LUT4 #(
		.INIT('h0008)
	) name26514 (
		_w32199_,
		_w32200_,
		_w32201_,
		_w32202_,
		_w32341_
	);
	LUT3 #(
		.INIT('h01)
	) name26515 (
		_w32209_,
		_w32301_,
		_w32341_,
		_w32342_
	);
	LUT3 #(
		.INIT('h10)
	) name26516 (
		_w32340_,
		_w32339_,
		_w32342_,
		_w32343_
	);
	LUT2 #(
		.INIT('h8)
	) name26517 (
		_w32199_,
		_w32205_,
		_w32344_
	);
	LUT2 #(
		.INIT('h8)
	) name26518 (
		_w32302_,
		_w32344_,
		_w32345_
	);
	LUT4 #(
		.INIT('h0040)
	) name26519 (
		_w32199_,
		_w32200_,
		_w32202_,
		_w32205_,
		_w32346_
	);
	LUT3 #(
		.INIT('h80)
	) name26520 (
		_w32200_,
		_w32202_,
		_w32209_,
		_w32347_
	);
	LUT3 #(
		.INIT('h23)
	) name26521 (
		_w32215_,
		_w32346_,
		_w32347_,
		_w32348_
	);
	LUT2 #(
		.INIT('h4)
	) name26522 (
		_w32345_,
		_w32348_,
		_w32349_
	);
	LUT4 #(
		.INIT('h56aa)
	) name26523 (
		\u0_L2_reg[30]/NET0131 ,
		_w32337_,
		_w32343_,
		_w32349_,
		_w32350_
	);
	LUT3 #(
		.INIT('h1b)
	) name26524 (
		_w31824_,
		_w31825_,
		_w31827_,
		_w32351_
	);
	LUT3 #(
		.INIT('h51)
	) name26525 (
		_w31822_,
		_w31824_,
		_w31825_,
		_w32352_
	);
	LUT4 #(
		.INIT('hdffc)
	) name26526 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w32353_
	);
	LUT4 #(
		.INIT('h1d00)
	) name26527 (
		_w31834_,
		_w32351_,
		_w32352_,
		_w32353_,
		_w32354_
	);
	LUT4 #(
		.INIT('h3400)
	) name26528 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31827_,
		_w32355_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name26529 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w32356_
	);
	LUT4 #(
		.INIT('h153f)
	) name26530 (
		_w31822_,
		_w31823_,
		_w31825_,
		_w31827_,
		_w32357_
	);
	LUT3 #(
		.INIT('h15)
	) name26531 (
		_w32355_,
		_w32356_,
		_w32357_,
		_w32358_
	);
	LUT4 #(
		.INIT('h0040)
	) name26532 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31827_,
		_w32359_
	);
	LUT4 #(
		.INIT('h77ef)
	) name26533 (
		_w31822_,
		_w31823_,
		_w31824_,
		_w31825_,
		_w32360_
	);
	LUT3 #(
		.INIT('h31)
	) name26534 (
		_w31827_,
		_w32359_,
		_w32360_,
		_w32361_
	);
	LUT4 #(
		.INIT('hd800)
	) name26535 (
		_w31821_,
		_w32358_,
		_w32354_,
		_w32361_,
		_w32362_
	);
	LUT2 #(
		.INIT('h9)
	) name26536 (
		\u0_L2_reg[18]/NET0131 ,
		_w32362_,
		_w32363_
	);
	LUT4 #(
		.INIT('hc693)
	) name26537 (
		decrypt_pad,
		\u0_R1_reg[28]/NET0131 ,
		\u0_uk_K_r1_reg[14]/NET0131 ,
		\u0_uk_K_r1_reg[8]/NET0131 ,
		_w32364_
	);
	LUT4 #(
		.INIT('hc963)
	) name26538 (
		decrypt_pad,
		\u0_R1_reg[27]/NET0131 ,
		\u0_uk_K_r1_reg[21]/NET0131 ,
		\u0_uk_K_r1_reg[31]/NET0131 ,
		_w32365_
	);
	LUT4 #(
		.INIT('hc963)
	) name26539 (
		decrypt_pad,
		\u0_R1_reg[26]/NET0131 ,
		\u0_uk_K_r1_reg[43]/NET0131 ,
		\u0_uk_K_r1_reg[49]/NET0131 ,
		_w32366_
	);
	LUT4 #(
		.INIT('hc963)
	) name26540 (
		decrypt_pad,
		\u0_R1_reg[24]/NET0131 ,
		\u0_uk_K_r1_reg[23]/NET0131 ,
		\u0_uk_K_r1_reg[29]/NET0131 ,
		_w32367_
	);
	LUT4 #(
		.INIT('hc963)
	) name26541 (
		decrypt_pad,
		\u0_R1_reg[25]/NET0131 ,
		\u0_uk_K_r1_reg[31]/NET0131 ,
		\u0_uk_K_r1_reg[9]/NET0131 ,
		_w32368_
	);
	LUT4 #(
		.INIT('hc963)
	) name26542 (
		decrypt_pad,
		\u0_R1_reg[29]/NET0131 ,
		\u0_uk_K_r1_reg[0]/NET0131 ,
		\u0_uk_K_r1_reg[37]/NET0131 ,
		_w32369_
	);
	LUT4 #(
		.INIT('h0004)
	) name26543 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32370_
	);
	LUT4 #(
		.INIT('h6659)
	) name26544 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32371_
	);
	LUT4 #(
		.INIT('h0008)
	) name26545 (
		_w32365_,
		_w32367_,
		_w32366_,
		_w32368_,
		_w32372_
	);
	LUT2 #(
		.INIT('h6)
	) name26546 (
		_w32367_,
		_w32366_,
		_w32373_
	);
	LUT4 #(
		.INIT('h9000)
	) name26547 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32374_
	);
	LUT4 #(
		.INIT('h0302)
	) name26548 (
		_w32365_,
		_w32372_,
		_w32374_,
		_w32371_,
		_w32375_
	);
	LUT2 #(
		.INIT('h1)
	) name26549 (
		_w32364_,
		_w32375_,
		_w32376_
	);
	LUT4 #(
		.INIT('h0200)
	) name26550 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32377_
	);
	LUT4 #(
		.INIT('hadff)
	) name26551 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32378_
	);
	LUT2 #(
		.INIT('h1)
	) name26552 (
		_w32365_,
		_w32378_,
		_w32379_
	);
	LUT3 #(
		.INIT('h15)
	) name26553 (
		_w32366_,
		_w32368_,
		_w32369_,
		_w32380_
	);
	LUT4 #(
		.INIT('h0888)
	) name26554 (
		_w32365_,
		_w32367_,
		_w32366_,
		_w32368_,
		_w32381_
	);
	LUT4 #(
		.INIT('h0400)
	) name26555 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32382_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name26556 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32383_
	);
	LUT3 #(
		.INIT('hb0)
	) name26557 (
		_w32380_,
		_w32381_,
		_w32383_,
		_w32384_
	);
	LUT4 #(
		.INIT('h4100)
	) name26558 (
		_w32365_,
		_w32367_,
		_w32366_,
		_w32368_,
		_w32385_
	);
	LUT4 #(
		.INIT('h0040)
	) name26559 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32386_
	);
	LUT4 #(
		.INIT('hfbb4)
	) name26560 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32387_
	);
	LUT3 #(
		.INIT('h31)
	) name26561 (
		_w32365_,
		_w32385_,
		_w32387_,
		_w32388_
	);
	LUT4 #(
		.INIT('h7500)
	) name26562 (
		_w32364_,
		_w32379_,
		_w32384_,
		_w32388_,
		_w32389_
	);
	LUT3 #(
		.INIT('h65)
	) name26563 (
		\u0_L1_reg[22]/NET0131 ,
		_w32376_,
		_w32389_,
		_w32390_
	);
	LUT4 #(
		.INIT('hc963)
	) name26564 (
		decrypt_pad,
		\u0_R1_reg[3]/NET0131 ,
		\u0_uk_K_r1_reg[24]/NET0131 ,
		\u0_uk_K_r1_reg[32]/NET0131 ,
		_w32391_
	);
	LUT4 #(
		.INIT('hc963)
	) name26565 (
		decrypt_pad,
		\u0_R1_reg[2]/NET0131 ,
		\u0_uk_K_r1_reg[47]/NET0131 ,
		\u0_uk_K_r1_reg[55]/NET0131 ,
		_w32392_
	);
	LUT4 #(
		.INIT('hc693)
	) name26566 (
		decrypt_pad,
		\u0_R1_reg[5]/NET0131 ,
		\u0_uk_K_r1_reg[13]/NET0131 ,
		\u0_uk_K_r1_reg[5]/NET0131 ,
		_w32393_
	);
	LUT2 #(
		.INIT('h9)
	) name26567 (
		_w32392_,
		_w32393_,
		_w32394_
	);
	LUT4 #(
		.INIT('hc963)
	) name26568 (
		decrypt_pad,
		\u0_R1_reg[32]/NET0131 ,
		\u0_uk_K_r1_reg[11]/NET0131 ,
		\u0_uk_K_r1_reg[19]/NET0131 ,
		_w32395_
	);
	LUT4 #(
		.INIT('hc963)
	) name26569 (
		decrypt_pad,
		\u0_R1_reg[1]/NET0131 ,
		\u0_uk_K_r1_reg[32]/NET0131 ,
		\u0_uk_K_r1_reg[40]/NET0131 ,
		_w32396_
	);
	LUT2 #(
		.INIT('h1)
	) name26570 (
		_w32396_,
		_w32393_,
		_w32397_
	);
	LUT2 #(
		.INIT('h8)
	) name26571 (
		_w32396_,
		_w32393_,
		_w32398_
	);
	LUT2 #(
		.INIT('h6)
	) name26572 (
		_w32396_,
		_w32393_,
		_w32399_
	);
	LUT4 #(
		.INIT('h100c)
	) name26573 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32400_
	);
	LUT3 #(
		.INIT('hb8)
	) name26574 (
		_w32395_,
		_w32396_,
		_w32393_,
		_w32401_
	);
	LUT4 #(
		.INIT('hc693)
	) name26575 (
		decrypt_pad,
		\u0_R1_reg[4]/NET0131 ,
		\u0_uk_K_r1_reg[10]/P0001 ,
		\u0_uk_K_r1_reg[34]/NET0131 ,
		_w32402_
	);
	LUT2 #(
		.INIT('h9)
	) name26576 (
		_w32395_,
		_w32392_,
		_w32403_
	);
	LUT3 #(
		.INIT('h09)
	) name26577 (
		_w32395_,
		_w32392_,
		_w32402_,
		_w32404_
	);
	LUT3 #(
		.INIT('h80)
	) name26578 (
		_w32396_,
		_w32392_,
		_w32393_,
		_w32405_
	);
	LUT4 #(
		.INIT('h8000)
	) name26579 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32406_
	);
	LUT4 #(
		.INIT('h000b)
	) name26580 (
		_w32401_,
		_w32404_,
		_w32406_,
		_w32400_,
		_w32407_
	);
	LUT2 #(
		.INIT('h1)
	) name26581 (
		_w32391_,
		_w32407_,
		_w32408_
	);
	LUT2 #(
		.INIT('h4)
	) name26582 (
		_w32391_,
		_w32396_,
		_w32409_
	);
	LUT4 #(
		.INIT('h4340)
	) name26583 (
		_w32391_,
		_w32395_,
		_w32396_,
		_w32392_,
		_w32410_
	);
	LUT4 #(
		.INIT('h0002)
	) name26584 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32411_
	);
	LUT3 #(
		.INIT('h10)
	) name26585 (
		_w32411_,
		_w32410_,
		_w32402_,
		_w32412_
	);
	LUT3 #(
		.INIT('h0b)
	) name26586 (
		_w32395_,
		_w32392_,
		_w32393_,
		_w32413_
	);
	LUT3 #(
		.INIT('h2a)
	) name26587 (
		_w32391_,
		_w32396_,
		_w32393_,
		_w32414_
	);
	LUT2 #(
		.INIT('h2)
	) name26588 (
		_w32391_,
		_w32392_,
		_w32415_
	);
	LUT3 #(
		.INIT('hc4)
	) name26589 (
		_w32391_,
		_w32396_,
		_w32392_,
		_w32416_
	);
	LUT2 #(
		.INIT('h4)
	) name26590 (
		_w32395_,
		_w32393_,
		_w32417_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name26591 (
		_w32413_,
		_w32414_,
		_w32416_,
		_w32417_,
		_w32418_
	);
	LUT2 #(
		.INIT('h8)
	) name26592 (
		_w32412_,
		_w32418_,
		_w32419_
	);
	LUT3 #(
		.INIT('h20)
	) name26593 (
		_w32395_,
		_w32392_,
		_w32393_,
		_w32420_
	);
	LUT3 #(
		.INIT('h23)
	) name26594 (
		_w32409_,
		_w32402_,
		_w32420_,
		_w32421_
	);
	LUT2 #(
		.INIT('h2)
	) name26595 (
		_w32396_,
		_w32393_,
		_w32422_
	);
	LUT3 #(
		.INIT('h80)
	) name26596 (
		_w32391_,
		_w32395_,
		_w32392_,
		_w32423_
	);
	LUT2 #(
		.INIT('h8)
	) name26597 (
		_w32422_,
		_w32423_,
		_w32424_
	);
	LUT4 #(
		.INIT('h0004)
	) name26598 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32425_
	);
	LUT3 #(
		.INIT('h20)
	) name26599 (
		_w32391_,
		_w32395_,
		_w32392_,
		_w32426_
	);
	LUT3 #(
		.INIT('h13)
	) name26600 (
		_w32398_,
		_w32425_,
		_w32426_,
		_w32427_
	);
	LUT3 #(
		.INIT('h40)
	) name26601 (
		_w32424_,
		_w32421_,
		_w32427_,
		_w32428_
	);
	LUT4 #(
		.INIT('h0008)
	) name26602 (
		_w32391_,
		_w32395_,
		_w32396_,
		_w32392_,
		_w32429_
	);
	LUT3 #(
		.INIT('h15)
	) name26603 (
		_w32429_,
		_w32397_,
		_w32426_,
		_w32430_
	);
	LUT4 #(
		.INIT('h0e00)
	) name26604 (
		_w32419_,
		_w32428_,
		_w32408_,
		_w32430_,
		_w32431_
	);
	LUT2 #(
		.INIT('h9)
	) name26605 (
		\u0_L1_reg[31]/NET0131 ,
		_w32431_,
		_w32432_
	);
	LUT4 #(
		.INIT('hc963)
	) name26606 (
		decrypt_pad,
		\u0_R1_reg[32]/NET0131 ,
		\u0_uk_K_r1_reg[28]/NET0131 ,
		\u0_uk_K_r1_reg[38]/NET0131 ,
		_w32433_
	);
	LUT4 #(
		.INIT('hc963)
	) name26607 (
		decrypt_pad,
		\u0_R1_reg[31]/NET0131 ,
		\u0_uk_K_r1_reg[22]/NET0131 ,
		\u0_uk_K_r1_reg[28]/NET0131 ,
		_w32434_
	);
	LUT4 #(
		.INIT('hc963)
	) name26608 (
		decrypt_pad,
		\u0_R1_reg[28]/NET0131 ,
		\u0_uk_K_r1_reg[37]/NET0131 ,
		\u0_uk_K_r1_reg[43]/NET0131 ,
		_w32435_
	);
	LUT4 #(
		.INIT('hc693)
	) name26609 (
		decrypt_pad,
		\u0_R1_reg[30]/NET0131 ,
		\u0_uk_K_r1_reg[16]/NET0131 ,
		\u0_uk_K_r1_reg[38]/NET0131 ,
		_w32436_
	);
	LUT4 #(
		.INIT('hc693)
	) name26610 (
		decrypt_pad,
		\u0_R1_reg[29]/NET0131 ,
		\u0_uk_K_r1_reg[15]/NET0131 ,
		\u0_uk_K_r1_reg[9]/NET0131 ,
		_w32437_
	);
	LUT3 #(
		.INIT('h01)
	) name26611 (
		_w32436_,
		_w32437_,
		_w32435_,
		_w32438_
	);
	LUT4 #(
		.INIT('hc693)
	) name26612 (
		decrypt_pad,
		\u0_R1_reg[1]/NET0131 ,
		\u0_uk_K_r1_reg[0]/NET0131 ,
		\u0_uk_K_r1_reg[49]/NET0131 ,
		_w32439_
	);
	LUT4 #(
		.INIT('h0400)
	) name26613 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32440_
	);
	LUT4 #(
		.INIT('h590c)
	) name26614 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32441_
	);
	LUT4 #(
		.INIT('h0080)
	) name26615 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32442_
	);
	LUT4 #(
		.INIT('h001b)
	) name26616 (
		_w32434_,
		_w32438_,
		_w32441_,
		_w32442_,
		_w32443_
	);
	LUT2 #(
		.INIT('h2)
	) name26617 (
		_w32433_,
		_w32443_,
		_w32444_
	);
	LUT4 #(
		.INIT('h2a35)
	) name26618 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32445_
	);
	LUT4 #(
		.INIT('hfdcf)
	) name26619 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32446_
	);
	LUT4 #(
		.INIT('h7bff)
	) name26620 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32447_
	);
	LUT4 #(
		.INIT('hb800)
	) name26621 (
		_w32446_,
		_w32434_,
		_w32445_,
		_w32447_,
		_w32448_
	);
	LUT4 #(
		.INIT('h1008)
	) name26622 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32449_
	);
	LUT4 #(
		.INIT('h0020)
	) name26623 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32450_
	);
	LUT4 #(
		.INIT('hffde)
	) name26624 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32451_
	);
	LUT3 #(
		.INIT('h20)
	) name26625 (
		_w32434_,
		_w32449_,
		_w32451_,
		_w32452_
	);
	LUT4 #(
		.INIT('h0800)
	) name26626 (
		_w32433_,
		_w32436_,
		_w32437_,
		_w32435_,
		_w32453_
	);
	LUT3 #(
		.INIT('h01)
	) name26627 (
		_w32434_,
		_w32440_,
		_w32453_,
		_w32454_
	);
	LUT4 #(
		.INIT('heee0)
	) name26628 (
		_w32433_,
		_w32448_,
		_w32452_,
		_w32454_,
		_w32455_
	);
	LUT3 #(
		.INIT('h9a)
	) name26629 (
		\u0_L1_reg[5]/NET0131 ,
		_w32444_,
		_w32455_,
		_w32456_
	);
	LUT4 #(
		.INIT('hc963)
	) name26630 (
		decrypt_pad,
		\u0_R1_reg[24]/NET0131 ,
		\u0_uk_K_r1_reg[1]/NET0131 ,
		\u0_uk_K_r1_reg[7]/P0001 ,
		_w32457_
	);
	LUT4 #(
		.INIT('hc693)
	) name26631 (
		decrypt_pad,
		\u0_R1_reg[22]/NET0131 ,
		\u0_uk_K_r1_reg[23]/NET0131 ,
		\u0_uk_K_r1_reg[45]/NET0131 ,
		_w32458_
	);
	LUT4 #(
		.INIT('hc693)
	) name26632 (
		decrypt_pad,
		\u0_R1_reg[21]/NET0131 ,
		\u0_uk_K_r1_reg[1]/NET0131 ,
		\u0_uk_K_r1_reg[50]/NET0131 ,
		_w32459_
	);
	LUT4 #(
		.INIT('hc963)
	) name26633 (
		decrypt_pad,
		\u0_R1_reg[20]/NET0131 ,
		\u0_uk_K_r1_reg[35]/NET0131 ,
		\u0_uk_K_r1_reg[45]/NET0131 ,
		_w32460_
	);
	LUT4 #(
		.INIT('hc693)
	) name26634 (
		decrypt_pad,
		\u0_R1_reg[25]/NET0131 ,
		\u0_uk_K_r1_reg[2]/NET0131 ,
		\u0_uk_K_r1_reg[51]/NET0131 ,
		_w32461_
	);
	LUT4 #(
		.INIT('he020)
	) name26635 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32462_
	);
	LUT4 #(
		.INIT('hc963)
	) name26636 (
		decrypt_pad,
		\u0_R1_reg[23]/NET0131 ,
		\u0_uk_K_r1_reg[30]/NET0131 ,
		\u0_uk_K_r1_reg[36]/NET0131 ,
		_w32463_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name26637 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32464_
	);
	LUT3 #(
		.INIT('h01)
	) name26638 (
		_w32463_,
		_w32464_,
		_w32462_,
		_w32465_
	);
	LUT4 #(
		.INIT('h0004)
	) name26639 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32466_
	);
	LUT4 #(
		.INIT('h57db)
	) name26640 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32467_
	);
	LUT2 #(
		.INIT('h1)
	) name26641 (
		_w32458_,
		_w32463_,
		_w32468_
	);
	LUT4 #(
		.INIT('h0200)
	) name26642 (
		_w32460_,
		_w32458_,
		_w32463_,
		_w32461_,
		_w32469_
	);
	LUT2 #(
		.INIT('h4)
	) name26643 (
		_w32459_,
		_w32469_,
		_w32470_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name26644 (
		_w32459_,
		_w32463_,
		_w32467_,
		_w32469_,
		_w32471_
	);
	LUT3 #(
		.INIT('h8a)
	) name26645 (
		_w32457_,
		_w32465_,
		_w32471_,
		_w32472_
	);
	LUT4 #(
		.INIT('h0028)
	) name26646 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32463_,
		_w32473_
	);
	LUT3 #(
		.INIT('hd0)
	) name26647 (
		_w32460_,
		_w32458_,
		_w32463_,
		_w32474_
	);
	LUT3 #(
		.INIT('h54)
	) name26648 (
		_w32459_,
		_w32460_,
		_w32461_,
		_w32475_
	);
	LUT2 #(
		.INIT('h8)
	) name26649 (
		_w32474_,
		_w32475_,
		_w32476_
	);
	LUT3 #(
		.INIT('hc4)
	) name26650 (
		_w32459_,
		_w32460_,
		_w32461_,
		_w32477_
	);
	LUT3 #(
		.INIT('h32)
	) name26651 (
		_w32460_,
		_w32458_,
		_w32463_,
		_w32478_
	);
	LUT4 #(
		.INIT('h0002)
	) name26652 (
		_w32460_,
		_w32458_,
		_w32463_,
		_w32461_,
		_w32479_
	);
	LUT4 #(
		.INIT('h4000)
	) name26653 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32480_
	);
	LUT4 #(
		.INIT('h000b)
	) name26654 (
		_w32477_,
		_w32478_,
		_w32479_,
		_w32480_,
		_w32481_
	);
	LUT4 #(
		.INIT('h00ef)
	) name26655 (
		_w32473_,
		_w32476_,
		_w32481_,
		_w32457_,
		_w32482_
	);
	LUT3 #(
		.INIT('h02)
	) name26656 (
		_w32459_,
		_w32458_,
		_w32461_,
		_w32483_
	);
	LUT4 #(
		.INIT('h33f5)
	) name26657 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32484_
	);
	LUT2 #(
		.INIT('h2)
	) name26658 (
		_w32474_,
		_w32484_,
		_w32485_
	);
	LUT3 #(
		.INIT('h01)
	) name26659 (
		_w32459_,
		_w32460_,
		_w32461_,
		_w32486_
	);
	LUT2 #(
		.INIT('h8)
	) name26660 (
		_w32468_,
		_w32486_,
		_w32487_
	);
	LUT4 #(
		.INIT('h0100)
	) name26661 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32488_
	);
	LUT3 #(
		.INIT('h08)
	) name26662 (
		_w32459_,
		_w32460_,
		_w32461_,
		_w32489_
	);
	LUT4 #(
		.INIT('h2e3f)
	) name26663 (
		_w32458_,
		_w32463_,
		_w32488_,
		_w32489_,
		_w32490_
	);
	LUT3 #(
		.INIT('h04)
	) name26664 (
		_w32487_,
		_w32490_,
		_w32485_,
		_w32491_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name26665 (
		\u0_L1_reg[11]/NET0131 ,
		_w32482_,
		_w32472_,
		_w32491_,
		_w32492_
	);
	LUT4 #(
		.INIT('hc693)
	) name26666 (
		decrypt_pad,
		\u0_R1_reg[16]/NET0131 ,
		\u0_uk_K_r1_reg[12]/NET0131 ,
		\u0_uk_K_r1_reg[4]/NET0131 ,
		_w32493_
	);
	LUT4 #(
		.INIT('hc693)
	) name26667 (
		decrypt_pad,
		\u0_R1_reg[15]/NET0131 ,
		\u0_uk_K_r1_reg[4]/NET0131 ,
		\u0_uk_K_r1_reg[53]/NET0131 ,
		_w32494_
	);
	LUT4 #(
		.INIT('hc963)
	) name26668 (
		decrypt_pad,
		\u0_R1_reg[13]/NET0131 ,
		\u0_uk_K_r1_reg[19]/NET0131 ,
		\u0_uk_K_r1_reg[27]/NET0131 ,
		_w32495_
	);
	LUT4 #(
		.INIT('hc693)
	) name26669 (
		decrypt_pad,
		\u0_R1_reg[17]/NET0131 ,
		\u0_uk_K_r1_reg[17]/NET0131 ,
		\u0_uk_K_r1_reg[41]/NET0131 ,
		_w32496_
	);
	LUT4 #(
		.INIT('hc963)
	) name26670 (
		decrypt_pad,
		\u0_R1_reg[12]/NET0131 ,
		\u0_uk_K_r1_reg[25]/NET0131 ,
		\u0_uk_K_r1_reg[33]/NET0131 ,
		_w32497_
	);
	LUT3 #(
		.INIT('h40)
	) name26671 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32498_
	);
	LUT4 #(
		.INIT('h4000)
	) name26672 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32494_,
		_w32499_
	);
	LUT4 #(
		.INIT('hc963)
	) name26673 (
		decrypt_pad,
		\u0_R1_reg[14]/NET0131 ,
		\u0_uk_K_r1_reg[20]/NET0131 ,
		\u0_uk_K_r1_reg[53]/NET0131 ,
		_w32500_
	);
	LUT2 #(
		.INIT('h2)
	) name26674 (
		_w32496_,
		_w32497_,
		_w32501_
	);
	LUT3 #(
		.INIT('h20)
	) name26675 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32502_
	);
	LUT4 #(
		.INIT('h0020)
	) name26676 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32503_
	);
	LUT2 #(
		.INIT('h1)
	) name26677 (
		_w32499_,
		_w32503_,
		_w32504_
	);
	LUT2 #(
		.INIT('h6)
	) name26678 (
		_w32496_,
		_w32494_,
		_w32505_
	);
	LUT4 #(
		.INIT('h1110)
	) name26679 (
		_w32497_,
		_w32495_,
		_w32494_,
		_w32500_,
		_w32506_
	);
	LUT4 #(
		.INIT('h0006)
	) name26680 (
		_w32497_,
		_w32495_,
		_w32494_,
		_w32500_,
		_w32507_
	);
	LUT4 #(
		.INIT('h8000)
	) name26681 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32508_
	);
	LUT4 #(
		.INIT('h1011)
	) name26682 (
		_w32507_,
		_w32508_,
		_w32505_,
		_w32506_,
		_w32509_
	);
	LUT3 #(
		.INIT('h2a)
	) name26683 (
		_w32493_,
		_w32504_,
		_w32509_,
		_w32510_
	);
	LUT4 #(
		.INIT('hfe00)
	) name26684 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32494_,
		_w32511_
	);
	LUT4 #(
		.INIT('h7e00)
	) name26685 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32494_,
		_w32512_
	);
	LUT3 #(
		.INIT('h40)
	) name26686 (
		_w32496_,
		_w32497_,
		_w32500_,
		_w32513_
	);
	LUT3 #(
		.INIT('h0d)
	) name26687 (
		_w32496_,
		_w32495_,
		_w32494_,
		_w32514_
	);
	LUT3 #(
		.INIT('h45)
	) name26688 (
		_w32512_,
		_w32513_,
		_w32514_,
		_w32515_
	);
	LUT4 #(
		.INIT('h1000)
	) name26689 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32516_
	);
	LUT4 #(
		.INIT('heffe)
	) name26690 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32517_
	);
	LUT2 #(
		.INIT('h8)
	) name26691 (
		_w32494_,
		_w32500_,
		_w32518_
	);
	LUT3 #(
		.INIT('h80)
	) name26692 (
		_w32495_,
		_w32494_,
		_w32500_,
		_w32519_
	);
	LUT4 #(
		.INIT('h4000)
	) name26693 (
		_w32497_,
		_w32495_,
		_w32494_,
		_w32500_,
		_w32520_
	);
	LUT4 #(
		.INIT('h0008)
	) name26694 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32521_
	);
	LUT3 #(
		.INIT('h10)
	) name26695 (
		_w32520_,
		_w32521_,
		_w32517_,
		_w32522_
	);
	LUT3 #(
		.INIT('h45)
	) name26696 (
		_w32493_,
		_w32515_,
		_w32522_,
		_w32523_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name26697 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32524_
	);
	LUT2 #(
		.INIT('h2)
	) name26698 (
		_w32494_,
		_w32524_,
		_w32525_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26699 (
		_w32494_,
		_w32500_,
		_w32502_,
		_w32498_,
		_w32526_
	);
	LUT2 #(
		.INIT('h4)
	) name26700 (
		_w32525_,
		_w32526_,
		_w32527_
	);
	LUT4 #(
		.INIT('h5655)
	) name26701 (
		\u0_L1_reg[20]/NET0131 ,
		_w32523_,
		_w32510_,
		_w32527_,
		_w32528_
	);
	LUT4 #(
		.INIT('hc963)
	) name26702 (
		decrypt_pad,
		\u0_R1_reg[19]/NET0131 ,
		\u0_uk_K_r1_reg[29]/NET0131 ,
		\u0_uk_K_r1_reg[35]/NET0131 ,
		_w32529_
	);
	LUT4 #(
		.INIT('hc963)
	) name26703 (
		decrypt_pad,
		\u0_R1_reg[16]/NET0131 ,
		\u0_uk_K_r1_reg[2]/NET0131 ,
		\u0_uk_K_r1_reg[8]/NET0131 ,
		_w32530_
	);
	LUT4 #(
		.INIT('hc963)
	) name26704 (
		decrypt_pad,
		\u0_R1_reg[21]/NET0131 ,
		\u0_uk_K_r1_reg[14]/NET0131 ,
		\u0_uk_K_r1_reg[51]/NET0131 ,
		_w32531_
	);
	LUT4 #(
		.INIT('hc963)
	) name26705 (
		decrypt_pad,
		\u0_R1_reg[18]/NET0131 ,
		\u0_uk_K_r1_reg[42]/NET0131 ,
		\u0_uk_K_r1_reg[52]/NET0131 ,
		_w32532_
	);
	LUT4 #(
		.INIT('hc693)
	) name26706 (
		decrypt_pad,
		\u0_R1_reg[17]/NET0131 ,
		\u0_uk_K_r1_reg[30]/NET0131 ,
		\u0_uk_K_r1_reg[52]/NET0131 ,
		_w32533_
	);
	LUT4 #(
		.INIT('h0800)
	) name26707 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32534_
	);
	LUT4 #(
		.INIT('h0002)
	) name26708 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32535_
	);
	LUT4 #(
		.INIT('hc7b9)
	) name26709 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32536_
	);
	LUT3 #(
		.INIT('h10)
	) name26710 (
		_w32530_,
		_w32532_,
		_w32533_,
		_w32537_
	);
	LUT4 #(
		.INIT('h7a6e)
	) name26711 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32538_
	);
	LUT4 #(
		.INIT('h0080)
	) name26712 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32539_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name26713 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32540_
	);
	LUT4 #(
		.INIT('he400)
	) name26714 (
		_w32529_,
		_w32536_,
		_w32538_,
		_w32540_,
		_w32541_
	);
	LUT4 #(
		.INIT('hc963)
	) name26715 (
		decrypt_pad,
		\u0_R1_reg[20]/NET0131 ,
		\u0_uk_K_r1_reg[44]/P0001 ,
		\u0_uk_K_r1_reg[50]/NET0131 ,
		_w32542_
	);
	LUT2 #(
		.INIT('h1)
	) name26716 (
		_w32541_,
		_w32542_,
		_w32543_
	);
	LUT4 #(
		.INIT('h95b3)
	) name26717 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32544_
	);
	LUT2 #(
		.INIT('h2)
	) name26718 (
		_w32529_,
		_w32544_,
		_w32545_
	);
	LUT2 #(
		.INIT('h6)
	) name26719 (
		_w32532_,
		_w32533_,
		_w32546_
	);
	LUT4 #(
		.INIT('h0220)
	) name26720 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32547_
	);
	LUT3 #(
		.INIT('h40)
	) name26721 (
		_w32529_,
		_w32530_,
		_w32531_,
		_w32548_
	);
	LUT3 #(
		.INIT('h23)
	) name26722 (
		_w32546_,
		_w32547_,
		_w32548_,
		_w32549_
	);
	LUT3 #(
		.INIT('h8a)
	) name26723 (
		_w32542_,
		_w32545_,
		_w32549_,
		_w32550_
	);
	LUT4 #(
		.INIT('h1040)
	) name26724 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32551_
	);
	LUT3 #(
		.INIT('hbe)
	) name26725 (
		_w32530_,
		_w32531_,
		_w32533_,
		_w32552_
	);
	LUT2 #(
		.INIT('h4)
	) name26726 (
		_w32532_,
		_w32542_,
		_w32553_
	);
	LUT4 #(
		.INIT('h0045)
	) name26727 (
		_w32529_,
		_w32552_,
		_w32553_,
		_w32551_,
		_w32554_
	);
	LUT4 #(
		.INIT('h0200)
	) name26728 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32555_
	);
	LUT3 #(
		.INIT('h10)
	) name26729 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32556_
	);
	LUT4 #(
		.INIT('h0010)
	) name26730 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32557_
	);
	LUT3 #(
		.INIT('h02)
	) name26731 (
		_w32529_,
		_w32557_,
		_w32555_,
		_w32558_
	);
	LUT2 #(
		.INIT('h1)
	) name26732 (
		_w32554_,
		_w32558_,
		_w32559_
	);
	LUT4 #(
		.INIT('h5556)
	) name26733 (
		\u0_L1_reg[14]/NET0131 ,
		_w32543_,
		_w32550_,
		_w32559_,
		_w32560_
	);
	LUT4 #(
		.INIT('hefe7)
	) name26734 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32561_
	);
	LUT2 #(
		.INIT('h2)
	) name26735 (
		_w32494_,
		_w32561_,
		_w32562_
	);
	LUT4 #(
		.INIT('h7dff)
	) name26736 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32563_
	);
	LUT2 #(
		.INIT('h2)
	) name26737 (
		_w32496_,
		_w32500_,
		_w32564_
	);
	LUT4 #(
		.INIT('hbb1b)
	) name26738 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32565_
	);
	LUT3 #(
		.INIT('h08)
	) name26739 (
		_w32497_,
		_w32495_,
		_w32500_,
		_w32566_
	);
	LUT4 #(
		.INIT('h0f07)
	) name26740 (
		_w32497_,
		_w32495_,
		_w32494_,
		_w32500_,
		_w32567_
	);
	LUT3 #(
		.INIT('h8a)
	) name26741 (
		_w32563_,
		_w32565_,
		_w32567_,
		_w32568_
	);
	LUT3 #(
		.INIT('h8a)
	) name26742 (
		_w32493_,
		_w32562_,
		_w32568_,
		_w32569_
	);
	LUT4 #(
		.INIT('hdcfe)
	) name26743 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32494_,
		_w32570_
	);
	LUT2 #(
		.INIT('h1)
	) name26744 (
		_w32518_,
		_w32570_,
		_w32571_
	);
	LUT3 #(
		.INIT('h20)
	) name26745 (
		_w32497_,
		_w32495_,
		_w32494_,
		_w32572_
	);
	LUT2 #(
		.INIT('h4)
	) name26746 (
		_w32564_,
		_w32572_,
		_w32573_
	);
	LUT4 #(
		.INIT('h0008)
	) name26747 (
		_w32496_,
		_w32497_,
		_w32494_,
		_w32500_,
		_w32574_
	);
	LUT3 #(
		.INIT('h01)
	) name26748 (
		_w32516_,
		_w32574_,
		_w32566_,
		_w32575_
	);
	LUT4 #(
		.INIT('h5455)
	) name26749 (
		_w32493_,
		_w32571_,
		_w32573_,
		_w32575_,
		_w32576_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name26750 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32577_
	);
	LUT2 #(
		.INIT('h1)
	) name26751 (
		_w32494_,
		_w32577_,
		_w32578_
	);
	LUT3 #(
		.INIT('h23)
	) name26752 (
		_w32500_,
		_w32520_,
		_w32499_,
		_w32579_
	);
	LUT2 #(
		.INIT('h4)
	) name26753 (
		_w32578_,
		_w32579_,
		_w32580_
	);
	LUT4 #(
		.INIT('h5655)
	) name26754 (
		\u0_L1_reg[10]/NET0131 ,
		_w32576_,
		_w32569_,
		_w32580_,
		_w32581_
	);
	LUT4 #(
		.INIT('h5515)
	) name26755 (
		_w32529_,
		_w32530_,
		_w32531_,
		_w32533_,
		_w32582_
	);
	LUT2 #(
		.INIT('h4)
	) name26756 (
		_w32537_,
		_w32582_,
		_w32583_
	);
	LUT3 #(
		.INIT('ha8)
	) name26757 (
		_w32529_,
		_w32530_,
		_w32533_,
		_w32584_
	);
	LUT3 #(
		.INIT('h80)
	) name26758 (
		_w32530_,
		_w32531_,
		_w32533_,
		_w32585_
	);
	LUT4 #(
		.INIT('h77fc)
	) name26759 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32586_
	);
	LUT3 #(
		.INIT('h40)
	) name26760 (
		_w32556_,
		_w32584_,
		_w32586_,
		_w32587_
	);
	LUT4 #(
		.INIT('hd3ff)
	) name26761 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32588_
	);
	LUT4 #(
		.INIT('h02aa)
	) name26762 (
		_w32542_,
		_w32583_,
		_w32587_,
		_w32588_,
		_w32589_
	);
	LUT3 #(
		.INIT('h8a)
	) name26763 (
		_w32529_,
		_w32531_,
		_w32533_,
		_w32590_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name26764 (
		_w32529_,
		_w32530_,
		_w32532_,
		_w32533_,
		_w32591_
	);
	LUT2 #(
		.INIT('h4)
	) name26765 (
		_w32590_,
		_w32591_,
		_w32592_
	);
	LUT4 #(
		.INIT('h4000)
	) name26766 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32593_
	);
	LUT4 #(
		.INIT('hafdd)
	) name26767 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32594_
	);
	LUT3 #(
		.INIT('h32)
	) name26768 (
		_w32529_,
		_w32593_,
		_w32594_,
		_w32595_
	);
	LUT4 #(
		.INIT('hdfeb)
	) name26769 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32596_
	);
	LUT4 #(
		.INIT('h0040)
	) name26770 (
		_w32529_,
		_w32530_,
		_w32532_,
		_w32533_,
		_w32597_
	);
	LUT4 #(
		.INIT('h0031)
	) name26771 (
		_w32529_,
		_w32534_,
		_w32596_,
		_w32597_,
		_w32598_
	);
	LUT4 #(
		.INIT('hba00)
	) name26772 (
		_w32542_,
		_w32592_,
		_w32595_,
		_w32598_,
		_w32599_
	);
	LUT3 #(
		.INIT('h65)
	) name26773 (
		\u0_L1_reg[25]/NET0131 ,
		_w32589_,
		_w32599_,
		_w32600_
	);
	LUT4 #(
		.INIT('h0800)
	) name26774 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32601_
	);
	LUT4 #(
		.INIT('h0010)
	) name26775 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32602_
	);
	LUT3 #(
		.INIT('h41)
	) name26776 (
		_w32365_,
		_w32368_,
		_w32369_,
		_w32603_
	);
	LUT3 #(
		.INIT('h01)
	) name26777 (
		_w32602_,
		_w32603_,
		_w32601_,
		_w32604_
	);
	LUT3 #(
		.INIT('h14)
	) name26778 (
		_w32367_,
		_w32368_,
		_w32369_,
		_w32605_
	);
	LUT3 #(
		.INIT('h70)
	) name26779 (
		_w32365_,
		_w32367_,
		_w32366_,
		_w32606_
	);
	LUT2 #(
		.INIT('h4)
	) name26780 (
		_w32605_,
		_w32606_,
		_w32607_
	);
	LUT4 #(
		.INIT('h0200)
	) name26781 (
		_w32365_,
		_w32367_,
		_w32368_,
		_w32369_,
		_w32608_
	);
	LUT4 #(
		.INIT('h0002)
	) name26782 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32609_
	);
	LUT3 #(
		.INIT('h01)
	) name26783 (
		_w32364_,
		_w32608_,
		_w32609_,
		_w32610_
	);
	LUT3 #(
		.INIT('h40)
	) name26784 (
		_w32607_,
		_w32610_,
		_w32604_,
		_w32611_
	);
	LUT3 #(
		.INIT('h02)
	) name26785 (
		_w32364_,
		_w32377_,
		_w32386_,
		_w32612_
	);
	LUT4 #(
		.INIT('h5554)
	) name26786 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32613_
	);
	LUT3 #(
		.INIT('ha2)
	) name26787 (
		_w32365_,
		_w32367_,
		_w32368_,
		_w32614_
	);
	LUT2 #(
		.INIT('h4)
	) name26788 (
		_w32613_,
		_w32614_,
		_w32615_
	);
	LUT4 #(
		.INIT('h1008)
	) name26789 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32616_
	);
	LUT3 #(
		.INIT('h0b)
	) name26790 (
		_w32365_,
		_w32382_,
		_w32616_,
		_w32617_
	);
	LUT3 #(
		.INIT('h40)
	) name26791 (
		_w32615_,
		_w32612_,
		_w32617_,
		_w32618_
	);
	LUT3 #(
		.INIT('ha9)
	) name26792 (
		\u0_L1_reg[12]/NET0131 ,
		_w32611_,
		_w32618_,
		_w32619_
	);
	LUT3 #(
		.INIT('h20)
	) name26793 (
		_w32391_,
		_w32395_,
		_w32396_,
		_w32620_
	);
	LUT2 #(
		.INIT('h4)
	) name26794 (
		_w32394_,
		_w32620_,
		_w32621_
	);
	LUT4 #(
		.INIT('h1080)
	) name26795 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32622_
	);
	LUT4 #(
		.INIT('hddea)
	) name26796 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32623_
	);
	LUT4 #(
		.INIT('h8008)
	) name26797 (
		_w32391_,
		_w32395_,
		_w32396_,
		_w32393_,
		_w32624_
	);
	LUT4 #(
		.INIT('h0032)
	) name26798 (
		_w32391_,
		_w32402_,
		_w32623_,
		_w32624_,
		_w32625_
	);
	LUT4 #(
		.INIT('h0200)
	) name26799 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32626_
	);
	LUT4 #(
		.INIT('ha9ab)
	) name26800 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32627_
	);
	LUT2 #(
		.INIT('h2)
	) name26801 (
		_w32391_,
		_w32627_,
		_w32628_
	);
	LUT4 #(
		.INIT('h4401)
	) name26802 (
		_w32391_,
		_w32395_,
		_w32396_,
		_w32392_,
		_w32629_
	);
	LUT4 #(
		.INIT('h0008)
	) name26803 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32630_
	);
	LUT4 #(
		.INIT('h0002)
	) name26804 (
		_w32402_,
		_w32405_,
		_w32630_,
		_w32629_,
		_w32631_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name26805 (
		_w32622_,
		_w32625_,
		_w32628_,
		_w32631_,
		_w32632_
	);
	LUT3 #(
		.INIT('h56)
	) name26806 (
		\u0_L1_reg[17]/NET0131 ,
		_w32621_,
		_w32632_,
		_w32633_
	);
	LUT4 #(
		.INIT('hd76b)
	) name26807 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32494_,
		_w32634_
	);
	LUT2 #(
		.INIT('h1)
	) name26808 (
		_w32500_,
		_w32634_,
		_w32635_
	);
	LUT3 #(
		.INIT('h20)
	) name26809 (
		_w32496_,
		_w32497_,
		_w32500_,
		_w32636_
	);
	LUT2 #(
		.INIT('h2)
	) name26810 (
		_w32511_,
		_w32636_,
		_w32637_
	);
	LUT3 #(
		.INIT('h80)
	) name26811 (
		_w32496_,
		_w32497_,
		_w32500_,
		_w32638_
	);
	LUT4 #(
		.INIT('h0002)
	) name26812 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32639_
	);
	LUT3 #(
		.INIT('h01)
	) name26813 (
		_w32494_,
		_w32639_,
		_w32638_,
		_w32640_
	);
	LUT4 #(
		.INIT('h6000)
	) name26814 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32641_
	);
	LUT4 #(
		.INIT('h0010)
	) name26815 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32642_
	);
	LUT3 #(
		.INIT('h02)
	) name26816 (
		_w32493_,
		_w32641_,
		_w32642_,
		_w32643_
	);
	LUT3 #(
		.INIT('he0)
	) name26817 (
		_w32637_,
		_w32640_,
		_w32643_,
		_w32644_
	);
	LUT2 #(
		.INIT('h2)
	) name26818 (
		_w32519_,
		_w32501_,
		_w32645_
	);
	LUT3 #(
		.INIT('h8a)
	) name26819 (
		_w32496_,
		_w32497_,
		_w32500_,
		_w32646_
	);
	LUT2 #(
		.INIT('h1)
	) name26820 (
		_w32495_,
		_w32494_,
		_w32647_
	);
	LUT4 #(
		.INIT('h5551)
	) name26821 (
		_w32493_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32648_
	);
	LUT3 #(
		.INIT('hb0)
	) name26822 (
		_w32646_,
		_w32647_,
		_w32648_,
		_w32649_
	);
	LUT3 #(
		.INIT('h20)
	) name26823 (
		_w32504_,
		_w32645_,
		_w32649_,
		_w32650_
	);
	LUT4 #(
		.INIT('h6665)
	) name26824 (
		\u0_L1_reg[26]/NET0131 ,
		_w32635_,
		_w32644_,
		_w32650_,
		_w32651_
	);
	LUT4 #(
		.INIT('hc693)
	) name26825 (
		decrypt_pad,
		\u0_R1_reg[8]/NET0131 ,
		\u0_uk_K_r1_reg[11]/NET0131 ,
		\u0_uk_K_r1_reg[3]/NET0131 ,
		_w32652_
	);
	LUT4 #(
		.INIT('hc963)
	) name26826 (
		decrypt_pad,
		\u0_R1_reg[7]/NET0131 ,
		\u0_uk_K_r1_reg[12]/NET0131 ,
		\u0_uk_K_r1_reg[20]/NET0131 ,
		_w32653_
	);
	LUT4 #(
		.INIT('hc963)
	) name26827 (
		decrypt_pad,
		\u0_R1_reg[6]/NET0131 ,
		\u0_uk_K_r1_reg[18]/NET0131 ,
		\u0_uk_K_r1_reg[26]/NET0131 ,
		_w32654_
	);
	LUT4 #(
		.INIT('hc963)
	) name26828 (
		decrypt_pad,
		\u0_R1_reg[5]/NET0131 ,
		\u0_uk_K_r1_reg[27]/NET0131 ,
		\u0_uk_K_r1_reg[3]/NET0131 ,
		_w32655_
	);
	LUT4 #(
		.INIT('hc693)
	) name26829 (
		decrypt_pad,
		\u0_R1_reg[4]/NET0131 ,
		\u0_uk_K_r1_reg[24]/NET0131 ,
		\u0_uk_K_r1_reg[48]/NET0131 ,
		_w32656_
	);
	LUT4 #(
		.INIT('hc963)
	) name26830 (
		decrypt_pad,
		\u0_R1_reg[9]/NET0131 ,
		\u0_uk_K_r1_reg[40]/NET0131 ,
		\u0_uk_K_r1_reg[48]/NET0131 ,
		_w32657_
	);
	LUT2 #(
		.INIT('h2)
	) name26831 (
		_w32655_,
		_w32657_,
		_w32658_
	);
	LUT4 #(
		.INIT('h3fc7)
	) name26832 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32659_
	);
	LUT2 #(
		.INIT('h2)
	) name26833 (
		_w32653_,
		_w32659_,
		_w32660_
	);
	LUT4 #(
		.INIT('hf3fa)
	) name26834 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32661_
	);
	LUT2 #(
		.INIT('h1)
	) name26835 (
		_w32653_,
		_w32661_,
		_w32662_
	);
	LUT2 #(
		.INIT('h4)
	) name26836 (
		_w32654_,
		_w32656_,
		_w32663_
	);
	LUT3 #(
		.INIT('h0b)
	) name26837 (
		_w32655_,
		_w32657_,
		_w32653_,
		_w32664_
	);
	LUT4 #(
		.INIT('h0200)
	) name26838 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32665_
	);
	LUT3 #(
		.INIT('h0d)
	) name26839 (
		_w32663_,
		_w32664_,
		_w32665_,
		_w32666_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name26840 (
		_w32652_,
		_w32662_,
		_w32660_,
		_w32666_,
		_w32667_
	);
	LUT4 #(
		.INIT('hfd7d)
	) name26841 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32668_
	);
	LUT2 #(
		.INIT('h1)
	) name26842 (
		_w32668_,
		_w32653_,
		_w32669_
	);
	LUT2 #(
		.INIT('h8)
	) name26843 (
		_w32653_,
		_w32661_,
		_w32670_
	);
	LUT3 #(
		.INIT('h10)
	) name26844 (
		_w32655_,
		_w32656_,
		_w32657_,
		_w32671_
	);
	LUT3 #(
		.INIT('h07)
	) name26845 (
		_w32655_,
		_w32656_,
		_w32653_,
		_w32672_
	);
	LUT3 #(
		.INIT('h04)
	) name26846 (
		_w32654_,
		_w32656_,
		_w32657_,
		_w32673_
	);
	LUT3 #(
		.INIT('h02)
	) name26847 (
		_w32672_,
		_w32673_,
		_w32671_,
		_w32674_
	);
	LUT2 #(
		.INIT('h6)
	) name26848 (
		_w32656_,
		_w32657_,
		_w32675_
	);
	LUT4 #(
		.INIT('hdf7d)
	) name26849 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32676_
	);
	LUT4 #(
		.INIT('h0155)
	) name26850 (
		_w32652_,
		_w32670_,
		_w32674_,
		_w32676_,
		_w32677_
	);
	LUT4 #(
		.INIT('h5556)
	) name26851 (
		\u0_L1_reg[28]/NET0131 ,
		_w32669_,
		_w32677_,
		_w32667_,
		_w32678_
	);
	LUT4 #(
		.INIT('h33cb)
	) name26852 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32679_
	);
	LUT4 #(
		.INIT('h0100)
	) name26853 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32680_
	);
	LUT4 #(
		.INIT('h5504)
	) name26854 (
		_w32433_,
		_w32434_,
		_w32679_,
		_w32680_,
		_w32681_
	);
	LUT4 #(
		.INIT('h0008)
	) name26855 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32682_
	);
	LUT4 #(
		.INIT('hddb6)
	) name26856 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32683_
	);
	LUT2 #(
		.INIT('h1)
	) name26857 (
		_w32434_,
		_w32683_,
		_w32684_
	);
	LUT3 #(
		.INIT('h40)
	) name26858 (
		_w32436_,
		_w32437_,
		_w32435_,
		_w32685_
	);
	LUT4 #(
		.INIT('h0020)
	) name26859 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32434_,
		_w32686_
	);
	LUT3 #(
		.INIT('h01)
	) name26860 (
		_w32685_,
		_w32682_,
		_w32686_,
		_w32687_
	);
	LUT4 #(
		.INIT('h0100)
	) name26861 (
		_w32437_,
		_w32439_,
		_w32435_,
		_w32434_,
		_w32688_
	);
	LUT4 #(
		.INIT('h2000)
	) name26862 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32689_
	);
	LUT2 #(
		.INIT('h1)
	) name26863 (
		_w32688_,
		_w32689_,
		_w32690_
	);
	LUT4 #(
		.INIT('h0010)
	) name26864 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32691_
	);
	LUT4 #(
		.INIT('hff6f)
	) name26865 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32692_
	);
	LUT4 #(
		.INIT('h0010)
	) name26866 (
		_w32433_,
		_w32437_,
		_w32435_,
		_w32434_,
		_w32693_
	);
	LUT3 #(
		.INIT('h0d)
	) name26867 (
		_w32434_,
		_w32692_,
		_w32693_,
		_w32694_
	);
	LUT4 #(
		.INIT('hd500)
	) name26868 (
		_w32433_,
		_w32687_,
		_w32690_,
		_w32694_,
		_w32695_
	);
	LUT4 #(
		.INIT('h5655)
	) name26869 (
		\u0_L1_reg[15]/P0001 ,
		_w32681_,
		_w32684_,
		_w32695_,
		_w32696_
	);
	LUT4 #(
		.INIT('hbc77)
	) name26870 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32697_
	);
	LUT2 #(
		.INIT('h2)
	) name26871 (
		_w32463_,
		_w32697_,
		_w32698_
	);
	LUT4 #(
		.INIT('h1000)
	) name26872 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32699_
	);
	LUT4 #(
		.INIT('hefdd)
	) name26873 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32700_
	);
	LUT4 #(
		.INIT('h0302)
	) name26874 (
		_w32463_,
		_w32466_,
		_w32469_,
		_w32700_,
		_w32701_
	);
	LUT3 #(
		.INIT('h45)
	) name26875 (
		_w32457_,
		_w32698_,
		_w32701_,
		_w32702_
	);
	LUT2 #(
		.INIT('h4)
	) name26876 (
		_w32477_,
		_w32468_,
		_w32703_
	);
	LUT4 #(
		.INIT('h0002)
	) name26877 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32704_
	);
	LUT4 #(
		.INIT('h2000)
	) name26878 (
		_w32460_,
		_w32458_,
		_w32463_,
		_w32461_,
		_w32705_
	);
	LUT3 #(
		.INIT('h80)
	) name26879 (
		_w32459_,
		_w32458_,
		_w32461_,
		_w32706_
	);
	LUT3 #(
		.INIT('h01)
	) name26880 (
		_w32705_,
		_w32704_,
		_w32706_,
		_w32707_
	);
	LUT4 #(
		.INIT('hd060)
	) name26881 (
		_w32459_,
		_w32460_,
		_w32463_,
		_w32461_,
		_w32708_
	);
	LUT4 #(
		.INIT('h070b)
	) name26882 (
		_w32459_,
		_w32460_,
		_w32463_,
		_w32461_,
		_w32709_
	);
	LUT4 #(
		.INIT('h0001)
	) name26883 (
		_w32460_,
		_w32458_,
		_w32463_,
		_w32461_,
		_w32710_
	);
	LUT4 #(
		.INIT('h00fd)
	) name26884 (
		_w32458_,
		_w32709_,
		_w32708_,
		_w32710_,
		_w32711_
	);
	LUT4 #(
		.INIT('h7500)
	) name26885 (
		_w32457_,
		_w32703_,
		_w32707_,
		_w32711_,
		_w32712_
	);
	LUT3 #(
		.INIT('h65)
	) name26886 (
		\u0_L1_reg[4]/NET0131 ,
		_w32702_,
		_w32712_,
		_w32713_
	);
	LUT2 #(
		.INIT('h4)
	) name26887 (
		_w32437_,
		_w32434_,
		_w32714_
	);
	LUT3 #(
		.INIT('h40)
	) name26888 (
		_w32436_,
		_w32439_,
		_w32435_,
		_w32715_
	);
	LUT4 #(
		.INIT('hfdfe)
	) name26889 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32716_
	);
	LUT3 #(
		.INIT('hb0)
	) name26890 (
		_w32714_,
		_w32715_,
		_w32716_,
		_w32717_
	);
	LUT4 #(
		.INIT('hd1ff)
	) name26891 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32718_
	);
	LUT2 #(
		.INIT('h2)
	) name26892 (
		_w32434_,
		_w32718_,
		_w32719_
	);
	LUT4 #(
		.INIT('h5515)
	) name26893 (
		_w32433_,
		_w32436_,
		_w32437_,
		_w32435_,
		_w32720_
	);
	LUT4 #(
		.INIT('h0008)
	) name26894 (
		_w32436_,
		_w32439_,
		_w32435_,
		_w32434_,
		_w32721_
	);
	LUT4 #(
		.INIT('h0002)
	) name26895 (
		_w32437_,
		_w32439_,
		_w32435_,
		_w32434_,
		_w32722_
	);
	LUT3 #(
		.INIT('h10)
	) name26896 (
		_w32721_,
		_w32722_,
		_w32720_,
		_w32723_
	);
	LUT3 #(
		.INIT('h40)
	) name26897 (
		_w32719_,
		_w32723_,
		_w32717_,
		_w32724_
	);
	LUT4 #(
		.INIT('hf700)
	) name26898 (
		_w32437_,
		_w32439_,
		_w32435_,
		_w32434_,
		_w32725_
	);
	LUT4 #(
		.INIT('h67ef)
	) name26899 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32726_
	);
	LUT4 #(
		.INIT('h00ef)
	) name26900 (
		_w32436_,
		_w32439_,
		_w32435_,
		_w32434_,
		_w32727_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name26901 (
		_w32689_,
		_w32725_,
		_w32726_,
		_w32727_,
		_w32728_
	);
	LUT4 #(
		.INIT('h0802)
	) name26902 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32729_
	);
	LUT3 #(
		.INIT('h02)
	) name26903 (
		_w32433_,
		_w32691_,
		_w32729_,
		_w32730_
	);
	LUT2 #(
		.INIT('h4)
	) name26904 (
		_w32728_,
		_w32730_,
		_w32731_
	);
	LUT4 #(
		.INIT('hfe00)
	) name26905 (
		_w32436_,
		_w32437_,
		_w32435_,
		_w32434_,
		_w32732_
	);
	LUT4 #(
		.INIT('h4000)
	) name26906 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32733_
	);
	LUT3 #(
		.INIT('h32)
	) name26907 (
		_w32434_,
		_w32732_,
		_w32733_,
		_w32734_
	);
	LUT4 #(
		.INIT('h55a9)
	) name26908 (
		\u0_L1_reg[21]/NET0131 ,
		_w32724_,
		_w32731_,
		_w32734_,
		_w32735_
	);
	LUT4 #(
		.INIT('h779a)
	) name26909 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32736_
	);
	LUT4 #(
		.INIT('hf17d)
	) name26910 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32737_
	);
	LUT4 #(
		.INIT('h3120)
	) name26911 (
		_w32463_,
		_w32699_,
		_w32736_,
		_w32737_,
		_w32738_
	);
	LUT2 #(
		.INIT('h1)
	) name26912 (
		_w32457_,
		_w32738_,
		_w32739_
	);
	LUT4 #(
		.INIT('hdd7d)
	) name26913 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32740_
	);
	LUT2 #(
		.INIT('h2)
	) name26914 (
		_w32463_,
		_w32740_,
		_w32741_
	);
	LUT4 #(
		.INIT('h3fce)
	) name26915 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32742_
	);
	LUT2 #(
		.INIT('h1)
	) name26916 (
		_w32463_,
		_w32742_,
		_w32743_
	);
	LUT4 #(
		.INIT('h0010)
	) name26917 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32744_
	);
	LUT4 #(
		.INIT('h0001)
	) name26918 (
		_w32479_,
		_w32480_,
		_w32488_,
		_w32744_,
		_w32745_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name26919 (
		_w32457_,
		_w32743_,
		_w32741_,
		_w32745_,
		_w32746_
	);
	LUT4 #(
		.INIT('h2000)
	) name26920 (
		_w32459_,
		_w32458_,
		_w32463_,
		_w32461_,
		_w32747_
	);
	LUT2 #(
		.INIT('h1)
	) name26921 (
		_w32466_,
		_w32747_,
		_w32748_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name26922 (
		\u0_L1_reg[29]/NET0131 ,
		_w32746_,
		_w32739_,
		_w32748_,
		_w32749_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name26923 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32750_
	);
	LUT3 #(
		.INIT('h40)
	) name26924 (
		_w32655_,
		_w32656_,
		_w32657_,
		_w32751_
	);
	LUT4 #(
		.INIT('h00bf)
	) name26925 (
		_w32655_,
		_w32656_,
		_w32657_,
		_w32653_,
		_w32752_
	);
	LUT2 #(
		.INIT('h4)
	) name26926 (
		_w32750_,
		_w32752_,
		_w32753_
	);
	LUT2 #(
		.INIT('h8)
	) name26927 (
		_w32654_,
		_w32653_,
		_w32754_
	);
	LUT3 #(
		.INIT('h15)
	) name26928 (
		_w32652_,
		_w32751_,
		_w32754_,
		_w32755_
	);
	LUT4 #(
		.INIT('h0010)
	) name26929 (
		_w32654_,
		_w32655_,
		_w32657_,
		_w32653_,
		_w32756_
	);
	LUT4 #(
		.INIT('h0800)
	) name26930 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32757_
	);
	LUT4 #(
		.INIT('h0144)
	) name26931 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32758_
	);
	LUT3 #(
		.INIT('h01)
	) name26932 (
		_w32756_,
		_w32757_,
		_w32758_,
		_w32759_
	);
	LUT3 #(
		.INIT('h40)
	) name26933 (
		_w32753_,
		_w32755_,
		_w32759_,
		_w32760_
	);
	LUT4 #(
		.INIT('h002a)
	) name26934 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32653_,
		_w32761_
	);
	LUT2 #(
		.INIT('h4)
	) name26935 (
		_w32675_,
		_w32761_,
		_w32762_
	);
	LUT4 #(
		.INIT('hc400)
	) name26936 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32653_,
		_w32763_
	);
	LUT4 #(
		.INIT('h4010)
	) name26937 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32764_
	);
	LUT4 #(
		.INIT('h0001)
	) name26938 (
		_w32655_,
		_w32656_,
		_w32657_,
		_w32653_,
		_w32765_
	);
	LUT4 #(
		.INIT('h0002)
	) name26939 (
		_w32652_,
		_w32764_,
		_w32763_,
		_w32765_,
		_w32766_
	);
	LUT2 #(
		.INIT('h4)
	) name26940 (
		_w32762_,
		_w32766_,
		_w32767_
	);
	LUT4 #(
		.INIT('h0002)
	) name26941 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32768_
	);
	LUT4 #(
		.INIT('hbfbd)
	) name26942 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32769_
	);
	LUT2 #(
		.INIT('h9)
	) name26943 (
		_w32654_,
		_w32655_,
		_w32770_
	);
	LUT3 #(
		.INIT('h04)
	) name26944 (
		_w32656_,
		_w32657_,
		_w32653_,
		_w32771_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name26945 (
		_w32653_,
		_w32769_,
		_w32770_,
		_w32771_,
		_w32772_
	);
	LUT4 #(
		.INIT('ha955)
	) name26946 (
		\u0_L1_reg[2]/NET0131 ,
		_w32760_,
		_w32767_,
		_w32772_,
		_w32773_
	);
	LUT4 #(
		.INIT('hf5f1)
	) name26947 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32774_
	);
	LUT4 #(
		.INIT('h6dff)
	) name26948 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32775_
	);
	LUT4 #(
		.INIT('h08cc)
	) name26949 (
		_w32493_,
		_w32494_,
		_w32774_,
		_w32775_,
		_w32776_
	);
	LUT4 #(
		.INIT('hfbee)
	) name26950 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32777_
	);
	LUT2 #(
		.INIT('h2)
	) name26951 (
		_w32494_,
		_w32777_,
		_w32778_
	);
	LUT4 #(
		.INIT('h0060)
	) name26952 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32779_
	);
	LUT3 #(
		.INIT('hd8)
	) name26953 (
		_w32496_,
		_w32495_,
		_w32500_,
		_w32780_
	);
	LUT2 #(
		.INIT('h2)
	) name26954 (
		_w32497_,
		_w32494_,
		_w32781_
	);
	LUT4 #(
		.INIT('h0045)
	) name26955 (
		_w32508_,
		_w32780_,
		_w32781_,
		_w32779_,
		_w32782_
	);
	LUT3 #(
		.INIT('h54)
	) name26956 (
		_w32493_,
		_w32496_,
		_w32494_,
		_w32783_
	);
	LUT4 #(
		.INIT('h4300)
	) name26957 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32784_
	);
	LUT4 #(
		.INIT('hdf0f)
	) name26958 (
		_w32496_,
		_w32497_,
		_w32495_,
		_w32500_,
		_w32785_
	);
	LUT4 #(
		.INIT('h008a)
	) name26959 (
		_w32493_,
		_w32496_,
		_w32497_,
		_w32494_,
		_w32786_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name26960 (
		_w32783_,
		_w32784_,
		_w32785_,
		_w32786_,
		_w32787_
	);
	LUT4 #(
		.INIT('hba00)
	) name26961 (
		_w32493_,
		_w32778_,
		_w32782_,
		_w32787_,
		_w32788_
	);
	LUT3 #(
		.INIT('h65)
	) name26962 (
		\u0_L1_reg[1]/NET0131 ,
		_w32776_,
		_w32788_,
		_w32789_
	);
	LUT3 #(
		.INIT('h13)
	) name26963 (
		_w32459_,
		_w32463_,
		_w32461_,
		_w32790_
	);
	LUT4 #(
		.INIT('hc4e6)
	) name26964 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32791_
	);
	LUT4 #(
		.INIT('h0201)
	) name26965 (
		_w32459_,
		_w32460_,
		_w32463_,
		_w32461_,
		_w32792_
	);
	LUT4 #(
		.INIT('h1011)
	) name26966 (
		_w32457_,
		_w32792_,
		_w32790_,
		_w32791_,
		_w32793_
	);
	LUT4 #(
		.INIT('h2010)
	) name26967 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32461_,
		_w32794_
	);
	LUT3 #(
		.INIT('h02)
	) name26968 (
		_w32457_,
		_w32488_,
		_w32483_,
		_w32795_
	);
	LUT4 #(
		.INIT('h0800)
	) name26969 (
		_w32459_,
		_w32460_,
		_w32458_,
		_w32463_,
		_w32796_
	);
	LUT4 #(
		.INIT('h1404)
	) name26970 (
		_w32459_,
		_w32460_,
		_w32463_,
		_w32461_,
		_w32797_
	);
	LUT2 #(
		.INIT('h1)
	) name26971 (
		_w32796_,
		_w32797_,
		_w32798_
	);
	LUT4 #(
		.INIT('h4555)
	) name26972 (
		_w32793_,
		_w32794_,
		_w32795_,
		_w32798_,
		_w32799_
	);
	LUT2 #(
		.INIT('h2)
	) name26973 (
		_w32490_,
		_w32470_,
		_w32800_
	);
	LUT3 #(
		.INIT('h65)
	) name26974 (
		\u0_L1_reg[19]/NET0131 ,
		_w32799_,
		_w32800_,
		_w32801_
	);
	LUT4 #(
		.INIT('h0102)
	) name26975 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32802_
	);
	LUT4 #(
		.INIT('h5545)
	) name26976 (
		_w32365_,
		_w32367_,
		_w32368_,
		_w32369_,
		_w32803_
	);
	LUT3 #(
		.INIT('h10)
	) name26977 (
		_w32601_,
		_w32802_,
		_w32803_,
		_w32804_
	);
	LUT4 #(
		.INIT('h3088)
	) name26978 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32805_
	);
	LUT4 #(
		.INIT('haaa8)
	) name26979 (
		_w32365_,
		_w32367_,
		_w32368_,
		_w32369_,
		_w32806_
	);
	LUT2 #(
		.INIT('h4)
	) name26980 (
		_w32805_,
		_w32806_,
		_w32807_
	);
	LUT4 #(
		.INIT('h0080)
	) name26981 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32808_
	);
	LUT4 #(
		.INIT('haa02)
	) name26982 (
		_w32364_,
		_w32804_,
		_w32807_,
		_w32808_,
		_w32809_
	);
	LUT4 #(
		.INIT('h8040)
	) name26983 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32810_
	);
	LUT3 #(
		.INIT('h02)
	) name26984 (
		_w32367_,
		_w32366_,
		_w32369_,
		_w32811_
	);
	LUT3 #(
		.INIT('h31)
	) name26985 (
		_w32603_,
		_w32810_,
		_w32811_,
		_w32812_
	);
	LUT4 #(
		.INIT('hf5dd)
	) name26986 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32813_
	);
	LUT4 #(
		.INIT('h0420)
	) name26987 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32814_
	);
	LUT3 #(
		.INIT('h0d)
	) name26988 (
		_w32365_,
		_w32813_,
		_w32814_,
		_w32815_
	);
	LUT4 #(
		.INIT('h5010)
	) name26989 (
		_w32365_,
		_w32367_,
		_w32368_,
		_w32369_,
		_w32816_
	);
	LUT4 #(
		.INIT('h135f)
	) name26990 (
		_w32365_,
		_w32373_,
		_w32382_,
		_w32816_,
		_w32817_
	);
	LUT4 #(
		.INIT('hea00)
	) name26991 (
		_w32364_,
		_w32812_,
		_w32815_,
		_w32817_,
		_w32818_
	);
	LUT3 #(
		.INIT('h65)
	) name26992 (
		\u0_L1_reg[32]/NET0131 ,
		_w32809_,
		_w32818_,
		_w32819_
	);
	LUT4 #(
		.INIT('hae16)
	) name26993 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32820_
	);
	LUT4 #(
		.INIT('h4880)
	) name26994 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32821_
	);
	LUT4 #(
		.INIT('h2210)
	) name26995 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32822_
	);
	LUT4 #(
		.INIT('h1032)
	) name26996 (
		_w32365_,
		_w32821_,
		_w32820_,
		_w32822_,
		_w32823_
	);
	LUT2 #(
		.INIT('h2)
	) name26997 (
		_w32364_,
		_w32823_,
		_w32824_
	);
	LUT4 #(
		.INIT('h4080)
	) name26998 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32825_
	);
	LUT4 #(
		.INIT('h2a11)
	) name26999 (
		_w32367_,
		_w32366_,
		_w32368_,
		_w32369_,
		_w32826_
	);
	LUT4 #(
		.INIT('h3332)
	) name27000 (
		_w32364_,
		_w32370_,
		_w32826_,
		_w32825_,
		_w32827_
	);
	LUT4 #(
		.INIT('h5150)
	) name27001 (
		_w32364_,
		_w32365_,
		_w32370_,
		_w32822_,
		_w32828_
	);
	LUT4 #(
		.INIT('h00b1)
	) name27002 (
		_w32365_,
		_w32821_,
		_w32827_,
		_w32828_,
		_w32829_
	);
	LUT3 #(
		.INIT('h65)
	) name27003 (
		\u0_L1_reg[7]/NET0131 ,
		_w32824_,
		_w32829_,
		_w32830_
	);
	LUT4 #(
		.INIT('hc963)
	) name27004 (
		decrypt_pad,
		\u0_R1_reg[11]/NET0131 ,
		\u0_uk_K_r1_reg[55]/NET0131 ,
		\u0_uk_K_r1_reg[6]/NET0131 ,
		_w32831_
	);
	LUT4 #(
		.INIT('hc963)
	) name27005 (
		decrypt_pad,
		\u0_R1_reg[12]/NET0131 ,
		\u0_uk_K_r1_reg[13]/NET0131 ,
		\u0_uk_K_r1_reg[46]/NET0131 ,
		_w32832_
	);
	LUT4 #(
		.INIT('hc963)
	) name27006 (
		decrypt_pad,
		\u0_R1_reg[9]/NET0131 ,
		\u0_uk_K_r1_reg[46]/NET0131 ,
		\u0_uk_K_r1_reg[54]/NET0131 ,
		_w32833_
	);
	LUT4 #(
		.INIT('hc963)
	) name27007 (
		decrypt_pad,
		\u0_R1_reg[13]/NET0131 ,
		\u0_uk_K_r1_reg[26]/NET0131 ,
		\u0_uk_K_r1_reg[34]/NET0131 ,
		_w32834_
	);
	LUT4 #(
		.INIT('hc963)
	) name27008 (
		decrypt_pad,
		\u0_R1_reg[10]/NET0131 ,
		\u0_uk_K_r1_reg[54]/NET0131 ,
		\u0_uk_K_r1_reg[5]/NET0131 ,
		_w32835_
	);
	LUT4 #(
		.INIT('hc963)
	) name27009 (
		decrypt_pad,
		\u0_R1_reg[8]/NET0131 ,
		\u0_uk_K_r1_reg[17]/NET0131 ,
		\u0_uk_K_r1_reg[25]/NET0131 ,
		_w32836_
	);
	LUT4 #(
		.INIT('hc34f)
	) name27010 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32837_
	);
	LUT2 #(
		.INIT('h1)
	) name27011 (
		_w32835_,
		_w32833_,
		_w32838_
	);
	LUT4 #(
		.INIT('h0001)
	) name27012 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32839_
	);
	LUT4 #(
		.INIT('hdfde)
	) name27013 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32840_
	);
	LUT4 #(
		.INIT('h08cc)
	) name27014 (
		_w32832_,
		_w32831_,
		_w32837_,
		_w32840_,
		_w32841_
	);
	LUT2 #(
		.INIT('h9)
	) name27015 (
		_w32835_,
		_w32833_,
		_w32842_
	);
	LUT2 #(
		.INIT('h6)
	) name27016 (
		_w32834_,
		_w32836_,
		_w32843_
	);
	LUT3 #(
		.INIT('h46)
	) name27017 (
		_w32834_,
		_w32836_,
		_w32831_,
		_w32844_
	);
	LUT4 #(
		.INIT('h0400)
	) name27018 (
		_w32835_,
		_w32833_,
		_w32836_,
		_w32831_,
		_w32845_
	);
	LUT4 #(
		.INIT('h1054)
	) name27019 (
		_w32845_,
		_w32842_,
		_w32843_,
		_w32844_,
		_w32846_
	);
	LUT2 #(
		.INIT('h8)
	) name27020 (
		_w32832_,
		_w32835_,
		_w32847_
	);
	LUT3 #(
		.INIT('h02)
	) name27021 (
		_w32833_,
		_w32834_,
		_w32836_,
		_w32848_
	);
	LUT4 #(
		.INIT('h30bb)
	) name27022 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32849_
	);
	LUT3 #(
		.INIT('h0d)
	) name27023 (
		_w32833_,
		_w32834_,
		_w32831_,
		_w32850_
	);
	LUT4 #(
		.INIT('h00a2)
	) name27024 (
		_w32832_,
		_w32833_,
		_w32834_,
		_w32831_,
		_w32851_
	);
	LUT4 #(
		.INIT('h7077)
	) name27025 (
		_w32847_,
		_w32848_,
		_w32849_,
		_w32851_,
		_w32852_
	);
	LUT4 #(
		.INIT('h3200)
	) name27026 (
		_w32832_,
		_w32841_,
		_w32846_,
		_w32852_,
		_w32853_
	);
	LUT2 #(
		.INIT('h9)
	) name27027 (
		\u0_L1_reg[6]/NET0131 ,
		_w32853_,
		_w32854_
	);
	LUT4 #(
		.INIT('hc004)
	) name27028 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32855_
	);
	LUT3 #(
		.INIT('hd7)
	) name27029 (
		_w32437_,
		_w32439_,
		_w32435_,
		_w32856_
	);
	LUT4 #(
		.INIT('he4f5)
	) name27030 (
		_w32434_,
		_w32438_,
		_w32855_,
		_w32856_,
		_w32857_
	);
	LUT4 #(
		.INIT('hed6f)
	) name27031 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32858_
	);
	LUT3 #(
		.INIT('h8a)
	) name27032 (
		_w32433_,
		_w32857_,
		_w32858_,
		_w32859_
	);
	LUT4 #(
		.INIT('hf700)
	) name27033 (
		_w32436_,
		_w32437_,
		_w32435_,
		_w32434_,
		_w32860_
	);
	LUT3 #(
		.INIT('h4b)
	) name27034 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32861_
	);
	LUT2 #(
		.INIT('h8)
	) name27035 (
		_w32860_,
		_w32861_,
		_w32862_
	);
	LUT4 #(
		.INIT('h0080)
	) name27036 (
		_w32436_,
		_w32439_,
		_w32435_,
		_w32434_,
		_w32863_
	);
	LUT3 #(
		.INIT('h01)
	) name27037 (
		_w32450_,
		_w32722_,
		_w32863_,
		_w32864_
	);
	LUT4 #(
		.INIT('hebf7)
	) name27038 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32435_,
		_w32865_
	);
	LUT4 #(
		.INIT('h0200)
	) name27039 (
		_w32436_,
		_w32437_,
		_w32439_,
		_w32434_,
		_w32866_
	);
	LUT3 #(
		.INIT('h0e)
	) name27040 (
		_w32434_,
		_w32865_,
		_w32866_,
		_w32867_
	);
	LUT4 #(
		.INIT('hba00)
	) name27041 (
		_w32433_,
		_w32862_,
		_w32864_,
		_w32867_,
		_w32868_
	);
	LUT3 #(
		.INIT('h65)
	) name27042 (
		\u0_L1_reg[27]/NET0131 ,
		_w32859_,
		_w32868_,
		_w32869_
	);
	LUT3 #(
		.INIT('h8c)
	) name27043 (
		_w32426_,
		_w32394_,
		_w32399_,
		_w32870_
	);
	LUT4 #(
		.INIT('h4440)
	) name27044 (
		_w32391_,
		_w32395_,
		_w32396_,
		_w32392_,
		_w32871_
	);
	LUT4 #(
		.INIT('h0020)
	) name27045 (
		_w32391_,
		_w32395_,
		_w32396_,
		_w32393_,
		_w32872_
	);
	LUT4 #(
		.INIT('h0203)
	) name27046 (
		_w32397_,
		_w32402_,
		_w32872_,
		_w32871_,
		_w32873_
	);
	LUT4 #(
		.INIT('h002a)
	) name27047 (
		_w32402_,
		_w32422_,
		_w32423_,
		_w32626_,
		_w32874_
	);
	LUT4 #(
		.INIT('h2000)
	) name27048 (
		_w32391_,
		_w32395_,
		_w32396_,
		_w32393_,
		_w32875_
	);
	LUT3 #(
		.INIT('h07)
	) name27049 (
		_w32397_,
		_w32426_,
		_w32875_,
		_w32876_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name27050 (
		_w32870_,
		_w32873_,
		_w32874_,
		_w32876_,
		_w32877_
	);
	LUT4 #(
		.INIT('h7ef7)
	) name27051 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32878_
	);
	LUT2 #(
		.INIT('h1)
	) name27052 (
		_w32391_,
		_w32878_,
		_w32879_
	);
	LUT3 #(
		.INIT('h96)
	) name27053 (
		_w32395_,
		_w32396_,
		_w32393_,
		_w32880_
	);
	LUT3 #(
		.INIT('ha2)
	) name27054 (
		_w32395_,
		_w32392_,
		_w32393_,
		_w32881_
	);
	LUT2 #(
		.INIT('h4)
	) name27055 (
		_w32391_,
		_w32402_,
		_w32882_
	);
	LUT3 #(
		.INIT('h20)
	) name27056 (
		_w32880_,
		_w32881_,
		_w32882_,
		_w32883_
	);
	LUT3 #(
		.INIT('h13)
	) name27057 (
		_w32391_,
		_w32429_,
		_w32425_,
		_w32884_
	);
	LUT3 #(
		.INIT('h10)
	) name27058 (
		_w32879_,
		_w32883_,
		_w32884_,
		_w32885_
	);
	LUT3 #(
		.INIT('h9a)
	) name27059 (
		\u0_L1_reg[23]/NET0131 ,
		_w32877_,
		_w32885_,
		_w32886_
	);
	LUT4 #(
		.INIT('hfde3)
	) name27060 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32887_
	);
	LUT2 #(
		.INIT('h1)
	) name27061 (
		_w32653_,
		_w32887_,
		_w32888_
	);
	LUT4 #(
		.INIT('h8b00)
	) name27062 (
		_w32654_,
		_w32656_,
		_w32657_,
		_w32653_,
		_w32889_
	);
	LUT4 #(
		.INIT('h87df)
	) name27063 (
		_w32655_,
		_w32656_,
		_w32657_,
		_w32653_,
		_w32890_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name27064 (
		_w32654_,
		_w32658_,
		_w32889_,
		_w32890_,
		_w32891_
	);
	LUT3 #(
		.INIT('h45)
	) name27065 (
		_w32652_,
		_w32888_,
		_w32891_,
		_w32892_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name27066 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32893_
	);
	LUT2 #(
		.INIT('h1)
	) name27067 (
		_w32653_,
		_w32893_,
		_w32894_
	);
	LUT3 #(
		.INIT('h02)
	) name27068 (
		_w32654_,
		_w32655_,
		_w32657_,
		_w32895_
	);
	LUT3 #(
		.INIT('h01)
	) name27069 (
		_w32654_,
		_w32655_,
		_w32657_,
		_w32896_
	);
	LUT4 #(
		.INIT('hdf00)
	) name27070 (
		_w32654_,
		_w32656_,
		_w32657_,
		_w32653_,
		_w32897_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name27071 (
		_w32752_,
		_w32895_,
		_w32896_,
		_w32897_,
		_w32898_
	);
	LUT4 #(
		.INIT('hbf7b)
	) name27072 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w32899_
	);
	LUT3 #(
		.INIT('h10)
	) name27073 (
		_w32756_,
		_w32757_,
		_w32899_,
		_w32900_
	);
	LUT4 #(
		.INIT('h1311)
	) name27074 (
		_w32652_,
		_w32894_,
		_w32898_,
		_w32900_,
		_w32901_
	);
	LUT3 #(
		.INIT('h9a)
	) name27075 (
		\u0_L1_reg[13]/NET0131 ,
		_w32892_,
		_w32901_,
		_w32902_
	);
	LUT4 #(
		.INIT('h0001)
	) name27076 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32903_
	);
	LUT4 #(
		.INIT('hff76)
	) name27077 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32904_
	);
	LUT3 #(
		.INIT('h04)
	) name27078 (
		_w32529_,
		_w32530_,
		_w32532_,
		_w32905_
	);
	LUT4 #(
		.INIT('h0031)
	) name27079 (
		_w32529_,
		_w32551_,
		_w32904_,
		_w32905_,
		_w32906_
	);
	LUT2 #(
		.INIT('h2)
	) name27080 (
		_w32542_,
		_w32906_,
		_w32907_
	);
	LUT3 #(
		.INIT('h02)
	) name27081 (
		_w32529_,
		_w32535_,
		_w32585_,
		_w32908_
	);
	LUT4 #(
		.INIT('h4404)
	) name27082 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32909_
	);
	LUT2 #(
		.INIT('h2)
	) name27083 (
		_w32582_,
		_w32909_,
		_w32910_
	);
	LUT4 #(
		.INIT('hdaef)
	) name27084 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32911_
	);
	LUT4 #(
		.INIT('h0155)
	) name27085 (
		_w32542_,
		_w32908_,
		_w32910_,
		_w32911_,
		_w32912_
	);
	LUT4 #(
		.INIT('hcbbf)
	) name27086 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32913_
	);
	LUT4 #(
		.INIT('hcf45)
	) name27087 (
		_w32529_,
		_w32531_,
		_w32597_,
		_w32913_,
		_w32914_
	);
	LUT4 #(
		.INIT('h5655)
	) name27088 (
		\u0_L1_reg[8]/NET0131 ,
		_w32912_,
		_w32907_,
		_w32914_,
		_w32915_
	);
	LUT3 #(
		.INIT('h20)
	) name27089 (
		_w32835_,
		_w32833_,
		_w32836_,
		_w32916_
	);
	LUT4 #(
		.INIT('h0200)
	) name27090 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32917_
	);
	LUT4 #(
		.INIT('hdda1)
	) name27091 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32918_
	);
	LUT4 #(
		.INIT('h5054)
	) name27092 (
		_w32832_,
		_w32831_,
		_w32917_,
		_w32918_,
		_w32919_
	);
	LUT4 #(
		.INIT('h665e)
	) name27093 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32920_
	);
	LUT2 #(
		.INIT('h2)
	) name27094 (
		_w32831_,
		_w32920_,
		_w32921_
	);
	LUT3 #(
		.INIT('h0e)
	) name27095 (
		_w32835_,
		_w32833_,
		_w32831_,
		_w32922_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name27096 (
		_w32838_,
		_w32843_,
		_w32844_,
		_w32922_,
		_w32923_
	);
	LUT3 #(
		.INIT('h8a)
	) name27097 (
		_w32832_,
		_w32921_,
		_w32923_,
		_w32924_
	);
	LUT4 #(
		.INIT('h1001)
	) name27098 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32925_
	);
	LUT4 #(
		.INIT('he35e)
	) name27099 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32926_
	);
	LUT2 #(
		.INIT('h1)
	) name27100 (
		_w32832_,
		_w32831_,
		_w32927_
	);
	LUT2 #(
		.INIT('h4)
	) name27101 (
		_w32926_,
		_w32927_,
		_w32928_
	);
	LUT3 #(
		.INIT('h10)
	) name27102 (
		_w32835_,
		_w32834_,
		_w32836_,
		_w32929_
	);
	LUT2 #(
		.INIT('h4)
	) name27103 (
		_w32833_,
		_w32831_,
		_w32930_
	);
	LUT2 #(
		.INIT('h8)
	) name27104 (
		_w32929_,
		_w32930_,
		_w32931_
	);
	LUT3 #(
		.INIT('h80)
	) name27105 (
		_w32833_,
		_w32834_,
		_w32836_,
		_w32932_
	);
	LUT2 #(
		.INIT('h2)
	) name27106 (
		_w32835_,
		_w32831_,
		_w32933_
	);
	LUT4 #(
		.INIT('h0777)
	) name27107 (
		_w32834_,
		_w32845_,
		_w32932_,
		_w32933_,
		_w32934_
	);
	LUT3 #(
		.INIT('h10)
	) name27108 (
		_w32931_,
		_w32928_,
		_w32934_,
		_w32935_
	);
	LUT4 #(
		.INIT('h5655)
	) name27109 (
		\u0_L1_reg[24]/NET0131 ,
		_w32924_,
		_w32919_,
		_w32935_,
		_w32936_
	);
	LUT4 #(
		.INIT('h59fb)
	) name27110 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32937_
	);
	LUT2 #(
		.INIT('h2)
	) name27111 (
		_w32831_,
		_w32937_,
		_w32938_
	);
	LUT3 #(
		.INIT('h5c)
	) name27112 (
		_w32835_,
		_w32833_,
		_w32836_,
		_w32939_
	);
	LUT2 #(
		.INIT('h8)
	) name27113 (
		_w32850_,
		_w32939_,
		_w32940_
	);
	LUT4 #(
		.INIT('h0020)
	) name27114 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32941_
	);
	LUT3 #(
		.INIT('h01)
	) name27115 (
		_w32832_,
		_w32925_,
		_w32941_,
		_w32942_
	);
	LUT3 #(
		.INIT('h10)
	) name27116 (
		_w32938_,
		_w32940_,
		_w32942_,
		_w32943_
	);
	LUT4 #(
		.INIT('h55f3)
	) name27117 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32944_
	);
	LUT2 #(
		.INIT('h1)
	) name27118 (
		_w32831_,
		_w32944_,
		_w32945_
	);
	LUT4 #(
		.INIT('h0600)
	) name27119 (
		_w32835_,
		_w32834_,
		_w32836_,
		_w32831_,
		_w32946_
	);
	LUT4 #(
		.INIT('h002a)
	) name27120 (
		_w32832_,
		_w32929_,
		_w32930_,
		_w32946_,
		_w32947_
	);
	LUT2 #(
		.INIT('h4)
	) name27121 (
		_w32945_,
		_w32947_,
		_w32948_
	);
	LUT3 #(
		.INIT('h2a)
	) name27122 (
		_w32833_,
		_w32834_,
		_w32836_,
		_w32949_
	);
	LUT4 #(
		.INIT('hbf00)
	) name27123 (
		_w32833_,
		_w32834_,
		_w32836_,
		_w32831_,
		_w32950_
	);
	LUT4 #(
		.INIT('haa08)
	) name27124 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32831_,
		_w32951_
	);
	LUT4 #(
		.INIT('h7077)
	) name27125 (
		_w32847_,
		_w32949_,
		_w32950_,
		_w32951_,
		_w32952_
	);
	LUT4 #(
		.INIT('h56aa)
	) name27126 (
		\u0_L1_reg[30]/NET0131 ,
		_w32943_,
		_w32948_,
		_w32952_,
		_w32953_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name27127 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32954_
	);
	LUT2 #(
		.INIT('h2)
	) name27128 (
		_w32529_,
		_w32954_,
		_w32955_
	);
	LUT4 #(
		.INIT('h2e26)
	) name27129 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32956_
	);
	LUT4 #(
		.INIT('h00d0)
	) name27130 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32957_
	);
	LUT4 #(
		.INIT('h0032)
	) name27131 (
		_w32529_,
		_w32542_,
		_w32956_,
		_w32957_,
		_w32958_
	);
	LUT4 #(
		.INIT('he6f7)
	) name27132 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32959_
	);
	LUT2 #(
		.INIT('h2)
	) name27133 (
		_w32529_,
		_w32959_,
		_w32960_
	);
	LUT4 #(
		.INIT('h0020)
	) name27134 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32961_
	);
	LUT4 #(
		.INIT('h1000)
	) name27135 (
		_w32529_,
		_w32530_,
		_w32531_,
		_w32533_,
		_w32962_
	);
	LUT4 #(
		.INIT('h0004)
	) name27136 (
		_w32534_,
		_w32542_,
		_w32961_,
		_w32962_,
		_w32963_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name27137 (
		_w32955_,
		_w32958_,
		_w32960_,
		_w32963_,
		_w32964_
	);
	LUT4 #(
		.INIT('h0040)
	) name27138 (
		_w32530_,
		_w32531_,
		_w32532_,
		_w32533_,
		_w32965_
	);
	LUT3 #(
		.INIT('h02)
	) name27139 (
		_w32529_,
		_w32535_,
		_w32965_,
		_w32966_
	);
	LUT4 #(
		.INIT('h0001)
	) name27140 (
		_w32529_,
		_w32539_,
		_w32555_,
		_w32903_,
		_w32967_
	);
	LUT2 #(
		.INIT('h1)
	) name27141 (
		_w32966_,
		_w32967_,
		_w32968_
	);
	LUT3 #(
		.INIT('h56)
	) name27142 (
		\u0_L1_reg[3]/NET0131 ,
		_w32964_,
		_w32968_,
		_w32969_
	);
	LUT4 #(
		.INIT('h696b)
	) name27143 (
		_w32833_,
		_w32834_,
		_w32836_,
		_w32831_,
		_w32970_
	);
	LUT4 #(
		.INIT('h0080)
	) name27144 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32971_
	);
	LUT4 #(
		.INIT('h0012)
	) name27145 (
		_w32835_,
		_w32834_,
		_w32836_,
		_w32831_,
		_w32972_
	);
	LUT4 #(
		.INIT('h0032)
	) name27146 (
		_w32835_,
		_w32971_,
		_w32970_,
		_w32972_,
		_w32973_
	);
	LUT2 #(
		.INIT('h2)
	) name27147 (
		_w32832_,
		_w32973_,
		_w32974_
	);
	LUT4 #(
		.INIT('h3fca)
	) name27148 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32975_
	);
	LUT4 #(
		.INIT('h3031)
	) name27149 (
		_w32832_,
		_w32831_,
		_w32916_,
		_w32975_,
		_w32976_
	);
	LUT3 #(
		.INIT('h04)
	) name27150 (
		_w32832_,
		_w32839_,
		_w32975_,
		_w32977_
	);
	LUT4 #(
		.INIT('h0802)
	) name27151 (
		_w32835_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32978_
	);
	LUT4 #(
		.INIT('h1440)
	) name27152 (
		_w32832_,
		_w32833_,
		_w32834_,
		_w32836_,
		_w32979_
	);
	LUT3 #(
		.INIT('ha8)
	) name27153 (
		_w32831_,
		_w32978_,
		_w32979_,
		_w32980_
	);
	LUT3 #(
		.INIT('h01)
	) name27154 (
		_w32977_,
		_w32980_,
		_w32976_,
		_w32981_
	);
	LUT3 #(
		.INIT('h65)
	) name27155 (
		\u0_L1_reg[16]/NET0131 ,
		_w32974_,
		_w32981_,
		_w32982_
	);
	LUT4 #(
		.INIT('h2810)
	) name27156 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32983_
	);
	LUT3 #(
		.INIT('h02)
	) name27157 (
		_w32395_,
		_w32392_,
		_w32393_,
		_w32984_
	);
	LUT3 #(
		.INIT('h28)
	) name27158 (
		_w32391_,
		_w32396_,
		_w32393_,
		_w32985_
	);
	LUT3 #(
		.INIT('h43)
	) name27159 (
		_w32395_,
		_w32396_,
		_w32393_,
		_w32986_
	);
	LUT4 #(
		.INIT('h1005)
	) name27160 (
		_w32391_,
		_w32395_,
		_w32396_,
		_w32393_,
		_w32987_
	);
	LUT4 #(
		.INIT('h1011)
	) name27161 (
		_w32402_,
		_w32987_,
		_w32984_,
		_w32985_,
		_w32988_
	);
	LUT4 #(
		.INIT('h9060)
	) name27162 (
		_w32395_,
		_w32396_,
		_w32392_,
		_w32393_,
		_w32989_
	);
	LUT4 #(
		.INIT('h020a)
	) name27163 (
		_w32402_,
		_w32415_,
		_w32630_,
		_w32986_,
		_w32990_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name27164 (
		_w32983_,
		_w32988_,
		_w32989_,
		_w32990_,
		_w32991_
	);
	LUT3 #(
		.INIT('h40)
	) name27165 (
		_w32391_,
		_w32396_,
		_w32393_,
		_w32992_
	);
	LUT2 #(
		.INIT('h4)
	) name27166 (
		_w32403_,
		_w32992_,
		_w32993_
	);
	LUT3 #(
		.INIT('h56)
	) name27167 (
		\u0_L1_reg[9]/NET0131 ,
		_w32991_,
		_w32993_,
		_w32994_
	);
	LUT4 #(
		.INIT('h1a00)
	) name27168 (
		_w32655_,
		_w32656_,
		_w32657_,
		_w32653_,
		_w32995_
	);
	LUT3 #(
		.INIT('hac)
	) name27169 (
		_w32654_,
		_w32655_,
		_w32657_,
		_w32996_
	);
	LUT2 #(
		.INIT('h2)
	) name27170 (
		_w32656_,
		_w32653_,
		_w32997_
	);
	LUT4 #(
		.INIT('h2022)
	) name27171 (
		_w32652_,
		_w32768_,
		_w32996_,
		_w32997_,
		_w32998_
	);
	LUT4 #(
		.INIT('h8000)
	) name27172 (
		_w32655_,
		_w32656_,
		_w32657_,
		_w32653_,
		_w32999_
	);
	LUT4 #(
		.INIT('h00fe)
	) name27173 (
		_w32654_,
		_w32655_,
		_w32657_,
		_w32652_,
		_w33000_
	);
	LUT4 #(
		.INIT('h2080)
	) name27174 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32657_,
		_w33001_
	);
	LUT4 #(
		.INIT('h0109)
	) name27175 (
		_w32654_,
		_w32655_,
		_w32656_,
		_w32653_,
		_w33002_
	);
	LUT4 #(
		.INIT('h0100)
	) name27176 (
		_w32999_,
		_w33001_,
		_w33002_,
		_w33000_,
		_w33003_
	);
	LUT3 #(
		.INIT('h0b)
	) name27177 (
		_w32654_,
		_w32655_,
		_w32657_,
		_w33004_
	);
	LUT4 #(
		.INIT('h0020)
	) name27178 (
		_w32655_,
		_w32656_,
		_w32657_,
		_w32653_,
		_w33005_
	);
	LUT3 #(
		.INIT('h0d)
	) name27179 (
		_w32889_,
		_w33004_,
		_w33005_,
		_w33006_
	);
	LUT4 #(
		.INIT('hf400)
	) name27180 (
		_w32995_,
		_w32998_,
		_w33003_,
		_w33006_,
		_w33007_
	);
	LUT2 #(
		.INIT('h9)
	) name27181 (
		\u0_L1_reg[18]/NET0131 ,
		_w33007_,
		_w33008_
	);
	LUT4 #(
		.INIT('hc963)
	) name27182 (
		decrypt_pad,
		\u0_R0_reg[4]/NET0131 ,
		\u0_uk_K_r0_reg[20]/NET0131 ,
		\u0_uk_K_r0_reg[24]/P0001 ,
		_w33009_
	);
	LUT4 #(
		.INIT('hc963)
	) name27183 (
		decrypt_pad,
		\u0_R0_reg[1]/NET0131 ,
		\u0_uk_K_r0_reg[18]/NET0131 ,
		\u0_uk_K_r0_reg[54]/NET0131 ,
		_w33010_
	);
	LUT4 #(
		.INIT('hc693)
	) name27184 (
		decrypt_pad,
		\u0_R0_reg[32]/NET0131 ,
		\u0_uk_K_r0_reg[33]/NET0131 ,
		\u0_uk_K_r0_reg[54]/NET0131 ,
		_w33011_
	);
	LUT4 #(
		.INIT('hc693)
	) name27185 (
		decrypt_pad,
		\u0_R0_reg[2]/NET0131 ,
		\u0_uk_K_r0_reg[12]/NET0131 ,
		\u0_uk_K_r0_reg[33]/NET0131 ,
		_w33012_
	);
	LUT4 #(
		.INIT('hc963)
	) name27186 (
		decrypt_pad,
		\u0_R0_reg[3]/NET0131 ,
		\u0_uk_K_r0_reg[10]/NET0131 ,
		\u0_uk_K_r0_reg[46]/NET0131 ,
		_w33013_
	);
	LUT3 #(
		.INIT('h40)
	) name27187 (
		_w33011_,
		_w33012_,
		_w33013_,
		_w33014_
	);
	LUT4 #(
		.INIT('hc693)
	) name27188 (
		decrypt_pad,
		\u0_R0_reg[5]/NET0131 ,
		\u0_uk_K_r0_reg[27]/NET0131 ,
		\u0_uk_K_r0_reg[48]/NET0131 ,
		_w33015_
	);
	LUT4 #(
		.INIT('h4000)
	) name27189 (
		_w33011_,
		_w33012_,
		_w33013_,
		_w33015_,
		_w33016_
	);
	LUT4 #(
		.INIT('hbfee)
	) name27190 (
		_w33011_,
		_w33012_,
		_w33013_,
		_w33015_,
		_w33017_
	);
	LUT2 #(
		.INIT('h2)
	) name27191 (
		_w33010_,
		_w33017_,
		_w33018_
	);
	LUT2 #(
		.INIT('h9)
	) name27192 (
		_w33011_,
		_w33012_,
		_w33019_
	);
	LUT3 #(
		.INIT('h09)
	) name27193 (
		_w33011_,
		_w33012_,
		_w33013_,
		_w33020_
	);
	LUT3 #(
		.INIT('h47)
	) name27194 (
		_w33011_,
		_w33010_,
		_w33015_,
		_w33021_
	);
	LUT2 #(
		.INIT('h8)
	) name27195 (
		_w33020_,
		_w33021_,
		_w33022_
	);
	LUT4 #(
		.INIT('h0080)
	) name27196 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33023_
	);
	LUT4 #(
		.INIT('hdd7f)
	) name27197 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33024_
	);
	LUT4 #(
		.INIT('h0200)
	) name27198 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33025_
	);
	LUT3 #(
		.INIT('h0d)
	) name27199 (
		_w33013_,
		_w33024_,
		_w33025_,
		_w33026_
	);
	LUT4 #(
		.INIT('h5455)
	) name27200 (
		_w33009_,
		_w33022_,
		_w33018_,
		_w33026_,
		_w33027_
	);
	LUT4 #(
		.INIT('hf0bb)
	) name27201 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33028_
	);
	LUT2 #(
		.INIT('h2)
	) name27202 (
		_w33013_,
		_w33028_,
		_w33029_
	);
	LUT2 #(
		.INIT('h4)
	) name27203 (
		_w33012_,
		_w33013_,
		_w33030_
	);
	LUT3 #(
		.INIT('hb0)
	) name27204 (
		_w33012_,
		_w33013_,
		_w33010_,
		_w33031_
	);
	LUT2 #(
		.INIT('h4)
	) name27205 (
		_w33011_,
		_w33015_,
		_w33032_
	);
	LUT2 #(
		.INIT('h4)
	) name27206 (
		_w33013_,
		_w33010_,
		_w33033_
	);
	LUT4 #(
		.INIT('h0a44)
	) name27207 (
		_w33011_,
		_w33012_,
		_w33013_,
		_w33010_,
		_w33034_
	);
	LUT2 #(
		.INIT('h1)
	) name27208 (
		_w33010_,
		_w33015_,
		_w33035_
	);
	LUT4 #(
		.INIT('h0002)
	) name27209 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33036_
	);
	LUT4 #(
		.INIT('h1011)
	) name27210 (
		_w33034_,
		_w33036_,
		_w33031_,
		_w33032_,
		_w33037_
	);
	LUT3 #(
		.INIT('h8a)
	) name27211 (
		_w33009_,
		_w33029_,
		_w33037_,
		_w33038_
	);
	LUT3 #(
		.INIT('h80)
	) name27212 (
		_w33011_,
		_w33012_,
		_w33015_,
		_w33039_
	);
	LUT4 #(
		.INIT('h0400)
	) name27213 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33040_
	);
	LUT4 #(
		.INIT('h7bcf)
	) name27214 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33041_
	);
	LUT2 #(
		.INIT('h1)
	) name27215 (
		_w33013_,
		_w33041_,
		_w33042_
	);
	LUT4 #(
		.INIT('h0020)
	) name27216 (
		_w33011_,
		_w33012_,
		_w33013_,
		_w33010_,
		_w33043_
	);
	LUT3 #(
		.INIT('h07)
	) name27217 (
		_w33014_,
		_w33035_,
		_w33043_,
		_w33044_
	);
	LUT2 #(
		.INIT('h4)
	) name27218 (
		_w33042_,
		_w33044_,
		_w33045_
	);
	LUT4 #(
		.INIT('h5655)
	) name27219 (
		\u0_L0_reg[31]/NET0131 ,
		_w33027_,
		_w33038_,
		_w33045_,
		_w33046_
	);
	LUT4 #(
		.INIT('hc693)
	) name27220 (
		decrypt_pad,
		\u0_R0_reg[24]/NET0131 ,
		\u0_uk_K_r0_reg[21]/NET0131 ,
		\u0_uk_K_r0_reg[42]/NET0131 ,
		_w33047_
	);
	LUT4 #(
		.INIT('hc963)
	) name27221 (
		decrypt_pad,
		\u0_R0_reg[22]/NET0131 ,
		\u0_uk_K_r0_reg[31]/NET0131 ,
		\u0_uk_K_r0_reg[37]/NET0131 ,
		_w33048_
	);
	LUT4 #(
		.INIT('hc693)
	) name27222 (
		decrypt_pad,
		\u0_R0_reg[21]/NET0131 ,
		\u0_uk_K_r0_reg[15]/NET0131 ,
		\u0_uk_K_r0_reg[36]/NET0131 ,
		_w33049_
	);
	LUT4 #(
		.INIT('hc693)
	) name27223 (
		decrypt_pad,
		\u0_R0_reg[20]/NET0131 ,
		\u0_uk_K_r0_reg[0]/NET0131 ,
		\u0_uk_K_r0_reg[21]/NET0131 ,
		_w33050_
	);
	LUT4 #(
		.INIT('hc693)
	) name27224 (
		decrypt_pad,
		\u0_R0_reg[25]/NET0131 ,
		\u0_uk_K_r0_reg[16]/NET0131 ,
		\u0_uk_K_r0_reg[37]/NET0131 ,
		_w33051_
	);
	LUT4 #(
		.INIT('he020)
	) name27225 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33052_
	);
	LUT4 #(
		.INIT('hc963)
	) name27226 (
		decrypt_pad,
		\u0_R0_reg[23]/NET0131 ,
		\u0_uk_K_r0_reg[16]/NET0131 ,
		\u0_uk_K_r0_reg[50]/NET0131 ,
		_w33053_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name27227 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33054_
	);
	LUT3 #(
		.INIT('h01)
	) name27228 (
		_w33053_,
		_w33054_,
		_w33052_,
		_w33055_
	);
	LUT4 #(
		.INIT('h0004)
	) name27229 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33056_
	);
	LUT4 #(
		.INIT('h57db)
	) name27230 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33057_
	);
	LUT2 #(
		.INIT('h1)
	) name27231 (
		_w33048_,
		_w33053_,
		_w33058_
	);
	LUT4 #(
		.INIT('h0200)
	) name27232 (
		_w33050_,
		_w33048_,
		_w33053_,
		_w33051_,
		_w33059_
	);
	LUT2 #(
		.INIT('h4)
	) name27233 (
		_w33049_,
		_w33059_,
		_w33060_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name27234 (
		_w33049_,
		_w33053_,
		_w33057_,
		_w33059_,
		_w33061_
	);
	LUT3 #(
		.INIT('h8a)
	) name27235 (
		_w33047_,
		_w33055_,
		_w33061_,
		_w33062_
	);
	LUT4 #(
		.INIT('h0028)
	) name27236 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33053_,
		_w33063_
	);
	LUT3 #(
		.INIT('hd0)
	) name27237 (
		_w33050_,
		_w33048_,
		_w33053_,
		_w33064_
	);
	LUT3 #(
		.INIT('h54)
	) name27238 (
		_w33049_,
		_w33050_,
		_w33051_,
		_w33065_
	);
	LUT2 #(
		.INIT('h8)
	) name27239 (
		_w33064_,
		_w33065_,
		_w33066_
	);
	LUT3 #(
		.INIT('hc4)
	) name27240 (
		_w33049_,
		_w33050_,
		_w33051_,
		_w33067_
	);
	LUT3 #(
		.INIT('h32)
	) name27241 (
		_w33050_,
		_w33048_,
		_w33053_,
		_w33068_
	);
	LUT4 #(
		.INIT('h0002)
	) name27242 (
		_w33050_,
		_w33048_,
		_w33053_,
		_w33051_,
		_w33069_
	);
	LUT4 #(
		.INIT('h4000)
	) name27243 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33070_
	);
	LUT4 #(
		.INIT('h000b)
	) name27244 (
		_w33067_,
		_w33068_,
		_w33069_,
		_w33070_,
		_w33071_
	);
	LUT4 #(
		.INIT('h00ef)
	) name27245 (
		_w33063_,
		_w33066_,
		_w33071_,
		_w33047_,
		_w33072_
	);
	LUT3 #(
		.INIT('h02)
	) name27246 (
		_w33049_,
		_w33048_,
		_w33051_,
		_w33073_
	);
	LUT4 #(
		.INIT('h33f5)
	) name27247 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33074_
	);
	LUT2 #(
		.INIT('h2)
	) name27248 (
		_w33064_,
		_w33074_,
		_w33075_
	);
	LUT3 #(
		.INIT('h01)
	) name27249 (
		_w33049_,
		_w33050_,
		_w33051_,
		_w33076_
	);
	LUT2 #(
		.INIT('h8)
	) name27250 (
		_w33058_,
		_w33076_,
		_w33077_
	);
	LUT4 #(
		.INIT('h0100)
	) name27251 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33078_
	);
	LUT3 #(
		.INIT('h08)
	) name27252 (
		_w33049_,
		_w33050_,
		_w33051_,
		_w33079_
	);
	LUT4 #(
		.INIT('h2e3f)
	) name27253 (
		_w33048_,
		_w33053_,
		_w33078_,
		_w33079_,
		_w33080_
	);
	LUT3 #(
		.INIT('h04)
	) name27254 (
		_w33077_,
		_w33080_,
		_w33075_,
		_w33081_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name27255 (
		\u0_L0_reg[11]/NET0131 ,
		_w33072_,
		_w33062_,
		_w33081_,
		_w33082_
	);
	LUT4 #(
		.INIT('hc693)
	) name27256 (
		decrypt_pad,
		\u0_R0_reg[28]/NET0131 ,
		\u0_uk_K_r0_reg[28]/NET0131 ,
		\u0_uk_K_r0_reg[49]/NET0131 ,
		_w33083_
	);
	LUT4 #(
		.INIT('hc693)
	) name27257 (
		decrypt_pad,
		\u0_R0_reg[27]/NET0131 ,
		\u0_uk_K_r0_reg[45]/NET0131 ,
		\u0_uk_K_r0_reg[7]/NET0131 ,
		_w33084_
	);
	LUT4 #(
		.INIT('hc963)
	) name27258 (
		decrypt_pad,
		\u0_R0_reg[26]/NET0131 ,
		\u0_uk_K_r0_reg[29]/NET0131 ,
		\u0_uk_K_r0_reg[8]/NET0131 ,
		_w33085_
	);
	LUT4 #(
		.INIT('hc693)
	) name27259 (
		decrypt_pad,
		\u0_R0_reg[24]/NET0131 ,
		\u0_uk_K_r0_reg[43]/NET0131 ,
		\u0_uk_K_r0_reg[9]/NET0131 ,
		_w33086_
	);
	LUT4 #(
		.INIT('hc963)
	) name27260 (
		decrypt_pad,
		\u0_R0_reg[29]/NET0131 ,
		\u0_uk_K_r0_reg[45]/NET0131 ,
		\u0_uk_K_r0_reg[51]/NET0131 ,
		_w33087_
	);
	LUT4 #(
		.INIT('hc693)
	) name27261 (
		decrypt_pad,
		\u0_R0_reg[25]/NET0131 ,
		\u0_uk_K_r0_reg[23]/NET0131 ,
		\u0_uk_K_r0_reg[44]/NET0131 ,
		_w33088_
	);
	LUT4 #(
		.INIT('h737d)
	) name27262 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33089_
	);
	LUT2 #(
		.INIT('h1)
	) name27263 (
		_w33084_,
		_w33089_,
		_w33090_
	);
	LUT4 #(
		.INIT('h9000)
	) name27264 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33091_
	);
	LUT4 #(
		.INIT('hf5b9)
	) name27265 (
		_w33086_,
		_w33087_,
		_w33088_,
		_w33084_,
		_w33092_
	);
	LUT3 #(
		.INIT('h32)
	) name27266 (
		_w33085_,
		_w33091_,
		_w33092_,
		_w33093_
	);
	LUT3 #(
		.INIT('h45)
	) name27267 (
		_w33083_,
		_w33090_,
		_w33093_,
		_w33094_
	);
	LUT4 #(
		.INIT('h0040)
	) name27268 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33095_
	);
	LUT4 #(
		.INIT('hcfbf)
	) name27269 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33096_
	);
	LUT2 #(
		.INIT('h1)
	) name27270 (
		_w33084_,
		_w33096_,
		_w33097_
	);
	LUT2 #(
		.INIT('h6)
	) name27271 (
		_w33085_,
		_w33088_,
		_w33098_
	);
	LUT2 #(
		.INIT('h8)
	) name27272 (
		_w33086_,
		_w33084_,
		_w33099_
	);
	LUT4 #(
		.INIT('hc800)
	) name27273 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33084_,
		_w33100_
	);
	LUT2 #(
		.INIT('h2)
	) name27274 (
		_w33085_,
		_w33088_,
		_w33101_
	);
	LUT4 #(
		.INIT('hffde)
	) name27275 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33102_
	);
	LUT3 #(
		.INIT('h70)
	) name27276 (
		_w33098_,
		_w33100_,
		_w33102_,
		_w33103_
	);
	LUT4 #(
		.INIT('h0200)
	) name27277 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33104_
	);
	LUT4 #(
		.INIT('hfdd3)
	) name27278 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33105_
	);
	LUT4 #(
		.INIT('h0090)
	) name27279 (
		_w33085_,
		_w33086_,
		_w33088_,
		_w33084_,
		_w33106_
	);
	LUT4 #(
		.INIT('h0100)
	) name27280 (
		_w33085_,
		_w33087_,
		_w33088_,
		_w33084_,
		_w33107_
	);
	LUT4 #(
		.INIT('h0031)
	) name27281 (
		_w33084_,
		_w33106_,
		_w33105_,
		_w33107_,
		_w33108_
	);
	LUT4 #(
		.INIT('h7500)
	) name27282 (
		_w33083_,
		_w33097_,
		_w33103_,
		_w33108_,
		_w33109_
	);
	LUT3 #(
		.INIT('h65)
	) name27283 (
		\u0_L0_reg[22]/NET0131 ,
		_w33094_,
		_w33109_,
		_w33110_
	);
	LUT2 #(
		.INIT('h9)
	) name27284 (
		_w33012_,
		_w33015_,
		_w33111_
	);
	LUT3 #(
		.INIT('h40)
	) name27285 (
		_w33011_,
		_w33013_,
		_w33010_,
		_w33112_
	);
	LUT2 #(
		.INIT('h4)
	) name27286 (
		_w33111_,
		_w33112_,
		_w33113_
	);
	LUT4 #(
		.INIT('h0809)
	) name27287 (
		_w33011_,
		_w33012_,
		_w33013_,
		_w33010_,
		_w33114_
	);
	LUT4 #(
		.INIT('ha9ab)
	) name27288 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33115_
	);
	LUT4 #(
		.INIT('hc020)
	) name27289 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33116_
	);
	LUT4 #(
		.INIT('h00c4)
	) name27290 (
		_w33013_,
		_w33009_,
		_w33115_,
		_w33116_,
		_w33117_
	);
	LUT4 #(
		.INIT('hf5ea)
	) name27291 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33118_
	);
	LUT2 #(
		.INIT('h1)
	) name27292 (
		_w33013_,
		_w33118_,
		_w33119_
	);
	LUT4 #(
		.INIT('h8008)
	) name27293 (
		_w33011_,
		_w33013_,
		_w33010_,
		_w33015_,
		_w33120_
	);
	LUT4 #(
		.INIT('h0001)
	) name27294 (
		_w33009_,
		_w33023_,
		_w33040_,
		_w33120_,
		_w33121_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name27295 (
		_w33114_,
		_w33117_,
		_w33119_,
		_w33121_,
		_w33122_
	);
	LUT3 #(
		.INIT('h56)
	) name27296 (
		\u0_L0_reg[17]/NET0131 ,
		_w33113_,
		_w33122_,
		_w33123_
	);
	LUT4 #(
		.INIT('hbc77)
	) name27297 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33124_
	);
	LUT2 #(
		.INIT('h2)
	) name27298 (
		_w33053_,
		_w33124_,
		_w33125_
	);
	LUT4 #(
		.INIT('h1000)
	) name27299 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33126_
	);
	LUT4 #(
		.INIT('hefdd)
	) name27300 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33127_
	);
	LUT4 #(
		.INIT('h0302)
	) name27301 (
		_w33053_,
		_w33056_,
		_w33059_,
		_w33127_,
		_w33128_
	);
	LUT3 #(
		.INIT('h45)
	) name27302 (
		_w33047_,
		_w33125_,
		_w33128_,
		_w33129_
	);
	LUT2 #(
		.INIT('h4)
	) name27303 (
		_w33067_,
		_w33058_,
		_w33130_
	);
	LUT4 #(
		.INIT('h0002)
	) name27304 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33131_
	);
	LUT4 #(
		.INIT('h2000)
	) name27305 (
		_w33050_,
		_w33048_,
		_w33053_,
		_w33051_,
		_w33132_
	);
	LUT3 #(
		.INIT('h80)
	) name27306 (
		_w33049_,
		_w33048_,
		_w33051_,
		_w33133_
	);
	LUT3 #(
		.INIT('h01)
	) name27307 (
		_w33132_,
		_w33131_,
		_w33133_,
		_w33134_
	);
	LUT4 #(
		.INIT('hd060)
	) name27308 (
		_w33049_,
		_w33050_,
		_w33053_,
		_w33051_,
		_w33135_
	);
	LUT4 #(
		.INIT('h070b)
	) name27309 (
		_w33049_,
		_w33050_,
		_w33053_,
		_w33051_,
		_w33136_
	);
	LUT4 #(
		.INIT('h0001)
	) name27310 (
		_w33050_,
		_w33048_,
		_w33053_,
		_w33051_,
		_w33137_
	);
	LUT4 #(
		.INIT('h00fd)
	) name27311 (
		_w33048_,
		_w33136_,
		_w33135_,
		_w33137_,
		_w33138_
	);
	LUT4 #(
		.INIT('h7500)
	) name27312 (
		_w33047_,
		_w33130_,
		_w33134_,
		_w33138_,
		_w33139_
	);
	LUT3 #(
		.INIT('h65)
	) name27313 (
		\u0_L0_reg[4]/NET0131 ,
		_w33129_,
		_w33139_,
		_w33140_
	);
	LUT4 #(
		.INIT('hc693)
	) name27314 (
		decrypt_pad,
		\u0_R0_reg[15]/NET0131 ,
		\u0_uk_K_r0_reg[18]/NET0131 ,
		\u0_uk_K_r0_reg[39]/NET0131 ,
		_w33141_
	);
	LUT4 #(
		.INIT('hc963)
	) name27315 (
		decrypt_pad,
		\u0_R0_reg[17]/NET0131 ,
		\u0_uk_K_r0_reg[27]/NET0131 ,
		\u0_uk_K_r0_reg[6]/NET0131 ,
		_w33142_
	);
	LUT4 #(
		.INIT('hc693)
	) name27316 (
		decrypt_pad,
		\u0_R0_reg[14]/NET0131 ,
		\u0_uk_K_r0_reg[10]/NET0131 ,
		\u0_uk_K_r0_reg[6]/NET0131 ,
		_w33143_
	);
	LUT4 #(
		.INIT('hc963)
	) name27317 (
		decrypt_pad,
		\u0_R0_reg[12]/NET0131 ,
		\u0_uk_K_r0_reg[11]/NET0131 ,
		\u0_uk_K_r0_reg[47]/NET0131 ,
		_w33144_
	);
	LUT4 #(
		.INIT('hc693)
	) name27318 (
		decrypt_pad,
		\u0_R0_reg[13]/NET0131 ,
		\u0_uk_K_r0_reg[41]/NET0131 ,
		\u0_uk_K_r0_reg[5]/NET0131 ,
		_w33145_
	);
	LUT2 #(
		.INIT('h4)
	) name27319 (
		_w33144_,
		_w33145_,
		_w33146_
	);
	LUT4 #(
		.INIT('hfec3)
	) name27320 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33147_
	);
	LUT2 #(
		.INIT('h1)
	) name27321 (
		_w33141_,
		_w33147_,
		_w33148_
	);
	LUT4 #(
		.INIT('h0020)
	) name27322 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33149_
	);
	LUT4 #(
		.INIT('h4000)
	) name27323 (
		_w33142_,
		_w33144_,
		_w33141_,
		_w33145_,
		_w33150_
	);
	LUT2 #(
		.INIT('h1)
	) name27324 (
		_w33149_,
		_w33150_,
		_w33151_
	);
	LUT4 #(
		.INIT('h8000)
	) name27325 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33152_
	);
	LUT4 #(
		.INIT('h0020)
	) name27326 (
		_w33142_,
		_w33144_,
		_w33141_,
		_w33145_,
		_w33153_
	);
	LUT4 #(
		.INIT('hc693)
	) name27327 (
		decrypt_pad,
		\u0_R0_reg[16]/NET0131 ,
		\u0_uk_K_r0_reg[26]/NET0131 ,
		\u0_uk_K_r0_reg[47]/NET0131 ,
		_w33154_
	);
	LUT3 #(
		.INIT('h10)
	) name27328 (
		_w33153_,
		_w33152_,
		_w33154_,
		_w33155_
	);
	LUT3 #(
		.INIT('h20)
	) name27329 (
		_w33151_,
		_w33148_,
		_w33155_,
		_w33156_
	);
	LUT4 #(
		.INIT('h0008)
	) name27330 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33157_
	);
	LUT4 #(
		.INIT('h1000)
	) name27331 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33158_
	);
	LUT4 #(
		.INIT('heff6)
	) name27332 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33159_
	);
	LUT4 #(
		.INIT('hb1f5)
	) name27333 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33160_
	);
	LUT2 #(
		.INIT('h1)
	) name27334 (
		_w33141_,
		_w33160_,
		_w33161_
	);
	LUT2 #(
		.INIT('h2)
	) name27335 (
		_w33141_,
		_w33145_,
		_w33162_
	);
	LUT4 #(
		.INIT('h0010)
	) name27336 (
		_w33142_,
		_w33144_,
		_w33141_,
		_w33145_,
		_w33163_
	);
	LUT4 #(
		.INIT('h8000)
	) name27337 (
		_w33142_,
		_w33144_,
		_w33141_,
		_w33145_,
		_w33164_
	);
	LUT2 #(
		.INIT('h8)
	) name27338 (
		_w33141_,
		_w33143_,
		_w33165_
	);
	LUT4 #(
		.INIT('h4000)
	) name27339 (
		_w33144_,
		_w33141_,
		_w33145_,
		_w33143_,
		_w33166_
	);
	LUT4 #(
		.INIT('h0001)
	) name27340 (
		_w33154_,
		_w33163_,
		_w33164_,
		_w33166_,
		_w33167_
	);
	LUT3 #(
		.INIT('h40)
	) name27341 (
		_w33161_,
		_w33167_,
		_w33159_,
		_w33168_
	);
	LUT3 #(
		.INIT('hbe)
	) name27342 (
		_w33142_,
		_w33144_,
		_w33143_,
		_w33169_
	);
	LUT2 #(
		.INIT('h2)
	) name27343 (
		_w33162_,
		_w33169_,
		_w33170_
	);
	LUT2 #(
		.INIT('h2)
	) name27344 (
		_w33142_,
		_w33143_,
		_w33171_
	);
	LUT3 #(
		.INIT('h02)
	) name27345 (
		_w33142_,
		_w33141_,
		_w33143_,
		_w33172_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name27346 (
		_w33143_,
		_w33150_,
		_w33146_,
		_w33172_,
		_w33173_
	);
	LUT2 #(
		.INIT('h4)
	) name27347 (
		_w33170_,
		_w33173_,
		_w33174_
	);
	LUT4 #(
		.INIT('ha955)
	) name27348 (
		\u0_L0_reg[20]/NET0131 ,
		_w33156_,
		_w33168_,
		_w33174_,
		_w33175_
	);
	LUT4 #(
		.INIT('h779a)
	) name27349 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33176_
	);
	LUT4 #(
		.INIT('hf17d)
	) name27350 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33177_
	);
	LUT4 #(
		.INIT('h3120)
	) name27351 (
		_w33053_,
		_w33126_,
		_w33176_,
		_w33177_,
		_w33178_
	);
	LUT2 #(
		.INIT('h1)
	) name27352 (
		_w33047_,
		_w33178_,
		_w33179_
	);
	LUT4 #(
		.INIT('hdd7d)
	) name27353 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33180_
	);
	LUT2 #(
		.INIT('h2)
	) name27354 (
		_w33053_,
		_w33180_,
		_w33181_
	);
	LUT4 #(
		.INIT('h3fce)
	) name27355 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33182_
	);
	LUT2 #(
		.INIT('h1)
	) name27356 (
		_w33053_,
		_w33182_,
		_w33183_
	);
	LUT4 #(
		.INIT('h0010)
	) name27357 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33184_
	);
	LUT4 #(
		.INIT('h0001)
	) name27358 (
		_w33069_,
		_w33070_,
		_w33078_,
		_w33184_,
		_w33185_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name27359 (
		_w33047_,
		_w33183_,
		_w33181_,
		_w33185_,
		_w33186_
	);
	LUT4 #(
		.INIT('h2000)
	) name27360 (
		_w33049_,
		_w33048_,
		_w33053_,
		_w33051_,
		_w33187_
	);
	LUT2 #(
		.INIT('h1)
	) name27361 (
		_w33056_,
		_w33187_,
		_w33188_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name27362 (
		\u0_L0_reg[29]/NET0131 ,
		_w33186_,
		_w33179_,
		_w33188_,
		_w33189_
	);
	LUT4 #(
		.INIT('hc693)
	) name27363 (
		decrypt_pad,
		\u0_R0_reg[7]/NET0131 ,
		\u0_uk_K_r0_reg[34]/NET0131 ,
		\u0_uk_K_r0_reg[55]/NET0131 ,
		_w33190_
	);
	LUT4 #(
		.INIT('hc963)
	) name27364 (
		decrypt_pad,
		\u0_R0_reg[5]/NET0131 ,
		\u0_uk_K_r0_reg[13]/NET0131 ,
		\u0_uk_K_r0_reg[17]/NET0131 ,
		_w33191_
	);
	LUT4 #(
		.INIT('hc693)
	) name27365 (
		decrypt_pad,
		\u0_R0_reg[6]/NET0131 ,
		\u0_uk_K_r0_reg[40]/NET0131 ,
		\u0_uk_K_r0_reg[4]/NET0131 ,
		_w33192_
	);
	LUT4 #(
		.INIT('hc963)
	) name27366 (
		decrypt_pad,
		\u0_R0_reg[9]/NET0131 ,
		\u0_uk_K_r0_reg[26]/NET0131 ,
		\u0_uk_K_r0_reg[5]/NET0131 ,
		_w33193_
	);
	LUT4 #(
		.INIT('hc693)
	) name27367 (
		decrypt_pad,
		\u0_R0_reg[4]/NET0131 ,
		\u0_uk_K_r0_reg[13]/NET0131 ,
		\u0_uk_K_r0_reg[34]/NET0131 ,
		_w33194_
	);
	LUT4 #(
		.INIT('h2000)
	) name27368 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33195_
	);
	LUT2 #(
		.INIT('h8)
	) name27369 (
		_w33190_,
		_w33195_,
		_w33196_
	);
	LUT4 #(
		.INIT('h0080)
	) name27370 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33197_
	);
	LUT4 #(
		.INIT('h0004)
	) name27371 (
		_w33190_,
		_w33193_,
		_w33191_,
		_w33192_,
		_w33198_
	);
	LUT4 #(
		.INIT('hc693)
	) name27372 (
		decrypt_pad,
		\u0_R0_reg[8]/NET0131 ,
		\u0_uk_K_r0_reg[25]/P0001 ,
		\u0_uk_K_r0_reg[46]/NET0131 ,
		_w33199_
	);
	LUT3 #(
		.INIT('h01)
	) name27373 (
		_w33197_,
		_w33198_,
		_w33199_,
		_w33200_
	);
	LUT3 #(
		.INIT('h02)
	) name27374 (
		_w33193_,
		_w33191_,
		_w33194_,
		_w33201_
	);
	LUT4 #(
		.INIT('h2fdd)
	) name27375 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33202_
	);
	LUT4 #(
		.INIT('h0406)
	) name27376 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33203_
	);
	LUT3 #(
		.INIT('h0e)
	) name27377 (
		_w33190_,
		_w33202_,
		_w33203_,
		_w33204_
	);
	LUT2 #(
		.INIT('h1)
	) name27378 (
		_w33193_,
		_w33192_,
		_w33205_
	);
	LUT4 #(
		.INIT('h0100)
	) name27379 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33206_
	);
	LUT2 #(
		.INIT('h4)
	) name27380 (
		_w33192_,
		_w33194_,
		_w33207_
	);
	LUT4 #(
		.INIT('h0800)
	) name27381 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33208_
	);
	LUT4 #(
		.INIT('h8808)
	) name27382 (
		_w33190_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33209_
	);
	LUT4 #(
		.INIT('h0002)
	) name27383 (
		_w33199_,
		_w33208_,
		_w33206_,
		_w33209_,
		_w33210_
	);
	LUT4 #(
		.INIT('h00bf)
	) name27384 (
		_w33196_,
		_w33200_,
		_w33204_,
		_w33210_,
		_w33211_
	);
	LUT4 #(
		.INIT('h0010)
	) name27385 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33212_
	);
	LUT4 #(
		.INIT('hf3ef)
	) name27386 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33213_
	);
	LUT2 #(
		.INIT('h2)
	) name27387 (
		_w33190_,
		_w33213_,
		_w33214_
	);
	LUT4 #(
		.INIT('h008a)
	) name27388 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33215_
	);
	LUT3 #(
		.INIT('hb0)
	) name27389 (
		_w33191_,
		_w33192_,
		_w33194_,
		_w33216_
	);
	LUT3 #(
		.INIT('h90)
	) name27390 (
		_w33193_,
		_w33194_,
		_w33199_,
		_w33217_
	);
	LUT3 #(
		.INIT('h51)
	) name27391 (
		_w33190_,
		_w33191_,
		_w33192_,
		_w33218_
	);
	LUT4 #(
		.INIT('hba00)
	) name27392 (
		_w33215_,
		_w33216_,
		_w33217_,
		_w33218_,
		_w33219_
	);
	LUT2 #(
		.INIT('h1)
	) name27393 (
		_w33214_,
		_w33219_,
		_w33220_
	);
	LUT3 #(
		.INIT('h65)
	) name27394 (
		\u0_L0_reg[2]/NET0131 ,
		_w33211_,
		_w33220_,
		_w33221_
	);
	LUT4 #(
		.INIT('hc963)
	) name27395 (
		decrypt_pad,
		\u0_R0_reg[32]/NET0131 ,
		\u0_uk_K_r0_reg[14]/NET0131 ,
		\u0_uk_K_r0_reg[52]/NET0131 ,
		_w33222_
	);
	LUT4 #(
		.INIT('hc693)
	) name27396 (
		decrypt_pad,
		\u0_R0_reg[31]/NET0131 ,
		\u0_uk_K_r0_reg[42]/NET0131 ,
		\u0_uk_K_r0_reg[8]/NET0131 ,
		_w33223_
	);
	LUT4 #(
		.INIT('hc693)
	) name27397 (
		decrypt_pad,
		\u0_R0_reg[30]/NET0131 ,
		\u0_uk_K_r0_reg[30]/NET0131 ,
		\u0_uk_K_r0_reg[51]/NET0131 ,
		_w33224_
	);
	LUT4 #(
		.INIT('hc963)
	) name27398 (
		decrypt_pad,
		\u0_R0_reg[28]/NET0131 ,
		\u0_uk_K_r0_reg[23]/NET0131 ,
		\u0_uk_K_r0_reg[2]/NET0131 ,
		_w33225_
	);
	LUT4 #(
		.INIT('hc693)
	) name27399 (
		decrypt_pad,
		\u0_R0_reg[1]/NET0131 ,
		\u0_uk_K_r0_reg[14]/NET0131 ,
		\u0_uk_K_r0_reg[35]/NET0131 ,
		_w33226_
	);
	LUT4 #(
		.INIT('hc693)
	) name27400 (
		decrypt_pad,
		\u0_R0_reg[29]/NET0131 ,
		\u0_uk_K_r0_reg[29]/NET0131 ,
		\u0_uk_K_r0_reg[50]/NET0131 ,
		_w33227_
	);
	LUT4 #(
		.INIT('h23a5)
	) name27401 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33228_
	);
	LUT4 #(
		.INIT('h0020)
	) name27402 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33229_
	);
	LUT4 #(
		.INIT('hfcdf)
	) name27403 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33230_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name27404 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33231_
	);
	LUT4 #(
		.INIT('he400)
	) name27405 (
		_w33223_,
		_w33228_,
		_w33230_,
		_w33231_,
		_w33232_
	);
	LUT3 #(
		.INIT('h01)
	) name27406 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33233_
	);
	LUT4 #(
		.INIT('h509c)
	) name27407 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33234_
	);
	LUT4 #(
		.INIT('h0800)
	) name27408 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33235_
	);
	LUT4 #(
		.INIT('h001d)
	) name27409 (
		_w33233_,
		_w33223_,
		_w33234_,
		_w33235_,
		_w33236_
	);
	LUT4 #(
		.INIT('h0009)
	) name27410 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33237_
	);
	LUT4 #(
		.INIT('hedf6)
	) name27411 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33238_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name27412 (
		_w33224_,
		_w33227_,
		_w33226_,
		_w33222_,
		_w33239_
	);
	LUT4 #(
		.INIT('hf3d1)
	) name27413 (
		_w33225_,
		_w33223_,
		_w33238_,
		_w33239_,
		_w33240_
	);
	LUT4 #(
		.INIT('hb800)
	) name27414 (
		_w33236_,
		_w33222_,
		_w33232_,
		_w33240_,
		_w33241_
	);
	LUT2 #(
		.INIT('h6)
	) name27415 (
		\u0_L0_reg[5]/NET0131 ,
		_w33241_,
		_w33242_
	);
	LUT4 #(
		.INIT('h9d81)
	) name27416 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33243_
	);
	LUT4 #(
		.INIT('h6000)
	) name27417 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33244_
	);
	LUT3 #(
		.INIT('h04)
	) name27418 (
		_w33224_,
		_w33225_,
		_w33226_,
		_w33245_
	);
	LUT4 #(
		.INIT('hddd8)
	) name27419 (
		_w33223_,
		_w33243_,
		_w33244_,
		_w33245_,
		_w33246_
	);
	LUT4 #(
		.INIT('h0082)
	) name27420 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33247_
	);
	LUT4 #(
		.INIT('h0100)
	) name27421 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33248_
	);
	LUT3 #(
		.INIT('h02)
	) name27422 (
		_w33222_,
		_w33247_,
		_w33248_,
		_w33249_
	);
	LUT2 #(
		.INIT('h4)
	) name27423 (
		_w33246_,
		_w33249_,
		_w33250_
	);
	LUT4 #(
		.INIT('hde1e)
	) name27424 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33251_
	);
	LUT2 #(
		.INIT('h2)
	) name27425 (
		_w33223_,
		_w33251_,
		_w33252_
	);
	LUT4 #(
		.INIT('hf3ee)
	) name27426 (
		_w33227_,
		_w33225_,
		_w33223_,
		_w33226_,
		_w33253_
	);
	LUT2 #(
		.INIT('h1)
	) name27427 (
		_w33224_,
		_w33253_,
		_w33254_
	);
	LUT4 #(
		.INIT('h00f7)
	) name27428 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33222_,
		_w33255_
	);
	LUT4 #(
		.INIT('h0200)
	) name27429 (
		_w33224_,
		_w33225_,
		_w33223_,
		_w33226_,
		_w33256_
	);
	LUT4 #(
		.INIT('h0002)
	) name27430 (
		_w33227_,
		_w33225_,
		_w33223_,
		_w33226_,
		_w33257_
	);
	LUT4 #(
		.INIT('h4000)
	) name27431 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33258_
	);
	LUT4 #(
		.INIT('h0001)
	) name27432 (
		_w33229_,
		_w33256_,
		_w33257_,
		_w33258_,
		_w33259_
	);
	LUT4 #(
		.INIT('h1000)
	) name27433 (
		_w33254_,
		_w33252_,
		_w33255_,
		_w33259_,
		_w33260_
	);
	LUT3 #(
		.INIT('ha9)
	) name27434 (
		\u0_L0_reg[21]/NET0131 ,
		_w33250_,
		_w33260_,
		_w33261_
	);
	LUT4 #(
		.INIT('h1000)
	) name27435 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33262_
	);
	LUT4 #(
		.INIT('h0002)
	) name27436 (
		_w33083_,
		_w33095_,
		_w33104_,
		_w33262_,
		_w33263_
	);
	LUT3 #(
		.INIT('hd9)
	) name27437 (
		_w33086_,
		_w33087_,
		_w33084_,
		_w33264_
	);
	LUT4 #(
		.INIT('h33fe)
	) name27438 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33265_
	);
	LUT4 #(
		.INIT('hf351)
	) name27439 (
		_w33084_,
		_w33101_,
		_w33264_,
		_w33265_,
		_w33266_
	);
	LUT2 #(
		.INIT('h8)
	) name27440 (
		_w33263_,
		_w33266_,
		_w33267_
	);
	LUT3 #(
		.INIT('h15)
	) name27441 (
		_w33086_,
		_w33087_,
		_w33088_,
		_w33268_
	);
	LUT4 #(
		.INIT('ha200)
	) name27442 (
		_w33086_,
		_w33087_,
		_w33088_,
		_w33084_,
		_w33269_
	);
	LUT3 #(
		.INIT('h02)
	) name27443 (
		_w33085_,
		_w33269_,
		_w33268_,
		_w33270_
	);
	LUT4 #(
		.INIT('h0400)
	) name27444 (
		_w33086_,
		_w33087_,
		_w33088_,
		_w33084_,
		_w33271_
	);
	LUT4 #(
		.INIT('h0004)
	) name27445 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33272_
	);
	LUT3 #(
		.INIT('h01)
	) name27446 (
		_w33083_,
		_w33272_,
		_w33271_,
		_w33273_
	);
	LUT3 #(
		.INIT('h09)
	) name27447 (
		_w33087_,
		_w33088_,
		_w33084_,
		_w33274_
	);
	LUT4 #(
		.INIT('h0102)
	) name27448 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33275_
	);
	LUT2 #(
		.INIT('h1)
	) name27449 (
		_w33274_,
		_w33275_,
		_w33276_
	);
	LUT3 #(
		.INIT('h40)
	) name27450 (
		_w33270_,
		_w33273_,
		_w33276_,
		_w33277_
	);
	LUT3 #(
		.INIT('ha9)
	) name27451 (
		\u0_L0_reg[12]/NET0131 ,
		_w33267_,
		_w33277_,
		_w33278_
	);
	LUT4 #(
		.INIT('h575f)
	) name27452 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33279_
	);
	LUT2 #(
		.INIT('h1)
	) name27453 (
		_w33013_,
		_w33279_,
		_w33280_
	);
	LUT4 #(
		.INIT('h0040)
	) name27454 (
		_w33011_,
		_w33013_,
		_w33010_,
		_w33015_,
		_w33281_
	);
	LUT3 #(
		.INIT('h81)
	) name27455 (
		_w33012_,
		_w33010_,
		_w33015_,
		_w33282_
	);
	LUT4 #(
		.INIT('h0001)
	) name27456 (
		_w33009_,
		_w33016_,
		_w33281_,
		_w33282_,
		_w33283_
	);
	LUT2 #(
		.INIT('h4)
	) name27457 (
		_w33280_,
		_w33283_,
		_w33284_
	);
	LUT3 #(
		.INIT('h48)
	) name27458 (
		_w33011_,
		_w33010_,
		_w33015_,
		_w33285_
	);
	LUT3 #(
		.INIT('h96)
	) name27459 (
		_w33011_,
		_w33010_,
		_w33015_,
		_w33286_
	);
	LUT4 #(
		.INIT('h050d)
	) name27460 (
		_w33011_,
		_w33012_,
		_w33013_,
		_w33015_,
		_w33287_
	);
	LUT2 #(
		.INIT('h8)
	) name27461 (
		_w33286_,
		_w33287_,
		_w33288_
	);
	LUT3 #(
		.INIT('hd0)
	) name27462 (
		_w33011_,
		_w33012_,
		_w33013_,
		_w33289_
	);
	LUT2 #(
		.INIT('h8)
	) name27463 (
		_w33285_,
		_w33289_,
		_w33290_
	);
	LUT4 #(
		.INIT('h0070)
	) name27464 (
		_w33014_,
		_w33035_,
		_w33009_,
		_w33025_,
		_w33291_
	);
	LUT3 #(
		.INIT('h10)
	) name27465 (
		_w33288_,
		_w33290_,
		_w33291_,
		_w33292_
	);
	LUT4 #(
		.INIT('hfe9f)
	) name27466 (
		_w33011_,
		_w33013_,
		_w33010_,
		_w33015_,
		_w33293_
	);
	LUT2 #(
		.INIT('h1)
	) name27467 (
		_w33012_,
		_w33293_,
		_w33294_
	);
	LUT3 #(
		.INIT('h15)
	) name27468 (
		_w33043_,
		_w33033_,
		_w33039_,
		_w33295_
	);
	LUT2 #(
		.INIT('h4)
	) name27469 (
		_w33294_,
		_w33295_,
		_w33296_
	);
	LUT4 #(
		.INIT('h56aa)
	) name27470 (
		\u0_L0_reg[23]/NET0131 ,
		_w33284_,
		_w33292_,
		_w33296_,
		_w33297_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name27471 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33298_
	);
	LUT4 #(
		.INIT('h4010)
	) name27472 (
		_w33142_,
		_w33144_,
		_w33141_,
		_w33143_,
		_w33299_
	);
	LUT2 #(
		.INIT('h4)
	) name27473 (
		_w33298_,
		_w33299_,
		_w33300_
	);
	LUT3 #(
		.INIT('h73)
	) name27474 (
		_w33142_,
		_w33144_,
		_w33143_,
		_w33301_
	);
	LUT2 #(
		.INIT('h1)
	) name27475 (
		_w33141_,
		_w33145_,
		_w33302_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name27476 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33303_
	);
	LUT3 #(
		.INIT('hb0)
	) name27477 (
		_w33301_,
		_w33302_,
		_w33303_,
		_w33304_
	);
	LUT3 #(
		.INIT('h45)
	) name27478 (
		_w33154_,
		_w33300_,
		_w33304_,
		_w33305_
	);
	LUT4 #(
		.INIT('hdf4f)
	) name27479 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33306_
	);
	LUT4 #(
		.INIT('hbcff)
	) name27480 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33307_
	);
	LUT4 #(
		.INIT('h04cc)
	) name27481 (
		_w33141_,
		_w33154_,
		_w33306_,
		_w33307_,
		_w33308_
	);
	LUT4 #(
		.INIT('h7dff)
	) name27482 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33309_
	);
	LUT4 #(
		.INIT('h6dff)
	) name27483 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33310_
	);
	LUT2 #(
		.INIT('h2)
	) name27484 (
		_w33141_,
		_w33310_,
		_w33311_
	);
	LUT4 #(
		.INIT('hbeff)
	) name27485 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33312_
	);
	LUT4 #(
		.INIT('hf5f1)
	) name27486 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33313_
	);
	LUT4 #(
		.INIT('hfa72)
	) name27487 (
		_w33141_,
		_w33154_,
		_w33312_,
		_w33313_,
		_w33314_
	);
	LUT3 #(
		.INIT('h10)
	) name27488 (
		_w33311_,
		_w33308_,
		_w33314_,
		_w33315_
	);
	LUT3 #(
		.INIT('h65)
	) name27489 (
		\u0_L0_reg[1]/NET0131 ,
		_w33305_,
		_w33315_,
		_w33316_
	);
	LUT4 #(
		.INIT('h008d)
	) name27490 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33317_
	);
	LUT2 #(
		.INIT('h2)
	) name27491 (
		_w33190_,
		_w33317_,
		_w33318_
	);
	LUT4 #(
		.INIT('hcd00)
	) name27492 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33319_
	);
	LUT4 #(
		.INIT('h5545)
	) name27493 (
		_w33190_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33320_
	);
	LUT3 #(
		.INIT('h04)
	) name27494 (
		_w33201_,
		_w33320_,
		_w33319_,
		_w33321_
	);
	LUT3 #(
		.INIT('h21)
	) name27495 (
		_w33193_,
		_w33191_,
		_w33194_,
		_w33322_
	);
	LUT4 #(
		.INIT('h6010)
	) name27496 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33323_
	);
	LUT2 #(
		.INIT('h1)
	) name27497 (
		_w33199_,
		_w33323_,
		_w33324_
	);
	LUT3 #(
		.INIT('he0)
	) name27498 (
		_w33318_,
		_w33321_,
		_w33324_,
		_w33325_
	);
	LUT3 #(
		.INIT('hb0)
	) name27499 (
		_w33193_,
		_w33191_,
		_w33194_,
		_w33326_
	);
	LUT3 #(
		.INIT('h90)
	) name27500 (
		_w33193_,
		_w33191_,
		_w33194_,
		_w33327_
	);
	LUT4 #(
		.INIT('h0040)
	) name27501 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33328_
	);
	LUT3 #(
		.INIT('h02)
	) name27502 (
		_w33190_,
		_w33328_,
		_w33327_,
		_w33329_
	);
	LUT4 #(
		.INIT('h4000)
	) name27503 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33330_
	);
	LUT3 #(
		.INIT('h04)
	) name27504 (
		_w33317_,
		_w33320_,
		_w33330_,
		_w33331_
	);
	LUT3 #(
		.INIT('h51)
	) name27505 (
		_w33190_,
		_w33193_,
		_w33191_,
		_w33332_
	);
	LUT4 #(
		.INIT('h0020)
	) name27506 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33333_
	);
	LUT4 #(
		.INIT('h00c4)
	) name27507 (
		_w33207_,
		_w33199_,
		_w33332_,
		_w33333_,
		_w33334_
	);
	LUT3 #(
		.INIT('he0)
	) name27508 (
		_w33329_,
		_w33331_,
		_w33334_,
		_w33335_
	);
	LUT3 #(
		.INIT('ha9)
	) name27509 (
		\u0_L0_reg[28]/NET0131 ,
		_w33325_,
		_w33335_,
		_w33336_
	);
	LUT4 #(
		.INIT('h3c3b)
	) name27510 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33337_
	);
	LUT4 #(
		.INIT('h0010)
	) name27511 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33338_
	);
	LUT4 #(
		.INIT('h0301)
	) name27512 (
		_w33223_,
		_w33222_,
		_w33338_,
		_w33337_,
		_w33339_
	);
	LUT4 #(
		.INIT('hdfdd)
	) name27513 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33223_,
		_w33340_
	);
	LUT2 #(
		.INIT('h2)
	) name27514 (
		_w33226_,
		_w33340_,
		_w33341_
	);
	LUT4 #(
		.INIT('h0008)
	) name27515 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33342_
	);
	LUT4 #(
		.INIT('h0010)
	) name27516 (
		_w33227_,
		_w33225_,
		_w33223_,
		_w33226_,
		_w33343_
	);
	LUT4 #(
		.INIT('hbf00)
	) name27517 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33222_,
		_w33344_
	);
	LUT3 #(
		.INIT('h10)
	) name27518 (
		_w33343_,
		_w33342_,
		_w33344_,
		_w33345_
	);
	LUT3 #(
		.INIT('h45)
	) name27519 (
		_w33339_,
		_w33341_,
		_w33345_,
		_w33346_
	);
	LUT4 #(
		.INIT('h2030)
	) name27520 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33222_,
		_w33347_
	);
	LUT4 #(
		.INIT('h0400)
	) name27521 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33348_
	);
	LUT4 #(
		.INIT('h0001)
	) name27522 (
		_w33223_,
		_w33237_,
		_w33348_,
		_w33347_,
		_w33349_
	);
	LUT3 #(
		.INIT('h02)
	) name27523 (
		_w33223_,
		_w33235_,
		_w33248_,
		_w33350_
	);
	LUT2 #(
		.INIT('h1)
	) name27524 (
		_w33349_,
		_w33350_,
		_w33351_
	);
	LUT3 #(
		.INIT('h56)
	) name27525 (
		\u0_L0_reg[15]/P0001 ,
		_w33346_,
		_w33351_,
		_w33352_
	);
	LUT4 #(
		.INIT('hc963)
	) name27526 (
		decrypt_pad,
		\u0_R0_reg[12]/NET0131 ,
		\u0_uk_K_r0_reg[24]/P0001 ,
		\u0_uk_K_r0_reg[3]/NET0131 ,
		_w33353_
	);
	LUT4 #(
		.INIT('hc693)
	) name27527 (
		decrypt_pad,
		\u0_R0_reg[9]/NET0131 ,
		\u0_uk_K_r0_reg[11]/NET0131 ,
		\u0_uk_K_r0_reg[32]/NET0131 ,
		_w33354_
	);
	LUT4 #(
		.INIT('hc693)
	) name27528 (
		decrypt_pad,
		\u0_R0_reg[8]/NET0131 ,
		\u0_uk_K_r0_reg[39]/NET0131 ,
		\u0_uk_K_r0_reg[3]/NET0131 ,
		_w33355_
	);
	LUT4 #(
		.INIT('hc693)
	) name27529 (
		decrypt_pad,
		\u0_R0_reg[10]/NET0131 ,
		\u0_uk_K_r0_reg[19]/NET0131 ,
		\u0_uk_K_r0_reg[40]/NET0131 ,
		_w33356_
	);
	LUT4 #(
		.INIT('hc963)
	) name27530 (
		decrypt_pad,
		\u0_R0_reg[13]/NET0131 ,
		\u0_uk_K_r0_reg[12]/NET0131 ,
		\u0_uk_K_r0_reg[48]/NET0131 ,
		_w33357_
	);
	LUT4 #(
		.INIT('h0010)
	) name27531 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33358_
	);
	LUT2 #(
		.INIT('h4)
	) name27532 (
		_w33355_,
		_w33357_,
		_w33359_
	);
	LUT3 #(
		.INIT('h10)
	) name27533 (
		_w33356_,
		_w33355_,
		_w33357_,
		_w33360_
	);
	LUT4 #(
		.INIT('hc693)
	) name27534 (
		decrypt_pad,
		\u0_R0_reg[11]/NET0131 ,
		\u0_uk_K_r0_reg[20]/NET0131 ,
		\u0_uk_K_r0_reg[41]/NET0131 ,
		_w33361_
	);
	LUT2 #(
		.INIT('h1)
	) name27535 (
		_w33354_,
		_w33361_,
		_w33362_
	);
	LUT3 #(
		.INIT('h15)
	) name27536 (
		_w33358_,
		_w33360_,
		_w33362_,
		_w33363_
	);
	LUT2 #(
		.INIT('h1)
	) name27537 (
		_w33355_,
		_w33357_,
		_w33364_
	);
	LUT2 #(
		.INIT('h8)
	) name27538 (
		_w33355_,
		_w33357_,
		_w33365_
	);
	LUT4 #(
		.INIT('he00e)
	) name27539 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33366_
	);
	LUT4 #(
		.INIT('h6006)
	) name27540 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33367_
	);
	LUT4 #(
		.INIT('h0800)
	) name27541 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33368_
	);
	LUT4 #(
		.INIT('h0080)
	) name27542 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33369_
	);
	LUT4 #(
		.INIT('h0200)
	) name27543 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33361_,
		_w33370_
	);
	LUT4 #(
		.INIT('h000b)
	) name27544 (
		_w33361_,
		_w33368_,
		_w33369_,
		_w33370_,
		_w33371_
	);
	LUT4 #(
		.INIT('h4555)
	) name27545 (
		_w33353_,
		_w33367_,
		_w33363_,
		_w33371_,
		_w33372_
	);
	LUT4 #(
		.INIT('ha25f)
	) name27546 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33373_
	);
	LUT2 #(
		.INIT('h8)
	) name27547 (
		_w33353_,
		_w33361_,
		_w33374_
	);
	LUT2 #(
		.INIT('h4)
	) name27548 (
		_w33373_,
		_w33374_,
		_w33375_
	);
	LUT3 #(
		.INIT('h0d)
	) name27549 (
		_w33354_,
		_w33357_,
		_w33361_,
		_w33376_
	);
	LUT3 #(
		.INIT('h0d)
	) name27550 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33377_
	);
	LUT3 #(
		.INIT('h8a)
	) name27551 (
		_w33353_,
		_w33354_,
		_w33357_,
		_w33378_
	);
	LUT3 #(
		.INIT('h40)
	) name27552 (
		_w33377_,
		_w33376_,
		_w33378_,
		_w33379_
	);
	LUT4 #(
		.INIT('h0001)
	) name27553 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33380_
	);
	LUT4 #(
		.INIT('hbbfe)
	) name27554 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33381_
	);
	LUT3 #(
		.INIT('h80)
	) name27555 (
		_w33353_,
		_w33354_,
		_w33356_,
		_w33382_
	);
	LUT4 #(
		.INIT('h51f3)
	) name27556 (
		_w33364_,
		_w33361_,
		_w33381_,
		_w33382_,
		_w33383_
	);
	LUT3 #(
		.INIT('h10)
	) name27557 (
		_w33379_,
		_w33375_,
		_w33383_,
		_w33384_
	);
	LUT3 #(
		.INIT('h65)
	) name27558 (
		\u0_L0_reg[6]/NET0131 ,
		_w33372_,
		_w33384_,
		_w33385_
	);
	LUT4 #(
		.INIT('hc963)
	) name27559 (
		decrypt_pad,
		\u0_R0_reg[20]/NET0131 ,
		\u0_uk_K_r0_reg[30]/NET0131 ,
		\u0_uk_K_r0_reg[9]/NET0131 ,
		_w33386_
	);
	LUT4 #(
		.INIT('hc963)
	) name27560 (
		decrypt_pad,
		\u0_R0_reg[18]/NET0131 ,
		\u0_uk_K_r0_reg[28]/NET0131 ,
		\u0_uk_K_r0_reg[7]/NET0131 ,
		_w33387_
	);
	LUT4 #(
		.INIT('hc963)
	) name27561 (
		decrypt_pad,
		\u0_R0_reg[21]/NET0131 ,
		\u0_uk_K_r0_reg[0]/NET0131 ,
		\u0_uk_K_r0_reg[38]/NET0131 ,
		_w33388_
	);
	LUT4 #(
		.INIT('hc963)
	) name27562 (
		decrypt_pad,
		\u0_R0_reg[19]/NET0131 ,
		\u0_uk_K_r0_reg[15]/NET0131 ,
		\u0_uk_K_r0_reg[49]/NET0131 ,
		_w33389_
	);
	LUT4 #(
		.INIT('hc963)
	) name27563 (
		decrypt_pad,
		\u0_R0_reg[17]/NET0131 ,
		\u0_uk_K_r0_reg[38]/NET0131 ,
		\u0_uk_K_r0_reg[44]/NET0131 ,
		_w33390_
	);
	LUT4 #(
		.INIT('hc693)
	) name27564 (
		decrypt_pad,
		\u0_R0_reg[16]/NET0131 ,
		\u0_uk_K_r0_reg[22]/NET0131 ,
		\u0_uk_K_r0_reg[43]/NET0131 ,
		_w33391_
	);
	LUT4 #(
		.INIT('h0020)
	) name27565 (
		_w33390_,
		_w33391_,
		_w33388_,
		_w33389_,
		_w33392_
	);
	LUT4 #(
		.INIT('hb796)
	) name27566 (
		_w33390_,
		_w33391_,
		_w33388_,
		_w33389_,
		_w33393_
	);
	LUT2 #(
		.INIT('h1)
	) name27567 (
		_w33387_,
		_w33393_,
		_w33394_
	);
	LUT3 #(
		.INIT('h80)
	) name27568 (
		_w33390_,
		_w33391_,
		_w33388_,
		_w33395_
	);
	LUT4 #(
		.INIT('hfb7b)
	) name27569 (
		_w33390_,
		_w33391_,
		_w33388_,
		_w33389_,
		_w33396_
	);
	LUT4 #(
		.INIT('ha43f)
	) name27570 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33397_
	);
	LUT4 #(
		.INIT('hf531)
	) name27571 (
		_w33387_,
		_w33389_,
		_w33396_,
		_w33397_,
		_w33398_
	);
	LUT3 #(
		.INIT('h8a)
	) name27572 (
		_w33386_,
		_w33394_,
		_w33398_,
		_w33399_
	);
	LUT4 #(
		.INIT('h0010)
	) name27573 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33400_
	);
	LUT4 #(
		.INIT('h4000)
	) name27574 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33401_
	);
	LUT4 #(
		.INIT('hbc67)
	) name27575 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33402_
	);
	LUT4 #(
		.INIT('h5bf8)
	) name27576 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33403_
	);
	LUT4 #(
		.INIT('h2000)
	) name27577 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33404_
	);
	LUT4 #(
		.INIT('hdffb)
	) name27578 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33405_
	);
	LUT4 #(
		.INIT('he400)
	) name27579 (
		_w33389_,
		_w33402_,
		_w33403_,
		_w33405_,
		_w33406_
	);
	LUT4 #(
		.INIT('h0208)
	) name27580 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33407_
	);
	LUT4 #(
		.INIT('h0040)
	) name27581 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33408_
	);
	LUT4 #(
		.INIT('hffbd)
	) name27582 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33409_
	);
	LUT3 #(
		.INIT('hb1)
	) name27583 (
		_w33389_,
		_w33407_,
		_w33409_,
		_w33410_
	);
	LUT3 #(
		.INIT('he0)
	) name27584 (
		_w33386_,
		_w33406_,
		_w33410_,
		_w33411_
	);
	LUT3 #(
		.INIT('h65)
	) name27585 (
		\u0_L0_reg[14]/NET0131 ,
		_w33399_,
		_w33411_,
		_w33412_
	);
	LUT3 #(
		.INIT('h13)
	) name27586 (
		_w33049_,
		_w33053_,
		_w33051_,
		_w33413_
	);
	LUT4 #(
		.INIT('hc4e6)
	) name27587 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33414_
	);
	LUT4 #(
		.INIT('h0201)
	) name27588 (
		_w33049_,
		_w33050_,
		_w33053_,
		_w33051_,
		_w33415_
	);
	LUT4 #(
		.INIT('h1011)
	) name27589 (
		_w33047_,
		_w33415_,
		_w33413_,
		_w33414_,
		_w33416_
	);
	LUT4 #(
		.INIT('h2010)
	) name27590 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33051_,
		_w33417_
	);
	LUT3 #(
		.INIT('h02)
	) name27591 (
		_w33047_,
		_w33078_,
		_w33073_,
		_w33418_
	);
	LUT4 #(
		.INIT('h0800)
	) name27592 (
		_w33049_,
		_w33050_,
		_w33048_,
		_w33053_,
		_w33419_
	);
	LUT4 #(
		.INIT('h1404)
	) name27593 (
		_w33049_,
		_w33050_,
		_w33053_,
		_w33051_,
		_w33420_
	);
	LUT2 #(
		.INIT('h1)
	) name27594 (
		_w33419_,
		_w33420_,
		_w33421_
	);
	LUT4 #(
		.INIT('h4555)
	) name27595 (
		_w33416_,
		_w33417_,
		_w33418_,
		_w33421_,
		_w33422_
	);
	LUT2 #(
		.INIT('h2)
	) name27596 (
		_w33080_,
		_w33060_,
		_w33423_
	);
	LUT3 #(
		.INIT('h65)
	) name27597 (
		\u0_L0_reg[19]/P0001 ,
		_w33422_,
		_w33423_,
		_w33424_
	);
	LUT4 #(
		.INIT('h3ce4)
	) name27598 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33425_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name27599 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33426_
	);
	LUT4 #(
		.INIT('hbb7f)
	) name27600 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33427_
	);
	LUT4 #(
		.INIT('he400)
	) name27601 (
		_w33389_,
		_w33426_,
		_w33425_,
		_w33427_,
		_w33428_
	);
	LUT2 #(
		.INIT('h2)
	) name27602 (
		_w33386_,
		_w33428_,
		_w33429_
	);
	LUT4 #(
		.INIT('hf5ee)
	) name27603 (
		_w33390_,
		_w33391_,
		_w33388_,
		_w33389_,
		_w33430_
	);
	LUT2 #(
		.INIT('h1)
	) name27604 (
		_w33387_,
		_w33430_,
		_w33431_
	);
	LUT4 #(
		.INIT('h0004)
	) name27605 (
		_w33390_,
		_w33391_,
		_w33388_,
		_w33389_,
		_w33432_
	);
	LUT2 #(
		.INIT('h4)
	) name27606 (
		_w33388_,
		_w33389_,
		_w33433_
	);
	LUT3 #(
		.INIT('h08)
	) name27607 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33434_
	);
	LUT3 #(
		.INIT('h45)
	) name27608 (
		_w33432_,
		_w33433_,
		_w33434_,
		_w33435_
	);
	LUT4 #(
		.INIT('hff7d)
	) name27609 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33436_
	);
	LUT4 #(
		.INIT('hfe7d)
	) name27610 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33437_
	);
	LUT4 #(
		.INIT('h0020)
	) name27611 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33389_,
		_w33438_
	);
	LUT4 #(
		.INIT('h0031)
	) name27612 (
		_w33389_,
		_w33401_,
		_w33437_,
		_w33438_,
		_w33439_
	);
	LUT4 #(
		.INIT('hba00)
	) name27613 (
		_w33386_,
		_w33431_,
		_w33435_,
		_w33439_,
		_w33440_
	);
	LUT3 #(
		.INIT('h65)
	) name27614 (
		\u0_L0_reg[25]/NET0131 ,
		_w33429_,
		_w33440_,
		_w33441_
	);
	LUT3 #(
		.INIT('hd0)
	) name27615 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33442_
	);
	LUT4 #(
		.INIT('h0094)
	) name27616 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33443_
	);
	LUT2 #(
		.INIT('h1)
	) name27617 (
		_w33142_,
		_w33145_,
		_w33444_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name27618 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33445_
	);
	LUT4 #(
		.INIT('h0054)
	) name27619 (
		_w33141_,
		_w33154_,
		_w33445_,
		_w33443_,
		_w33446_
	);
	LUT3 #(
		.INIT('h02)
	) name27620 (
		_w33141_,
		_w33149_,
		_w33157_,
		_w33447_
	);
	LUT2 #(
		.INIT('h1)
	) name27621 (
		_w33446_,
		_w33447_,
		_w33448_
	);
	LUT4 #(
		.INIT('h4010)
	) name27622 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33449_
	);
	LUT3 #(
		.INIT('h02)
	) name27623 (
		_w33154_,
		_w33163_,
		_w33449_,
		_w33450_
	);
	LUT4 #(
		.INIT('h77fd)
	) name27624 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w33451_
	);
	LUT4 #(
		.INIT('hdddf)
	) name27625 (
		_w33142_,
		_w33144_,
		_w33141_,
		_w33145_,
		_w33452_
	);
	LUT4 #(
		.INIT('hfa32)
	) name27626 (
		_w33141_,
		_w33143_,
		_w33451_,
		_w33452_,
		_w33453_
	);
	LUT4 #(
		.INIT('h00fd)
	) name27627 (
		_w33144_,
		_w33145_,
		_w33143_,
		_w33154_,
		_w33454_
	);
	LUT3 #(
		.INIT('h70)
	) name27628 (
		_w33165_,
		_w33442_,
		_w33454_,
		_w33455_
	);
	LUT4 #(
		.INIT('h153f)
	) name27629 (
		_w33151_,
		_w33450_,
		_w33453_,
		_w33455_,
		_w33456_
	);
	LUT3 #(
		.INIT('h56)
	) name27630 (
		\u0_L0_reg[26]/NET0131 ,
		_w33448_,
		_w33456_,
		_w33457_
	);
	LUT4 #(
		.INIT('hb000)
	) name27631 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33458_
	);
	LUT4 #(
		.INIT('h0400)
	) name27632 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33459_
	);
	LUT4 #(
		.INIT('h0002)
	) name27633 (
		_w33190_,
		_w33322_,
		_w33459_,
		_w33458_,
		_w33460_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name27634 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33461_
	);
	LUT4 #(
		.INIT('h5545)
	) name27635 (
		_w33190_,
		_w33193_,
		_w33191_,
		_w33194_,
		_w33462_
	);
	LUT4 #(
		.INIT('h1000)
	) name27636 (
		_w33206_,
		_w33333_,
		_w33461_,
		_w33462_,
		_w33463_
	);
	LUT2 #(
		.INIT('h1)
	) name27637 (
		_w33190_,
		_w33191_,
		_w33464_
	);
	LUT3 #(
		.INIT('h02)
	) name27638 (
		_w33193_,
		_w33192_,
		_w33194_,
		_w33465_
	);
	LUT3 #(
		.INIT('h45)
	) name27639 (
		_w33199_,
		_w33464_,
		_w33465_,
		_w33466_
	);
	LUT3 #(
		.INIT('he0)
	) name27640 (
		_w33460_,
		_w33463_,
		_w33466_,
		_w33467_
	);
	LUT3 #(
		.INIT('h10)
	) name27641 (
		_w33197_,
		_w33198_,
		_w33199_,
		_w33468_
	);
	LUT4 #(
		.INIT('h0004)
	) name27642 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33469_
	);
	LUT3 #(
		.INIT('he4)
	) name27643 (
		_w33193_,
		_w33192_,
		_w33194_,
		_w33470_
	);
	LUT3 #(
		.INIT('h13)
	) name27644 (
		_w33464_,
		_w33469_,
		_w33470_,
		_w33471_
	);
	LUT4 #(
		.INIT('hfe5e)
	) name27645 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33472_
	);
	LUT3 #(
		.INIT('hc4)
	) name27646 (
		_w33190_,
		_w33461_,
		_w33472_,
		_w33473_
	);
	LUT3 #(
		.INIT('h80)
	) name27647 (
		_w33468_,
		_w33471_,
		_w33473_,
		_w33474_
	);
	LUT3 #(
		.INIT('h56)
	) name27648 (
		\u0_L0_reg[13]/NET0131 ,
		_w33467_,
		_w33474_,
		_w33475_
	);
	LUT4 #(
		.INIT('h0001)
	) name27649 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33476_
	);
	LUT4 #(
		.INIT('hcffe)
	) name27650 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33477_
	);
	LUT4 #(
		.INIT('haa8a)
	) name27651 (
		_w33386_,
		_w33387_,
		_w33391_,
		_w33389_,
		_w33478_
	);
	LUT4 #(
		.INIT('h3100)
	) name27652 (
		_w33389_,
		_w33407_,
		_w33477_,
		_w33478_,
		_w33479_
	);
	LUT3 #(
		.INIT('h02)
	) name27653 (
		_w33389_,
		_w33400_,
		_w33395_,
		_w33480_
	);
	LUT4 #(
		.INIT('h0d00)
	) name27654 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33481_
	);
	LUT4 #(
		.INIT('h00bf)
	) name27655 (
		_w33390_,
		_w33391_,
		_w33388_,
		_w33389_,
		_w33482_
	);
	LUT2 #(
		.INIT('h4)
	) name27656 (
		_w33481_,
		_w33482_,
		_w33483_
	);
	LUT4 #(
		.INIT('h5545)
	) name27657 (
		_w33386_,
		_w33387_,
		_w33390_,
		_w33391_,
		_w33484_
	);
	LUT2 #(
		.INIT('h8)
	) name27658 (
		_w33436_,
		_w33484_,
		_w33485_
	);
	LUT4 #(
		.INIT('h0155)
	) name27659 (
		_w33479_,
		_w33480_,
		_w33483_,
		_w33485_,
		_w33486_
	);
	LUT4 #(
		.INIT('hf977)
	) name27660 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33487_
	);
	LUT4 #(
		.INIT('haf23)
	) name27661 (
		_w33388_,
		_w33389_,
		_w33438_,
		_w33487_,
		_w33488_
	);
	LUT3 #(
		.INIT('h65)
	) name27662 (
		\u0_L0_reg[8]/NET0131 ,
		_w33486_,
		_w33488_,
		_w33489_
	);
	LUT3 #(
		.INIT('h80)
	) name27663 (
		_w33354_,
		_w33355_,
		_w33357_,
		_w33490_
	);
	LUT4 #(
		.INIT('h696b)
	) name27664 (
		_w33354_,
		_w33355_,
		_w33357_,
		_w33361_,
		_w33491_
	);
	LUT2 #(
		.INIT('h1)
	) name27665 (
		_w33356_,
		_w33491_,
		_w33492_
	);
	LUT4 #(
		.INIT('h0006)
	) name27666 (
		_w33356_,
		_w33355_,
		_w33357_,
		_w33361_,
		_w33493_
	);
	LUT3 #(
		.INIT('h02)
	) name27667 (
		_w33353_,
		_w33368_,
		_w33493_,
		_w33494_
	);
	LUT4 #(
		.INIT('h5afc)
	) name27668 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33495_
	);
	LUT2 #(
		.INIT('h1)
	) name27669 (
		_w33361_,
		_w33495_,
		_w33496_
	);
	LUT4 #(
		.INIT('h6800)
	) name27670 (
		_w33354_,
		_w33355_,
		_w33357_,
		_w33361_,
		_w33497_
	);
	LUT3 #(
		.INIT('h01)
	) name27671 (
		_w33353_,
		_w33380_,
		_w33497_,
		_w33498_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name27672 (
		_w33492_,
		_w33494_,
		_w33496_,
		_w33498_,
		_w33499_
	);
	LUT3 #(
		.INIT('h40)
	) name27673 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33500_
	);
	LUT4 #(
		.INIT('h00bf)
	) name27674 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33361_,
		_w33501_
	);
	LUT4 #(
		.INIT('h0004)
	) name27675 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33502_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name27676 (
		_w33361_,
		_w33369_,
		_w33501_,
		_w33502_,
		_w33503_
	);
	LUT3 #(
		.INIT('h56)
	) name27677 (
		\u0_L0_reg[16]/NET0131 ,
		_w33499_,
		_w33503_,
		_w33504_
	);
	LUT4 #(
		.INIT('hc1e6)
	) name27678 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33505_
	);
	LUT4 #(
		.INIT('h2880)
	) name27679 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33506_
	);
	LUT4 #(
		.INIT('h4140)
	) name27680 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33507_
	);
	LUT4 #(
		.INIT('h1032)
	) name27681 (
		_w33084_,
		_w33506_,
		_w33505_,
		_w33507_,
		_w33508_
	);
	LUT2 #(
		.INIT('h2)
	) name27682 (
		_w33083_,
		_w33508_,
		_w33509_
	);
	LUT2 #(
		.INIT('h2)
	) name27683 (
		_w33083_,
		_w33084_,
		_w33510_
	);
	LUT4 #(
		.INIT('h0002)
	) name27684 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33511_
	);
	LUT4 #(
		.INIT('h0f04)
	) name27685 (
		_w33084_,
		_w33507_,
		_w33510_,
		_w33511_,
		_w33512_
	);
	LUT2 #(
		.INIT('h4)
	) name27686 (
		_w33084_,
		_w33506_,
		_w33513_
	);
	LUT4 #(
		.INIT('h41c1)
	) name27687 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33514_
	);
	LUT4 #(
		.INIT('h2800)
	) name27688 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33515_
	);
	LUT2 #(
		.INIT('h4)
	) name27689 (
		_w33083_,
		_w33084_,
		_w33516_
	);
	LUT3 #(
		.INIT('h10)
	) name27690 (
		_w33515_,
		_w33514_,
		_w33516_,
		_w33517_
	);
	LUT3 #(
		.INIT('h01)
	) name27691 (
		_w33513_,
		_w33512_,
		_w33517_,
		_w33518_
	);
	LUT3 #(
		.INIT('h65)
	) name27692 (
		\u0_L0_reg[7]/NET0131 ,
		_w33509_,
		_w33518_,
		_w33519_
	);
	LUT4 #(
		.INIT('h2804)
	) name27693 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33520_
	);
	LUT3 #(
		.INIT('h20)
	) name27694 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33521_
	);
	LUT3 #(
		.INIT('h28)
	) name27695 (
		_w33013_,
		_w33010_,
		_w33015_,
		_w33522_
	);
	LUT3 #(
		.INIT('h43)
	) name27696 (
		_w33011_,
		_w33010_,
		_w33015_,
		_w33523_
	);
	LUT4 #(
		.INIT('h1003)
	) name27697 (
		_w33011_,
		_w33013_,
		_w33010_,
		_w33015_,
		_w33524_
	);
	LUT4 #(
		.INIT('h1011)
	) name27698 (
		_w33009_,
		_w33524_,
		_w33521_,
		_w33522_,
		_w33525_
	);
	LUT4 #(
		.INIT('h8448)
	) name27699 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33526_
	);
	LUT4 #(
		.INIT('h0020)
	) name27700 (
		_w33011_,
		_w33012_,
		_w33010_,
		_w33015_,
		_w33527_
	);
	LUT4 #(
		.INIT('h002a)
	) name27701 (
		_w33009_,
		_w33030_,
		_w33523_,
		_w33527_,
		_w33528_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name27702 (
		_w33520_,
		_w33525_,
		_w33526_,
		_w33528_,
		_w33529_
	);
	LUT3 #(
		.INIT('h40)
	) name27703 (
		_w33013_,
		_w33010_,
		_w33015_,
		_w33530_
	);
	LUT2 #(
		.INIT('h4)
	) name27704 (
		_w33019_,
		_w33530_,
		_w33531_
	);
	LUT3 #(
		.INIT('h56)
	) name27705 (
		\u0_L0_reg[9]/NET0131 ,
		_w33529_,
		_w33531_,
		_w33532_
	);
	LUT4 #(
		.INIT('hc043)
	) name27706 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33533_
	);
	LUT4 #(
		.INIT('h3c28)
	) name27707 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33534_
	);
	LUT3 #(
		.INIT('h01)
	) name27708 (
		_w33084_,
		_w33533_,
		_w33534_,
		_w33535_
	);
	LUT4 #(
		.INIT('h0800)
	) name27709 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33536_
	);
	LUT3 #(
		.INIT('he2)
	) name27710 (
		_w33085_,
		_w33087_,
		_w33088_,
		_w33537_
	);
	LUT4 #(
		.INIT('ha7f4)
	) name27711 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33538_
	);
	LUT3 #(
		.INIT('h31)
	) name27712 (
		_w33084_,
		_w33536_,
		_w33538_,
		_w33539_
	);
	LUT3 #(
		.INIT('h8a)
	) name27713 (
		_w33083_,
		_w33535_,
		_w33539_,
		_w33540_
	);
	LUT3 #(
		.INIT('h04)
	) name27714 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33541_
	);
	LUT2 #(
		.INIT('h2)
	) name27715 (
		_w33274_,
		_w33541_,
		_w33542_
	);
	LUT4 #(
		.INIT('h79df)
	) name27716 (
		_w33085_,
		_w33086_,
		_w33087_,
		_w33088_,
		_w33543_
	);
	LUT3 #(
		.INIT('hd0)
	) name27717 (
		_w33099_,
		_w33537_,
		_w33543_,
		_w33544_
	);
	LUT4 #(
		.INIT('h00e0)
	) name27718 (
		_w33085_,
		_w33087_,
		_w33088_,
		_w33084_,
		_w33545_
	);
	LUT4 #(
		.INIT('h195f)
	) name27719 (
		_w33085_,
		_w33086_,
		_w33271_,
		_w33545_,
		_w33546_
	);
	LUT4 #(
		.INIT('hba00)
	) name27720 (
		_w33083_,
		_w33542_,
		_w33544_,
		_w33546_,
		_w33547_
	);
	LUT3 #(
		.INIT('h65)
	) name27721 (
		\u0_L0_reg[32]/NET0131 ,
		_w33540_,
		_w33547_,
		_w33548_
	);
	LUT4 #(
		.INIT('hc004)
	) name27722 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33549_
	);
	LUT3 #(
		.INIT('h28)
	) name27723 (
		_w33227_,
		_w33225_,
		_w33226_,
		_w33550_
	);
	LUT4 #(
		.INIT('hf3e2)
	) name27724 (
		_w33233_,
		_w33223_,
		_w33549_,
		_w33550_,
		_w33551_
	);
	LUT3 #(
		.INIT('h10)
	) name27725 (
		_w33224_,
		_w33227_,
		_w33226_,
		_w33552_
	);
	LUT4 #(
		.INIT('h0004)
	) name27726 (
		_w33235_,
		_w33222_,
		_w33229_,
		_w33552_,
		_w33553_
	);
	LUT4 #(
		.INIT('hf700)
	) name27727 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33223_,
		_w33554_
	);
	LUT3 #(
		.INIT('h4b)
	) name27728 (
		_w33224_,
		_w33227_,
		_w33226_,
		_w33555_
	);
	LUT2 #(
		.INIT('h8)
	) name27729 (
		_w33554_,
		_w33555_,
		_w33556_
	);
	LUT4 #(
		.INIT('he2ff)
	) name27730 (
		_w33227_,
		_w33225_,
		_w33223_,
		_w33226_,
		_w33557_
	);
	LUT4 #(
		.INIT('h0301)
	) name27731 (
		_w33224_,
		_w33222_,
		_w33257_,
		_w33557_,
		_w33558_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name27732 (
		_w33551_,
		_w33553_,
		_w33556_,
		_w33558_,
		_w33559_
	);
	LUT4 #(
		.INIT('hefb7)
	) name27733 (
		_w33224_,
		_w33227_,
		_w33225_,
		_w33226_,
		_w33560_
	);
	LUT4 #(
		.INIT('h0020)
	) name27734 (
		_w33224_,
		_w33227_,
		_w33223_,
		_w33226_,
		_w33561_
	);
	LUT3 #(
		.INIT('h0e)
	) name27735 (
		_w33223_,
		_w33560_,
		_w33561_,
		_w33562_
	);
	LUT3 #(
		.INIT('h65)
	) name27736 (
		\u0_L0_reg[27]/NET0131 ,
		_w33559_,
		_w33562_,
		_w33563_
	);
	LUT4 #(
		.INIT('h3f9d)
	) name27737 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33564_
	);
	LUT2 #(
		.INIT('h2)
	) name27738 (
		_w33361_,
		_w33564_,
		_w33565_
	);
	LUT3 #(
		.INIT('h3a)
	) name27739 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33566_
	);
	LUT4 #(
		.INIT('hebfe)
	) name27740 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33567_
	);
	LUT4 #(
		.INIT('h1500)
	) name27741 (
		_w33353_,
		_w33376_,
		_w33566_,
		_w33567_,
		_w33568_
	);
	LUT4 #(
		.INIT('hfce3)
	) name27742 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33569_
	);
	LUT4 #(
		.INIT('h3f35)
	) name27743 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33570_
	);
	LUT4 #(
		.INIT('ha820)
	) name27744 (
		_w33353_,
		_w33361_,
		_w33570_,
		_w33569_,
		_w33571_
	);
	LUT3 #(
		.INIT('h0b)
	) name27745 (
		_w33565_,
		_w33568_,
		_w33571_,
		_w33572_
	);
	LUT2 #(
		.INIT('h8)
	) name27746 (
		_w33357_,
		_w33361_,
		_w33573_
	);
	LUT2 #(
		.INIT('h8)
	) name27747 (
		_w33500_,
		_w33573_,
		_w33574_
	);
	LUT2 #(
		.INIT('h2)
	) name27748 (
		_w33356_,
		_w33361_,
		_w33575_
	);
	LUT4 #(
		.INIT('h0008)
	) name27749 (
		_w33354_,
		_w33356_,
		_w33357_,
		_w33361_,
		_w33576_
	);
	LUT3 #(
		.INIT('h0b)
	) name27750 (
		_w33365_,
		_w33382_,
		_w33576_,
		_w33577_
	);
	LUT2 #(
		.INIT('h4)
	) name27751 (
		_w33574_,
		_w33577_,
		_w33578_
	);
	LUT3 #(
		.INIT('h9a)
	) name27752 (
		\u0_L0_reg[30]/P0001 ,
		_w33572_,
		_w33578_,
		_w33579_
	);
	LUT4 #(
		.INIT('h2028)
	) name27753 (
		_w33190_,
		_w33193_,
		_w33191_,
		_w33194_,
		_w33580_
	);
	LUT3 #(
		.INIT('h15)
	) name27754 (
		_w33190_,
		_w33193_,
		_w33192_,
		_w33581_
	);
	LUT4 #(
		.INIT('h0105)
	) name27755 (
		_w33212_,
		_w33326_,
		_w33580_,
		_w33581_,
		_w33582_
	);
	LUT2 #(
		.INIT('h2)
	) name27756 (
		_w33199_,
		_w33582_,
		_w33583_
	);
	LUT3 #(
		.INIT('h07)
	) name27757 (
		_w33190_,
		_w33191_,
		_w33194_,
		_w33584_
	);
	LUT2 #(
		.INIT('h9)
	) name27758 (
		_w33191_,
		_w33192_,
		_w33585_
	);
	LUT3 #(
		.INIT('he0)
	) name27759 (
		_w33205_,
		_w33584_,
		_w33585_,
		_w33586_
	);
	LUT4 #(
		.INIT('h8000)
	) name27760 (
		_w33190_,
		_w33193_,
		_w33191_,
		_w33194_,
		_w33587_
	);
	LUT3 #(
		.INIT('h01)
	) name27761 (
		_w33195_,
		_w33330_,
		_w33587_,
		_w33588_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name27762 (
		_w33193_,
		_w33191_,
		_w33192_,
		_w33194_,
		_w33589_
	);
	LUT4 #(
		.INIT('h0040)
	) name27763 (
		_w33190_,
		_w33193_,
		_w33191_,
		_w33194_,
		_w33590_
	);
	LUT3 #(
		.INIT('h0d)
	) name27764 (
		_w33190_,
		_w33589_,
		_w33590_,
		_w33591_
	);
	LUT4 #(
		.INIT('hba00)
	) name27765 (
		_w33199_,
		_w33586_,
		_w33588_,
		_w33591_,
		_w33592_
	);
	LUT3 #(
		.INIT('h65)
	) name27766 (
		\u0_L0_reg[18]/NET0131 ,
		_w33583_,
		_w33592_,
		_w33593_
	);
	LUT4 #(
		.INIT('h0040)
	) name27767 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33594_
	);
	LUT4 #(
		.INIT('hbcb1)
	) name27768 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33595_
	);
	LUT4 #(
		.INIT('h5054)
	) name27769 (
		_w33353_,
		_w33361_,
		_w33594_,
		_w33595_,
		_w33596_
	);
	LUT3 #(
		.INIT('h10)
	) name27770 (
		_w33354_,
		_w33356_,
		_w33361_,
		_w33597_
	);
	LUT2 #(
		.INIT('h4)
	) name27771 (
		_w33359_,
		_w33597_,
		_w33598_
	);
	LUT4 #(
		.INIT('h737f)
	) name27772 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33599_
	);
	LUT3 #(
		.INIT('hd1)
	) name27773 (
		_w33366_,
		_w33361_,
		_w33599_,
		_w33600_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name27774 (
		_w33353_,
		_w33363_,
		_w33598_,
		_w33600_,
		_w33601_
	);
	LUT4 #(
		.INIT('he35e)
	) name27775 (
		_w33354_,
		_w33356_,
		_w33355_,
		_w33357_,
		_w33602_
	);
	LUT2 #(
		.INIT('h1)
	) name27776 (
		_w33353_,
		_w33361_,
		_w33603_
	);
	LUT2 #(
		.INIT('h4)
	) name27777 (
		_w33602_,
		_w33603_,
		_w33604_
	);
	LUT2 #(
		.INIT('h8)
	) name27778 (
		_w33361_,
		_w33358_,
		_w33605_
	);
	LUT4 #(
		.INIT('h0777)
	) name27779 (
		_w33357_,
		_w33370_,
		_w33490_,
		_w33575_,
		_w33606_
	);
	LUT3 #(
		.INIT('h10)
	) name27780 (
		_w33604_,
		_w33605_,
		_w33606_,
		_w33607_
	);
	LUT4 #(
		.INIT('h5655)
	) name27781 (
		\u0_L0_reg[24]/NET0131 ,
		_w33601_,
		_w33596_,
		_w33607_,
		_w33608_
	);
	LUT4 #(
		.INIT('haff3)
	) name27782 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33609_
	);
	LUT2 #(
		.INIT('h2)
	) name27783 (
		_w33389_,
		_w33609_,
		_w33610_
	);
	LUT4 #(
		.INIT('h0020)
	) name27784 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33611_
	);
	LUT3 #(
		.INIT('h01)
	) name27785 (
		_w33401_,
		_w33392_,
		_w33611_,
		_w33612_
	);
	LUT3 #(
		.INIT('h8a)
	) name27786 (
		_w33386_,
		_w33610_,
		_w33612_,
		_w33613_
	);
	LUT4 #(
		.INIT('hd83d)
	) name27787 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33614_
	);
	LUT2 #(
		.INIT('h1)
	) name27788 (
		_w33386_,
		_w33614_,
		_w33615_
	);
	LUT4 #(
		.INIT('h0200)
	) name27789 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33616_
	);
	LUT3 #(
		.INIT('h02)
	) name27790 (
		_w33389_,
		_w33400_,
		_w33616_,
		_w33617_
	);
	LUT4 #(
		.INIT('h45f0)
	) name27791 (
		_w33387_,
		_w33390_,
		_w33391_,
		_w33388_,
		_w33618_
	);
	LUT3 #(
		.INIT('h0d)
	) name27792 (
		_w33386_,
		_w33404_,
		_w33618_,
		_w33619_
	);
	LUT3 #(
		.INIT('h01)
	) name27793 (
		_w33389_,
		_w33408_,
		_w33476_,
		_w33620_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name27794 (
		_w33615_,
		_w33617_,
		_w33619_,
		_w33620_,
		_w33621_
	);
	LUT3 #(
		.INIT('h56)
	) name27795 (
		\u0_L0_reg[3]/NET0131 ,
		_w33613_,
		_w33621_,
		_w33622_
	);
	LUT4 #(
		.INIT('hc693)
	) name27796 (
		decrypt_pad,
		\u0_desIn_r_reg[25]/NET0131 ,
		\u0_key_r_reg[35]/P0001 ,
		\u0_key_r_reg[42]/P0001 ,
		_w33623_
	);
	LUT4 #(
		.INIT('hc693)
	) name27797 (
		decrypt_pad,
		\u0_desIn_r_reg[9]/NET0131 ,
		\u0_key_r_reg[15]/NET0131 ,
		\u0_key_r_reg[22]/NET0131 ,
		_w33624_
	);
	LUT4 #(
		.INIT('hc963)
	) name27798 (
		decrypt_pad,
		\u0_desIn_r_reg[59]/NET0131 ,
		\u0_key_r_reg[2]/NET0131 ,
		\u0_key_r_reg[50]/NET0131 ,
		_w33625_
	);
	LUT4 #(
		.INIT('hc693)
	) name27799 (
		decrypt_pad,
		\u0_desIn_r_reg[33]/NET0131 ,
		\u0_key_r_reg[31]/NET0131 ,
		\u0_key_r_reg[38]/NET0131 ,
		_w33626_
	);
	LUT4 #(
		.INIT('hc693)
	) name27800 (
		decrypt_pad,
		\u0_desIn_r_reg[1]/NET0131 ,
		\u0_key_r_reg[30]/NET0131 ,
		\u0_key_r_reg[37]/NET0131 ,
		_w33627_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name27801 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33628_
	);
	LUT4 #(
		.INIT('hc963)
	) name27802 (
		decrypt_pad,
		\u0_desIn_r_reg[17]/NET0131 ,
		\u0_key_r_reg[0]/NET0131 ,
		\u0_key_r_reg[52]/NET0131 ,
		_w33629_
	);
	LUT4 #(
		.INIT('h0408)
	) name27803 (
		_w33625_,
		_w33626_,
		_w33629_,
		_w33627_,
		_w33630_
	);
	LUT2 #(
		.INIT('h4)
	) name27804 (
		_w33628_,
		_w33630_,
		_w33631_
	);
	LUT4 #(
		.INIT('h0800)
	) name27805 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33632_
	);
	LUT4 #(
		.INIT('hf75f)
	) name27806 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33633_
	);
	LUT4 #(
		.INIT('h0040)
	) name27807 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33634_
	);
	LUT4 #(
		.INIT('hffbe)
	) name27808 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33635_
	);
	LUT3 #(
		.INIT('hd0)
	) name27809 (
		_w33629_,
		_w33633_,
		_w33635_,
		_w33636_
	);
	LUT3 #(
		.INIT('h8a)
	) name27810 (
		_w33623_,
		_w33631_,
		_w33636_,
		_w33637_
	);
	LUT4 #(
		.INIT('h0010)
	) name27811 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33638_
	);
	LUT4 #(
		.INIT('h5d6f)
	) name27812 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33639_
	);
	LUT2 #(
		.INIT('h1)
	) name27813 (
		_w33629_,
		_w33639_,
		_w33640_
	);
	LUT2 #(
		.INIT('h2)
	) name27814 (
		_w33626_,
		_w33629_,
		_w33641_
	);
	LUT3 #(
		.INIT('h02)
	) name27815 (
		_w33625_,
		_w33624_,
		_w33627_,
		_w33642_
	);
	LUT2 #(
		.INIT('h1)
	) name27816 (
		_w33629_,
		_w33624_,
		_w33643_
	);
	LUT4 #(
		.INIT('h0004)
	) name27817 (
		_w33625_,
		_w33626_,
		_w33629_,
		_w33624_,
		_w33644_
	);
	LUT4 #(
		.INIT('h8400)
	) name27818 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33645_
	);
	LUT4 #(
		.INIT('h1011)
	) name27819 (
		_w33644_,
		_w33645_,
		_w33641_,
		_w33642_,
		_w33646_
	);
	LUT4 #(
		.INIT('hef9c)
	) name27820 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33647_
	);
	LUT4 #(
		.INIT('h2100)
	) name27821 (
		_w33625_,
		_w33629_,
		_w33624_,
		_w33627_,
		_w33648_
	);
	LUT3 #(
		.INIT('h0d)
	) name27822 (
		_w33629_,
		_w33647_,
		_w33648_,
		_w33649_
	);
	LUT4 #(
		.INIT('hba00)
	) name27823 (
		_w33623_,
		_w33640_,
		_w33646_,
		_w33649_,
		_w33650_
	);
	LUT3 #(
		.INIT('h65)
	) name27824 (
		\u0_desIn_r_reg[42]/NET0131 ,
		_w33637_,
		_w33650_,
		_w33651_
	);
	LUT4 #(
		.INIT('hc693)
	) name27825 (
		decrypt_pad,
		\u0_desIn_r_reg[57]/NET0131 ,
		\u0_key_r_reg[40]/NET0131 ,
		\u0_key_r_reg[47]/NET0131 ,
		_w33652_
	);
	LUT4 #(
		.INIT('hc963)
	) name27826 (
		decrypt_pad,
		\u0_desIn_r_reg[23]/NET0131 ,
		\u0_key_r_reg[3]/NET0131 ,
		\u0_key_r_reg[53]/NET0131 ,
		_w33653_
	);
	LUT4 #(
		.INIT('hc963)
	) name27827 (
		decrypt_pad,
		\u0_desIn_r_reg[7]/NET0131 ,
		\u0_key_r_reg[11]/NET0131 ,
		\u0_key_r_reg[4]/NET0131 ,
		_w33654_
	);
	LUT4 #(
		.INIT('hc693)
	) name27828 (
		decrypt_pad,
		\u0_desIn_r_reg[39]/NET0131 ,
		\u0_key_r_reg[34]/NET0131 ,
		\u0_key_r_reg[41]/NET0131 ,
		_w33655_
	);
	LUT4 #(
		.INIT('hc693)
	) name27829 (
		decrypt_pad,
		\u0_desIn_r_reg[15]/NET0131 ,
		\u0_key_r_reg[19]/NET0131 ,
		\u0_key_r_reg[26]/NET0131 ,
		_w33656_
	);
	LUT4 #(
		.INIT('hafac)
	) name27830 (
		_w33653_,
		_w33656_,
		_w33654_,
		_w33655_,
		_w33657_
	);
	LUT2 #(
		.INIT('h2)
	) name27831 (
		_w33652_,
		_w33657_,
		_w33658_
	);
	LUT4 #(
		.INIT('hccf5)
	) name27832 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w33659_
	);
	LUT2 #(
		.INIT('h2)
	) name27833 (
		_w33653_,
		_w33659_,
		_w33660_
	);
	LUT4 #(
		.INIT('hc963)
	) name27834 (
		decrypt_pad,
		\u0_desIn_r_reg[31]/NET0131 ,
		\u0_key_r_reg[13]/NET0131 ,
		\u0_key_r_reg[6]/NET0131 ,
		_w33661_
	);
	LUT2 #(
		.INIT('h2)
	) name27835 (
		_w33653_,
		_w33656_,
		_w33662_
	);
	LUT3 #(
		.INIT('hd0)
	) name27836 (
		_w33653_,
		_w33656_,
		_w33654_,
		_w33663_
	);
	LUT3 #(
		.INIT('hcd)
	) name27837 (
		_w33656_,
		_w33652_,
		_w33655_,
		_w33664_
	);
	LUT3 #(
		.INIT('ha8)
	) name27838 (
		_w33661_,
		_w33663_,
		_w33664_,
		_w33665_
	);
	LUT3 #(
		.INIT('h10)
	) name27839 (
		_w33660_,
		_w33658_,
		_w33665_,
		_w33666_
	);
	LUT4 #(
		.INIT('h4ff3)
	) name27840 (
		_w33653_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w33667_
	);
	LUT2 #(
		.INIT('h1)
	) name27841 (
		_w33656_,
		_w33667_,
		_w33668_
	);
	LUT3 #(
		.INIT('h08)
	) name27842 (
		_w33653_,
		_w33656_,
		_w33652_,
		_w33669_
	);
	LUT2 #(
		.INIT('h8)
	) name27843 (
		_w33654_,
		_w33655_,
		_w33670_
	);
	LUT2 #(
		.INIT('h8)
	) name27844 (
		_w33669_,
		_w33670_,
		_w33671_
	);
	LUT4 #(
		.INIT('h0080)
	) name27845 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w33672_
	);
	LUT3 #(
		.INIT('h13)
	) name27846 (
		_w33653_,
		_w33661_,
		_w33672_,
		_w33673_
	);
	LUT3 #(
		.INIT('h10)
	) name27847 (
		_w33668_,
		_w33671_,
		_w33673_,
		_w33674_
	);
	LUT2 #(
		.INIT('h1)
	) name27848 (
		_w33654_,
		_w33655_,
		_w33675_
	);
	LUT4 #(
		.INIT('hfbda)
	) name27849 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w33676_
	);
	LUT4 #(
		.INIT('h0200)
	) name27850 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w33677_
	);
	LUT4 #(
		.INIT('h7dbb)
	) name27851 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w33678_
	);
	LUT4 #(
		.INIT('h0155)
	) name27852 (
		_w33653_,
		_w33676_,
		_w33661_,
		_w33678_,
		_w33679_
	);
	LUT4 #(
		.INIT('h0200)
	) name27853 (
		_w33653_,
		_w33656_,
		_w33654_,
		_w33652_,
		_w33680_
	);
	LUT3 #(
		.INIT('h15)
	) name27854 (
		_w33680_,
		_w33675_,
		_w33669_,
		_w33681_
	);
	LUT2 #(
		.INIT('h4)
	) name27855 (
		_w33679_,
		_w33681_,
		_w33682_
	);
	LUT4 #(
		.INIT('ha955)
	) name27856 (
		\u0_desIn_r_reg[48]/NET0131 ,
		_w33666_,
		_w33674_,
		_w33682_,
		_w33683_
	);
	LUT4 #(
		.INIT('hc963)
	) name27857 (
		decrypt_pad,
		\u0_desIn_r_reg[29]/NET0131 ,
		\u0_key_r_reg[4]/NET0131 ,
		\u0_key_r_reg[54]/NET0131 ,
		_w33684_
	);
	LUT4 #(
		.INIT('hc693)
	) name27858 (
		decrypt_pad,
		\u0_desIn_r_reg[3]/NET0131 ,
		\u0_key_r_reg[13]/NET0131 ,
		\u0_key_r_reg[20]/NET0131 ,
		_w33685_
	);
	LUT4 #(
		.INIT('hc693)
	) name27859 (
		decrypt_pad,
		\u0_desIn_r_reg[37]/NET0131 ,
		\u0_key_r_reg[48]/NET0131 ,
		\u0_key_r_reg[55]/NET0131 ,
		_w33686_
	);
	LUT4 #(
		.INIT('hc693)
	) name27860 (
		decrypt_pad,
		\u0_desIn_r_reg[45]/NET0131 ,
		\u0_key_r_reg[17]/NET0131 ,
		\u0_key_r_reg[24]/NET0131 ,
		_w33687_
	);
	LUT4 #(
		.INIT('h0040)
	) name27861 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33688_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name27862 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33689_
	);
	LUT4 #(
		.INIT('hc693)
	) name27863 (
		decrypt_pad,
		\u0_desIn_r_reg[53]/NET0131 ,
		\u0_key_r_reg[25]/NET0131 ,
		\u0_key_r_reg[32]/NET0131 ,
		_w33690_
	);
	LUT2 #(
		.INIT('h8)
	) name27864 (
		_w33690_,
		_w33686_,
		_w33691_
	);
	LUT4 #(
		.INIT('h2000)
	) name27865 (
		_w33684_,
		_w33685_,
		_w33690_,
		_w33686_,
		_w33692_
	);
	LUT2 #(
		.INIT('h2)
	) name27866 (
		_w33690_,
		_w33686_,
		_w33693_
	);
	LUT4 #(
		.INIT('h0040)
	) name27867 (
		_w33684_,
		_w33685_,
		_w33690_,
		_w33686_,
		_w33694_
	);
	LUT4 #(
		.INIT('hc693)
	) name27868 (
		decrypt_pad,
		\u0_desIn_r_reg[61]/NET0131 ,
		\u0_key_r_reg[33]/NET0131 ,
		\u0_key_r_reg[40]/NET0131 ,
		_w33695_
	);
	LUT3 #(
		.INIT('h10)
	) name27869 (
		_w33694_,
		_w33692_,
		_w33695_,
		_w33696_
	);
	LUT4 #(
		.INIT('h0012)
	) name27870 (
		_w33684_,
		_w33690_,
		_w33686_,
		_w33687_,
		_w33697_
	);
	LUT2 #(
		.INIT('h4)
	) name27871 (
		_w33690_,
		_w33687_,
		_w33698_
	);
	LUT3 #(
		.INIT('h01)
	) name27872 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33699_
	);
	LUT3 #(
		.INIT('h15)
	) name27873 (
		_w33697_,
		_w33698_,
		_w33699_,
		_w33700_
	);
	LUT3 #(
		.INIT('h80)
	) name27874 (
		_w33689_,
		_w33696_,
		_w33700_,
		_w33701_
	);
	LUT4 #(
		.INIT('h0008)
	) name27875 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33702_
	);
	LUT3 #(
		.INIT('h27)
	) name27876 (
		_w33684_,
		_w33685_,
		_w33687_,
		_w33703_
	);
	LUT3 #(
		.INIT('h10)
	) name27877 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33704_
	);
	LUT4 #(
		.INIT('h1000)
	) name27878 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33705_
	);
	LUT4 #(
		.INIT('h000d)
	) name27879 (
		_w33691_,
		_w33703_,
		_w33705_,
		_w33702_,
		_w33706_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name27880 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33707_
	);
	LUT2 #(
		.INIT('h1)
	) name27881 (
		_w33690_,
		_w33707_,
		_w33708_
	);
	LUT3 #(
		.INIT('h0b)
	) name27882 (
		_w33698_,
		_w33699_,
		_w33695_,
		_w33709_
	);
	LUT3 #(
		.INIT('h40)
	) name27883 (
		_w33708_,
		_w33709_,
		_w33706_,
		_w33710_
	);
	LUT4 #(
		.INIT('h0020)
	) name27884 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33711_
	);
	LUT3 #(
		.INIT('he4)
	) name27885 (
		_w33690_,
		_w33688_,
		_w33711_,
		_w33712_
	);
	LUT3 #(
		.INIT('h01)
	) name27886 (
		_w33684_,
		_w33685_,
		_w33687_,
		_w33713_
	);
	LUT3 #(
		.INIT('hde)
	) name27887 (
		_w33684_,
		_w33685_,
		_w33687_,
		_w33714_
	);
	LUT2 #(
		.INIT('h2)
	) name27888 (
		_w33693_,
		_w33714_,
		_w33715_
	);
	LUT2 #(
		.INIT('h1)
	) name27889 (
		_w33712_,
		_w33715_,
		_w33716_
	);
	LUT4 #(
		.INIT('ha955)
	) name27890 (
		\u0_desIn_r_reg[26]/NET0131 ,
		_w33701_,
		_w33710_,
		_w33716_,
		_w33717_
	);
	LUT4 #(
		.INIT('hc963)
	) name27891 (
		decrypt_pad,
		\u0_desIn_r_reg[25]/NET0131 ,
		\u0_key_r_reg[16]/NET0131 ,
		\u0_key_r_reg[9]/NET0131 ,
		_w33718_
	);
	LUT4 #(
		.INIT('hc693)
	) name27892 (
		decrypt_pad,
		\u0_desIn_r_reg[7]/NET0131 ,
		\u0_key_r_reg[21]/NET0131 ,
		\u0_key_r_reg[28]/NET0131 ,
		_w33719_
	);
	LUT4 #(
		.INIT('hc693)
	) name27893 (
		decrypt_pad,
		\u0_desIn_r_reg[33]/NET0131 ,
		\u0_key_r_reg[36]/NET0131 ,
		\u0_key_r_reg[43]/NET0131 ,
		_w33720_
	);
	LUT4 #(
		.INIT('hc693)
	) name27894 (
		decrypt_pad,
		\u0_desIn_r_reg[41]/NET0131 ,
		\u0_key_r_reg[37]/NET0131 ,
		\u0_key_r_reg[44]/NET0131 ,
		_w33721_
	);
	LUT4 #(
		.INIT('hc963)
	) name27895 (
		decrypt_pad,
		\u0_desIn_r_reg[49]/NET0131 ,
		\u0_key_r_reg[1]/NET0131 ,
		\u0_key_r_reg[49]/NET0131 ,
		_w33722_
	);
	LUT4 #(
		.INIT('h7b70)
	) name27896 (
		_w33719_,
		_w33720_,
		_w33721_,
		_w33722_,
		_w33723_
	);
	LUT2 #(
		.INIT('h2)
	) name27897 (
		_w33718_,
		_w33723_,
		_w33724_
	);
	LUT4 #(
		.INIT('hf9fb)
	) name27898 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w33725_
	);
	LUT2 #(
		.INIT('h4)
	) name27899 (
		_w33725_,
		_w33722_,
		_w33726_
	);
	LUT4 #(
		.INIT('hc693)
	) name27900 (
		decrypt_pad,
		\u0_desIn_r_reg[57]/NET0131 ,
		\u0_key_r_reg[0]/NET0131 ,
		\u0_key_r_reg[7]/NET0131 ,
		_w33727_
	);
	LUT3 #(
		.INIT('h0d)
	) name27901 (
		_w33719_,
		_w33720_,
		_w33722_,
		_w33728_
	);
	LUT3 #(
		.INIT('hdc)
	) name27902 (
		_w33718_,
		_w33719_,
		_w33721_,
		_w33729_
	);
	LUT3 #(
		.INIT('h15)
	) name27903 (
		_w33727_,
		_w33728_,
		_w33729_,
		_w33730_
	);
	LUT3 #(
		.INIT('h10)
	) name27904 (
		_w33726_,
		_w33724_,
		_w33730_,
		_w33731_
	);
	LUT4 #(
		.INIT('h0020)
	) name27905 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w33732_
	);
	LUT4 #(
		.INIT('hcf45)
	) name27906 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w33733_
	);
	LUT3 #(
		.INIT('h02)
	) name27907 (
		_w33722_,
		_w33733_,
		_w33732_,
		_w33734_
	);
	LUT4 #(
		.INIT('h0001)
	) name27908 (
		_w33718_,
		_w33720_,
		_w33721_,
		_w33722_,
		_w33735_
	);
	LUT4 #(
		.INIT('h4000)
	) name27909 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w33736_
	);
	LUT3 #(
		.INIT('h02)
	) name27910 (
		_w33727_,
		_w33736_,
		_w33735_,
		_w33737_
	);
	LUT2 #(
		.INIT('h4)
	) name27911 (
		_w33734_,
		_w33737_,
		_w33738_
	);
	LUT4 #(
		.INIT('h0001)
	) name27912 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w33739_
	);
	LUT4 #(
		.INIT('h0400)
	) name27913 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w33740_
	);
	LUT4 #(
		.INIT('hebf7)
	) name27914 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w33741_
	);
	LUT3 #(
		.INIT('h20)
	) name27915 (
		_w33722_,
		_w33739_,
		_w33741_,
		_w33742_
	);
	LUT4 #(
		.INIT('h0800)
	) name27916 (
		_w33727_,
		_w33718_,
		_w33720_,
		_w33721_,
		_w33743_
	);
	LUT3 #(
		.INIT('h01)
	) name27917 (
		_w33722_,
		_w33732_,
		_w33743_,
		_w33744_
	);
	LUT2 #(
		.INIT('h1)
	) name27918 (
		_w33742_,
		_w33744_,
		_w33745_
	);
	LUT4 #(
		.INIT('haa56)
	) name27919 (
		\u0_desIn_r_reg[38]/NET0131 ,
		_w33731_,
		_w33738_,
		_w33745_,
		_w33746_
	);
	LUT4 #(
		.INIT('hc693)
	) name27920 (
		decrypt_pad,
		\u0_desIn_r_reg[29]/NET0131 ,
		\u0_key_r_reg[10]/P0001 ,
		\u0_key_r_reg[17]/NET0131 ,
		_w33747_
	);
	LUT4 #(
		.INIT('hc693)
	) name27921 (
		decrypt_pad,
		\u0_desIn_r_reg[37]/NET0131 ,
		\u0_key_r_reg[55]/NET0131 ,
		\u0_key_r_reg[5]/NET0131 ,
		_w33748_
	);
	LUT4 #(
		.INIT('hc693)
	) name27922 (
		decrypt_pad,
		\u0_desIn_r_reg[63]/NET0131 ,
		\u0_key_r_reg[46]/NET0131 ,
		\u0_key_r_reg[53]/NET0131 ,
		_w33749_
	);
	LUT2 #(
		.INIT('h2)
	) name27923 (
		_w33748_,
		_w33749_,
		_w33750_
	);
	LUT4 #(
		.INIT('hc693)
	) name27924 (
		decrypt_pad,
		\u0_desIn_r_reg[13]/NET0131 ,
		\u0_key_r_reg[26]/NET0131 ,
		\u0_key_r_reg[33]/NET0131 ,
		_w33751_
	);
	LUT4 #(
		.INIT('hc693)
	) name27925 (
		decrypt_pad,
		\u0_desIn_r_reg[5]/NET0131 ,
		\u0_key_r_reg[18]/NET0131 ,
		\u0_key_r_reg[25]/NET0131 ,
		_w33752_
	);
	LUT4 #(
		.INIT('h2000)
	) name27926 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w33753_
	);
	LUT4 #(
		.INIT('hc693)
	) name27927 (
		decrypt_pad,
		\u0_desIn_r_reg[21]/NET0131 ,
		\u0_key_r_reg[27]/NET0131 ,
		\u0_key_r_reg[34]/NET0131 ,
		_w33754_
	);
	LUT2 #(
		.INIT('h6)
	) name27928 (
		_w33748_,
		_w33749_,
		_w33755_
	);
	LUT4 #(
		.INIT('hbf6f)
	) name27929 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w33756_
	);
	LUT3 #(
		.INIT('hd0)
	) name27930 (
		_w33753_,
		_w33754_,
		_w33756_,
		_w33757_
	);
	LUT2 #(
		.INIT('h8)
	) name27931 (
		_w33748_,
		_w33754_,
		_w33758_
	);
	LUT3 #(
		.INIT('h46)
	) name27932 (
		_w33748_,
		_w33749_,
		_w33754_,
		_w33759_
	);
	LUT2 #(
		.INIT('h4)
	) name27933 (
		_w33751_,
		_w33752_,
		_w33760_
	);
	LUT2 #(
		.INIT('h1)
	) name27934 (
		_w33751_,
		_w33752_,
		_w33761_
	);
	LUT2 #(
		.INIT('h8)
	) name27935 (
		_w33759_,
		_w33761_,
		_w33762_
	);
	LUT3 #(
		.INIT('heb)
	) name27936 (
		_w33751_,
		_w33752_,
		_w33759_,
		_w33763_
	);
	LUT3 #(
		.INIT('h15)
	) name27937 (
		_w33747_,
		_w33757_,
		_w33763_,
		_w33764_
	);
	LUT2 #(
		.INIT('h4)
	) name27938 (
		_w33748_,
		_w33749_,
		_w33765_
	);
	LUT4 #(
		.INIT('h9b55)
	) name27939 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w33766_
	);
	LUT2 #(
		.INIT('h8)
	) name27940 (
		_w33747_,
		_w33754_,
		_w33767_
	);
	LUT2 #(
		.INIT('h4)
	) name27941 (
		_w33766_,
		_w33767_,
		_w33768_
	);
	LUT4 #(
		.INIT('h0001)
	) name27942 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w33769_
	);
	LUT4 #(
		.INIT('hff5e)
	) name27943 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w33770_
	);
	LUT2 #(
		.INIT('h2)
	) name27944 (
		_w33754_,
		_w33770_,
		_w33771_
	);
	LUT3 #(
		.INIT('h10)
	) name27945 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33772_
	);
	LUT2 #(
		.INIT('h8)
	) name27946 (
		_w33747_,
		_w33752_,
		_w33773_
	);
	LUT3 #(
		.INIT('h45)
	) name27947 (
		_w33749_,
		_w33751_,
		_w33752_,
		_w33774_
	);
	LUT2 #(
		.INIT('h2)
	) name27948 (
		_w33747_,
		_w33754_,
		_w33775_
	);
	LUT4 #(
		.INIT('h0082)
	) name27949 (
		_w33747_,
		_w33748_,
		_w33752_,
		_w33754_,
		_w33776_
	);
	LUT4 #(
		.INIT('h7077)
	) name27950 (
		_w33772_,
		_w33773_,
		_w33774_,
		_w33776_,
		_w33777_
	);
	LUT3 #(
		.INIT('h10)
	) name27951 (
		_w33771_,
		_w33768_,
		_w33777_,
		_w33778_
	);
	LUT3 #(
		.INIT('h65)
	) name27952 (
		\u0_desIn_r_reg[46]/NET0131 ,
		_w33764_,
		_w33778_,
		_w33779_
	);
	LUT4 #(
		.INIT('hc693)
	) name27953 (
		decrypt_pad,
		\u0_desIn_r_reg[59]/NET0131 ,
		\u0_key_r_reg[28]/NET0131 ,
		\u0_key_r_reg[35]/P0001 ,
		_w33780_
	);
	LUT4 #(
		.INIT('hc693)
	) name27954 (
		decrypt_pad,
		\u0_desIn_r_reg[51]/NET0131 ,
		\u0_key_r_reg[2]/NET0131 ,
		\u0_key_r_reg[9]/NET0131 ,
		_w33781_
	);
	LUT4 #(
		.INIT('hc693)
	) name27955 (
		decrypt_pad,
		\u0_desIn_r_reg[35]/NET0131 ,
		\u0_key_r_reg[22]/NET0131 ,
		\u0_key_r_reg[29]/NET0131 ,
		_w33782_
	);
	LUT4 #(
		.INIT('hc963)
	) name27956 (
		decrypt_pad,
		\u0_desIn_r_reg[27]/NET0131 ,
		\u0_key_r_reg[14]/NET0131 ,
		\u0_key_r_reg[7]/NET0131 ,
		_w33783_
	);
	LUT4 #(
		.INIT('hc693)
	) name27957 (
		decrypt_pad,
		\u0_desIn_r_reg[1]/NET0131 ,
		\u0_key_r_reg[23]/NET0131 ,
		\u0_key_r_reg[30]/NET0131 ,
		_w33784_
	);
	LUT4 #(
		.INIT('hc693)
	) name27958 (
		decrypt_pad,
		\u0_desIn_r_reg[43]/NET0131 ,
		\u0_key_r_reg[44]/NET0131 ,
		\u0_key_r_reg[51]/NET0131 ,
		_w33785_
	);
	LUT4 #(
		.INIT('he65f)
	) name27959 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33786_
	);
	LUT2 #(
		.INIT('h2)
	) name27960 (
		_w33781_,
		_w33786_,
		_w33787_
	);
	LUT4 #(
		.INIT('h0400)
	) name27961 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33788_
	);
	LUT4 #(
		.INIT('hfbaf)
	) name27962 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33789_
	);
	LUT2 #(
		.INIT('h1)
	) name27963 (
		_w33785_,
		_w33781_,
		_w33790_
	);
	LUT4 #(
		.INIT('h0020)
	) name27964 (
		_w33783_,
		_w33785_,
		_w33784_,
		_w33781_,
		_w33791_
	);
	LUT4 #(
		.INIT('h0002)
	) name27965 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33792_
	);
	LUT4 #(
		.INIT('h0032)
	) name27966 (
		_w33781_,
		_w33791_,
		_w33789_,
		_w33792_,
		_w33793_
	);
	LUT3 #(
		.INIT('h45)
	) name27967 (
		_w33780_,
		_w33787_,
		_w33793_,
		_w33794_
	);
	LUT4 #(
		.INIT('heece)
	) name27968 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33795_
	);
	LUT4 #(
		.INIT('h2000)
	) name27969 (
		_w33783_,
		_w33785_,
		_w33784_,
		_w33781_,
		_w33796_
	);
	LUT4 #(
		.INIT('hc010)
	) name27970 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33797_
	);
	LUT4 #(
		.INIT('h000e)
	) name27971 (
		_w33795_,
		_w33781_,
		_w33796_,
		_w33797_,
		_w33798_
	);
	LUT3 #(
		.INIT('h01)
	) name27972 (
		_w33783_,
		_w33782_,
		_w33784_,
		_w33799_
	);
	LUT3 #(
		.INIT('hb6)
	) name27973 (
		_w33783_,
		_w33782_,
		_w33784_,
		_w33800_
	);
	LUT2 #(
		.INIT('h8)
	) name27974 (
		_w33785_,
		_w33781_,
		_w33801_
	);
	LUT4 #(
		.INIT('h4cc4)
	) name27975 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33802_
	);
	LUT4 #(
		.INIT('h00cd)
	) name27976 (
		_w33783_,
		_w33785_,
		_w33784_,
		_w33781_,
		_w33803_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name27977 (
		_w33800_,
		_w33801_,
		_w33802_,
		_w33803_,
		_w33804_
	);
	LUT3 #(
		.INIT('hb0)
	) name27978 (
		_w33798_,
		_w33780_,
		_w33804_,
		_w33805_
	);
	LUT3 #(
		.INIT('h65)
	) name27979 (
		\u0_desIn_r_reg[30]/NET0131 ,
		_w33794_,
		_w33805_,
		_w33806_
	);
	LUT4 #(
		.INIT('hc693)
	) name27980 (
		decrypt_pad,
		\u0_desIn_r_reg[19]/NET0131 ,
		\u0_key_r_reg[1]/NET0131 ,
		\u0_key_r_reg[8]/NET0131 ,
		_w33807_
	);
	LUT4 #(
		.INIT('hc693)
	) name27981 (
		decrypt_pad,
		\u0_desIn_r_reg[61]/NET0131 ,
		\u0_key_r_reg[29]/NET0131 ,
		\u0_key_r_reg[36]/NET0131 ,
		_w33808_
	);
	LUT4 #(
		.INIT('hc693)
	) name27982 (
		decrypt_pad,
		\u0_desIn_r_reg[35]/NET0131 ,
		\u0_key_r_reg[45]/NET0131 ,
		\u0_key_r_reg[52]/NET0131 ,
		_w33809_
	);
	LUT4 #(
		.INIT('hc963)
	) name27983 (
		decrypt_pad,
		\u0_desIn_r_reg[3]/NET0131 ,
		\u0_key_r_reg[31]/NET0131 ,
		\u0_key_r_reg[51]/NET0131 ,
		_w33810_
	);
	LUT4 #(
		.INIT('hc693)
	) name27984 (
		decrypt_pad,
		\u0_desIn_r_reg[11]/NET0131 ,
		\u0_key_r_reg[14]/NET0131 ,
		\u0_key_r_reg[21]/NET0131 ,
		_w33811_
	);
	LUT4 #(
		.INIT('h0800)
	) name27985 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33812_
	);
	LUT4 #(
		.INIT('h0100)
	) name27986 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33813_
	);
	LUT4 #(
		.INIT('hb69d)
	) name27987 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33814_
	);
	LUT3 #(
		.INIT('h02)
	) name27988 (
		_w33810_,
		_w33811_,
		_w33808_,
		_w33815_
	);
	LUT4 #(
		.INIT('h5fe2)
	) name27989 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33816_
	);
	LUT4 #(
		.INIT('h2000)
	) name27990 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33817_
	);
	LUT4 #(
		.INIT('hdffb)
	) name27991 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33818_
	);
	LUT4 #(
		.INIT('he400)
	) name27992 (
		_w33807_,
		_w33814_,
		_w33816_,
		_w33818_,
		_w33819_
	);
	LUT4 #(
		.INIT('hc693)
	) name27993 (
		decrypt_pad,
		\u0_desIn_r_reg[27]/NET0131 ,
		\u0_key_r_reg[16]/NET0131 ,
		\u0_key_r_reg[23]/NET0131 ,
		_w33820_
	);
	LUT2 #(
		.INIT('h1)
	) name27994 (
		_w33819_,
		_w33820_,
		_w33821_
	);
	LUT4 #(
		.INIT('hb15d)
	) name27995 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33822_
	);
	LUT2 #(
		.INIT('h2)
	) name27996 (
		_w33807_,
		_w33822_,
		_w33823_
	);
	LUT2 #(
		.INIT('h1)
	) name27997 (
		_w33807_,
		_w33811_,
		_w33824_
	);
	LUT3 #(
		.INIT('h08)
	) name27998 (
		_w33809_,
		_w33810_,
		_w33808_,
		_w33825_
	);
	LUT3 #(
		.INIT('hf6)
	) name27999 (
		_w33809_,
		_w33810_,
		_w33808_,
		_w33826_
	);
	LUT2 #(
		.INIT('h2)
	) name28000 (
		_w33824_,
		_w33826_,
		_w33827_
	);
	LUT2 #(
		.INIT('h9)
	) name28001 (
		_w33810_,
		_w33811_,
		_w33828_
	);
	LUT4 #(
		.INIT('h1400)
	) name28002 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33829_
	);
	LUT4 #(
		.INIT('h4c00)
	) name28003 (
		_w33807_,
		_w33809_,
		_w33810_,
		_w33808_,
		_w33830_
	);
	LUT3 #(
		.INIT('h13)
	) name28004 (
		_w33828_,
		_w33829_,
		_w33830_,
		_w33831_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name28005 (
		_w33820_,
		_w33823_,
		_w33827_,
		_w33831_,
		_w33832_
	);
	LUT4 #(
		.INIT('hfbef)
	) name28006 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33833_
	);
	LUT4 #(
		.INIT('h0020)
	) name28007 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33834_
	);
	LUT4 #(
		.INIT('hff9f)
	) name28008 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33835_
	);
	LUT3 #(
		.INIT('hd8)
	) name28009 (
		_w33807_,
		_w33833_,
		_w33835_,
		_w33836_
	);
	LUT4 #(
		.INIT('h5655)
	) name28010 (
		\u0_desIn_r_reg[44]/NET0131 ,
		_w33821_,
		_w33832_,
		_w33836_,
		_w33837_
	);
	LUT4 #(
		.INIT('heb73)
	) name28011 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33838_
	);
	LUT2 #(
		.INIT('h1)
	) name28012 (
		_w33781_,
		_w33838_,
		_w33839_
	);
	LUT4 #(
		.INIT('h1fbd)
	) name28013 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33840_
	);
	LUT2 #(
		.INIT('h4)
	) name28014 (
		_w33782_,
		_w33791_,
		_w33841_
	);
	LUT4 #(
		.INIT('haf23)
	) name28015 (
		_w33782_,
		_w33781_,
		_w33791_,
		_w33840_,
		_w33842_
	);
	LUT3 #(
		.INIT('h8a)
	) name28016 (
		_w33780_,
		_w33839_,
		_w33842_,
		_w33843_
	);
	LUT4 #(
		.INIT('h1960)
	) name28017 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33781_,
		_w33844_
	);
	LUT4 #(
		.INIT('h0002)
	) name28018 (
		_w33783_,
		_w33785_,
		_w33784_,
		_w33781_,
		_w33845_
	);
	LUT4 #(
		.INIT('h0800)
	) name28019 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33846_
	);
	LUT4 #(
		.INIT('h1000)
	) name28020 (
		_w33783_,
		_w33782_,
		_w33784_,
		_w33781_,
		_w33847_
	);
	LUT4 #(
		.INIT('h0020)
	) name28021 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33848_
	);
	LUT4 #(
		.INIT('h0001)
	) name28022 (
		_w33847_,
		_w33845_,
		_w33846_,
		_w33848_,
		_w33849_
	);
	LUT3 #(
		.INIT('h45)
	) name28023 (
		_w33780_,
		_w33844_,
		_w33849_,
		_w33850_
	);
	LUT4 #(
		.INIT('h23af)
	) name28024 (
		_w33785_,
		_w33782_,
		_w33847_,
		_w33845_,
		_w33851_
	);
	LUT4 #(
		.INIT('h45cf)
	) name28025 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33852_
	);
	LUT4 #(
		.INIT('hcd00)
	) name28026 (
		_w33783_,
		_w33785_,
		_w33784_,
		_w33781_,
		_w33853_
	);
	LUT4 #(
		.INIT('h7077)
	) name28027 (
		_w33799_,
		_w33790_,
		_w33852_,
		_w33853_,
		_w33854_
	);
	LUT2 #(
		.INIT('h8)
	) name28028 (
		_w33851_,
		_w33854_,
		_w33855_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name28029 (
		\u0_desIn_r_reg[20]/NET0131 ,
		_w33850_,
		_w33843_,
		_w33855_,
		_w33856_
	);
	LUT3 #(
		.INIT('h02)
	) name28030 (
		_w33690_,
		_w33704_,
		_w33702_,
		_w33857_
	);
	LUT4 #(
		.INIT('h2202)
	) name28031 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33858_
	);
	LUT3 #(
		.INIT('h01)
	) name28032 (
		_w33690_,
		_w33688_,
		_w33858_,
		_w33859_
	);
	LUT3 #(
		.INIT('h90)
	) name28033 (
		_w33684_,
		_w33686_,
		_w33687_,
		_w33860_
	);
	LUT4 #(
		.INIT('h8400)
	) name28034 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33861_
	);
	LUT4 #(
		.INIT('haa02)
	) name28035 (
		_w33695_,
		_w33857_,
		_w33859_,
		_w33861_,
		_w33862_
	);
	LUT3 #(
		.INIT('hd1)
	) name28036 (
		_w33690_,
		_w33686_,
		_w33687_,
		_w33863_
	);
	LUT4 #(
		.INIT('haaa2)
	) name28037 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33864_
	);
	LUT2 #(
		.INIT('h4)
	) name28038 (
		_w33863_,
		_w33864_,
		_w33865_
	);
	LUT2 #(
		.INIT('h8)
	) name28039 (
		_w33690_,
		_w33687_,
		_w33866_
	);
	LUT4 #(
		.INIT('hbfae)
	) name28040 (
		_w33684_,
		_w33685_,
		_w33690_,
		_w33686_,
		_w33867_
	);
	LUT4 #(
		.INIT('h0008)
	) name28041 (
		_w33684_,
		_w33685_,
		_w33690_,
		_w33687_,
		_w33868_
	);
	LUT4 #(
		.INIT('h0054)
	) name28042 (
		_w33705_,
		_w33866_,
		_w33867_,
		_w33868_,
		_w33869_
	);
	LUT3 #(
		.INIT('h45)
	) name28043 (
		_w33695_,
		_w33865_,
		_w33869_,
		_w33870_
	);
	LUT4 #(
		.INIT('h4000)
	) name28044 (
		_w33684_,
		_w33690_,
		_w33686_,
		_w33687_,
		_w33871_
	);
	LUT4 #(
		.INIT('h0001)
	) name28045 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33872_
	);
	LUT4 #(
		.INIT('hddd8)
	) name28046 (
		_w33690_,
		_w33711_,
		_w33861_,
		_w33872_,
		_w33873_
	);
	LUT2 #(
		.INIT('h1)
	) name28047 (
		_w33871_,
		_w33873_,
		_w33874_
	);
	LUT4 #(
		.INIT('h5655)
	) name28048 (
		\u0_desIn_r_reg[12]/NET0131 ,
		_w33862_,
		_w33870_,
		_w33874_,
		_w33875_
	);
	LUT4 #(
		.INIT('hdd75)
	) name28049 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33876_
	);
	LUT3 #(
		.INIT('h32)
	) name28050 (
		_w33807_,
		_w33815_,
		_w33876_,
		_w33877_
	);
	LUT4 #(
		.INIT('h76ff)
	) name28051 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33878_
	);
	LUT4 #(
		.INIT('hbfef)
	) name28052 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33879_
	);
	LUT3 #(
		.INIT('hd0)
	) name28053 (
		_w33807_,
		_w33878_,
		_w33879_,
		_w33880_
	);
	LUT3 #(
		.INIT('h15)
	) name28054 (
		_w33820_,
		_w33877_,
		_w33880_,
		_w33881_
	);
	LUT4 #(
		.INIT('hddfe)
	) name28055 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33882_
	);
	LUT3 #(
		.INIT('h10)
	) name28056 (
		_w33807_,
		_w33811_,
		_w33808_,
		_w33883_
	);
	LUT4 #(
		.INIT('h00c4)
	) name28057 (
		_w33807_,
		_w33835_,
		_w33882_,
		_w33883_,
		_w33884_
	);
	LUT3 #(
		.INIT('h40)
	) name28058 (
		_w33810_,
		_w33811_,
		_w33808_,
		_w33885_
	);
	LUT4 #(
		.INIT('hbf97)
	) name28059 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33886_
	);
	LUT4 #(
		.INIT('hef45)
	) name28060 (
		_w33807_,
		_w33809_,
		_w33885_,
		_w33886_,
		_w33887_
	);
	LUT3 #(
		.INIT('hd0)
	) name28061 (
		_w33820_,
		_w33884_,
		_w33887_,
		_w33888_
	);
	LUT3 #(
		.INIT('h65)
	) name28062 (
		\u0_desIn_r_reg[62]/NET0131 ,
		_w33881_,
		_w33888_,
		_w33889_
	);
	LUT3 #(
		.INIT('h02)
	) name28063 (
		_w33690_,
		_w33688_,
		_w33702_,
		_w33890_
	);
	LUT4 #(
		.INIT('h0092)
	) name28064 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33891_
	);
	LUT3 #(
		.INIT('h8c)
	) name28065 (
		_w33684_,
		_w33685_,
		_w33687_,
		_w33892_
	);
	LUT2 #(
		.INIT('h1)
	) name28066 (
		_w33686_,
		_w33695_,
		_w33893_
	);
	LUT4 #(
		.INIT('h0045)
	) name28067 (
		_w33690_,
		_w33892_,
		_w33893_,
		_w33891_,
		_w33894_
	);
	LUT2 #(
		.INIT('h1)
	) name28068 (
		_w33890_,
		_w33894_,
		_w33895_
	);
	LUT3 #(
		.INIT('hb0)
	) name28069 (
		_w33684_,
		_w33685_,
		_w33687_,
		_w33896_
	);
	LUT2 #(
		.INIT('h8)
	) name28070 (
		_w33691_,
		_w33896_,
		_w33897_
	);
	LUT3 #(
		.INIT('h02)
	) name28071 (
		_w33684_,
		_w33686_,
		_w33687_,
		_w33898_
	);
	LUT3 #(
		.INIT('h01)
	) name28072 (
		_w33688_,
		_w33692_,
		_w33898_,
		_w33899_
	);
	LUT3 #(
		.INIT('h45)
	) name28073 (
		_w33695_,
		_w33897_,
		_w33899_,
		_w33900_
	);
	LUT4 #(
		.INIT('h7773)
	) name28074 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w33901_
	);
	LUT2 #(
		.INIT('h1)
	) name28075 (
		_w33690_,
		_w33901_,
		_w33902_
	);
	LUT3 #(
		.INIT('h0b)
	) name28076 (
		_w33684_,
		_w33690_,
		_w33686_,
		_w33903_
	);
	LUT3 #(
		.INIT('h01)
	) name28077 (
		_w33705_,
		_w33892_,
		_w33903_,
		_w33904_
	);
	LUT3 #(
		.INIT('hd0)
	) name28078 (
		_w33684_,
		_w33687_,
		_w33695_,
		_w33905_
	);
	LUT3 #(
		.INIT('he0)
	) name28079 (
		_w33902_,
		_w33904_,
		_w33905_,
		_w33906_
	);
	LUT4 #(
		.INIT('h5556)
	) name28080 (
		\u0_desIn_r_reg[8]/NET0131 ,
		_w33895_,
		_w33900_,
		_w33906_,
		_w33907_
	);
	LUT4 #(
		.INIT('hc693)
	) name28081 (
		decrypt_pad,
		\u0_desIn_r_reg[55]/NET0131 ,
		\u0_key_r_reg[41]/NET0131 ,
		\u0_key_r_reg[48]/NET0131 ,
		_w33908_
	);
	LUT4 #(
		.INIT('hc693)
	) name28082 (
		decrypt_pad,
		\u0_desIn_r_reg[39]/NET0131 ,
		\u0_key_r_reg[24]/NET0131 ,
		\u0_key_r_reg[6]/NET0131 ,
		_w33909_
	);
	LUT4 #(
		.INIT('hc693)
	) name28083 (
		decrypt_pad,
		\u0_desIn_r_reg[5]/NET0131 ,
		\u0_key_r_reg[12]/NET0131 ,
		\u0_key_r_reg[19]/NET0131 ,
		_w33910_
	);
	LUT4 #(
		.INIT('hc693)
	) name28084 (
		decrypt_pad,
		\u0_desIn_r_reg[47]/NET0131 ,
		\u0_key_r_reg[47]/NET0131 ,
		\u0_key_r_reg[54]/NET0131 ,
		_w33911_
	);
	LUT4 #(
		.INIT('h0004)
	) name28085 (
		_w33908_,
		_w33910_,
		_w33909_,
		_w33911_,
		_w33912_
	);
	LUT4 #(
		.INIT('hc693)
	) name28086 (
		decrypt_pad,
		\u0_desIn_r_reg[31]/NET0131 ,
		\u0_key_r_reg[20]/NET0131 ,
		\u0_key_r_reg[27]/NET0131 ,
		_w33913_
	);
	LUT2 #(
		.INIT('h2)
	) name28087 (
		_w33910_,
		_w33913_,
		_w33914_
	);
	LUT4 #(
		.INIT('h0800)
	) name28088 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33915_
	);
	LUT2 #(
		.INIT('h1)
	) name28089 (
		_w33912_,
		_w33915_,
		_w33916_
	);
	LUT4 #(
		.INIT('hc693)
	) name28090 (
		decrypt_pad,
		\u0_desIn_r_reg[63]/NET0131 ,
		\u0_key_r_reg[32]/NET0131 ,
		\u0_key_r_reg[39]/P0001 ,
		_w33917_
	);
	LUT2 #(
		.INIT('h2)
	) name28091 (
		_w33910_,
		_w33909_,
		_w33918_
	);
	LUT3 #(
		.INIT('h80)
	) name28092 (
		_w33908_,
		_w33913_,
		_w33911_,
		_w33919_
	);
	LUT3 #(
		.INIT('h15)
	) name28093 (
		_w33917_,
		_w33918_,
		_w33919_,
		_w33920_
	);
	LUT2 #(
		.INIT('h4)
	) name28094 (
		_w33910_,
		_w33909_,
		_w33921_
	);
	LUT4 #(
		.INIT('h0046)
	) name28095 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33922_
	);
	LUT4 #(
		.INIT('h5155)
	) name28096 (
		_w33908_,
		_w33910_,
		_w33909_,
		_w33913_,
		_w33923_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name28097 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33924_
	);
	LUT3 #(
		.INIT('h51)
	) name28098 (
		_w33922_,
		_w33923_,
		_w33924_,
		_w33925_
	);
	LUT3 #(
		.INIT('h80)
	) name28099 (
		_w33916_,
		_w33920_,
		_w33925_,
		_w33926_
	);
	LUT2 #(
		.INIT('h4)
	) name28100 (
		_w33908_,
		_w33911_,
		_w33927_
	);
	LUT3 #(
		.INIT('hda)
	) name28101 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33928_
	);
	LUT2 #(
		.INIT('h2)
	) name28102 (
		_w33927_,
		_w33928_,
		_w33929_
	);
	LUT4 #(
		.INIT('h8088)
	) name28103 (
		_w33908_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33930_
	);
	LUT4 #(
		.INIT('h0001)
	) name28104 (
		_w33908_,
		_w33910_,
		_w33909_,
		_w33913_,
		_w33931_
	);
	LUT2 #(
		.INIT('h2)
	) name28105 (
		_w33913_,
		_w33911_,
		_w33932_
	);
	LUT3 #(
		.INIT('h04)
	) name28106 (
		_w33910_,
		_w33913_,
		_w33911_,
		_w33933_
	);
	LUT4 #(
		.INIT('h0010)
	) name28107 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33934_
	);
	LUT4 #(
		.INIT('hff6f)
	) name28108 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33935_
	);
	LUT4 #(
		.INIT('h0200)
	) name28109 (
		_w33917_,
		_w33931_,
		_w33930_,
		_w33935_,
		_w33936_
	);
	LUT2 #(
		.INIT('h4)
	) name28110 (
		_w33929_,
		_w33936_,
		_w33937_
	);
	LUT4 #(
		.INIT('h0100)
	) name28111 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33938_
	);
	LUT4 #(
		.INIT('hfe3f)
	) name28112 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33939_
	);
	LUT3 #(
		.INIT('hae)
	) name28113 (
		_w33908_,
		_w33909_,
		_w33911_,
		_w33940_
	);
	LUT4 #(
		.INIT('h080a)
	) name28114 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33941_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name28115 (
		_w33908_,
		_w33939_,
		_w33940_,
		_w33941_,
		_w33942_
	);
	LUT4 #(
		.INIT('ha955)
	) name28116 (
		\u0_desIn_r_reg[14]/NET0131 ,
		_w33926_,
		_w33937_,
		_w33942_,
		_w33943_
	);
	LUT4 #(
		.INIT('hf7f2)
	) name28117 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33944_
	);
	LUT4 #(
		.INIT('h0551)
	) name28118 (
		_w33908_,
		_w33910_,
		_w33909_,
		_w33913_,
		_w33945_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name28119 (
		_w33908_,
		_w33933_,
		_w33944_,
		_w33945_,
		_w33946_
	);
	LUT4 #(
		.INIT('h9eff)
	) name28120 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33947_
	);
	LUT3 #(
		.INIT('h45)
	) name28121 (
		_w33917_,
		_w33946_,
		_w33947_,
		_w33948_
	);
	LUT3 #(
		.INIT('hb0)
	) name28122 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33949_
	);
	LUT3 #(
		.INIT('h04)
	) name28123 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33950_
	);
	LUT4 #(
		.INIT('h6b6f)
	) name28124 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33951_
	);
	LUT2 #(
		.INIT('h2)
	) name28125 (
		_w33908_,
		_w33951_,
		_w33952_
	);
	LUT2 #(
		.INIT('h1)
	) name28126 (
		_w33908_,
		_w33944_,
		_w33953_
	);
	LUT3 #(
		.INIT('h51)
	) name28127 (
		_w33908_,
		_w33910_,
		_w33909_,
		_w33954_
	);
	LUT4 #(
		.INIT('h0200)
	) name28128 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w33955_
	);
	LUT3 #(
		.INIT('h0d)
	) name28129 (
		_w33932_,
		_w33954_,
		_w33955_,
		_w33956_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name28130 (
		_w33917_,
		_w33953_,
		_w33952_,
		_w33956_,
		_w33957_
	);
	LUT3 #(
		.INIT('h23)
	) name28131 (
		_w33909_,
		_w33913_,
		_w33911_,
		_w33958_
	);
	LUT3 #(
		.INIT('h51)
	) name28132 (
		_w33908_,
		_w33913_,
		_w33911_,
		_w33959_
	);
	LUT3 #(
		.INIT('h10)
	) name28133 (
		_w33949_,
		_w33958_,
		_w33959_,
		_w33960_
	);
	LUT4 #(
		.INIT('h5556)
	) name28134 (
		\u0_desIn_r_reg[24]/NET0131 ,
		_w33957_,
		_w33960_,
		_w33948_,
		_w33961_
	);
	LUT4 #(
		.INIT('h768c)
	) name28135 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33962_
	);
	LUT4 #(
		.INIT('hddf3)
	) name28136 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33963_
	);
	LUT4 #(
		.INIT('hb7f7)
	) name28137 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33964_
	);
	LUT4 #(
		.INIT('he400)
	) name28138 (
		_w33807_,
		_w33963_,
		_w33962_,
		_w33964_,
		_w33965_
	);
	LUT2 #(
		.INIT('h2)
	) name28139 (
		_w33820_,
		_w33965_,
		_w33966_
	);
	LUT3 #(
		.INIT('h8a)
	) name28140 (
		_w33807_,
		_w33809_,
		_w33810_,
		_w33967_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name28141 (
		_w33807_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33968_
	);
	LUT2 #(
		.INIT('h4)
	) name28142 (
		_w33967_,
		_w33968_,
		_w33969_
	);
	LUT4 #(
		.INIT('h0080)
	) name28143 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33970_
	);
	LUT3 #(
		.INIT('h23)
	) name28144 (
		_w33809_,
		_w33810_,
		_w33808_,
		_w33971_
	);
	LUT4 #(
		.INIT('h1151)
	) name28145 (
		_w33807_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33972_
	);
	LUT3 #(
		.INIT('h45)
	) name28146 (
		_w33970_,
		_w33971_,
		_w33972_,
		_w33973_
	);
	LUT4 #(
		.INIT('hbfed)
	) name28147 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w33974_
	);
	LUT4 #(
		.INIT('h2301)
	) name28148 (
		_w33807_,
		_w33812_,
		_w33885_,
		_w33974_,
		_w33975_
	);
	LUT4 #(
		.INIT('hba00)
	) name28149 (
		_w33820_,
		_w33969_,
		_w33973_,
		_w33975_,
		_w33976_
	);
	LUT3 #(
		.INIT('h65)
	) name28150 (
		\u0_desIn_r_reg[0]/NET0131 ,
		_w33966_,
		_w33976_,
		_w33977_
	);
	LUT4 #(
		.INIT('h55fe)
	) name28151 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33978_
	);
	LUT2 #(
		.INIT('h2)
	) name28152 (
		_w33629_,
		_w33978_,
		_w33979_
	);
	LUT3 #(
		.INIT('h40)
	) name28153 (
		_w33625_,
		_w33624_,
		_w33627_,
		_w33980_
	);
	LUT4 #(
		.INIT('h1020)
	) name28154 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33981_
	);
	LUT2 #(
		.INIT('h2)
	) name28155 (
		_w33623_,
		_w33981_,
		_w33982_
	);
	LUT4 #(
		.INIT('h0408)
	) name28156 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33983_
	);
	LUT3 #(
		.INIT('h0b)
	) name28157 (
		_w33629_,
		_w33634_,
		_w33983_,
		_w33984_
	);
	LUT3 #(
		.INIT('h40)
	) name28158 (
		_w33979_,
		_w33982_,
		_w33984_,
		_w33985_
	);
	LUT4 #(
		.INIT('h4000)
	) name28159 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33986_
	);
	LUT4 #(
		.INIT('h0040)
	) name28160 (
		_w33625_,
		_w33626_,
		_w33629_,
		_w33627_,
		_w33987_
	);
	LUT4 #(
		.INIT('h0012)
	) name28161 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33988_
	);
	LUT4 #(
		.INIT('h0001)
	) name28162 (
		_w33623_,
		_w33986_,
		_w33987_,
		_w33988_,
		_w33989_
	);
	LUT4 #(
		.INIT('h0180)
	) name28163 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33990_
	);
	LUT2 #(
		.INIT('h6)
	) name28164 (
		_w33626_,
		_w33627_,
		_w33991_
	);
	LUT4 #(
		.INIT('h134c)
	) name28165 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w33992_
	);
	LUT3 #(
		.INIT('h32)
	) name28166 (
		_w33629_,
		_w33990_,
		_w33992_,
		_w33993_
	);
	LUT2 #(
		.INIT('h8)
	) name28167 (
		_w33989_,
		_w33993_,
		_w33994_
	);
	LUT3 #(
		.INIT('ha9)
	) name28168 (
		\u0_desIn_r_reg[28]/NET0131 ,
		_w33985_,
		_w33994_,
		_w33995_
	);
	LUT4 #(
		.INIT('haf6f)
	) name28169 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33996_
	);
	LUT2 #(
		.INIT('h2)
	) name28170 (
		_w33781_,
		_w33996_,
		_w33997_
	);
	LUT4 #(
		.INIT('h77ba)
	) name28171 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w33998_
	);
	LUT2 #(
		.INIT('h1)
	) name28172 (
		_w33781_,
		_w33998_,
		_w33999_
	);
	LUT4 #(
		.INIT('h0104)
	) name28173 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w34000_
	);
	LUT3 #(
		.INIT('h01)
	) name28174 (
		_w33845_,
		_w33846_,
		_w34000_,
		_w34001_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name28175 (
		_w33780_,
		_w33997_,
		_w33999_,
		_w34001_,
		_w34002_
	);
	LUT4 #(
		.INIT('hcd6f)
	) name28176 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w34003_
	);
	LUT4 #(
		.INIT('h5fb4)
	) name28177 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w34004_
	);
	LUT4 #(
		.INIT('h3120)
	) name28178 (
		_w33781_,
		_w33788_,
		_w34004_,
		_w34003_,
		_w34005_
	);
	LUT4 #(
		.INIT('h4000)
	) name28179 (
		_w33785_,
		_w33782_,
		_w33784_,
		_w33781_,
		_w34006_
	);
	LUT2 #(
		.INIT('h1)
	) name28180 (
		_w33792_,
		_w34006_,
		_w34007_
	);
	LUT3 #(
		.INIT('he0)
	) name28181 (
		_w33780_,
		_w34005_,
		_w34007_,
		_w34008_
	);
	LUT3 #(
		.INIT('h9a)
	) name28182 (
		\u0_desIn_r_reg[32]/NET0131 ,
		_w34002_,
		_w34008_,
		_w34009_
	);
	LUT4 #(
		.INIT('h082a)
	) name28183 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w34010_
	);
	LUT4 #(
		.INIT('h0200)
	) name28184 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w34011_
	);
	LUT4 #(
		.INIT('hfad8)
	) name28185 (
		_w33690_,
		_w33713_,
		_w34010_,
		_w34011_,
		_w34012_
	);
	LUT4 #(
		.INIT('h7f9f)
	) name28186 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w34013_
	);
	LUT3 #(
		.INIT('h45)
	) name28187 (
		_w33695_,
		_w34012_,
		_w34013_,
		_w34014_
	);
	LUT4 #(
		.INIT('h9400)
	) name28188 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w34015_
	);
	LUT4 #(
		.INIT('hf3f1)
	) name28189 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w34016_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name28190 (
		_w33690_,
		_w33695_,
		_w34015_,
		_w34016_,
		_w34017_
	);
	LUT4 #(
		.INIT('h2500)
	) name28191 (
		_w33684_,
		_w33685_,
		_w33686_,
		_w33687_,
		_w34018_
	);
	LUT4 #(
		.INIT('h0d00)
	) name28192 (
		_w33684_,
		_w33685_,
		_w33690_,
		_w33686_,
		_w34019_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name28193 (
		_w33695_,
		_w33896_,
		_w34018_,
		_w34019_,
		_w34020_
	);
	LUT2 #(
		.INIT('h1)
	) name28194 (
		_w33685_,
		_w33690_,
		_w34021_
	);
	LUT2 #(
		.INIT('h8)
	) name28195 (
		_w33860_,
		_w34021_,
		_w34022_
	);
	LUT3 #(
		.INIT('h01)
	) name28196 (
		_w34017_,
		_w34020_,
		_w34022_,
		_w34023_
	);
	LUT3 #(
		.INIT('h65)
	) name28197 (
		\u0_desIn_r_reg[6]/NET0131 ,
		_w34014_,
		_w34023_,
		_w34024_
	);
	LUT4 #(
		.INIT('h1000)
	) name28198 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34025_
	);
	LUT4 #(
		.INIT('he1f1)
	) name28199 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34026_
	);
	LUT2 #(
		.INIT('h2)
	) name28200 (
		_w33653_,
		_w34026_,
		_w34027_
	);
	LUT4 #(
		.INIT('h0040)
	) name28201 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34028_
	);
	LUT4 #(
		.INIT('h4401)
	) name28202 (
		_w33653_,
		_w33656_,
		_w33654_,
		_w33652_,
		_w34029_
	);
	LUT3 #(
		.INIT('h80)
	) name28203 (
		_w33656_,
		_w33654_,
		_w33655_,
		_w34030_
	);
	LUT4 #(
		.INIT('h0002)
	) name28204 (
		_w33661_,
		_w34028_,
		_w34029_,
		_w34030_,
		_w34031_
	);
	LUT4 #(
		.INIT('h0408)
	) name28205 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34032_
	);
	LUT2 #(
		.INIT('h9)
	) name28206 (
		_w33654_,
		_w33655_,
		_w34033_
	);
	LUT4 #(
		.INIT('h2a8a)
	) name28207 (
		_w33653_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34034_
	);
	LUT3 #(
		.INIT('h41)
	) name28208 (
		_w33654_,
		_w33652_,
		_w33655_,
		_w34035_
	);
	LUT4 #(
		.INIT('h5554)
	) name28209 (
		_w33653_,
		_w33656_,
		_w33652_,
		_w33655_,
		_w34036_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name28210 (
		_w34032_,
		_w34034_,
		_w34035_,
		_w34036_,
		_w34037_
	);
	LUT3 #(
		.INIT('h01)
	) name28211 (
		_w33677_,
		_w33661_,
		_w33672_,
		_w34038_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name28212 (
		_w34027_,
		_w34031_,
		_w34037_,
		_w34038_,
		_w34039_
	);
	LUT2 #(
		.INIT('h6)
	) name28213 (
		\u0_desIn_r_reg[2]/NET0131 ,
		_w34039_,
		_w34040_
	);
	LUT3 #(
		.INIT('h0e)
	) name28214 (
		_w33908_,
		_w33909_,
		_w33911_,
		_w34041_
	);
	LUT4 #(
		.INIT('h51f3)
	) name28215 (
		_w33914_,
		_w33919_,
		_w33921_,
		_w34041_,
		_w34042_
	);
	LUT2 #(
		.INIT('h1)
	) name28216 (
		_w33908_,
		_w33917_,
		_w34043_
	);
	LUT4 #(
		.INIT('h0100)
	) name28217 (
		_w33934_,
		_w33950_,
		_w33955_,
		_w34043_,
		_w34044_
	);
	LUT3 #(
		.INIT('h10)
	) name28218 (
		_w33910_,
		_w33909_,
		_w33911_,
		_w34045_
	);
	LUT3 #(
		.INIT('h20)
	) name28219 (
		_w33910_,
		_w33913_,
		_w33911_,
		_w34046_
	);
	LUT4 #(
		.INIT('haaa8)
	) name28220 (
		_w33908_,
		_w33910_,
		_w33909_,
		_w33911_,
		_w34047_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name28221 (
		_w33923_,
		_w34045_,
		_w34046_,
		_w34047_,
		_w34048_
	);
	LUT4 #(
		.INIT('h0004)
	) name28222 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w34049_
	);
	LUT4 #(
		.INIT('h0010)
	) name28223 (
		_w33912_,
		_w33915_,
		_w33917_,
		_w34049_,
		_w34050_
	);
	LUT4 #(
		.INIT('h7077)
	) name28224 (
		_w34042_,
		_w34044_,
		_w34048_,
		_w34050_,
		_w34051_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name28225 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w34052_
	);
	LUT3 #(
		.INIT('h21)
	) name28226 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w34053_
	);
	LUT4 #(
		.INIT('h0040)
	) name28227 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w34054_
	);
	LUT2 #(
		.INIT('h2)
	) name28228 (
		_w33908_,
		_w33917_,
		_w34055_
	);
	LUT2 #(
		.INIT('h4)
	) name28229 (
		_w34054_,
		_w34055_,
		_w34056_
	);
	LUT3 #(
		.INIT('h20)
	) name28230 (
		_w34042_,
		_w34053_,
		_w34056_,
		_w34057_
	);
	LUT4 #(
		.INIT('h559a)
	) name28231 (
		\u0_desIn_r_reg[36]/NET0131 ,
		_w34051_,
		_w34052_,
		_w34057_,
		_w34058_
	);
	LUT4 #(
		.INIT('h0041)
	) name28232 (
		_w33783_,
		_w33782_,
		_w33784_,
		_w33781_,
		_w34059_
	);
	LUT4 #(
		.INIT('h7525)
	) name28233 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w34060_
	);
	LUT4 #(
		.INIT('h8000)
	) name28234 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w34061_
	);
	LUT4 #(
		.INIT('h0301)
	) name28235 (
		_w33781_,
		_w33780_,
		_w34061_,
		_w34060_,
		_w34062_
	);
	LUT4 #(
		.INIT('hfb00)
	) name28236 (
		_w33785_,
		_w33782_,
		_w33784_,
		_w33780_,
		_w34063_
	);
	LUT4 #(
		.INIT('hefdd)
	) name28237 (
		_w33783_,
		_w33782_,
		_w33784_,
		_w33781_,
		_w34064_
	);
	LUT4 #(
		.INIT('h2000)
	) name28238 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33781_,
		_w34065_
	);
	LUT4 #(
		.INIT('hbefb)
	) name28239 (
		_w33783_,
		_w33785_,
		_w33782_,
		_w33784_,
		_w34066_
	);
	LUT4 #(
		.INIT('h4000)
	) name28240 (
		_w34065_,
		_w34063_,
		_w34064_,
		_w34066_,
		_w34067_
	);
	LUT3 #(
		.INIT('h0b)
	) name28241 (
		_w34059_,
		_w34062_,
		_w34067_,
		_w34068_
	);
	LUT2 #(
		.INIT('h2)
	) name28242 (
		_w33851_,
		_w33841_,
		_w34069_
	);
	LUT3 #(
		.INIT('h65)
	) name28243 (
		\u0_desIn_r_reg[18]/NET0131 ,
		_w34068_,
		_w34069_,
		_w34070_
	);
	LUT4 #(
		.INIT('h1f3f)
	) name28244 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34071_
	);
	LUT2 #(
		.INIT('h1)
	) name28245 (
		_w33653_,
		_w34071_,
		_w34072_
	);
	LUT4 #(
		.INIT('h0800)
	) name28246 (
		_w33653_,
		_w33656_,
		_w33652_,
		_w33655_,
		_w34073_
	);
	LUT4 #(
		.INIT('h0008)
	) name28247 (
		_w33653_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34074_
	);
	LUT3 #(
		.INIT('h7e)
	) name28248 (
		_w33656_,
		_w33654_,
		_w33655_,
		_w34075_
	);
	LUT3 #(
		.INIT('h10)
	) name28249 (
		_w34074_,
		_w34073_,
		_w34075_,
		_w34076_
	);
	LUT3 #(
		.INIT('h45)
	) name28250 (
		_w33661_,
		_w34072_,
		_w34076_,
		_w34077_
	);
	LUT4 #(
		.INIT('hfcd3)
	) name28251 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34078_
	);
	LUT4 #(
		.INIT('h7ebf)
	) name28252 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34079_
	);
	LUT4 #(
		.INIT('h0455)
	) name28253 (
		_w33653_,
		_w33661_,
		_w34078_,
		_w34079_,
		_w34080_
	);
	LUT3 #(
		.INIT('hb9)
	) name28254 (
		_w33654_,
		_w33652_,
		_w33655_,
		_w34081_
	);
	LUT2 #(
		.INIT('h2)
	) name28255 (
		_w33662_,
		_w34081_,
		_w34082_
	);
	LUT4 #(
		.INIT('h0a08)
	) name28256 (
		_w33653_,
		_w33656_,
		_w33652_,
		_w33655_,
		_w34083_
	);
	LUT2 #(
		.INIT('h8)
	) name28257 (
		_w34033_,
		_w34083_,
		_w34084_
	);
	LUT3 #(
		.INIT('h07)
	) name28258 (
		_w33653_,
		_w33672_,
		_w34025_,
		_w34085_
	);
	LUT4 #(
		.INIT('h1311)
	) name28259 (
		_w33661_,
		_w34082_,
		_w34084_,
		_w34085_,
		_w34086_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name28260 (
		\u0_desIn_r_reg[50]/NET0131 ,
		_w34080_,
		_w34077_,
		_w34086_,
		_w34087_
	);
	LUT4 #(
		.INIT('h0800)
	) name28261 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34088_
	);
	LUT4 #(
		.INIT('hf7dd)
	) name28262 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34089_
	);
	LUT4 #(
		.INIT('h1fb3)
	) name28263 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34090_
	);
	LUT4 #(
		.INIT('h0004)
	) name28264 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34091_
	);
	LUT4 #(
		.INIT('hdefb)
	) name28265 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34092_
	);
	LUT4 #(
		.INIT('hd800)
	) name28266 (
		_w33722_,
		_w34090_,
		_w34089_,
		_w34092_,
		_w34093_
	);
	LUT2 #(
		.INIT('h2)
	) name28267 (
		_w33727_,
		_w34093_,
		_w34094_
	);
	LUT4 #(
		.INIT('hd5df)
	) name28268 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34095_
	);
	LUT2 #(
		.INIT('h2)
	) name28269 (
		_w33722_,
		_w34095_,
		_w34096_
	);
	LUT4 #(
		.INIT('hadff)
	) name28270 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34097_
	);
	LUT2 #(
		.INIT('h2)
	) name28271 (
		_w33720_,
		_w33722_,
		_w34098_
	);
	LUT4 #(
		.INIT('h0010)
	) name28272 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33722_,
		_w34099_
	);
	LUT4 #(
		.INIT('h0040)
	) name28273 (
		_w33718_,
		_w33719_,
		_w33721_,
		_w33722_,
		_w34100_
	);
	LUT3 #(
		.INIT('h10)
	) name28274 (
		_w34099_,
		_w34100_,
		_w34097_,
		_w34101_
	);
	LUT2 #(
		.INIT('h4)
	) name28275 (
		_w33720_,
		_w33722_,
		_w34102_
	);
	LUT3 #(
		.INIT('h08)
	) name28276 (
		_w33718_,
		_w33719_,
		_w33721_,
		_w34103_
	);
	LUT3 #(
		.INIT('h45)
	) name28277 (
		_w33739_,
		_w34102_,
		_w34103_,
		_w34104_
	);
	LUT4 #(
		.INIT('h4555)
	) name28278 (
		_w33727_,
		_w34096_,
		_w34101_,
		_w34104_,
		_w34105_
	);
	LUT4 #(
		.INIT('h0100)
	) name28279 (
		_w33718_,
		_w33720_,
		_w33721_,
		_w33722_,
		_w34106_
	);
	LUT3 #(
		.INIT('h07)
	) name28280 (
		_w34098_,
		_w34103_,
		_w34106_,
		_w34107_
	);
	LUT4 #(
		.INIT('h5655)
	) name28281 (
		\u0_desIn_r_reg[34]/NET0131 ,
		_w34105_,
		_w34094_,
		_w34107_,
		_w34108_
	);
	LUT3 #(
		.INIT('h80)
	) name28282 (
		_w33748_,
		_w33749_,
		_w33752_,
		_w34109_
	);
	LUT4 #(
		.INIT('h6979)
	) name28283 (
		_w33748_,
		_w33749_,
		_w33752_,
		_w33754_,
		_w34110_
	);
	LUT4 #(
		.INIT('h0014)
	) name28284 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33754_,
		_w34111_
	);
	LUT4 #(
		.INIT('h0032)
	) name28285 (
		_w33751_,
		_w33753_,
		_w34110_,
		_w34111_,
		_w34112_
	);
	LUT4 #(
		.INIT('h76dc)
	) name28286 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w34113_
	);
	LUT3 #(
		.INIT('he0)
	) name28287 (
		_w33748_,
		_w33749_,
		_w33754_,
		_w34114_
	);
	LUT4 #(
		.INIT('h6800)
	) name28288 (
		_w33748_,
		_w33749_,
		_w33752_,
		_w33754_,
		_w34115_
	);
	LUT4 #(
		.INIT('h0032)
	) name28289 (
		_w33754_,
		_w33769_,
		_w34113_,
		_w34115_,
		_w34116_
	);
	LUT2 #(
		.INIT('h2)
	) name28290 (
		_w33751_,
		_w33754_,
		_w34117_
	);
	LUT4 #(
		.INIT('h0008)
	) name28291 (
		_w33749_,
		_w33751_,
		_w33752_,
		_w33754_,
		_w34118_
	);
	LUT4 #(
		.INIT('hbfef)
	) name28292 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w34119_
	);
	LUT3 #(
		.INIT('h31)
	) name28293 (
		_w33754_,
		_w34118_,
		_w34119_,
		_w34120_
	);
	LUT4 #(
		.INIT('hd800)
	) name28294 (
		_w33747_,
		_w34112_,
		_w34116_,
		_w34120_,
		_w34121_
	);
	LUT2 #(
		.INIT('h9)
	) name28295 (
		\u0_desIn_r_reg[60]/NET0131 ,
		_w34121_,
		_w34122_
	);
	LUT4 #(
		.INIT('h1f1a)
	) name28296 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34123_
	);
	LUT3 #(
		.INIT('h07)
	) name28297 (
		_w33718_,
		_w33719_,
		_w33722_,
		_w34124_
	);
	LUT2 #(
		.INIT('h4)
	) name28298 (
		_w34123_,
		_w34124_,
		_w34125_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name28299 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34126_
	);
	LUT3 #(
		.INIT('hd0)
	) name28300 (
		_w33718_,
		_w33719_,
		_w33722_,
		_w34127_
	);
	LUT4 #(
		.INIT('hbdf3)
	) name28301 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34128_
	);
	LUT3 #(
		.INIT('h70)
	) name28302 (
		_w34126_,
		_w34127_,
		_w34128_,
		_w34129_
	);
	LUT3 #(
		.INIT('h8a)
	) name28303 (
		_w33727_,
		_w34125_,
		_w34129_,
		_w34130_
	);
	LUT4 #(
		.INIT('hbf00)
	) name28304 (
		_w33718_,
		_w33720_,
		_w33721_,
		_w33722_,
		_w34131_
	);
	LUT3 #(
		.INIT('h59)
	) name28305 (
		_w33719_,
		_w33720_,
		_w33721_,
		_w34132_
	);
	LUT2 #(
		.INIT('h8)
	) name28306 (
		_w34131_,
		_w34132_,
		_w34133_
	);
	LUT4 #(
		.INIT('h0080)
	) name28307 (
		_w33718_,
		_w33719_,
		_w33721_,
		_w33722_,
		_w34134_
	);
	LUT3 #(
		.INIT('h01)
	) name28308 (
		_w33740_,
		_w34099_,
		_w34134_,
		_w34135_
	);
	LUT4 #(
		.INIT('hefd7)
	) name28309 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34136_
	);
	LUT4 #(
		.INIT('h1000)
	) name28310 (
		_w33719_,
		_w33720_,
		_w33721_,
		_w33722_,
		_w34137_
	);
	LUT3 #(
		.INIT('h0e)
	) name28311 (
		_w33722_,
		_w34136_,
		_w34137_,
		_w34138_
	);
	LUT4 #(
		.INIT('hba00)
	) name28312 (
		_w33727_,
		_w34133_,
		_w34135_,
		_w34138_,
		_w34139_
	);
	LUT3 #(
		.INIT('h65)
	) name28313 (
		\u0_desIn_r_reg[16]/NET0131 ,
		_w34130_,
		_w34139_,
		_w34140_
	);
	LUT4 #(
		.INIT('hee79)
	) name28314 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w34141_
	);
	LUT4 #(
		.INIT('h2000)
	) name28315 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w34142_
	);
	LUT4 #(
		.INIT('hd3ce)
	) name28316 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w34143_
	);
	LUT4 #(
		.INIT('h3120)
	) name28317 (
		_w33629_,
		_w34142_,
		_w34143_,
		_w34141_,
		_w34144_
	);
	LUT2 #(
		.INIT('h2)
	) name28318 (
		_w33623_,
		_w34144_,
		_w34145_
	);
	LUT4 #(
		.INIT('h318c)
	) name28319 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w34146_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name28320 (
		_w33625_,
		_w33626_,
		_w33629_,
		_w33624_,
		_w34147_
	);
	LUT3 #(
		.INIT('h32)
	) name28321 (
		_w33991_,
		_w34146_,
		_w34147_,
		_w34148_
	);
	LUT4 #(
		.INIT('hfd75)
	) name28322 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w34149_
	);
	LUT4 #(
		.INIT('h9000)
	) name28323 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w34150_
	);
	LUT3 #(
		.INIT('h0d)
	) name28324 (
		_w33629_,
		_w34149_,
		_w34150_,
		_w34151_
	);
	LUT4 #(
		.INIT('hddd8)
	) name28325 (
		_w33629_,
		_w33634_,
		_w33632_,
		_w33980_,
		_w34152_
	);
	LUT4 #(
		.INIT('h00ba)
	) name28326 (
		_w33623_,
		_w34148_,
		_w34151_,
		_w34152_,
		_w34153_
	);
	LUT3 #(
		.INIT('h65)
	) name28327 (
		\u0_desIn_r_reg[56]/NET0131 ,
		_w34145_,
		_w34153_,
		_w34154_
	);
	LUT4 #(
		.INIT('h5d0a)
	) name28328 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w34155_
	);
	LUT4 #(
		.INIT('h2030)
	) name28329 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w34156_
	);
	LUT4 #(
		.INIT('hbbf5)
	) name28330 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w34157_
	);
	LUT4 #(
		.INIT('h3120)
	) name28331 (
		_w33807_,
		_w34156_,
		_w34157_,
		_w34155_,
		_w34158_
	);
	LUT2 #(
		.INIT('h1)
	) name28332 (
		_w33820_,
		_w34158_,
		_w34159_
	);
	LUT4 #(
		.INIT('hf5bb)
	) name28333 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w34160_
	);
	LUT4 #(
		.INIT('he7ff)
	) name28334 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w34161_
	);
	LUT4 #(
		.INIT('hb100)
	) name28335 (
		_w33807_,
		_w33825_,
		_w34160_,
		_w34161_,
		_w34162_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name28336 (
		_w33809_,
		_w33810_,
		_w33811_,
		_w33808_,
		_w34163_
	);
	LUT3 #(
		.INIT('h10)
	) name28337 (
		_w33807_,
		_w33817_,
		_w34163_,
		_w34164_
	);
	LUT3 #(
		.INIT('h02)
	) name28338 (
		_w33807_,
		_w33813_,
		_w33834_,
		_w34165_
	);
	LUT4 #(
		.INIT('hddd0)
	) name28339 (
		_w33820_,
		_w34162_,
		_w34164_,
		_w34165_,
		_w34166_
	);
	LUT3 #(
		.INIT('h65)
	) name28340 (
		\u0_desIn_r_reg[22]/NET0131 ,
		_w34159_,
		_w34166_,
		_w34167_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name28341 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w34168_
	);
	LUT4 #(
		.INIT('hbf00)
	) name28342 (
		_w33748_,
		_w33751_,
		_w33752_,
		_w33754_,
		_w34169_
	);
	LUT3 #(
		.INIT('h0e)
	) name28343 (
		_w33749_,
		_w33752_,
		_w33754_,
		_w34170_
	);
	LUT4 #(
		.INIT('hffd6)
	) name28344 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w34171_
	);
	LUT4 #(
		.INIT('h1b00)
	) name28345 (
		_w34168_,
		_w34169_,
		_w34170_,
		_w34171_,
		_w34172_
	);
	LUT2 #(
		.INIT('h1)
	) name28346 (
		_w33747_,
		_w34172_,
		_w34173_
	);
	LUT4 #(
		.INIT('h1200)
	) name28347 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33754_,
		_w34174_
	);
	LUT3 #(
		.INIT('h10)
	) name28348 (
		_w33751_,
		_w33752_,
		_w33754_,
		_w34175_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name28349 (
		_w33747_,
		_w33765_,
		_w34174_,
		_w34175_,
		_w34176_
	);
	LUT4 #(
		.INIT('h2e3f)
	) name28350 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w34177_
	);
	LUT2 #(
		.INIT('h2)
	) name28351 (
		_w33775_,
		_w34177_,
		_w34178_
	);
	LUT3 #(
		.INIT('h70)
	) name28352 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w34179_
	);
	LUT2 #(
		.INIT('h8)
	) name28353 (
		_w33773_,
		_w34179_,
		_w34180_
	);
	LUT3 #(
		.INIT('h08)
	) name28354 (
		_w33749_,
		_w33751_,
		_w33752_,
		_w34181_
	);
	LUT4 #(
		.INIT('h0040)
	) name28355 (
		_w33748_,
		_w33751_,
		_w33752_,
		_w33754_,
		_w34182_
	);
	LUT3 #(
		.INIT('h07)
	) name28356 (
		_w33758_,
		_w34181_,
		_w34182_,
		_w34183_
	);
	LUT4 #(
		.INIT('h0100)
	) name28357 (
		_w34176_,
		_w34178_,
		_w34180_,
		_w34183_,
		_w34184_
	);
	LUT3 #(
		.INIT('h9a)
	) name28358 (
		\u0_desIn_r_reg[40]/NET0131 ,
		_w34173_,
		_w34184_,
		_w34185_
	);
	LUT4 #(
		.INIT('h89da)
	) name28359 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w34186_
	);
	LUT2 #(
		.INIT('h1)
	) name28360 (
		_w33629_,
		_w34186_,
		_w34187_
	);
	LUT4 #(
		.INIT('h6080)
	) name28361 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w34188_
	);
	LUT3 #(
		.INIT('h98)
	) name28362 (
		_w33625_,
		_w33626_,
		_w33627_,
		_w34189_
	);
	LUT2 #(
		.INIT('h2)
	) name28363 (
		_w33629_,
		_w33624_,
		_w34190_
	);
	LUT3 #(
		.INIT('h15)
	) name28364 (
		_w34188_,
		_w34189_,
		_w34190_,
		_w34191_
	);
	LUT3 #(
		.INIT('h8a)
	) name28365 (
		_w33623_,
		_w34187_,
		_w34191_,
		_w34192_
	);
	LUT4 #(
		.INIT('h6989)
	) name28366 (
		_w33625_,
		_w33626_,
		_w33624_,
		_w33627_,
		_w34193_
	);
	LUT4 #(
		.INIT('h00c4)
	) name28367 (
		_w33623_,
		_w33629_,
		_w33638_,
		_w34193_,
		_w34194_
	);
	LUT2 #(
		.INIT('h4)
	) name28368 (
		_w33629_,
		_w34188_,
		_w34195_
	);
	LUT4 #(
		.INIT('h5450)
	) name28369 (
		_w33623_,
		_w33643_,
		_w33638_,
		_w34189_,
		_w34196_
	);
	LUT3 #(
		.INIT('h01)
	) name28370 (
		_w34195_,
		_w34196_,
		_w34194_,
		_w34197_
	);
	LUT3 #(
		.INIT('h65)
	) name28371 (
		\u0_desIn_r_reg[54]/NET0131 ,
		_w34192_,
		_w34197_,
		_w34198_
	);
	LUT4 #(
		.INIT('h6002)
	) name28372 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34199_
	);
	LUT4 #(
		.INIT('h4440)
	) name28373 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34200_
	);
	LUT3 #(
		.INIT('h28)
	) name28374 (
		_w33653_,
		_w33654_,
		_w33655_,
		_w34201_
	);
	LUT3 #(
		.INIT('h25)
	) name28375 (
		_w33654_,
		_w33652_,
		_w33655_,
		_w34202_
	);
	LUT4 #(
		.INIT('h0411)
	) name28376 (
		_w33653_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34203_
	);
	LUT4 #(
		.INIT('h1011)
	) name28377 (
		_w33661_,
		_w34203_,
		_w34200_,
		_w34201_,
		_w34204_
	);
	LUT4 #(
		.INIT('h8228)
	) name28378 (
		_w33656_,
		_w33654_,
		_w33652_,
		_w33655_,
		_w34205_
	);
	LUT4 #(
		.INIT('h040c)
	) name28379 (
		_w33662_,
		_w33661_,
		_w34028_,
		_w34202_,
		_w34206_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name28380 (
		_w34199_,
		_w34204_,
		_w34205_,
		_w34206_,
		_w34207_
	);
	LUT3 #(
		.INIT('he0)
	) name28381 (
		_w33656_,
		_w33652_,
		_w33655_,
		_w34208_
	);
	LUT4 #(
		.INIT('h1050)
	) name28382 (
		_w33653_,
		_w33656_,
		_w33654_,
		_w33652_,
		_w34209_
	);
	LUT2 #(
		.INIT('h8)
	) name28383 (
		_w34208_,
		_w34209_,
		_w34210_
	);
	LUT3 #(
		.INIT('h56)
	) name28384 (
		\u0_desIn_r_reg[4]/NET0131 ,
		_w34207_,
		_w34210_,
		_w34211_
	);
	LUT4 #(
		.INIT('h5b4b)
	) name28385 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34212_
	);
	LUT4 #(
		.INIT('h0002)
	) name28386 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34213_
	);
	LUT4 #(
		.INIT('h5504)
	) name28387 (
		_w33727_,
		_w33722_,
		_w34212_,
		_w34213_,
		_w34214_
	);
	LUT4 #(
		.INIT('h00df)
	) name28388 (
		_w33718_,
		_w33720_,
		_w33721_,
		_w33722_,
		_w34215_
	);
	LUT3 #(
		.INIT('h04)
	) name28389 (
		_w33727_,
		_w33718_,
		_w33720_,
		_w34216_
	);
	LUT4 #(
		.INIT('h0040)
	) name28390 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34217_
	);
	LUT4 #(
		.INIT('h1000)
	) name28391 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34218_
	);
	LUT4 #(
		.INIT('heffe)
	) name28392 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33721_,
		_w34219_
	);
	LUT4 #(
		.INIT('h1000)
	) name28393 (
		_w34216_,
		_w34217_,
		_w34215_,
		_w34219_,
		_w34220_
	);
	LUT3 #(
		.INIT('h02)
	) name28394 (
		_w33722_,
		_w33736_,
		_w34091_,
		_w34221_
	);
	LUT2 #(
		.INIT('h1)
	) name28395 (
		_w34220_,
		_w34221_,
		_w34222_
	);
	LUT3 #(
		.INIT('h08)
	) name28396 (
		_w33718_,
		_w33720_,
		_w33721_,
		_w34223_
	);
	LUT4 #(
		.INIT('h0020)
	) name28397 (
		_w33719_,
		_w33720_,
		_w33721_,
		_w33722_,
		_w34224_
	);
	LUT3 #(
		.INIT('h01)
	) name28398 (
		_w34088_,
		_w34223_,
		_w34224_,
		_w34225_
	);
	LUT4 #(
		.INIT('h0100)
	) name28399 (
		_w33718_,
		_w33719_,
		_w33720_,
		_w33722_,
		_w34226_
	);
	LUT2 #(
		.INIT('h1)
	) name28400 (
		_w34218_,
		_w34226_,
		_w34227_
	);
	LUT3 #(
		.INIT('h2a)
	) name28401 (
		_w33727_,
		_w34225_,
		_w34227_,
		_w34228_
	);
	LUT4 #(
		.INIT('h5556)
	) name28402 (
		\u0_desIn_r_reg[52]/NET0131 ,
		_w34214_,
		_w34222_,
		_w34228_,
		_w34229_
	);
	LUT3 #(
		.INIT('he4)
	) name28403 (
		decrypt_pad,
		\key1[51]_pad ,
		\key3[51]_pad ,
		_w34230_
	);
	LUT3 #(
		.INIT('hd8)
	) name28404 (
		decrypt_pad,
		\key1[33]_pad ,
		\key3[33]_pad ,
		_w34231_
	);
	LUT3 #(
		.INIT('hd8)
	) name28405 (
		decrypt_pad,
		\key1[35]_pad ,
		\key3[35]_pad ,
		_w34232_
	);
	LUT3 #(
		.INIT('hd8)
	) name28406 (
		decrypt_pad,
		\key1[45]_pad ,
		\key3[45]_pad ,
		_w34233_
	);
	LUT3 #(
		.INIT('hd8)
	) name28407 (
		decrypt_pad,
		\key1[7]_pad ,
		\key3[7]_pad ,
		_w34234_
	);
	LUT3 #(
		.INIT('hd8)
	) name28408 (
		decrypt_pad,
		\key1[38]_pad ,
		\key3[38]_pad ,
		_w34235_
	);
	LUT3 #(
		.INIT('he4)
	) name28409 (
		decrypt_pad,
		\key1[23]_pad ,
		\key3[23]_pad ,
		_w34236_
	);
	LUT3 #(
		.INIT('hd8)
	) name28410 (
		decrypt_pad,
		\key1[11]_pad ,
		\key3[11]_pad ,
		_w34237_
	);
	LUT3 #(
		.INIT('hd8)
	) name28411 (
		decrypt_pad,
		\key1[27]_pad ,
		\key3[27]_pad ,
		_w34238_
	);
	LUT3 #(
		.INIT('hd8)
	) name28412 (
		decrypt_pad,
		\key1[32]_pad ,
		\key3[32]_pad ,
		_w34239_
	);
	LUT3 #(
		.INIT('he4)
	) name28413 (
		decrypt_pad,
		\key1[10]_pad ,
		\key3[10]_pad ,
		_w34240_
	);
	LUT3 #(
		.INIT('he4)
	) name28414 (
		decrypt_pad,
		\key1[19]_pad ,
		\key3[19]_pad ,
		_w34241_
	);
	LUT3 #(
		.INIT('he4)
	) name28415 (
		decrypt_pad,
		\key1[14]_pad ,
		\key3[14]_pad ,
		_w34242_
	);
	LUT3 #(
		.INIT('he4)
	) name28416 (
		decrypt_pad,
		\key1[12]_pad ,
		\key3[12]_pad ,
		_w34243_
	);
	LUT3 #(
		.INIT('he4)
	) name28417 (
		decrypt_pad,
		\key1[30]_pad ,
		\key3[30]_pad ,
		_w34244_
	);
	LUT3 #(
		.INIT('he4)
	) name28418 (
		decrypt_pad,
		\key1[17]_pad ,
		\key3[17]_pad ,
		_w34245_
	);
	LUT3 #(
		.INIT('he4)
	) name28419 (
		decrypt_pad,
		\key1[2]_pad ,
		\key3[2]_pad ,
		_w34246_
	);
	LUT3 #(
		.INIT('hd8)
	) name28420 (
		decrypt_pad,
		\key1[10]_pad ,
		\key3[10]_pad ,
		_w34247_
	);
	LUT3 #(
		.INIT('he4)
	) name28421 (
		decrypt_pad,
		\key1[3]_pad ,
		\key3[3]_pad ,
		_w34248_
	);
	LUT3 #(
		.INIT('hd8)
	) name28422 (
		decrypt_pad,
		\key1[37]_pad ,
		\key3[37]_pad ,
		_w34249_
	);
	LUT3 #(
		.INIT('hd8)
	) name28423 (
		decrypt_pad,
		\key1[40]_pad ,
		\key3[40]_pad ,
		_w34250_
	);
	LUT3 #(
		.INIT('he4)
	) name28424 (
		decrypt_pad,
		\key1[33]_pad ,
		\key3[33]_pad ,
		_w34251_
	);
	LUT3 #(
		.INIT('hd8)
	) name28425 (
		decrypt_pad,
		\key1[6]_pad ,
		\key3[6]_pad ,
		_w34252_
	);
	LUT3 #(
		.INIT('hd8)
	) name28426 (
		decrypt_pad,
		\key1[53]_pad ,
		\key3[53]_pad ,
		_w34253_
	);
	LUT3 #(
		.INIT('he4)
	) name28427 (
		decrypt_pad,
		\key1[24]_pad ,
		\key3[24]_pad ,
		_w34254_
	);
	LUT3 #(
		.INIT('hd8)
	) name28428 (
		decrypt_pad,
		\key1[34]_pad ,
		\key3[34]_pad ,
		_w34255_
	);
	LUT3 #(
		.INIT('he4)
	) name28429 (
		decrypt_pad,
		\key1[49]_pad ,
		\key3[49]_pad ,
		_w34256_
	);
	LUT3 #(
		.INIT('hd8)
	) name28430 (
		decrypt_pad,
		\key1[14]_pad ,
		\key3[14]_pad ,
		_w34257_
	);
	LUT3 #(
		.INIT('hd8)
	) name28431 (
		decrypt_pad,
		\key1[29]_pad ,
		\key3[29]_pad ,
		_w34258_
	);
	LUT3 #(
		.INIT('hd8)
	) name28432 (
		decrypt_pad,
		\key1[21]_pad ,
		\key3[21]_pad ,
		_w34259_
	);
	LUT3 #(
		.INIT('he4)
	) name28433 (
		decrypt_pad,
		\key1[4]_pad ,
		\key3[4]_pad ,
		_w34260_
	);
	LUT3 #(
		.INIT('he4)
	) name28434 (
		decrypt_pad,
		\key1[37]_pad ,
		\key3[37]_pad ,
		_w34261_
	);
	LUT3 #(
		.INIT('he4)
	) name28435 (
		decrypt_pad,
		\key1[53]_pad ,
		\key3[53]_pad ,
		_w34262_
	);
	LUT3 #(
		.INIT('he4)
	) name28436 (
		decrypt_pad,
		\key1[31]_pad ,
		\key3[31]_pad ,
		_w34263_
	);
	LUT3 #(
		.INIT('hd8)
	) name28437 (
		decrypt_pad,
		\key1[42]_pad ,
		\key3[42]_pad ,
		_w34264_
	);
	LUT3 #(
		.INIT('he4)
	) name28438 (
		decrypt_pad,
		\key1[43]_pad ,
		\key3[43]_pad ,
		_w34265_
	);
	LUT3 #(
		.INIT('hd8)
	) name28439 (
		decrypt_pad,
		\key1[55]_pad ,
		\key3[55]_pad ,
		_w34266_
	);
	LUT3 #(
		.INIT('he4)
	) name28440 (
		decrypt_pad,
		\key1[20]_pad ,
		\key3[20]_pad ,
		_w34267_
	);
	LUT3 #(
		.INIT('he4)
	) name28441 (
		decrypt_pad,
		\key1[36]_pad ,
		\key3[36]_pad ,
		_w34268_
	);
	LUT3 #(
		.INIT('hd8)
	) name28442 (
		decrypt_pad,
		\key1[22]_pad ,
		\key3[22]_pad ,
		_w34269_
	);
	LUT3 #(
		.INIT('he4)
	) name28443 (
		decrypt_pad,
		\key1[55]_pad ,
		\key3[55]_pad ,
		_w34270_
	);
	LUT3 #(
		.INIT('he4)
	) name28444 (
		decrypt_pad,
		\key1[15]_pad ,
		\key3[15]_pad ,
		_w34271_
	);
	LUT3 #(
		.INIT('he4)
	) name28445 (
		decrypt_pad,
		\key1[40]_pad ,
		\key3[40]_pad ,
		_w34272_
	);
	LUT3 #(
		.INIT('he4)
	) name28446 (
		decrypt_pad,
		\key1[8]_pad ,
		\key3[8]_pad ,
		_w34273_
	);
	LUT3 #(
		.INIT('hd8)
	) name28447 (
		decrypt_pad,
		\key1[16]_pad ,
		\key3[16]_pad ,
		_w34274_
	);
	LUT3 #(
		.INIT('he4)
	) name28448 (
		decrypt_pad,
		\key1[22]_pad ,
		\key3[22]_pad ,
		_w34275_
	);
	LUT3 #(
		.INIT('he4)
	) name28449 (
		decrypt_pad,
		\key1[27]_pad ,
		\key3[27]_pad ,
		_w34276_
	);
	LUT3 #(
		.INIT('hd8)
	) name28450 (
		decrypt_pad,
		\key1[31]_pad ,
		\key3[31]_pad ,
		_w34277_
	);
	LUT3 #(
		.INIT('hd8)
	) name28451 (
		decrypt_pad,
		\key1[46]_pad ,
		\key3[46]_pad ,
		_w34278_
	);
	LUT3 #(
		.INIT('he4)
	) name28452 (
		decrypt_pad,
		\key1[26]_pad ,
		\key3[26]_pad ,
		_w34279_
	);
	LUT3 #(
		.INIT('hd8)
	) name28453 (
		decrypt_pad,
		\key1[24]_pad ,
		\key3[24]_pad ,
		_w34280_
	);
	LUT3 #(
		.INIT('he4)
	) name28454 (
		decrypt_pad,
		\key1[35]_pad ,
		\key3[35]_pad ,
		_w34281_
	);
	LUT3 #(
		.INIT('he4)
	) name28455 (
		decrypt_pad,
		\key1[28]_pad ,
		\key3[28]_pad ,
		_w34282_
	);
	LUT3 #(
		.INIT('he4)
	) name28456 (
		decrypt_pad,
		\key1[48]_pad ,
		\key3[48]_pad ,
		_w34283_
	);
	LUT3 #(
		.INIT('hd8)
	) name28457 (
		decrypt_pad,
		\key1[15]_pad ,
		\key3[15]_pad ,
		_w34284_
	);
	LUT3 #(
		.INIT('he4)
	) name28458 (
		decrypt_pad,
		\key1[38]_pad ,
		\key3[38]_pad ,
		_w34285_
	);
	LUT3 #(
		.INIT('he4)
	) name28459 (
		decrypt_pad,
		\key1[45]_pad ,
		\key3[45]_pad ,
		_w34286_
	);
	LUT3 #(
		.INIT('hd8)
	) name28460 (
		decrypt_pad,
		\key1[50]_pad ,
		\key3[50]_pad ,
		_w34287_
	);
	LUT3 #(
		.INIT('hd8)
	) name28461 (
		decrypt_pad,
		\key1[26]_pad ,
		\key3[26]_pad ,
		_w34288_
	);
	LUT3 #(
		.INIT('he4)
	) name28462 (
		decrypt_pad,
		\key1[9]_pad ,
		\key3[9]_pad ,
		_w34289_
	);
	LUT3 #(
		.INIT('hd8)
	) name28463 (
		decrypt_pad,
		\key1[39]_pad ,
		\key3[39]_pad ,
		_w34290_
	);
	LUT3 #(
		.INIT('he4)
	) name28464 (
		decrypt_pad,
		\key1[54]_pad ,
		\key3[54]_pad ,
		_w34291_
	);
	LUT3 #(
		.INIT('he4)
	) name28465 (
		decrypt_pad,
		\key1[25]_pad ,
		\key3[25]_pad ,
		_w34292_
	);
	LUT3 #(
		.INIT('hd8)
	) name28466 (
		decrypt_pad,
		\key1[8]_pad ,
		\key3[8]_pad ,
		_w34293_
	);
	LUT3 #(
		.INIT('hd8)
	) name28467 (
		decrypt_pad,
		\key1[0]_pad ,
		\key3[0]_pad ,
		_w34294_
	);
	LUT3 #(
		.INIT('hd8)
	) name28468 (
		decrypt_pad,
		\key1[20]_pad ,
		\key3[20]_pad ,
		_w34295_
	);
	LUT3 #(
		.INIT('he4)
	) name28469 (
		decrypt_pad,
		\key1[46]_pad ,
		\key3[46]_pad ,
		_w34296_
	);
	LUT3 #(
		.INIT('hd8)
	) name28470 (
		decrypt_pad,
		\key1[25]_pad ,
		\key3[25]_pad ,
		_w34297_
	);
	LUT3 #(
		.INIT('hd8)
	) name28471 (
		decrypt_pad,
		\key1[44]_pad ,
		\key3[44]_pad ,
		_w34298_
	);
	LUT3 #(
		.INIT('hd8)
	) name28472 (
		decrypt_pad,
		\key1[51]_pad ,
		\key3[51]_pad ,
		_w34299_
	);
	LUT3 #(
		.INIT('he4)
	) name28473 (
		decrypt_pad,
		\key1[50]_pad ,
		\key3[50]_pad ,
		_w34300_
	);
	LUT3 #(
		.INIT('he4)
	) name28474 (
		decrypt_pad,
		\key1[32]_pad ,
		\key3[32]_pad ,
		_w34301_
	);
	LUT3 #(
		.INIT('hd8)
	) name28475 (
		decrypt_pad,
		\key1[43]_pad ,
		\key3[43]_pad ,
		_w34302_
	);
	LUT3 #(
		.INIT('hd8)
	) name28476 (
		decrypt_pad,
		\key1[3]_pad ,
		\key3[3]_pad ,
		_w34303_
	);
	LUT3 #(
		.INIT('he4)
	) name28477 (
		decrypt_pad,
		\key1[7]_pad ,
		\key3[7]_pad ,
		_w34304_
	);
	LUT3 #(
		.INIT('he4)
	) name28478 (
		decrypt_pad,
		\key1[44]_pad ,
		\key3[44]_pad ,
		_w34305_
	);
	LUT3 #(
		.INIT('hd8)
	) name28479 (
		decrypt_pad,
		\key1[54]_pad ,
		\key3[54]_pad ,
		_w34306_
	);
	LUT3 #(
		.INIT('hd8)
	) name28480 (
		decrypt_pad,
		\key1[30]_pad ,
		\key3[30]_pad ,
		_w34307_
	);
	LUT3 #(
		.INIT('he4)
	) name28481 (
		decrypt_pad,
		\key1[1]_pad ,
		\key3[1]_pad ,
		_w34308_
	);
	LUT3 #(
		.INIT('hd8)
	) name28482 (
		decrypt_pad,
		\key1[18]_pad ,
		\key3[18]_pad ,
		_w34309_
	);
	LUT3 #(
		.INIT('hd8)
	) name28483 (
		decrypt_pad,
		\key1[28]_pad ,
		\key3[28]_pad ,
		_w34310_
	);
	LUT3 #(
		.INIT('he4)
	) name28484 (
		decrypt_pad,
		\key1[39]_pad ,
		\key3[39]_pad ,
		_w34311_
	);
	LUT3 #(
		.INIT('hd8)
	) name28485 (
		decrypt_pad,
		\key1[17]_pad ,
		\key3[17]_pad ,
		_w34312_
	);
	LUT3 #(
		.INIT('hd8)
	) name28486 (
		decrypt_pad,
		\key1[1]_pad ,
		\key3[1]_pad ,
		_w34313_
	);
	LUT3 #(
		.INIT('he4)
	) name28487 (
		decrypt_pad,
		\key1[13]_pad ,
		\key3[13]_pad ,
		_w34314_
	);
	LUT3 #(
		.INIT('hd8)
	) name28488 (
		decrypt_pad,
		\key1[19]_pad ,
		\key3[19]_pad ,
		_w34315_
	);
	LUT3 #(
		.INIT('he4)
	) name28489 (
		decrypt_pad,
		\key1[6]_pad ,
		\key3[6]_pad ,
		_w34316_
	);
	LUT3 #(
		.INIT('hd8)
	) name28490 (
		decrypt_pad,
		\key1[47]_pad ,
		\key3[47]_pad ,
		_w34317_
	);
	LUT3 #(
		.INIT('hd8)
	) name28491 (
		decrypt_pad,
		\key1[23]_pad ,
		\key3[23]_pad ,
		_w34318_
	);
	LUT3 #(
		.INIT('hd8)
	) name28492 (
		decrypt_pad,
		\key1[12]_pad ,
		\key3[12]_pad ,
		_w34319_
	);
	LUT3 #(
		.INIT('he4)
	) name28493 (
		decrypt_pad,
		\key1[52]_pad ,
		\key3[52]_pad ,
		_w34320_
	);
	LUT3 #(
		.INIT('hd8)
	) name28494 (
		decrypt_pad,
		\key1[5]_pad ,
		\key3[5]_pad ,
		_w34321_
	);
	LUT3 #(
		.INIT('hd8)
	) name28495 (
		decrypt_pad,
		\key1[9]_pad ,
		\key3[9]_pad ,
		_w34322_
	);
	LUT3 #(
		.INIT('he4)
	) name28496 (
		decrypt_pad,
		\key1[0]_pad ,
		\key3[0]_pad ,
		_w34323_
	);
	LUT3 #(
		.INIT('hd8)
	) name28497 (
		decrypt_pad,
		\key1[4]_pad ,
		\key3[4]_pad ,
		_w34324_
	);
	LUT3 #(
		.INIT('he4)
	) name28498 (
		decrypt_pad,
		\key1[11]_pad ,
		\key3[11]_pad ,
		_w34325_
	);
	LUT3 #(
		.INIT('hd8)
	) name28499 (
		decrypt_pad,
		\key1[52]_pad ,
		\key3[52]_pad ,
		_w34326_
	);
	LUT3 #(
		.INIT('he4)
	) name28500 (
		decrypt_pad,
		\key1[18]_pad ,
		\key3[18]_pad ,
		_w34327_
	);
	LUT3 #(
		.INIT('hd8)
	) name28501 (
		decrypt_pad,
		\key1[36]_pad ,
		\key3[36]_pad ,
		_w34328_
	);
	LUT3 #(
		.INIT('he4)
	) name28502 (
		decrypt_pad,
		\key1[5]_pad ,
		\key3[5]_pad ,
		_w34329_
	);
	LUT3 #(
		.INIT('he4)
	) name28503 (
		decrypt_pad,
		\key1[42]_pad ,
		\key3[42]_pad ,
		_w34330_
	);
	LUT3 #(
		.INIT('hd8)
	) name28504 (
		decrypt_pad,
		\key1[2]_pad ,
		\key3[2]_pad ,
		_w34331_
	);
	LUT3 #(
		.INIT('hd8)
	) name28505 (
		decrypt_pad,
		\key1[48]_pad ,
		\key3[48]_pad ,
		_w34332_
	);
	LUT3 #(
		.INIT('he4)
	) name28506 (
		decrypt_pad,
		\key1[34]_pad ,
		\key3[34]_pad ,
		_w34333_
	);
	LUT3 #(
		.INIT('he4)
	) name28507 (
		decrypt_pad,
		\key1[21]_pad ,
		\key3[21]_pad ,
		_w34334_
	);
	LUT3 #(
		.INIT('hd8)
	) name28508 (
		decrypt_pad,
		\key1[49]_pad ,
		\key3[49]_pad ,
		_w34335_
	);
	LUT3 #(
		.INIT('he4)
	) name28509 (
		decrypt_pad,
		\key1[47]_pad ,
		\key3[47]_pad ,
		_w34336_
	);
	LUT3 #(
		.INIT('he4)
	) name28510 (
		decrypt_pad,
		\key1[29]_pad ,
		\key3[29]_pad ,
		_w34337_
	);
	LUT3 #(
		.INIT('hd8)
	) name28511 (
		decrypt_pad,
		\key1[13]_pad ,
		\key3[13]_pad ,
		_w34338_
	);
	LUT3 #(
		.INIT('hd8)
	) name28512 (
		decrypt_pad,
		\key1[41]_pad ,
		\key3[41]_pad ,
		_w34339_
	);
	LUT3 #(
		.INIT('he4)
	) name28513 (
		decrypt_pad,
		\key1[41]_pad ,
		\key3[41]_pad ,
		_w34340_
	);
	LUT3 #(
		.INIT('he4)
	) name28514 (
		decrypt_pad,
		\key1[16]_pad ,
		\key3[16]_pad ,
		_w34341_
	);
	LUT4 #(
		.INIT('h1000)
	) name28515 (
		_w23070_,
		_w23071_,
		_w23072_,
		_w23069_,
		_w34342_
	);
	LUT4 #(
		.INIT('h002a)
	) name28516 (
		_w23068_,
		_w23073_,
		_w23088_,
		_w23094_,
		_w34343_
	);
	LUT4 #(
		.INIT('h0014)
	) name28517 (
		_w23073_,
		_w23070_,
		_w23071_,
		_w23069_,
		_w34344_
	);
	LUT2 #(
		.INIT('h1)
	) name28518 (
		_w23179_,
		_w34344_,
		_w34345_
	);
	LUT3 #(
		.INIT('h40)
	) name28519 (
		_w34342_,
		_w34343_,
		_w34345_,
		_w34346_
	);
	LUT3 #(
		.INIT('h0b)
	) name28520 (
		_w23070_,
		_w23072_,
		_w23069_,
		_w34347_
	);
	LUT4 #(
		.INIT('h7e00)
	) name28521 (
		_w23070_,
		_w23071_,
		_w23072_,
		_w23069_,
		_w34348_
	);
	LUT3 #(
		.INIT('h0b)
	) name28522 (
		_w23170_,
		_w34347_,
		_w34348_,
		_w34349_
	);
	LUT4 #(
		.INIT('h0001)
	) name28523 (
		_w23068_,
		_w23084_,
		_w23096_,
		_w23074_,
		_w34350_
	);
	LUT2 #(
		.INIT('h4)
	) name28524 (
		_w34349_,
		_w34350_,
		_w34351_
	);
	LUT2 #(
		.INIT('h4)
	) name28525 (
		_w23070_,
		_w23069_,
		_w34352_
	);
	LUT2 #(
		.INIT('h4)
	) name28526 (
		_w23203_,
		_w34352_,
		_w34353_
	);
	LUT4 #(
		.INIT('h8caf)
	) name28527 (
		_w23073_,
		_w23069_,
		_w23094_,
		_w23207_,
		_w34354_
	);
	LUT2 #(
		.INIT('h4)
	) name28528 (
		_w34353_,
		_w34354_,
		_w34355_
	);
	LUT4 #(
		.INIT('ha955)
	) name28529 (
		\u1_L1_reg[20]/NET0131 ,
		_w34346_,
		_w34351_,
		_w34355_,
		_w34356_
	);
	LUT4 #(
		.INIT('hf04f)
	) name28530 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w34357_
	);
	LUT3 #(
		.INIT('hbc)
	) name28531 (
		_w27420_,
		_w27417_,
		_w27418_,
		_w34358_
	);
	LUT4 #(
		.INIT('hb7fd)
	) name28532 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w34359_
	);
	LUT4 #(
		.INIT('hd800)
	) name28533 (
		_w27416_,
		_w34357_,
		_w34358_,
		_w34359_,
		_w34360_
	);
	LUT4 #(
		.INIT('h9fff)
	) name28534 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w34361_
	);
	LUT2 #(
		.INIT('h1)
	) name28535 (
		_w27416_,
		_w34361_,
		_w34362_
	);
	LUT4 #(
		.INIT('h8228)
	) name28536 (
		_w27419_,
		_w27420_,
		_w27417_,
		_w27418_,
		_w34363_
	);
	LUT4 #(
		.INIT('h0031)
	) name28537 (
		_w27424_,
		_w27755_,
		_w34358_,
		_w34363_,
		_w34364_
	);
	LUT4 #(
		.INIT('h0e04)
	) name28538 (
		_w27415_,
		_w34360_,
		_w34362_,
		_w34364_,
		_w34365_
	);
	LUT2 #(
		.INIT('h9)
	) name28539 (
		\u0_L9_reg[9]/NET0131 ,
		_w34365_,
		_w34366_
	);
	LUT4 #(
		.INIT('hefe7)
	) name28540 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w34367_
	);
	LUT4 #(
		.INIT('hbbdb)
	) name28541 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w34368_
	);
	LUT4 #(
		.INIT('hc840)
	) name28542 (
		_w33141_,
		_w33309_,
		_w34368_,
		_w34367_,
		_w34369_
	);
	LUT2 #(
		.INIT('h2)
	) name28543 (
		_w33154_,
		_w34369_,
		_w34370_
	);
	LUT4 #(
		.INIT('hff0d)
	) name28544 (
		_w33142_,
		_w33141_,
		_w33145_,
		_w33143_,
		_w34371_
	);
	LUT2 #(
		.INIT('h2)
	) name28545 (
		_w33144_,
		_w34371_,
		_w34372_
	);
	LUT4 #(
		.INIT('h0020)
	) name28546 (
		_w33142_,
		_w33144_,
		_w33141_,
		_w33143_,
		_w34373_
	);
	LUT2 #(
		.INIT('h1)
	) name28547 (
		_w33158_,
		_w34373_,
		_w34374_
	);
	LUT3 #(
		.INIT('h15)
	) name28548 (
		_w33144_,
		_w33141_,
		_w33143_,
		_w34375_
	);
	LUT3 #(
		.INIT('h08)
	) name28549 (
		_w33144_,
		_w33141_,
		_w33145_,
		_w34376_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name28550 (
		_w33171_,
		_w33444_,
		_w34375_,
		_w34376_,
		_w34377_
	);
	LUT4 #(
		.INIT('h4555)
	) name28551 (
		_w33154_,
		_w34372_,
		_w34374_,
		_w34377_,
		_w34378_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name28552 (
		_w33142_,
		_w33144_,
		_w33145_,
		_w33143_,
		_w34379_
	);
	LUT2 #(
		.INIT('h1)
	) name28553 (
		_w33141_,
		_w34379_,
		_w34380_
	);
	LUT3 #(
		.INIT('h0b)
	) name28554 (
		_w33143_,
		_w33150_,
		_w33166_,
		_w34381_
	);
	LUT2 #(
		.INIT('h4)
	) name28555 (
		_w34380_,
		_w34381_,
		_w34382_
	);
	LUT4 #(
		.INIT('h5655)
	) name28556 (
		\u0_L0_reg[10]/NET0131 ,
		_w34378_,
		_w34370_,
		_w34382_,
		_w34383_
	);
	LUT4 #(
		.INIT('h4044)
	) name28557 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w34384_
	);
	LUT3 #(
		.INIT('h01)
	) name28558 (
		_w19283_,
		_w19306_,
		_w34384_,
		_w34385_
	);
	LUT3 #(
		.INIT('h02)
	) name28559 (
		_w19283_,
		_w19295_,
		_w19288_,
		_w34386_
	);
	LUT4 #(
		.INIT('h888a)
	) name28560 (
		_w19289_,
		_w19513_,
		_w34385_,
		_w34386_,
		_w34387_
	);
	LUT4 #(
		.INIT('h0008)
	) name28561 (
		_w19283_,
		_w19287_,
		_w19281_,
		_w19284_,
		_w34388_
	);
	LUT2 #(
		.INIT('h1)
	) name28562 (
		_w19301_,
		_w34388_,
		_w34389_
	);
	LUT3 #(
		.INIT('h0b)
	) name28563 (
		_w19283_,
		_w19287_,
		_w19282_,
		_w34390_
	);
	LUT3 #(
		.INIT('hf2)
	) name28564 (
		_w19287_,
		_w19284_,
		_w19282_,
		_w34391_
	);
	LUT4 #(
		.INIT('hf351)
	) name28565 (
		_w19307_,
		_w19581_,
		_w34390_,
		_w34391_,
		_w34392_
	);
	LUT4 #(
		.INIT('h1333)
	) name28566 (
		_w19296_,
		_w19289_,
		_w34389_,
		_w34392_,
		_w34393_
	);
	LUT4 #(
		.INIT('h7fde)
	) name28567 (
		_w19287_,
		_w19281_,
		_w19284_,
		_w19282_,
		_w34394_
	);
	LUT2 #(
		.INIT('h1)
	) name28568 (
		_w19283_,
		_w34394_,
		_w34395_
	);
	LUT3 #(
		.INIT('h0b)
	) name28569 (
		_w19284_,
		_w19308_,
		_w19286_,
		_w34396_
	);
	LUT2 #(
		.INIT('h4)
	) name28570 (
		_w34395_,
		_w34396_,
		_w34397_
	);
	LUT4 #(
		.INIT('h5655)
	) name28571 (
		\u1_L7_reg[10]/NET0131 ,
		_w34387_,
		_w34393_,
		_w34397_,
		_w34398_
	);
	LUT3 #(
		.INIT('h02)
	) name28572 (
		_w29976_,
		_w29980_,
		_w29992_,
		_w34399_
	);
	LUT4 #(
		.INIT('h4014)
	) name28573 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w34400_
	);
	LUT4 #(
		.INIT('hfdcc)
	) name28574 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w34401_
	);
	LUT4 #(
		.INIT('h0504)
	) name28575 (
		_w29976_,
		_w29984_,
		_w34400_,
		_w34401_,
		_w34402_
	);
	LUT2 #(
		.INIT('h1)
	) name28576 (
		_w34399_,
		_w34402_,
		_w34403_
	);
	LUT3 #(
		.INIT('h80)
	) name28577 (
		_w29971_,
		_w29973_,
		_w29974_,
		_w34404_
	);
	LUT4 #(
		.INIT('h0100)
	) name28578 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w34405_
	);
	LUT4 #(
		.INIT('h3332)
	) name28579 (
		_w29976_,
		_w29987_,
		_w34405_,
		_w34404_,
		_w34406_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name28580 (
		_w29976_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w34407_
	);
	LUT4 #(
		.INIT('h0084)
	) name28581 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29974_,
		_w34408_
	);
	LUT4 #(
		.INIT('h0c04)
	) name28582 (
		_w29971_,
		_w29984_,
		_w34408_,
		_w34407_,
		_w34409_
	);
	LUT2 #(
		.INIT('h4)
	) name28583 (
		_w29977_,
		_w29995_,
		_w34410_
	);
	LUT4 #(
		.INIT('h00ef)
	) name28584 (
		_w29971_,
		_w29972_,
		_w29973_,
		_w29984_,
		_w34411_
	);
	LUT3 #(
		.INIT('h10)
	) name28585 (
		_w29979_,
		_w29980_,
		_w34411_,
		_w34412_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name28586 (
		_w34406_,
		_w34409_,
		_w34410_,
		_w34412_,
		_w34413_
	);
	LUT3 #(
		.INIT('h56)
	) name28587 (
		\u0_L5_reg[26]/NET0131 ,
		_w34403_,
		_w34413_,
		_w34414_
	);
	LUT4 #(
		.INIT('h001d)
	) name28588 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w34415_
	);
	LUT4 #(
		.INIT('h6e00)
	) name28589 (
		_w31319_,
		_w31320_,
		_w31321_,
		_w31318_,
		_w34416_
	);
	LUT4 #(
		.INIT('h00fd)
	) name28590 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31318_,
		_w34417_
	);
	LUT4 #(
		.INIT('h8acf)
	) name28591 (
		_w31339_,
		_w34415_,
		_w34416_,
		_w34417_,
		_w34418_
	);
	LUT4 #(
		.INIT('hdd7f)
	) name28592 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w34419_
	);
	LUT3 #(
		.INIT('h8a)
	) name28593 (
		_w31317_,
		_w34418_,
		_w34419_,
		_w34420_
	);
	LUT4 #(
		.INIT('h7707)
	) name28594 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w34421_
	);
	LUT3 #(
		.INIT('h07)
	) name28595 (
		_w31319_,
		_w31320_,
		_w31318_,
		_w34422_
	);
	LUT2 #(
		.INIT('h4)
	) name28596 (
		_w34421_,
		_w34422_,
		_w34423_
	);
	LUT4 #(
		.INIT('h0200)
	) name28597 (
		_w31319_,
		_w31322_,
		_w31321_,
		_w31318_,
		_w34424_
	);
	LUT4 #(
		.INIT('h0001)
	) name28598 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31318_,
		_w34425_
	);
	LUT4 #(
		.INIT('h0800)
	) name28599 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w34426_
	);
	LUT3 #(
		.INIT('h01)
	) name28600 (
		_w34425_,
		_w34426_,
		_w34424_,
		_w34427_
	);
	LUT4 #(
		.INIT('hfe7b)
	) name28601 (
		_w31319_,
		_w31322_,
		_w31320_,
		_w31321_,
		_w34428_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name28602 (
		_w31319_,
		_w31322_,
		_w31321_,
		_w31318_,
		_w34429_
	);
	LUT4 #(
		.INIT('hf351)
	) name28603 (
		_w31320_,
		_w31318_,
		_w34428_,
		_w34429_,
		_w34430_
	);
	LUT4 #(
		.INIT('hba00)
	) name28604 (
		_w31317_,
		_w34423_,
		_w34427_,
		_w34430_,
		_w34431_
	);
	LUT3 #(
		.INIT('h65)
	) name28605 (
		\u0_L3_reg[25]/NET0131 ,
		_w34420_,
		_w34431_,
		_w34432_
	);
	LUT2 #(
		.INIT('h4)
	) name28606 (
		_w33750_,
		_w34175_,
		_w34433_
	);
	LUT3 #(
		.INIT('h0e)
	) name28607 (
		_w33751_,
		_w33752_,
		_w33754_,
		_w34434_
	);
	LUT3 #(
		.INIT('hc4)
	) name28608 (
		_w33749_,
		_w33751_,
		_w33752_,
		_w34435_
	);
	LUT4 #(
		.INIT('h23af)
	) name28609 (
		_w33755_,
		_w34114_,
		_w34434_,
		_w34435_,
		_w34436_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name28610 (
		_w33747_,
		_w33762_,
		_w34433_,
		_w34436_,
		_w34437_
	);
	LUT4 #(
		.INIT('hec2d)
	) name28611 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w34438_
	);
	LUT4 #(
		.INIT('h0040)
	) name28612 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w34439_
	);
	LUT4 #(
		.INIT('h5504)
	) name28613 (
		_w33747_,
		_w33754_,
		_w34438_,
		_w34439_,
		_w34440_
	);
	LUT4 #(
		.INIT('h9bd6)
	) name28614 (
		_w33748_,
		_w33749_,
		_w33751_,
		_w33752_,
		_w34441_
	);
	LUT2 #(
		.INIT('h1)
	) name28615 (
		_w33747_,
		_w33754_,
		_w34442_
	);
	LUT2 #(
		.INIT('h4)
	) name28616 (
		_w34441_,
		_w34442_,
		_w34443_
	);
	LUT3 #(
		.INIT('h20)
	) name28617 (
		_w33748_,
		_w33749_,
		_w33754_,
		_w34444_
	);
	LUT2 #(
		.INIT('h8)
	) name28618 (
		_w33760_,
		_w34444_,
		_w34445_
	);
	LUT4 #(
		.INIT('h153f)
	) name28619 (
		_w33765_,
		_w34117_,
		_w34109_,
		_w34175_,
		_w34446_
	);
	LUT4 #(
		.INIT('h0100)
	) name28620 (
		_w34440_,
		_w34445_,
		_w34443_,
		_w34446_,
		_w34447_
	);
	LUT3 #(
		.INIT('h65)
	) name28621 (
		\u0_desIn_r_reg[58]/NET0131 ,
		_w34437_,
		_w34447_,
		_w34448_
	);
	LUT4 #(
		.INIT('h1020)
	) name28622 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w34449_
	);
	LUT3 #(
		.INIT('h08)
	) name28623 (
		_w16226_,
		_w16223_,
		_w34449_,
		_w34450_
	);
	LUT4 #(
		.INIT('h2000)
	) name28624 (
		_w16216_,
		_w16217_,
		_w16220_,
		_w16235_,
		_w34451_
	);
	LUT3 #(
		.INIT('h01)
	) name28625 (
		_w16226_,
		_w16512_,
		_w34451_,
		_w34452_
	);
	LUT2 #(
		.INIT('h1)
	) name28626 (
		_w34450_,
		_w34452_,
		_w34453_
	);
	LUT4 #(
		.INIT('hef00)
	) name28627 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16226_,
		_w34454_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name28628 (
		_w16224_,
		_w16227_,
		_w16277_,
		_w34454_,
		_w34455_
	);
	LUT4 #(
		.INIT('h00ef)
	) name28629 (
		_w16216_,
		_w16219_,
		_w16220_,
		_w16226_,
		_w34456_
	);
	LUT3 #(
		.INIT('h23)
	) name28630 (
		_w16277_,
		_w34456_,
		_w34454_,
		_w34457_
	);
	LUT3 #(
		.INIT('hd0)
	) name28631 (
		_w16217_,
		_w16219_,
		_w16226_,
		_w34458_
	);
	LUT3 #(
		.INIT('h51)
	) name28632 (
		_w16235_,
		_w16236_,
		_w34458_,
		_w34459_
	);
	LUT3 #(
		.INIT('h10)
	) name28633 (
		_w34457_,
		_w34455_,
		_w34459_,
		_w34460_
	);
	LUT4 #(
		.INIT('h0ca6)
	) name28634 (
		_w16216_,
		_w16217_,
		_w16219_,
		_w16220_,
		_w34461_
	);
	LUT3 #(
		.INIT('h31)
	) name28635 (
		_w16226_,
		_w16500_,
		_w34461_,
		_w34462_
	);
	LUT2 #(
		.INIT('h4)
	) name28636 (
		_w16232_,
		_w16235_,
		_w34463_
	);
	LUT2 #(
		.INIT('h4)
	) name28637 (
		_w34462_,
		_w34463_,
		_w34464_
	);
	LUT4 #(
		.INIT('h999a)
	) name28638 (
		\u1_L12_reg[5]/NET0131 ,
		_w34453_,
		_w34460_,
		_w34464_,
		_w34465_
	);
	LUT4 #(
		.INIT('h70e0)
	) name28639 (
		_w28755_,
		_w28754_,
		_w28757_,
		_w28752_,
		_w34466_
	);
	LUT3 #(
		.INIT('h23)
	) name28640 (
		_w28754_,
		_w28757_,
		_w28752_,
		_w34467_
	);
	LUT3 #(
		.INIT('h23)
	) name28641 (
		_w28802_,
		_w34466_,
		_w34467_,
		_w34468_
	);
	LUT4 #(
		.INIT('h0001)
	) name28642 (
		_w28766_,
		_w28814_,
		_w28986_,
		_w28992_,
		_w34469_
	);
	LUT3 #(
		.INIT('h10)
	) name28643 (
		_w28989_,
		_w34468_,
		_w34469_,
		_w34470_
	);
	LUT4 #(
		.INIT('h0012)
	) name28644 (
		_w28755_,
		_w28753_,
		_w28754_,
		_w28757_,
		_w34471_
	);
	LUT4 #(
		.INIT('h1000)
	) name28645 (
		_w28755_,
		_w28754_,
		_w28757_,
		_w28752_,
		_w34472_
	);
	LUT4 #(
		.INIT('h0002)
	) name28646 (
		_w28766_,
		_w28773_,
		_w28775_,
		_w34472_,
		_w34473_
	);
	LUT3 #(
		.INIT('h07)
	) name28647 (
		_w28756_,
		_w28765_,
		_w28806_,
		_w34474_
	);
	LUT3 #(
		.INIT('h40)
	) name28648 (
		_w34471_,
		_w34473_,
		_w34474_,
		_w34475_
	);
	LUT3 #(
		.INIT('hf6)
	) name28649 (
		_w28755_,
		_w28753_,
		_w28752_,
		_w34476_
	);
	LUT2 #(
		.INIT('h2)
	) name28650 (
		_w28761_,
		_w34476_,
		_w34477_
	);
	LUT4 #(
		.INIT('h8caf)
	) name28651 (
		_w28753_,
		_w28757_,
		_w28773_,
		_w28775_,
		_w34478_
	);
	LUT2 #(
		.INIT('h4)
	) name28652 (
		_w34477_,
		_w34478_,
		_w34479_
	);
	LUT4 #(
		.INIT('ha955)
	) name28653 (
		\u0_L7_reg[20]/NET0131 ,
		_w34470_,
		_w34475_,
		_w34479_,
		_w34480_
	);
	LUT4 #(
		.INIT('h0403)
	) name28654 (
		_w33908_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w34481_
	);
	LUT3 #(
		.INIT('h47)
	) name28655 (
		_w33908_,
		_w33909_,
		_w33911_,
		_w34482_
	);
	LUT2 #(
		.INIT('h8)
	) name28656 (
		_w33910_,
		_w33913_,
		_w34483_
	);
	LUT4 #(
		.INIT('hbfee)
	) name28657 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w34484_
	);
	LUT4 #(
		.INIT('h0b00)
	) name28658 (
		_w34482_,
		_w34483_,
		_w34481_,
		_w34484_,
		_w34485_
	);
	LUT4 #(
		.INIT('h2028)
	) name28659 (
		_w33908_,
		_w33910_,
		_w33909_,
		_w33913_,
		_w34486_
	);
	LUT3 #(
		.INIT('he4)
	) name28660 (
		_w33910_,
		_w33909_,
		_w33911_,
		_w34487_
	);
	LUT2 #(
		.INIT('h4)
	) name28661 (
		_w33908_,
		_w33913_,
		_w34488_
	);
	LUT4 #(
		.INIT('h1011)
	) name28662 (
		_w33938_,
		_w34486_,
		_w34487_,
		_w34488_,
		_w34489_
	);
	LUT4 #(
		.INIT('h0040)
	) name28663 (
		_w33908_,
		_w33910_,
		_w33909_,
		_w33913_,
		_w34490_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name28664 (
		_w33910_,
		_w33909_,
		_w33913_,
		_w33911_,
		_w34491_
	);
	LUT3 #(
		.INIT('h31)
	) name28665 (
		_w33908_,
		_w34490_,
		_w34491_,
		_w34492_
	);
	LUT4 #(
		.INIT('hd800)
	) name28666 (
		_w33917_,
		_w34489_,
		_w34485_,
		_w34492_,
		_w34493_
	);
	LUT2 #(
		.INIT('h9)
	) name28667 (
		\u0_desIn_r_reg[10]/NET0131 ,
		_w34493_,
		_w34494_
	);
	LUT4 #(
		.INIT('h0008)
	) name28668 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w34495_
	);
	LUT4 #(
		.INIT('h0008)
	) name28669 (
		_w17540_,
		_w17546_,
		_w17749_,
		_w34495_,
		_w34496_
	);
	LUT4 #(
		.INIT('h0800)
	) name28670 (
		_w17534_,
		_w17536_,
		_w17537_,
		_w17542_,
		_w34497_
	);
	LUT3 #(
		.INIT('h01)
	) name28671 (
		_w17540_,
		_w17750_,
		_w34497_,
		_w34498_
	);
	LUT2 #(
		.INIT('h1)
	) name28672 (
		_w34496_,
		_w34498_,
		_w34499_
	);
	LUT4 #(
		.INIT('h8caf)
	) name28673 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w34500_
	);
	LUT3 #(
		.INIT('h02)
	) name28674 (
		_w17540_,
		_w17750_,
		_w34500_,
		_w34501_
	);
	LUT4 #(
		.INIT('h0001)
	) name28675 (
		_w17534_,
		_w17536_,
		_w17537_,
		_w17540_,
		_w34502_
	);
	LUT3 #(
		.INIT('h02)
	) name28676 (
		_w17542_,
		_w17557_,
		_w34502_,
		_w34503_
	);
	LUT2 #(
		.INIT('h4)
	) name28677 (
		_w34501_,
		_w34503_,
		_w34504_
	);
	LUT4 #(
		.INIT('hffd3)
	) name28678 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w34505_
	);
	LUT2 #(
		.INIT('h2)
	) name28679 (
		_w17540_,
		_w34505_,
		_w34506_
	);
	LUT4 #(
		.INIT('hefaa)
	) name28680 (
		_w17534_,
		_w17535_,
		_w17537_,
		_w17540_,
		_w34507_
	);
	LUT2 #(
		.INIT('h2)
	) name28681 (
		_w17536_,
		_w34507_,
		_w34508_
	);
	LUT3 #(
		.INIT('h4e)
	) name28682 (
		_w17535_,
		_w17536_,
		_w17537_,
		_w34509_
	);
	LUT3 #(
		.INIT('h0e)
	) name28683 (
		_w17534_,
		_w17535_,
		_w17540_,
		_w34510_
	);
	LUT4 #(
		.INIT('h8000)
	) name28684 (
		_w17534_,
		_w17535_,
		_w17536_,
		_w17537_,
		_w34511_
	);
	LUT4 #(
		.INIT('h1011)
	) name28685 (
		_w17542_,
		_w34511_,
		_w34509_,
		_w34510_,
		_w34512_
	);
	LUT3 #(
		.INIT('h10)
	) name28686 (
		_w34506_,
		_w34508_,
		_w34512_,
		_w34513_
	);
	LUT4 #(
		.INIT('h999a)
	) name28687 (
		\u1_L10_reg[5]/NET0131 ,
		_w34499_,
		_w34504_,
		_w34513_,
		_w34514_
	);
	LUT4 #(
		.INIT('hbf00)
	) name28688 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22916_,
		_w34515_
	);
	LUT3 #(
		.INIT('h51)
	) name28689 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w34516_
	);
	LUT4 #(
		.INIT('h8000)
	) name28690 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w34517_
	);
	LUT4 #(
		.INIT('h0041)
	) name28691 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w22916_,
		_w34518_
	);
	LUT4 #(
		.INIT('h0301)
	) name28692 (
		_w34515_,
		_w34517_,
		_w34518_,
		_w34516_,
		_w34519_
	);
	LUT4 #(
		.INIT('h400c)
	) name28693 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22916_,
		_w34520_
	);
	LUT4 #(
		.INIT('hdead)
	) name28694 (
		_w22913_,
		_w22910_,
		_w22911_,
		_w22912_,
		_w34521_
	);
	LUT3 #(
		.INIT('h10)
	) name28695 (
		_w22926_,
		_w34520_,
		_w34521_,
		_w34522_
	);
	LUT3 #(
		.INIT('hd7)
	) name28696 (
		_w22910_,
		_w22911_,
		_w22912_,
		_w34523_
	);
	LUT4 #(
		.INIT('hbfae)
	) name28697 (
		_w22913_,
		_w22916_,
		_w22925_,
		_w34523_,
		_w34524_
	);
	LUT4 #(
		.INIT('hd800)
	) name28698 (
		_w22909_,
		_w34522_,
		_w34519_,
		_w34524_,
		_w34525_
	);
	LUT2 #(
		.INIT('h9)
	) name28699 (
		\u1_L1_reg[19]/P0001 ,
		_w34525_,
		_w34526_
	);
	LUT4 #(
		.INIT('h3fef)
	) name28700 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w34527_
	);
	LUT2 #(
		.INIT('h1)
	) name28701 (
		_w26877_,
		_w34527_,
		_w34528_
	);
	LUT4 #(
		.INIT('h0002)
	) name28702 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w34529_
	);
	LUT3 #(
		.INIT('h04)
	) name28703 (
		_w26886_,
		_w26884_,
		_w34529_,
		_w34530_
	);
	LUT2 #(
		.INIT('h1)
	) name28704 (
		_w26877_,
		_w26878_,
		_w34531_
	);
	LUT3 #(
		.INIT('h40)
	) name28705 (
		_w26880_,
		_w26881_,
		_w26882_,
		_w34532_
	);
	LUT3 #(
		.INIT('h45)
	) name28706 (
		_w27089_,
		_w34531_,
		_w34532_,
		_w34533_
	);
	LUT3 #(
		.INIT('h40)
	) name28707 (
		_w34528_,
		_w34530_,
		_w34533_,
		_w34534_
	);
	LUT2 #(
		.INIT('h8)
	) name28708 (
		_w26879_,
		_w27086_,
		_w34535_
	);
	LUT4 #(
		.INIT('h00fb)
	) name28709 (
		_w26878_,
		_w26880_,
		_w26882_,
		_w26884_,
		_w34536_
	);
	LUT3 #(
		.INIT('h10)
	) name28710 (
		_w26895_,
		_w26900_,
		_w34536_,
		_w34537_
	);
	LUT2 #(
		.INIT('h4)
	) name28711 (
		_w34535_,
		_w34537_,
		_w34538_
	);
	LUT4 #(
		.INIT('h0086)
	) name28712 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w34539_
	);
	LUT4 #(
		.INIT('heafa)
	) name28713 (
		_w26878_,
		_w26880_,
		_w26881_,
		_w26882_,
		_w34540_
	);
	LUT4 #(
		.INIT('h0504)
	) name28714 (
		_w26877_,
		_w26884_,
		_w34539_,
		_w34540_,
		_w34541_
	);
	LUT3 #(
		.INIT('h02)
	) name28715 (
		_w26877_,
		_w26887_,
		_w26900_,
		_w34542_
	);
	LUT2 #(
		.INIT('h1)
	) name28716 (
		_w34541_,
		_w34542_,
		_w34543_
	);
	LUT4 #(
		.INIT('h55a9)
	) name28717 (
		\u0_L10_reg[26]/NET0131 ,
		_w34534_,
		_w34538_,
		_w34543_,
		_w34544_
	);
	LUT4 #(
		.INIT('h7776)
	) name28718 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w34545_
	);
	LUT2 #(
		.INIT('h2)
	) name28719 (
		_w31137_,
		_w34545_,
		_w34546_
	);
	LUT4 #(
		.INIT('h0660)
	) name28720 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w34547_
	);
	LUT4 #(
		.INIT('h008a)
	) name28721 (
		_w31136_,
		_w31137_,
		_w31157_,
		_w34547_,
		_w34548_
	);
	LUT3 #(
		.INIT('h27)
	) name28722 (
		_w31142_,
		_w31138_,
		_w31137_,
		_w34549_
	);
	LUT4 #(
		.INIT('h0002)
	) name28723 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w34550_
	);
	LUT4 #(
		.INIT('h0501)
	) name28724 (
		_w31136_,
		_w31141_,
		_w34550_,
		_w34549_,
		_w34551_
	);
	LUT4 #(
		.INIT('h134c)
	) name28725 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w34552_
	);
	LUT4 #(
		.INIT('h2014)
	) name28726 (
		_w31139_,
		_w31142_,
		_w31138_,
		_w31140_,
		_w34553_
	);
	LUT3 #(
		.INIT('h0e)
	) name28727 (
		_w31137_,
		_w34552_,
		_w34553_,
		_w34554_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name28728 (
		_w34546_,
		_w34548_,
		_w34551_,
		_w34554_,
		_w34555_
	);
	LUT2 #(
		.INIT('h6)
	) name28729 (
		\u0_L3_reg[12]/NET0131 ,
		_w34555_,
		_w34556_
	);
	LUT4 #(
		.INIT('haaa7)
	) name28730 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w34557_
	);
	LUT2 #(
		.INIT('h2)
	) name28731 (
		_w31165_,
		_w34557_,
		_w34558_
	);
	LUT4 #(
		.INIT('h00a1)
	) name28732 (
		_w31166_,
		_w31167_,
		_w31169_,
		_w31165_,
		_w34559_
	);
	LUT4 #(
		.INIT('h7f00)
	) name28733 (
		_w31168_,
		_w31167_,
		_w31169_,
		_w31164_,
		_w34560_
	);
	LUT3 #(
		.INIT('h10)
	) name28734 (
		_w31499_,
		_w34559_,
		_w34560_,
		_w34561_
	);
	LUT4 #(
		.INIT('h0919)
	) name28735 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w34562_
	);
	LUT4 #(
		.INIT('h1040)
	) name28736 (
		_w31166_,
		_w31168_,
		_w31167_,
		_w31169_,
		_w34563_
	);
	LUT4 #(
		.INIT('hfad8)
	) name28737 (
		_w31165_,
		_w31495_,
		_w34562_,
		_w34563_,
		_w34564_
	);
	LUT3 #(
		.INIT('h01)
	) name28738 (
		_w31164_,
		_w31170_,
		_w31188_,
		_w34565_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name28739 (
		_w34558_,
		_w34561_,
		_w34564_,
		_w34565_,
		_w34566_
	);
	LUT2 #(
		.INIT('h6)
	) name28740 (
		\u0_L3_reg[17]/NET0131 ,
		_w34566_,
		_w34567_
	);
	LUT4 #(
		.INIT('hfb9e)
	) name28741 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w34568_
	);
	LUT4 #(
		.INIT('hfd00)
	) name28742 (
		_w13040_,
		_w13218_,
		_w13216_,
		_w34568_,
		_w34569_
	);
	LUT2 #(
		.INIT('h2)
	) name28743 (
		_w13043_,
		_w34569_,
		_w34570_
	);
	LUT4 #(
		.INIT('hffa7)
	) name28744 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w34571_
	);
	LUT2 #(
		.INIT('h2)
	) name28745 (
		_w13043_,
		_w34571_,
		_w34572_
	);
	LUT4 #(
		.INIT('h0026)
	) name28746 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13043_,
		_w34573_
	);
	LUT3 #(
		.INIT('h70)
	) name28747 (
		_w13035_,
		_w13036_,
		_w13043_,
		_w34574_
	);
	LUT4 #(
		.INIT('h0301)
	) name28748 (
		_w13081_,
		_w13216_,
		_w34573_,
		_w34574_,
		_w34575_
	);
	LUT3 #(
		.INIT('h45)
	) name28749 (
		_w13040_,
		_w34572_,
		_w34575_,
		_w34576_
	);
	LUT4 #(
		.INIT('h0009)
	) name28750 (
		_w13035_,
		_w13036_,
		_w13038_,
		_w13043_,
		_w34577_
	);
	LUT3 #(
		.INIT('ha8)
	) name28751 (
		_w13040_,
		_w13058_,
		_w34577_,
		_w34578_
	);
	LUT2 #(
		.INIT('h1)
	) name28752 (
		_w13217_,
		_w34578_,
		_w34579_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name28753 (
		\u2_L2_reg[5]/NET0131 ,
		_w34576_,
		_w34570_,
		_w34579_,
		_w34580_
	);
	LUT3 #(
		.INIT('h15)
	) name28754 (
		_w17938_,
		_w17943_,
		_w17940_,
		_w34581_
	);
	LUT4 #(
		.INIT('h8008)
	) name28755 (
		_w17938_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w34582_
	);
	LUT4 #(
		.INIT('h0820)
	) name28756 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w34583_
	);
	LUT4 #(
		.INIT('h0103)
	) name28757 (
		_w18465_,
		_w34582_,
		_w34583_,
		_w34581_,
		_w34584_
	);
	LUT3 #(
		.INIT('hed)
	) name28758 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w34585_
	);
	LUT2 #(
		.INIT('h2)
	) name28759 (
		_w18328_,
		_w34585_,
		_w34586_
	);
	LUT4 #(
		.INIT('hcc9d)
	) name28760 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w34587_
	);
	LUT4 #(
		.INIT('h4041)
	) name28761 (
		_w17938_,
		_w17942_,
		_w17943_,
		_w17940_,
		_w34588_
	);
	LUT4 #(
		.INIT('h5bff)
	) name28762 (
		_w17942_,
		_w17943_,
		_w17939_,
		_w17940_,
		_w34589_
	);
	LUT4 #(
		.INIT('h0d00)
	) name28763 (
		_w17938_,
		_w34587_,
		_w34588_,
		_w34589_,
		_w34590_
	);
	LUT4 #(
		.INIT('h0e04)
	) name28764 (
		_w17937_,
		_w34584_,
		_w34586_,
		_w34590_,
		_w34591_
	);
	LUT2 #(
		.INIT('h9)
	) name28765 (
		\u1_L9_reg[17]/NET0131 ,
		_w34591_,
		_w34592_
	);
	LUT4 #(
		.INIT('h7c00)
	) name28766 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28255_,
		_w34593_
	);
	LUT4 #(
		.INIT('hfaee)
	) name28767 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w34594_
	);
	LUT4 #(
		.INIT('h00fd)
	) name28768 (
		_w28257_,
		_w28259_,
		_w28254_,
		_w28255_,
		_w34595_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name28769 (
		_w28433_,
		_w34593_,
		_w34594_,
		_w34595_,
		_w34596_
	);
	LUT4 #(
		.INIT('hbf77)
	) name28770 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w34597_
	);
	LUT3 #(
		.INIT('h8a)
	) name28771 (
		_w28270_,
		_w34596_,
		_w34597_,
		_w34598_
	);
	LUT4 #(
		.INIT('he3ef)
	) name28772 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w34599_
	);
	LUT2 #(
		.INIT('h4)
	) name28773 (
		_w28258_,
		_w28255_,
		_w34600_
	);
	LUT3 #(
		.INIT('hb0)
	) name28774 (
		_w28258_,
		_w28257_,
		_w28255_,
		_w34601_
	);
	LUT4 #(
		.INIT('h0f01)
	) name28775 (
		_w28257_,
		_w28259_,
		_w28254_,
		_w28255_,
		_w34602_
	);
	LUT4 #(
		.INIT('he0ee)
	) name28776 (
		_w34599_,
		_w34600_,
		_w34601_,
		_w34602_,
		_w34603_
	);
	LUT4 #(
		.INIT('hbefd)
	) name28777 (
		_w28258_,
		_w28257_,
		_w28259_,
		_w28254_,
		_w34604_
	);
	LUT4 #(
		.INIT('h0040)
	) name28778 (
		_w28257_,
		_w28259_,
		_w28254_,
		_w28255_,
		_w34605_
	);
	LUT4 #(
		.INIT('h0031)
	) name28779 (
		_w28255_,
		_w28275_,
		_w34604_,
		_w34605_,
		_w34606_
	);
	LUT3 #(
		.INIT('he0)
	) name28780 (
		_w28270_,
		_w34603_,
		_w34606_,
		_w34607_
	);
	LUT3 #(
		.INIT('h65)
	) name28781 (
		\u0_L8_reg[25]/NET0131 ,
		_w34598_,
		_w34607_,
		_w34608_
	);
	LUT4 #(
		.INIT('h3dc3)
	) name28782 (
		_w19030_,
		_w19031_,
		_w19034_,
		_w19032_,
		_w34609_
	);
	LUT4 #(
		.INIT('h0110)
	) name28783 (
		_w19030_,
		_w19031_,
		_w19034_,
		_w19033_,
		_w34610_
	);
	LUT4 #(
		.INIT('h0032)
	) name28784 (
		_w19033_,
		_w19049_,
		_w34609_,
		_w34610_,
		_w34611_
	);
	LUT4 #(
		.INIT('h76dc)
	) name28785 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w34612_
	);
	LUT4 #(
		.INIT('h2880)
	) name28786 (
		_w19030_,
		_w19031_,
		_w19034_,
		_w19032_,
		_w34613_
	);
	LUT4 #(
		.INIT('h00f2)
	) name28787 (
		_w19030_,
		_w19039_,
		_w34612_,
		_w34613_,
		_w34614_
	);
	LUT4 #(
		.INIT('h0040)
	) name28788 (
		_w19030_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w34615_
	);
	LUT4 #(
		.INIT('hbfef)
	) name28789 (
		_w19031_,
		_w19034_,
		_w19033_,
		_w19032_,
		_w34616_
	);
	LUT3 #(
		.INIT('h31)
	) name28790 (
		_w19030_,
		_w34615_,
		_w34616_,
		_w34617_
	);
	LUT4 #(
		.INIT('hd800)
	) name28791 (
		_w19038_,
		_w34611_,
		_w34614_,
		_w34617_,
		_w34618_
	);
	LUT2 #(
		.INIT('h9)
	) name28792 (
		\u1_L8_reg[16]/NET0131 ,
		_w34618_,
		_w34619_
	);
	LUT4 #(
		.INIT('hefcc)
	) name28793 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w34620_
	);
	LUT4 #(
		.INIT('h0806)
	) name28794 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w34621_
	);
	LUT4 #(
		.INIT('h5501)
	) name28795 (
		_w21765_,
		_w21761_,
		_w34620_,
		_w34621_,
		_w34622_
	);
	LUT4 #(
		.INIT('h0010)
	) name28796 (
		_w21762_,
		_w21764_,
		_w21765_,
		_w21763_,
		_w34623_
	);
	LUT4 #(
		.INIT('hff7b)
	) name28797 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w34624_
	);
	LUT2 #(
		.INIT('h4)
	) name28798 (
		_w34623_,
		_w34624_,
		_w34625_
	);
	LUT4 #(
		.INIT('habff)
	) name28799 (
		_w21762_,
		_w21764_,
		_w21765_,
		_w21763_,
		_w34626_
	);
	LUT4 #(
		.INIT('h5eff)
	) name28800 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w34627_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name28801 (
		_w21765_,
		_w21767_,
		_w34626_,
		_w34627_,
		_w34628_
	);
	LUT3 #(
		.INIT('h2a)
	) name28802 (
		_w21761_,
		_w34625_,
		_w34628_,
		_w34629_
	);
	LUT4 #(
		.INIT('hf9ff)
	) name28803 (
		_w21762_,
		_w21764_,
		_w21767_,
		_w21763_,
		_w34630_
	);
	LUT2 #(
		.INIT('h2)
	) name28804 (
		_w21765_,
		_w34630_,
		_w34631_
	);
	LUT3 #(
		.INIT('h80)
	) name28805 (
		_w21764_,
		_w21765_,
		_w21767_,
		_w34632_
	);
	LUT3 #(
		.INIT('h23)
	) name28806 (
		_w21768_,
		_w21893_,
		_w34632_,
		_w34633_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name28807 (
		_w21761_,
		_w21770_,
		_w34631_,
		_w34633_,
		_w34634_
	);
	LUT4 #(
		.INIT('h5655)
	) name28808 (
		\u1_L3_reg[26]/NET0131 ,
		_w34629_,
		_w34622_,
		_w34634_,
		_w34635_
	);
	LUT4 #(
		.INIT('hafab)
	) name28809 (
		_w21862_,
		_w21860_,
		_w21859_,
		_w21866_,
		_w34636_
	);
	LUT2 #(
		.INIT('h2)
	) name28810 (
		_w21861_,
		_w34636_,
		_w34637_
	);
	LUT3 #(
		.INIT('h01)
	) name28811 (
		_w21870_,
		_w21872_,
		_w22104_,
		_w34638_
	);
	LUT3 #(
		.INIT('he0)
	) name28812 (
		_w21861_,
		_w21859_,
		_w21866_,
		_w34639_
	);
	LUT3 #(
		.INIT('h15)
	) name28813 (
		_w21884_,
		_w22093_,
		_w34639_,
		_w34640_
	);
	LUT3 #(
		.INIT('h40)
	) name28814 (
		_w34637_,
		_w34638_,
		_w34640_,
		_w34641_
	);
	LUT4 #(
		.INIT('h00fb)
	) name28815 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21866_,
		_w34642_
	);
	LUT4 #(
		.INIT('hbf00)
	) name28816 (
		_w21862_,
		_w21860_,
		_w21859_,
		_w21866_,
		_w34643_
	);
	LUT4 #(
		.INIT('h77af)
	) name28817 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w34644_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name28818 (
		_w21965_,
		_w34642_,
		_w34643_,
		_w34644_,
		_w34645_
	);
	LUT4 #(
		.INIT('h0802)
	) name28819 (
		_w21861_,
		_w21862_,
		_w21860_,
		_w21859_,
		_w34646_
	);
	LUT3 #(
		.INIT('h02)
	) name28820 (
		_w21870_,
		_w21971_,
		_w34646_,
		_w34647_
	);
	LUT2 #(
		.INIT('h4)
	) name28821 (
		_w34645_,
		_w34647_,
		_w34648_
	);
	LUT4 #(
		.INIT('h0100)
	) name28822 (
		_w21861_,
		_w21862_,
		_w21859_,
		_w21866_,
		_w34649_
	);
	LUT3 #(
		.INIT('hd0)
	) name28823 (
		_w21859_,
		_w21866_,
		_w21870_,
		_w34650_
	);
	LUT3 #(
		.INIT('h45)
	) name28824 (
		_w21861_,
		_w21859_,
		_w21866_,
		_w34651_
	);
	LUT4 #(
		.INIT('h3133)
	) name28825 (
		_w22105_,
		_w34649_,
		_w34650_,
		_w34651_,
		_w34652_
	);
	LUT4 #(
		.INIT('ha955)
	) name28826 (
		\u1_L3_reg[21]/NET0131 ,
		_w34641_,
		_w34648_,
		_w34652_,
		_w34653_
	);
	LUT4 #(
		.INIT('haf84)
	) name28827 (
		_w26279_,
		_w26278_,
		_w26280_,
		_w26276_,
		_w34654_
	);
	LUT2 #(
		.INIT('h1)
	) name28828 (
		_w26277_,
		_w34654_,
		_w34655_
	);
	LUT3 #(
		.INIT('h0d)
	) name28829 (
		_w26289_,
		_w26314_,
		_w26333_,
		_w34656_
	);
	LUT3 #(
		.INIT('h45)
	) name28830 (
		_w26285_,
		_w34655_,
		_w34656_,
		_w34657_
	);
	LUT3 #(
		.INIT('h15)
	) name28831 (
		_w26284_,
		_w26294_,
		_w26339_,
		_w34658_
	);
	LUT4 #(
		.INIT('h0802)
	) name28832 (
		_w26277_,
		_w26279_,
		_w26278_,
		_w26280_,
		_w34659_
	);
	LUT4 #(
		.INIT('h0888)
	) name28833 (
		_w26279_,
		_w26278_,
		_w26280_,
		_w26276_,
		_w34660_
	);
	LUT3 #(
		.INIT('h23)
	) name28834 (
		_w26294_,
		_w34659_,
		_w34660_,
		_w34661_
	);
	LUT4 #(
		.INIT('h134c)
	) name28835 (
		_w26277_,
		_w26278_,
		_w26280_,
		_w26276_,
		_w34662_
	);
	LUT4 #(
		.INIT('ha521)
	) name28836 (
		_w26277_,
		_w26278_,
		_w26280_,
		_w26276_,
		_w34663_
	);
	LUT3 #(
		.INIT('h01)
	) name28837 (
		_w26279_,
		_w34663_,
		_w34662_,
		_w34664_
	);
	LUT4 #(
		.INIT('h00d5)
	) name28838 (
		_w26285_,
		_w34658_,
		_w34661_,
		_w34664_,
		_w34665_
	);
	LUT3 #(
		.INIT('h65)
	) name28839 (
		\u0_L11_reg[26]/NET0131 ,
		_w34657_,
		_w34665_,
		_w34666_
	);
	LUT4 #(
		.INIT('h3c3b)
	) name28840 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w34667_
	);
	LUT4 #(
		.INIT('h0010)
	) name28841 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w34668_
	);
	LUT4 #(
		.INIT('h3302)
	) name28842 (
		_w5950_,
		_w5962_,
		_w34667_,
		_w34668_,
		_w34669_
	);
	LUT4 #(
		.INIT('h0400)
	) name28843 (
		_w5950_,
		_w5951_,
		_w5952_,
		_w5956_,
		_w34670_
	);
	LUT4 #(
		.INIT('h0008)
	) name28844 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w34671_
	);
	LUT4 #(
		.INIT('hbfb7)
	) name28845 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w34672_
	);
	LUT4 #(
		.INIT('h0002)
	) name28846 (
		_w5950_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w34673_
	);
	LUT4 #(
		.INIT('h0100)
	) name28847 (
		_w6094_,
		_w34673_,
		_w34670_,
		_w34672_,
		_w34674_
	);
	LUT2 #(
		.INIT('h2)
	) name28848 (
		_w5962_,
		_w34674_,
		_w34675_
	);
	LUT4 #(
		.INIT('h2420)
	) name28849 (
		_w5951_,
		_w5952_,
		_w5953_,
		_w5956_,
		_w34676_
	);
	LUT4 #(
		.INIT('h0001)
	) name28850 (
		_w5950_,
		_w5964_,
		_w34676_,
		_w34671_,
		_w34677_
	);
	LUT3 #(
		.INIT('h02)
	) name28851 (
		_w5950_,
		_w5960_,
		_w6098_,
		_w34678_
	);
	LUT4 #(
		.INIT('h0010)
	) name28852 (
		_w5950_,
		_w5952_,
		_w5953_,
		_w5962_,
		_w34679_
	);
	LUT3 #(
		.INIT('h0e)
	) name28853 (
		_w34677_,
		_w34678_,
		_w34679_,
		_w34680_
	);
	LUT4 #(
		.INIT('h5655)
	) name28854 (
		\u2_L13_reg[15]/NET0131 ,
		_w34669_,
		_w34675_,
		_w34680_,
		_w34681_
	);
	LUT4 #(
		.INIT('hef11)
	) name28855 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w34682_
	);
	LUT4 #(
		.INIT('h5001)
	) name28856 (
		_w16681_,
		_w16682_,
		_w16684_,
		_w16685_,
		_w34683_
	);
	LUT4 #(
		.INIT('h7d7f)
	) name28857 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w34684_
	);
	LUT4 #(
		.INIT('h0d00)
	) name28858 (
		_w16681_,
		_w34682_,
		_w34683_,
		_w34684_,
		_w34685_
	);
	LUT4 #(
		.INIT('haff8)
	) name28859 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w34686_
	);
	LUT4 #(
		.INIT('h0840)
	) name28860 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w16685_,
		_w34687_
	);
	LUT4 #(
		.INIT('h8200)
	) name28861 (
		_w16681_,
		_w16682_,
		_w16683_,
		_w16685_,
		_w34688_
	);
	LUT4 #(
		.INIT('h0032)
	) name28862 (
		_w16681_,
		_w34687_,
		_w34686_,
		_w34688_,
		_w34689_
	);
	LUT3 #(
		.INIT('hd7)
	) name28863 (
		_w16682_,
		_w16684_,
		_w16683_,
		_w34690_
	);
	LUT2 #(
		.INIT('h2)
	) name28864 (
		_w16696_,
		_w34690_,
		_w34691_
	);
	LUT4 #(
		.INIT('h0e04)
	) name28865 (
		_w16693_,
		_w34689_,
		_w34691_,
		_w34685_,
		_w34692_
	);
	LUT2 #(
		.INIT('h9)
	) name28866 (
		\u1_L11_reg[17]/NET0131 ,
		_w34692_,
		_w34693_
	);
	LUT4 #(
		.INIT('hb8b3)
	) name28867 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w34694_
	);
	LUT2 #(
		.INIT('h2)
	) name28868 (
		_w18791_,
		_w18794_,
		_w34695_
	);
	LUT3 #(
		.INIT('h08)
	) name28869 (
		_w18791_,
		_w18792_,
		_w18794_,
		_w34696_
	);
	LUT4 #(
		.INIT('h0514)
	) name28870 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w34697_
	);
	LUT4 #(
		.INIT('h0031)
	) name28871 (
		_w18794_,
		_w34696_,
		_w34694_,
		_w34697_,
		_w34698_
	);
	LUT2 #(
		.INIT('h2)
	) name28872 (
		_w18800_,
		_w34698_,
		_w34699_
	);
	LUT3 #(
		.INIT('hbc)
	) name28873 (
		_w18791_,
		_w18792_,
		_w18790_,
		_w34700_
	);
	LUT3 #(
		.INIT('h0b)
	) name28874 (
		_w18791_,
		_w18789_,
		_w18794_,
		_w34701_
	);
	LUT2 #(
		.INIT('h4)
	) name28875 (
		_w34700_,
		_w34701_,
		_w34702_
	);
	LUT4 #(
		.INIT('hdfee)
	) name28876 (
		_w18789_,
		_w18792_,
		_w18794_,
		_w18790_,
		_w34703_
	);
	LUT2 #(
		.INIT('h2)
	) name28877 (
		_w18791_,
		_w34703_,
		_w34704_
	);
	LUT3 #(
		.INIT('h08)
	) name28878 (
		_w18789_,
		_w18792_,
		_w18790_,
		_w34705_
	);
	LUT4 #(
		.INIT('h7077)
	) name28879 (
		_w18806_,
		_w18985_,
		_w34695_,
		_w34705_,
		_w34706_
	);
	LUT4 #(
		.INIT('h5455)
	) name28880 (
		_w18800_,
		_w34704_,
		_w34702_,
		_w34706_,
		_w34707_
	);
	LUT4 #(
		.INIT('h7bdd)
	) name28881 (
		_w18791_,
		_w18789_,
		_w18792_,
		_w18790_,
		_w34708_
	);
	LUT2 #(
		.INIT('h1)
	) name28882 (
		_w18794_,
		_w34708_,
		_w34709_
	);
	LUT4 #(
		.INIT('h0040)
	) name28883 (
		_w18791_,
		_w18792_,
		_w18794_,
		_w18790_,
		_w34710_
	);
	LUT3 #(
		.INIT('h07)
	) name28884 (
		_w18986_,
		_w18987_,
		_w34710_,
		_w34711_
	);
	LUT2 #(
		.INIT('h4)
	) name28885 (
		_w34709_,
		_w34711_,
		_w34712_
	);
	LUT4 #(
		.INIT('h5655)
	) name28886 (
		\u1_L8_reg[31]/NET0131 ,
		_w34707_,
		_w34699_,
		_w34712_,
		_w34713_
	);
	LUT3 #(
		.INIT('h04)
	) name28887 (
		_w20125_,
		_w20128_,
		_w20127_,
		_w34714_
	);
	LUT4 #(
		.INIT('hdf00)
	) name28888 (
		_w20128_,
		_w20126_,
		_w20127_,
		_w20124_,
		_w34715_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name28889 (
		_w20134_,
		_w20380_,
		_w34714_,
		_w34715_,
		_w34716_
	);
	LUT4 #(
		.INIT('h0002)
	) name28890 (
		_w20123_,
		_w20166_,
		_w20167_,
		_w20387_,
		_w34717_
	);
	LUT4 #(
		.INIT('h021a)
	) name28891 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w34718_
	);
	LUT3 #(
		.INIT('h04)
	) name28892 (
		_w20135_,
		_w20162_,
		_w34718_,
		_w34719_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name28893 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w34720_
	);
	LUT4 #(
		.INIT('hf400)
	) name28894 (
		_w34716_,
		_w34717_,
		_w34719_,
		_w34720_,
		_w34721_
	);
	LUT4 #(
		.INIT('h1121)
	) name28895 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w34722_
	);
	LUT4 #(
		.INIT('hc244)
	) name28896 (
		_w20125_,
		_w20128_,
		_w20126_,
		_w20127_,
		_w34723_
	);
	LUT2 #(
		.INIT('h2)
	) name28897 (
		_w20124_,
		_w20123_,
		_w34724_
	);
	LUT3 #(
		.INIT('h10)
	) name28898 (
		_w34723_,
		_w34722_,
		_w34724_,
		_w34725_
	);
	LUT3 #(
		.INIT('h56)
	) name28899 (
		\u1_L6_reg[13]/NET0131 ,
		_w34721_,
		_w34725_,
		_w34726_
	);
	LUT4 #(
		.INIT('h0020)
	) name28900 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w34727_
	);
	LUT4 #(
		.INIT('h0009)
	) name28901 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w34728_
	);
	LUT4 #(
		.INIT('h0002)
	) name28902 (
		_w5984_,
		_w6123_,
		_w34728_,
		_w34727_,
		_w34729_
	);
	LUT3 #(
		.INIT('h06)
	) name28903 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w34730_
	);
	LUT3 #(
		.INIT('h01)
	) name28904 (
		_w5984_,
		_w5999_,
		_w34730_,
		_w34731_
	);
	LUT2 #(
		.INIT('h8)
	) name28905 (
		_w5983_,
		_w5993_,
		_w34732_
	);
	LUT4 #(
		.INIT('h1000)
	) name28906 (
		_w5985_,
		_w5987_,
		_w5986_,
		_w5984_,
		_w34733_
	);
	LUT4 #(
		.INIT('h0002)
	) name28907 (
		_w5982_,
		_w5999_,
		_w6080_,
		_w34733_,
		_w34734_
	);
	LUT4 #(
		.INIT('h0e00)
	) name28908 (
		_w34729_,
		_w34731_,
		_w34732_,
		_w34734_,
		_w34735_
	);
	LUT4 #(
		.INIT('hcc5f)
	) name28909 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w34736_
	);
	LUT3 #(
		.INIT('h10)
	) name28910 (
		_w5984_,
		_w5999_,
		_w34736_,
		_w34737_
	);
	LUT4 #(
		.INIT('h37ae)
	) name28911 (
		_w5985_,
		_w5987_,
		_w5983_,
		_w5986_,
		_w34738_
	);
	LUT4 #(
		.INIT('h0200)
	) name28912 (
		_w5984_,
		_w34728_,
		_w34727_,
		_w34738_,
		_w34739_
	);
	LUT3 #(
		.INIT('h04)
	) name28913 (
		_w5982_,
		_w5995_,
		_w6126_,
		_w34740_
	);
	LUT3 #(
		.INIT('he0)
	) name28914 (
		_w34737_,
		_w34739_,
		_w34740_,
		_w34741_
	);
	LUT3 #(
		.INIT('ha9)
	) name28915 (
		\u2_L13_reg[20]/NET0131 ,
		_w34735_,
		_w34741_,
		_w34742_
	);
	LUT3 #(
		.INIT('h40)
	) name28916 (
		_w24794_,
		_w24796_,
		_w24792_,
		_w34743_
	);
	LUT2 #(
		.INIT('h4)
	) name28917 (
		_w24795_,
		_w24796_,
		_w34744_
	);
	LUT4 #(
		.INIT('h8acf)
	) name28918 (
		_w24794_,
		_w24795_,
		_w24796_,
		_w24792_,
		_w34745_
	);
	LUT3 #(
		.INIT('h02)
	) name28919 (
		_w24793_,
		_w34745_,
		_w34743_,
		_w34746_
	);
	LUT4 #(
		.INIT('h0007)
	) name28920 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24792_,
		_w34747_
	);
	LUT3 #(
		.INIT('h45)
	) name28921 (
		_w24791_,
		_w34744_,
		_w34747_,
		_w34748_
	);
	LUT3 #(
		.INIT('h04)
	) name28922 (
		_w24795_,
		_w24793_,
		_w24796_,
		_w34749_
	);
	LUT4 #(
		.INIT('h00f7)
	) name28923 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24792_,
		_w34750_
	);
	LUT4 #(
		.INIT('h1105)
	) name28924 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w34751_
	);
	LUT3 #(
		.INIT('h80)
	) name28925 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w34752_
	);
	LUT4 #(
		.INIT('h7c00)
	) name28926 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24792_,
		_w34753_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name28927 (
		_w34749_,
		_w34750_,
		_w34751_,
		_w34753_,
		_w34754_
	);
	LUT4 #(
		.INIT('h4000)
	) name28928 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w34755_
	);
	LUT4 #(
		.INIT('haa2a)
	) name28929 (
		_w24791_,
		_w24794_,
		_w24793_,
		_w24796_,
		_w34756_
	);
	LUT2 #(
		.INIT('h4)
	) name28930 (
		_w34755_,
		_w34756_,
		_w34757_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name28931 (
		_w34746_,
		_w34748_,
		_w34754_,
		_w34757_,
		_w34758_
	);
	LUT4 #(
		.INIT('hf7c7)
	) name28932 (
		_w24794_,
		_w24793_,
		_w24796_,
		_w24792_,
		_w34759_
	);
	LUT4 #(
		.INIT('hbefd)
	) name28933 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w34760_
	);
	LUT4 #(
		.INIT('hf531)
	) name28934 (
		_w24795_,
		_w24792_,
		_w34759_,
		_w34760_,
		_w34761_
	);
	LUT3 #(
		.INIT('h65)
	) name28935 (
		\u0_L14_reg[25]/P0001 ,
		_w34758_,
		_w34761_,
		_w34762_
	);
	LUT4 #(
		.INIT('hc963)
	) name28936 (
		decrypt_pad,
		\u0_R14_reg[16]/NET0131 ,
		\u0_uk_K_r14_reg[33]/NET0131 ,
		\u0_uk_K_r14_reg[40]/NET0131 ,
		_w34763_
	);
	LUT4 #(
		.INIT('hc693)
	) name28937 (
		decrypt_pad,
		\u0_R14_reg[12]/NET0131 ,
		\u0_uk_K_r14_reg[4]/NET0131 ,
		\u0_uk_K_r14_reg[54]/NET0131 ,
		_w34764_
	);
	LUT4 #(
		.INIT('hc963)
	) name28938 (
		decrypt_pad,
		\u0_R14_reg[15]/NET0131 ,
		\u0_uk_K_r14_reg[25]/NET0131 ,
		\u0_uk_K_r14_reg[32]/NET0131 ,
		_w34765_
	);
	LUT4 #(
		.INIT('hc963)
	) name28939 (
		decrypt_pad,
		\u0_R14_reg[14]/NET0131 ,
		\u0_uk_K_r14_reg[17]/NET0131 ,
		\u0_uk_K_r14_reg[24]/NET0131 ,
		_w34766_
	);
	LUT4 #(
		.INIT('hc963)
	) name28940 (
		decrypt_pad,
		\u0_R14_reg[13]/NET0131 ,
		\u0_uk_K_r14_reg[48]/NET0131 ,
		\u0_uk_K_r14_reg[55]/NET0131 ,
		_w34767_
	);
	LUT4 #(
		.INIT('hc963)
	) name28941 (
		decrypt_pad,
		\u0_R14_reg[17]/NET0131 ,
		\u0_uk_K_r14_reg[13]/NET0131 ,
		\u0_uk_K_r14_reg[20]/NET0131 ,
		_w34768_
	);
	LUT2 #(
		.INIT('h1)
	) name28942 (
		_w34766_,
		_w34765_,
		_w34769_
	);
	LUT4 #(
		.INIT('hc2cd)
	) name28943 (
		_w34768_,
		_w34766_,
		_w34767_,
		_w34765_,
		_w34770_
	);
	LUT2 #(
		.INIT('h2)
	) name28944 (
		_w34764_,
		_w34770_,
		_w34771_
	);
	LUT4 #(
		.INIT('h1000)
	) name28945 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34772_
	);
	LUT3 #(
		.INIT('h01)
	) name28946 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34773_
	);
	LUT4 #(
		.INIT('h0001)
	) name28947 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34774_
	);
	LUT4 #(
		.INIT('heffe)
	) name28948 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34775_
	);
	LUT4 #(
		.INIT('h0001)
	) name28949 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w34765_,
		_w34776_
	);
	LUT2 #(
		.INIT('h4)
	) name28950 (
		_w34764_,
		_w34768_,
		_w34777_
	);
	LUT4 #(
		.INIT('h0400)
	) name28951 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34765_,
		_w34778_
	);
	LUT3 #(
		.INIT('h02)
	) name28952 (
		_w34775_,
		_w34776_,
		_w34778_,
		_w34779_
	);
	LUT3 #(
		.INIT('h45)
	) name28953 (
		_w34763_,
		_w34771_,
		_w34779_,
		_w34780_
	);
	LUT2 #(
		.INIT('h8)
	) name28954 (
		_w34764_,
		_w34768_,
		_w34781_
	);
	LUT4 #(
		.INIT('h8000)
	) name28955 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34782_
	);
	LUT3 #(
		.INIT('h04)
	) name28956 (
		_w34764_,
		_w34766_,
		_w34767_,
		_w34783_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name28957 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34784_
	);
	LUT4 #(
		.INIT('h2022)
	) name28958 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34785_
	);
	LUT4 #(
		.INIT('h0400)
	) name28959 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34786_
	);
	LUT3 #(
		.INIT('h01)
	) name28960 (
		_w34785_,
		_w34765_,
		_w34786_,
		_w34787_
	);
	LUT4 #(
		.INIT('h0008)
	) name28961 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34788_
	);
	LUT4 #(
		.INIT('hef00)
	) name28962 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w34765_,
		_w34789_
	);
	LUT2 #(
		.INIT('h4)
	) name28963 (
		_w34788_,
		_w34789_,
		_w34790_
	);
	LUT4 #(
		.INIT('h5700)
	) name28964 (
		_w34784_,
		_w34787_,
		_w34790_,
		_w34763_,
		_w34791_
	);
	LUT4 #(
		.INIT('h7fbe)
	) name28965 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34792_
	);
	LUT2 #(
		.INIT('h1)
	) name28966 (
		_w34765_,
		_w34792_,
		_w34793_
	);
	LUT3 #(
		.INIT('h80)
	) name28967 (
		_w34766_,
		_w34767_,
		_w34765_,
		_w34794_
	);
	LUT4 #(
		.INIT('h4000)
	) name28968 (
		_w34764_,
		_w34766_,
		_w34767_,
		_w34765_,
		_w34795_
	);
	LUT4 #(
		.INIT('h2000)
	) name28969 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w34765_,
		_w34796_
	);
	LUT2 #(
		.INIT('h4)
	) name28970 (
		_w34766_,
		_w34796_,
		_w34797_
	);
	LUT3 #(
		.INIT('h23)
	) name28971 (
		_w34766_,
		_w34795_,
		_w34796_,
		_w34798_
	);
	LUT2 #(
		.INIT('h4)
	) name28972 (
		_w34793_,
		_w34798_,
		_w34799_
	);
	LUT4 #(
		.INIT('h5655)
	) name28973 (
		\u0_L14_reg[10]/P0001 ,
		_w34791_,
		_w34780_,
		_w34799_,
		_w34800_
	);
	LUT4 #(
		.INIT('h0082)
	) name28974 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34801_
	);
	LUT3 #(
		.INIT('h5d)
	) name28975 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w34802_
	);
	LUT4 #(
		.INIT('h0b00)
	) name28976 (
		_w24834_,
		_w24835_,
		_w24832_,
		_w24836_,
		_w34803_
	);
	LUT2 #(
		.INIT('h8)
	) name28977 (
		_w34802_,
		_w34803_,
		_w34804_
	);
	LUT2 #(
		.INIT('h1)
	) name28978 (
		_w24833_,
		_w24832_,
		_w34805_
	);
	LUT4 #(
		.INIT('h0001)
	) name28979 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24832_,
		_w34806_
	);
	LUT2 #(
		.INIT('h8)
	) name28980 (
		_w24833_,
		_w24832_,
		_w34807_
	);
	LUT4 #(
		.INIT('h80c0)
	) name28981 (
		_w24834_,
		_w24833_,
		_w24832_,
		_w24836_,
		_w34808_
	);
	LUT3 #(
		.INIT('h02)
	) name28982 (
		_w24831_,
		_w34808_,
		_w34806_,
		_w34809_
	);
	LUT3 #(
		.INIT('h10)
	) name28983 (
		_w34801_,
		_w34804_,
		_w34809_,
		_w34810_
	);
	LUT4 #(
		.INIT('h59fb)
	) name28984 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34811_
	);
	LUT2 #(
		.INIT('h1)
	) name28985 (
		_w24832_,
		_w34811_,
		_w34812_
	);
	LUT3 #(
		.INIT('h13)
	) name28986 (
		_w24832_,
		_w24831_,
		_w24844_,
		_w34813_
	);
	LUT4 #(
		.INIT('h0034)
	) name28987 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34814_
	);
	LUT4 #(
		.INIT('h0002)
	) name28988 (
		_w24835_,
		_w24833_,
		_w24832_,
		_w24836_,
		_w34815_
	);
	LUT4 #(
		.INIT('h4000)
	) name28989 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34816_
	);
	LUT3 #(
		.INIT('h01)
	) name28990 (
		_w34814_,
		_w34815_,
		_w34816_,
		_w34817_
	);
	LUT3 #(
		.INIT('h40)
	) name28991 (
		_w34812_,
		_w34813_,
		_w34817_,
		_w34818_
	);
	LUT4 #(
		.INIT('h0004)
	) name28992 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34819_
	);
	LUT3 #(
		.INIT('h01)
	) name28993 (
		_w24832_,
		_w34816_,
		_w34819_,
		_w34820_
	);
	LUT4 #(
		.INIT('hf070)
	) name28994 (
		_w24834_,
		_w24833_,
		_w24832_,
		_w24836_,
		_w34821_
	);
	LUT2 #(
		.INIT('h4)
	) name28995 (
		_w24840_,
		_w34821_,
		_w34822_
	);
	LUT2 #(
		.INIT('h1)
	) name28996 (
		_w34820_,
		_w34822_,
		_w34823_
	);
	LUT4 #(
		.INIT('h55a9)
	) name28997 (
		\u0_L14_reg[2]/P0001 ,
		_w34810_,
		_w34818_,
		_w34823_,
		_w34824_
	);
	LUT4 #(
		.INIT('hc963)
	) name28998 (
		decrypt_pad,
		\u0_R14_reg[23]/NET0131 ,
		\u0_uk_K_r14_reg[2]/NET0131 ,
		\u0_uk_K_r14_reg[9]/NET0131 ,
		_w34825_
	);
	LUT4 #(
		.INIT('hc963)
	) name28999 (
		decrypt_pad,
		\u0_R14_reg[21]/NET0131 ,
		\u0_uk_K_r14_reg[22]/NET0131 ,
		\u0_uk_K_r14_reg[29]/NET0131 ,
		_w34826_
	);
	LUT4 #(
		.INIT('hc693)
	) name29000 (
		decrypt_pad,
		\u0_R14_reg[20]/NET0131 ,
		\u0_uk_K_r14_reg[14]/NET0131 ,
		\u0_uk_K_r14_reg[7]/NET0131 ,
		_w34827_
	);
	LUT4 #(
		.INIT('hc963)
	) name29001 (
		decrypt_pad,
		\u0_R14_reg[25]/NET0131 ,
		\u0_uk_K_r14_reg[23]/NET0131 ,
		\u0_uk_K_r14_reg[30]/NET0131 ,
		_w34828_
	);
	LUT4 #(
		.INIT('hc963)
	) name29002 (
		decrypt_pad,
		\u0_R14_reg[22]/P0001 ,
		\u0_uk_K_r14_reg[44]/NET0131 ,
		\u0_uk_K_r14_reg[51]/NET0131 ,
		_w34829_
	);
	LUT4 #(
		.INIT('h45e5)
	) name29003 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34830_
	);
	LUT2 #(
		.INIT('h2)
	) name29004 (
		_w34825_,
		_w34830_,
		_w34831_
	);
	LUT3 #(
		.INIT('h01)
	) name29005 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34832_
	);
	LUT4 #(
		.INIT('h1001)
	) name29006 (
		_w34825_,
		_w34827_,
		_w34828_,
		_w34826_,
		_w34833_
	);
	LUT4 #(
		.INIT('h8000)
	) name29007 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34834_
	);
	LUT4 #(
		.INIT('hc963)
	) name29008 (
		decrypt_pad,
		\u0_R14_reg[24]/NET0131 ,
		\u0_uk_K_r14_reg[28]/NET0131 ,
		\u0_uk_K_r14_reg[35]/P0001 ,
		_w34835_
	);
	LUT3 #(
		.INIT('h01)
	) name29009 (
		_w34834_,
		_w34833_,
		_w34835_,
		_w34836_
	);
	LUT3 #(
		.INIT('h04)
	) name29010 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34837_
	);
	LUT4 #(
		.INIT('hfb5b)
	) name29011 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34838_
	);
	LUT2 #(
		.INIT('h2)
	) name29012 (
		_w34825_,
		_w34838_,
		_w34839_
	);
	LUT4 #(
		.INIT('hfefb)
	) name29013 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34840_
	);
	LUT4 #(
		.INIT('hfb00)
	) name29014 (
		_w34828_,
		_w34826_,
		_w34829_,
		_w34835_,
		_w34841_
	);
	LUT3 #(
		.INIT('h04)
	) name29015 (
		_w34825_,
		_w34827_,
		_w34826_,
		_w34842_
	);
	LUT4 #(
		.INIT('h4000)
	) name29016 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34843_
	);
	LUT4 #(
		.INIT('h0200)
	) name29017 (
		_w34840_,
		_w34842_,
		_w34843_,
		_w34841_,
		_w34844_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name29018 (
		_w34831_,
		_w34836_,
		_w34839_,
		_w34844_,
		_w34845_
	);
	LUT4 #(
		.INIT('h0008)
	) name29019 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34846_
	);
	LUT2 #(
		.INIT('h4)
	) name29020 (
		_w34825_,
		_w34846_,
		_w34847_
	);
	LUT4 #(
		.INIT('h0020)
	) name29021 (
		_w34825_,
		_w34827_,
		_w34828_,
		_w34826_,
		_w34848_
	);
	LUT2 #(
		.INIT('h1)
	) name29022 (
		_w34825_,
		_w34829_,
		_w34849_
	);
	LUT3 #(
		.INIT('h20)
	) name29023 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34850_
	);
	LUT4 #(
		.INIT('hcedf)
	) name29024 (
		_w34825_,
		_w34829_,
		_w34837_,
		_w34850_,
		_w34851_
	);
	LUT2 #(
		.INIT('h4)
	) name29025 (
		_w34847_,
		_w34851_,
		_w34852_
	);
	LUT3 #(
		.INIT('h65)
	) name29026 (
		\u0_L14_reg[19]/P0001 ,
		_w34845_,
		_w34852_,
		_w34853_
	);
	LUT3 #(
		.INIT('h40)
	) name29027 (
		_w34827_,
		_w34826_,
		_w34829_,
		_w34854_
	);
	LUT4 #(
		.INIT('h2740)
	) name29028 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34855_
	);
	LUT3 #(
		.INIT('h01)
	) name29029 (
		_w34825_,
		_w34846_,
		_w34855_,
		_w34856_
	);
	LUT4 #(
		.INIT('h0002)
	) name29030 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34857_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name29031 (
		_w34825_,
		_w34827_,
		_w34828_,
		_w34826_,
		_w34858_
	);
	LUT3 #(
		.INIT('h10)
	) name29032 (
		_w34854_,
		_w34857_,
		_w34858_,
		_w34859_
	);
	LUT3 #(
		.INIT('ha8)
	) name29033 (
		_w34835_,
		_w34856_,
		_w34859_,
		_w34860_
	);
	LUT4 #(
		.INIT('h0020)
	) name29034 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34861_
	);
	LUT3 #(
		.INIT('h01)
	) name29035 (
		_w34835_,
		_w34848_,
		_w34861_,
		_w34862_
	);
	LUT4 #(
		.INIT('h0822)
	) name29036 (
		_w34825_,
		_w34827_,
		_w34826_,
		_w34829_,
		_w34863_
	);
	LUT4 #(
		.INIT('h0004)
	) name29037 (
		_w34825_,
		_w34827_,
		_w34828_,
		_w34829_,
		_w34864_
	);
	LUT4 #(
		.INIT('h0800)
	) name29038 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34865_
	);
	LUT4 #(
		.INIT('h1040)
	) name29039 (
		_w34825_,
		_w34827_,
		_w34826_,
		_w34829_,
		_w34866_
	);
	LUT4 #(
		.INIT('h0001)
	) name29040 (
		_w34864_,
		_w34865_,
		_w34866_,
		_w34863_,
		_w34867_
	);
	LUT2 #(
		.INIT('h8)
	) name29041 (
		_w34862_,
		_w34867_,
		_w34868_
	);
	LUT4 #(
		.INIT('h0010)
	) name29042 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34869_
	);
	LUT4 #(
		.INIT('h77ef)
	) name29043 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34870_
	);
	LUT2 #(
		.INIT('h2)
	) name29044 (
		_w34825_,
		_w34870_,
		_w34871_
	);
	LUT2 #(
		.INIT('h8)
	) name29045 (
		_w34832_,
		_w34849_,
		_w34872_
	);
	LUT3 #(
		.INIT('h02)
	) name29046 (
		_w34851_,
		_w34872_,
		_w34871_,
		_w34873_
	);
	LUT4 #(
		.INIT('h56aa)
	) name29047 (
		\u0_L14_reg[11]/P0001 ,
		_w34860_,
		_w34868_,
		_w34873_,
		_w34874_
	);
	LUT4 #(
		.INIT('hbfae)
	) name29048 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34875_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name29049 (
		_w24834_,
		_w24833_,
		_w24832_,
		_w24836_,
		_w34876_
	);
	LUT3 #(
		.INIT('h40)
	) name29050 (
		_w24845_,
		_w34876_,
		_w34875_,
		_w34877_
	);
	LUT4 #(
		.INIT('h1000)
	) name29051 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34878_
	);
	LUT4 #(
		.INIT('h7d00)
	) name29052 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24832_,
		_w34879_
	);
	LUT2 #(
		.INIT('h4)
	) name29053 (
		_w34878_,
		_w34879_,
		_w34880_
	);
	LUT4 #(
		.INIT('h0400)
	) name29054 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34881_
	);
	LUT4 #(
		.INIT('h0008)
	) name29055 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34882_
	);
	LUT4 #(
		.INIT('hf070)
	) name29056 (
		_w24834_,
		_w24832_,
		_w24831_,
		_w24836_,
		_w34883_
	);
	LUT3 #(
		.INIT('h10)
	) name29057 (
		_w34882_,
		_w34881_,
		_w34883_,
		_w34884_
	);
	LUT3 #(
		.INIT('he0)
	) name29058 (
		_w34877_,
		_w34880_,
		_w34884_,
		_w34885_
	);
	LUT3 #(
		.INIT('h02)
	) name29059 (
		_w24834_,
		_w24835_,
		_w24836_,
		_w34886_
	);
	LUT4 #(
		.INIT('h5b59)
	) name29060 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34887_
	);
	LUT4 #(
		.INIT('h4e5f)
	) name29061 (
		_w24832_,
		_w24839_,
		_w34875_,
		_w34887_,
		_w34888_
	);
	LUT3 #(
		.INIT('h0b)
	) name29062 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w34889_
	);
	LUT4 #(
		.INIT('h0900)
	) name29063 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w34890_
	);
	LUT3 #(
		.INIT('h01)
	) name29064 (
		_w24831_,
		_w24845_,
		_w34890_,
		_w34891_
	);
	LUT2 #(
		.INIT('h4)
	) name29065 (
		_w34888_,
		_w34891_,
		_w34892_
	);
	LUT3 #(
		.INIT('ha9)
	) name29066 (
		\u0_L14_reg[28]/P0001 ,
		_w34885_,
		_w34892_,
		_w34893_
	);
	LUT2 #(
		.INIT('h1)
	) name29067 (
		_w34763_,
		_w34795_,
		_w34894_
	);
	LUT4 #(
		.INIT('h0100)
	) name29068 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w34765_,
		_w34895_
	);
	LUT3 #(
		.INIT('h2e)
	) name29069 (
		_w34766_,
		_w34767_,
		_w34765_,
		_w34896_
	);
	LUT3 #(
		.INIT('h31)
	) name29070 (
		_w34781_,
		_w34895_,
		_w34896_,
		_w34897_
	);
	LUT4 #(
		.INIT('hdf13)
	) name29071 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34898_
	);
	LUT3 #(
		.INIT('hc8)
	) name29072 (
		_w34765_,
		_w34775_,
		_w34898_,
		_w34899_
	);
	LUT3 #(
		.INIT('h80)
	) name29073 (
		_w34894_,
		_w34897_,
		_w34899_,
		_w34900_
	);
	LUT2 #(
		.INIT('h4)
	) name29074 (
		_w34782_,
		_w34763_,
		_w34901_
	);
	LUT4 #(
		.INIT('h0400)
	) name29075 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w34765_,
		_w34902_
	);
	LUT3 #(
		.INIT('h01)
	) name29076 (
		_w34786_,
		_w34796_,
		_w34902_,
		_w34903_
	);
	LUT2 #(
		.INIT('h8)
	) name29077 (
		_w34766_,
		_w34776_,
		_w34904_
	);
	LUT3 #(
		.INIT('h02)
	) name29078 (
		_w34764_,
		_w34766_,
		_w34767_,
		_w34905_
	);
	LUT3 #(
		.INIT('hed)
	) name29079 (
		_w34764_,
		_w34766_,
		_w34767_,
		_w34906_
	);
	LUT4 #(
		.INIT('h0012)
	) name29080 (
		_w34764_,
		_w34766_,
		_w34767_,
		_w34765_,
		_w34907_
	);
	LUT3 #(
		.INIT('h07)
	) name29081 (
		_w34766_,
		_w34776_,
		_w34907_,
		_w34908_
	);
	LUT3 #(
		.INIT('h80)
	) name29082 (
		_w34901_,
		_w34903_,
		_w34908_,
		_w34909_
	);
	LUT4 #(
		.INIT('h0020)
	) name29083 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w34910_
	);
	LUT4 #(
		.INIT('heee4)
	) name29084 (
		_w34765_,
		_w34786_,
		_w34774_,
		_w34910_,
		_w34911_
	);
	LUT2 #(
		.INIT('h1)
	) name29085 (
		_w34797_,
		_w34911_,
		_w34912_
	);
	LUT4 #(
		.INIT('ha955)
	) name29086 (
		\u0_L14_reg[20]/P0001 ,
		_w34900_,
		_w34909_,
		_w34912_,
		_w34913_
	);
	LUT4 #(
		.INIT('hc693)
	) name29087 (
		decrypt_pad,
		\u0_R14_reg[24]/NET0131 ,
		\u0_uk_K_r14_reg[2]/NET0131 ,
		\u0_uk_K_r14_reg[50]/NET0131 ,
		_w34914_
	);
	LUT4 #(
		.INIT('hc963)
	) name29088 (
		decrypt_pad,
		\u0_R14_reg[25]/NET0131 ,
		\u0_uk_K_r14_reg[30]/NET0131 ,
		\u0_uk_K_r14_reg[37]/NET0131 ,
		_w34915_
	);
	LUT2 #(
		.INIT('h6)
	) name29089 (
		_w34914_,
		_w34915_,
		_w34916_
	);
	LUT4 #(
		.INIT('hc963)
	) name29090 (
		decrypt_pad,
		\u0_R14_reg[26]/P0001 ,
		\u0_uk_K_r14_reg[15]/NET0131 ,
		\u0_uk_K_r14_reg[22]/NET0131 ,
		_w34917_
	);
	LUT4 #(
		.INIT('hc693)
	) name29091 (
		decrypt_pad,
		\u0_R14_reg[27]/P0001 ,
		\u0_uk_K_r14_reg[0]/NET0131 ,
		\u0_uk_K_r14_reg[52]/NET0131 ,
		_w34918_
	);
	LUT4 #(
		.INIT('hc963)
	) name29092 (
		decrypt_pad,
		\u0_R14_reg[29]/NET0131 ,
		\u0_uk_K_r14_reg[31]/NET0131 ,
		\u0_uk_K_r14_reg[38]/NET0131 ,
		_w34919_
	);
	LUT2 #(
		.INIT('h2)
	) name29093 (
		_w34919_,
		_w34914_,
		_w34920_
	);
	LUT4 #(
		.INIT('hf100)
	) name29094 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34918_,
		_w34921_
	);
	LUT2 #(
		.INIT('h4)
	) name29095 (
		_w34916_,
		_w34921_,
		_w34922_
	);
	LUT4 #(
		.INIT('h0008)
	) name29096 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w34923_
	);
	LUT4 #(
		.INIT('h0660)
	) name29097 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w34924_
	);
	LUT4 #(
		.INIT('hc963)
	) name29098 (
		decrypt_pad,
		\u0_R14_reg[28]/NET0131 ,
		\u0_uk_K_r14_reg[35]/P0001 ,
		\u0_uk_K_r14_reg[42]/P0001 ,
		_w34925_
	);
	LUT4 #(
		.INIT('h5100)
	) name29099 (
		_w34924_,
		_w34923_,
		_w34918_,
		_w34925_,
		_w34926_
	);
	LUT2 #(
		.INIT('h4)
	) name29100 (
		_w34922_,
		_w34926_,
		_w34927_
	);
	LUT4 #(
		.INIT('hf632)
	) name29101 (
		_w34919_,
		_w34917_,
		_w34915_,
		_w34918_,
		_w34928_
	);
	LUT2 #(
		.INIT('h2)
	) name29102 (
		_w34914_,
		_w34928_,
		_w34929_
	);
	LUT3 #(
		.INIT('h47)
	) name29103 (
		_w34917_,
		_w34915_,
		_w34918_,
		_w34930_
	);
	LUT3 #(
		.INIT('h51)
	) name29104 (
		_w34925_,
		_w34920_,
		_w34930_,
		_w34931_
	);
	LUT3 #(
		.INIT('h09)
	) name29105 (
		_w34919_,
		_w34915_,
		_w34918_,
		_w34932_
	);
	LUT4 #(
		.INIT('h0104)
	) name29106 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w34933_
	);
	LUT2 #(
		.INIT('h1)
	) name29107 (
		_w34932_,
		_w34933_,
		_w34934_
	);
	LUT3 #(
		.INIT('h40)
	) name29108 (
		_w34929_,
		_w34931_,
		_w34934_,
		_w34935_
	);
	LUT3 #(
		.INIT('ha9)
	) name29109 (
		\u0_L14_reg[12]/P0001 ,
		_w34927_,
		_w34935_,
		_w34936_
	);
	LUT4 #(
		.INIT('hcc9d)
	) name29110 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w34937_
	);
	LUT2 #(
		.INIT('h2)
	) name29111 (
		_w24726_,
		_w34937_,
		_w34938_
	);
	LUT4 #(
		.INIT('h5001)
	) name29112 (
		_w24726_,
		_w24728_,
		_w24727_,
		_w24730_,
		_w34939_
	);
	LUT4 #(
		.INIT('h0002)
	) name29113 (
		_w24725_,
		_w24749_,
		_w24748_,
		_w34939_,
		_w34940_
	);
	LUT4 #(
		.INIT('h5554)
	) name29114 (
		_w24726_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w34941_
	);
	LUT4 #(
		.INIT('h0220)
	) name29115 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w34942_
	);
	LUT4 #(
		.INIT('h2a8a)
	) name29116 (
		_w24726_,
		_w24728_,
		_w24727_,
		_w24729_,
		_w34943_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name29117 (
		_w24822_,
		_w34941_,
		_w34942_,
		_w34943_,
		_w34944_
	);
	LUT4 #(
		.INIT('h1000)
	) name29118 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w34945_
	);
	LUT3 #(
		.INIT('h01)
	) name29119 (
		_w24725_,
		_w24731_,
		_w34945_,
		_w34946_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name29120 (
		_w34938_,
		_w34940_,
		_w34944_,
		_w34946_,
		_w34947_
	);
	LUT2 #(
		.INIT('h6)
	) name29121 (
		\u0_L14_reg[17]/P0001 ,
		_w34947_,
		_w34948_
	);
	LUT4 #(
		.INIT('hff8a)
	) name29122 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34949_
	);
	LUT2 #(
		.INIT('h1)
	) name29123 (
		_w34825_,
		_w34949_,
		_w34950_
	);
	LUT4 #(
		.INIT('h0080)
	) name29124 (
		_w34825_,
		_w34827_,
		_w34828_,
		_w34829_,
		_w34951_
	);
	LUT3 #(
		.INIT('h02)
	) name29125 (
		_w34835_,
		_w34869_,
		_w34951_,
		_w34952_
	);
	LUT4 #(
		.INIT('hd79b)
	) name29126 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34953_
	);
	LUT4 #(
		.INIT('h0301)
	) name29127 (
		_w34825_,
		_w34835_,
		_w34857_,
		_w34953_,
		_w34954_
	);
	LUT3 #(
		.INIT('h0b)
	) name29128 (
		_w34950_,
		_w34952_,
		_w34954_,
		_w34955_
	);
	LUT4 #(
		.INIT('h0400)
	) name29129 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34956_
	);
	LUT4 #(
		.INIT('heb67)
	) name29130 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34957_
	);
	LUT3 #(
		.INIT('h01)
	) name29131 (
		_w34827_,
		_w34828_,
		_w34829_,
		_w34958_
	);
	LUT4 #(
		.INIT('h5501)
	) name29132 (
		_w34825_,
		_w34835_,
		_w34957_,
		_w34958_,
		_w34959_
	);
	LUT4 #(
		.INIT('h2802)
	) name29133 (
		_w34825_,
		_w34827_,
		_w34828_,
		_w34826_,
		_w34960_
	);
	LUT4 #(
		.INIT('h4004)
	) name29134 (
		_w34825_,
		_w34827_,
		_w34828_,
		_w34826_,
		_w34961_
	);
	LUT3 #(
		.INIT('h80)
	) name29135 (
		_w34828_,
		_w34826_,
		_w34835_,
		_w34962_
	);
	LUT4 #(
		.INIT('haaa8)
	) name29136 (
		_w34829_,
		_w34961_,
		_w34960_,
		_w34962_,
		_w34963_
	);
	LUT2 #(
		.INIT('h1)
	) name29137 (
		_w34959_,
		_w34963_,
		_w34964_
	);
	LUT3 #(
		.INIT('h65)
	) name29138 (
		\u0_L14_reg[4]/P0001 ,
		_w34955_,
		_w34964_,
		_w34965_
	);
	LUT4 #(
		.INIT('h9faf)
	) name29139 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34966_
	);
	LUT2 #(
		.INIT('h2)
	) name29140 (
		_w34825_,
		_w34966_,
		_w34967_
	);
	LUT4 #(
		.INIT('h66fe)
	) name29141 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34968_
	);
	LUT2 #(
		.INIT('h1)
	) name29142 (
		_w34825_,
		_w34968_,
		_w34969_
	);
	LUT3 #(
		.INIT('h02)
	) name29143 (
		_w34840_,
		_w34864_,
		_w34865_,
		_w34970_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name29144 (
		_w34835_,
		_w34967_,
		_w34969_,
		_w34970_,
		_w34971_
	);
	LUT4 #(
		.INIT('h6d7c)
	) name29145 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34972_
	);
	LUT4 #(
		.INIT('h3032)
	) name29146 (
		_w34825_,
		_w34835_,
		_w34956_,
		_w34972_,
		_w34973_
	);
	LUT4 #(
		.INIT('hdf27)
	) name29147 (
		_w34827_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34974_
	);
	LUT2 #(
		.INIT('h1)
	) name29148 (
		_w34825_,
		_w34835_,
		_w34975_
	);
	LUT4 #(
		.INIT('h0080)
	) name29149 (
		_w34825_,
		_w34828_,
		_w34826_,
		_w34829_,
		_w34976_
	);
	LUT4 #(
		.INIT('h1011)
	) name29150 (
		_w34857_,
		_w34976_,
		_w34974_,
		_w34975_,
		_w34977_
	);
	LUT2 #(
		.INIT('h4)
	) name29151 (
		_w34973_,
		_w34977_,
		_w34978_
	);
	LUT3 #(
		.INIT('h9a)
	) name29152 (
		\u0_L14_reg[29]/P0001 ,
		_w34971_,
		_w34978_,
		_w34979_
	);
	LUT4 #(
		.INIT('h1fb3)
	) name29153 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w34980_
	);
	LUT2 #(
		.INIT('h2)
	) name29154 (
		_w24705_,
		_w34980_,
		_w34981_
	);
	LUT4 #(
		.INIT('hf7dd)
	) name29155 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w34982_
	);
	LUT2 #(
		.INIT('h1)
	) name29156 (
		_w24705_,
		_w34982_,
		_w34983_
	);
	LUT4 #(
		.INIT('h2100)
	) name29157 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w34984_
	);
	LUT4 #(
		.INIT('h0004)
	) name29158 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w34985_
	);
	LUT3 #(
		.INIT('h02)
	) name29159 (
		_w24712_,
		_w34985_,
		_w34984_,
		_w34986_
	);
	LUT3 #(
		.INIT('h10)
	) name29160 (
		_w34983_,
		_w34981_,
		_w34986_,
		_w34987_
	);
	LUT3 #(
		.INIT('h75)
	) name29161 (
		_w24700_,
		_w24697_,
		_w24705_,
		_w34988_
	);
	LUT2 #(
		.INIT('h2)
	) name29162 (
		_w24701_,
		_w24698_,
		_w34989_
	);
	LUT2 #(
		.INIT('h4)
	) name29163 (
		_w34988_,
		_w34989_,
		_w34990_
	);
	LUT4 #(
		.INIT('h00bf)
	) name29164 (
		_w24700_,
		_w24697_,
		_w24698_,
		_w24712_,
		_w34991_
	);
	LUT4 #(
		.INIT('h0040)
	) name29165 (
		_w24700_,
		_w24701_,
		_w24698_,
		_w24705_,
		_w34992_
	);
	LUT3 #(
		.INIT('h10)
	) name29166 (
		_w24783_,
		_w34992_,
		_w34991_,
		_w34993_
	);
	LUT4 #(
		.INIT('h0201)
	) name29167 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w34994_
	);
	LUT4 #(
		.INIT('hd5df)
	) name29168 (
		_w24700_,
		_w24701_,
		_w24697_,
		_w24698_,
		_w34995_
	);
	LUT3 #(
		.INIT('h31)
	) name29169 (
		_w24705_,
		_w34994_,
		_w34995_,
		_w34996_
	);
	LUT3 #(
		.INIT('h40)
	) name29170 (
		_w34990_,
		_w34993_,
		_w34996_,
		_w34997_
	);
	LUT4 #(
		.INIT('h0100)
	) name29171 (
		_w24700_,
		_w24697_,
		_w24698_,
		_w24705_,
		_w34998_
	);
	LUT3 #(
		.INIT('h07)
	) name29172 (
		_w24709_,
		_w24713_,
		_w34998_,
		_w34999_
	);
	LUT4 #(
		.INIT('ha955)
	) name29173 (
		\u0_L14_reg[21]/P0001 ,
		_w34987_,
		_w34997_,
		_w34999_,
		_w35000_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name29174 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w35001_
	);
	LUT4 #(
		.INIT('hebed)
	) name29175 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w35002_
	);
	LUT4 #(
		.INIT('h0515)
	) name29176 (
		_w24832_,
		_w24831_,
		_w35001_,
		_w35002_,
		_w35003_
	);
	LUT4 #(
		.INIT('h74f6)
	) name29177 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w35004_
	);
	LUT2 #(
		.INIT('h2)
	) name29178 (
		_w24832_,
		_w35004_,
		_w35005_
	);
	LUT3 #(
		.INIT('h04)
	) name29179 (
		_w24834_,
		_w24835_,
		_w24836_,
		_w35006_
	);
	LUT2 #(
		.INIT('h4)
	) name29180 (
		_w34805_,
		_w35006_,
		_w35007_
	);
	LUT3 #(
		.INIT('h15)
	) name29181 (
		_w24831_,
		_w34807_,
		_w34886_,
		_w35008_
	);
	LUT3 #(
		.INIT('h10)
	) name29182 (
		_w35005_,
		_w35007_,
		_w35008_,
		_w35009_
	);
	LUT3 #(
		.INIT('hcd)
	) name29183 (
		_w24835_,
		_w24832_,
		_w24836_,
		_w35010_
	);
	LUT4 #(
		.INIT('h2202)
	) name29184 (
		_w24831_,
		_w24849_,
		_w34889_,
		_w35010_,
		_w35011_
	);
	LUT4 #(
		.INIT('hbbfc)
	) name29185 (
		_w24834_,
		_w24835_,
		_w24833_,
		_w24836_,
		_w35012_
	);
	LUT2 #(
		.INIT('h2)
	) name29186 (
		_w24832_,
		_w35012_,
		_w35013_
	);
	LUT3 #(
		.INIT('h10)
	) name29187 (
		_w34815_,
		_w34816_,
		_w35001_,
		_w35014_
	);
	LUT3 #(
		.INIT('h40)
	) name29188 (
		_w35013_,
		_w35011_,
		_w35014_,
		_w35015_
	);
	LUT4 #(
		.INIT('h999a)
	) name29189 (
		\u0_L14_reg[13]/P0001 ,
		_w35003_,
		_w35009_,
		_w35015_,
		_w35016_
	);
	LUT4 #(
		.INIT('hcffb)
	) name29190 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34918_,
		_w35017_
	);
	LUT2 #(
		.INIT('h1)
	) name29191 (
		_w34915_,
		_w35017_,
		_w35018_
	);
	LUT2 #(
		.INIT('h9)
	) name29192 (
		_w34917_,
		_w34914_,
		_w35019_
	);
	LUT3 #(
		.INIT('h8a)
	) name29193 (
		_w34919_,
		_w34915_,
		_w34918_,
		_w35020_
	);
	LUT2 #(
		.INIT('h8)
	) name29194 (
		_w35019_,
		_w35020_,
		_w35021_
	);
	LUT3 #(
		.INIT('h2e)
	) name29195 (
		_w34919_,
		_w34917_,
		_w34915_,
		_w35022_
	);
	LUT2 #(
		.INIT('h2)
	) name29196 (
		_w34914_,
		_w34918_,
		_w35023_
	);
	LUT3 #(
		.INIT('h45)
	) name29197 (
		_w34925_,
		_w35022_,
		_w35023_,
		_w35024_
	);
	LUT3 #(
		.INIT('h10)
	) name29198 (
		_w35018_,
		_w35021_,
		_w35024_,
		_w35025_
	);
	LUT4 #(
		.INIT('h0009)
	) name29199 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35026_
	);
	LUT2 #(
		.INIT('h2)
	) name29200 (
		_w34925_,
		_w35026_,
		_w35027_
	);
	LUT3 #(
		.INIT('h8b)
	) name29201 (
		_w34917_,
		_w34914_,
		_w34915_,
		_w35028_
	);
	LUT4 #(
		.INIT('h002a)
	) name29202 (
		_w34919_,
		_w34914_,
		_w34915_,
		_w34918_,
		_w35029_
	);
	LUT4 #(
		.INIT('hc800)
	) name29203 (
		_w34917_,
		_w34914_,
		_w34915_,
		_w34918_,
		_w35030_
	);
	LUT4 #(
		.INIT('h45cf)
	) name29204 (
		_w35022_,
		_w35028_,
		_w35029_,
		_w35030_,
		_w35031_
	);
	LUT2 #(
		.INIT('h8)
	) name29205 (
		_w35027_,
		_w35031_,
		_w35032_
	);
	LUT4 #(
		.INIT('hfba7)
	) name29206 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35033_
	);
	LUT4 #(
		.INIT('h0090)
	) name29207 (
		_w34917_,
		_w34914_,
		_w34915_,
		_w34918_,
		_w35034_
	);
	LUT4 #(
		.INIT('h0100)
	) name29208 (
		_w34919_,
		_w34917_,
		_w34915_,
		_w34918_,
		_w35035_
	);
	LUT4 #(
		.INIT('h0301)
	) name29209 (
		_w34918_,
		_w35034_,
		_w35035_,
		_w35033_,
		_w35036_
	);
	LUT4 #(
		.INIT('ha955)
	) name29210 (
		\u0_L14_reg[22]/P0001 ,
		_w35025_,
		_w35032_,
		_w35036_,
		_w35037_
	);
	LUT4 #(
		.INIT('h9d35)
	) name29211 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35038_
	);
	LUT2 #(
		.INIT('h2)
	) name29212 (
		_w24792_,
		_w35038_,
		_w35039_
	);
	LUT4 #(
		.INIT('hf7d6)
	) name29213 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24792_,
		_w35040_
	);
	LUT2 #(
		.INIT('h1)
	) name29214 (
		_w24796_,
		_w35040_,
		_w35041_
	);
	LUT3 #(
		.INIT('h80)
	) name29215 (
		_w24794_,
		_w24795_,
		_w24796_,
		_w35042_
	);
	LUT4 #(
		.INIT('hfbbf)
	) name29216 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35043_
	);
	LUT3 #(
		.INIT('h70)
	) name29217 (
		_w24814_,
		_w35042_,
		_w35043_,
		_w35044_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name29218 (
		_w24791_,
		_w35041_,
		_w35039_,
		_w35044_,
		_w35045_
	);
	LUT4 #(
		.INIT('had79)
	) name29219 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35046_
	);
	LUT4 #(
		.INIT('h76ce)
	) name29220 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35047_
	);
	LUT4 #(
		.INIT('hf7ef)
	) name29221 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35048_
	);
	LUT4 #(
		.INIT('he400)
	) name29222 (
		_w24792_,
		_w35046_,
		_w35047_,
		_w35048_,
		_w35049_
	);
	LUT4 #(
		.INIT('h1200)
	) name29223 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35050_
	);
	LUT4 #(
		.INIT('hfebf)
	) name29224 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35051_
	);
	LUT3 #(
		.INIT('hb1)
	) name29225 (
		_w24792_,
		_w35050_,
		_w35051_,
		_w35052_
	);
	LUT3 #(
		.INIT('he0)
	) name29226 (
		_w24791_,
		_w35049_,
		_w35052_,
		_w35053_
	);
	LUT3 #(
		.INIT('h65)
	) name29227 (
		\u0_L14_reg[14]/P0001 ,
		_w35045_,
		_w35053_,
		_w35054_
	);
	LUT4 #(
		.INIT('h2814)
	) name29228 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w35055_
	);
	LUT3 #(
		.INIT('h01)
	) name29229 (
		_w24902_,
		_w24916_,
		_w35055_,
		_w35056_
	);
	LUT2 #(
		.INIT('h4)
	) name29230 (
		_w24860_,
		_w24909_,
		_w35057_
	);
	LUT4 #(
		.INIT('h5155)
	) name29231 (
		_w24854_,
		_w24891_,
		_w35057_,
		_w35056_,
		_w35058_
	);
	LUT4 #(
		.INIT('h995d)
	) name29232 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w35059_
	);
	LUT4 #(
		.INIT('hdfde)
	) name29233 (
		_w24857_,
		_w24855_,
		_w24856_,
		_w24858_,
		_w35060_
	);
	LUT4 #(
		.INIT('h08aa)
	) name29234 (
		_w24860_,
		_w24854_,
		_w35059_,
		_w35060_,
		_w35061_
	);
	LUT3 #(
		.INIT('h0d)
	) name29235 (
		_w24855_,
		_w24856_,
		_w24858_,
		_w35062_
	);
	LUT4 #(
		.INIT('h0900)
	) name29236 (
		_w24857_,
		_w24855_,
		_w24860_,
		_w24854_,
		_w35063_
	);
	LUT4 #(
		.INIT('h7077)
	) name29237 (
		_w24864_,
		_w24882_,
		_w35062_,
		_w35063_,
		_w35064_
	);
	LUT2 #(
		.INIT('h4)
	) name29238 (
		_w35061_,
		_w35064_,
		_w35065_
	);
	LUT3 #(
		.INIT('h65)
	) name29239 (
		\u0_L14_reg[6]/P0001 ,
		_w35058_,
		_w35065_,
		_w35066_
	);
	LUT3 #(
		.INIT('hbe)
	) name29240 (
		_w24727_,
		_w24729_,
		_w24730_,
		_w35067_
	);
	LUT3 #(
		.INIT('h02)
	) name29241 (
		_w24728_,
		_w34941_,
		_w35067_,
		_w35068_
	);
	LUT4 #(
		.INIT('hf73f)
	) name29242 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w35069_
	);
	LUT3 #(
		.INIT('h31)
	) name29243 (
		_w24726_,
		_w24736_,
		_w35069_,
		_w35070_
	);
	LUT3 #(
		.INIT('h45)
	) name29244 (
		_w24725_,
		_w35068_,
		_w35070_,
		_w35071_
	);
	LUT4 #(
		.INIT('hfbdc)
	) name29245 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w35072_
	);
	LUT4 #(
		.INIT('h6ff5)
	) name29246 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w35073_
	);
	LUT4 #(
		.INIT('h0133)
	) name29247 (
		_w24725_,
		_w24726_,
		_w35072_,
		_w35073_,
		_w35074_
	);
	LUT4 #(
		.INIT('hacaf)
	) name29248 (
		_w24728_,
		_w24727_,
		_w24729_,
		_w24730_,
		_w35075_
	);
	LUT2 #(
		.INIT('h2)
	) name29249 (
		_w24726_,
		_w35075_,
		_w35076_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name29250 (
		_w24726_,
		_w24728_,
		_w24729_,
		_w24730_,
		_w35077_
	);
	LUT2 #(
		.INIT('h2)
	) name29251 (
		_w24727_,
		_w35077_,
		_w35078_
	);
	LUT3 #(
		.INIT('h10)
	) name29252 (
		_w24728_,
		_w24727_,
		_w24730_,
		_w35079_
	);
	LUT3 #(
		.INIT('hc4)
	) name29253 (
		_w24726_,
		_w24728_,
		_w24730_,
		_w35080_
	);
	LUT3 #(
		.INIT('h31)
	) name29254 (
		_w24821_,
		_w35079_,
		_w35080_,
		_w35081_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name29255 (
		_w24725_,
		_w35078_,
		_w35076_,
		_w35081_,
		_w35082_
	);
	LUT3 #(
		.INIT('h13)
	) name29256 (
		_w24734_,
		_w24756_,
		_w24735_,
		_w35083_
	);
	LUT4 #(
		.INIT('h0100)
	) name29257 (
		_w35082_,
		_w35074_,
		_w35071_,
		_w35083_,
		_w35084_
	);
	LUT2 #(
		.INIT('h9)
	) name29258 (
		\u0_L14_reg[31]/P0001 ,
		_w35084_,
		_w35085_
	);
	LUT4 #(
		.INIT('h010c)
	) name29259 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35086_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name29260 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35087_
	);
	LUT3 #(
		.INIT('h01)
	) name29261 (
		_w34918_,
		_w35087_,
		_w35086_,
		_w35088_
	);
	LUT4 #(
		.INIT('h4800)
	) name29262 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35089_
	);
	LUT3 #(
		.INIT('h08)
	) name29263 (
		_w34919_,
		_w34914_,
		_w34915_,
		_w35090_
	);
	LUT4 #(
		.INIT('hb77f)
	) name29264 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35091_
	);
	LUT3 #(
		.INIT('h21)
	) name29265 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w35092_
	);
	LUT4 #(
		.INIT('h2120)
	) name29266 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35093_
	);
	LUT3 #(
		.INIT('h4c)
	) name29267 (
		_w34918_,
		_w35091_,
		_w35093_,
		_w35094_
	);
	LUT3 #(
		.INIT('h8a)
	) name29268 (
		_w34925_,
		_w35088_,
		_w35094_,
		_w35095_
	);
	LUT2 #(
		.INIT('h4)
	) name29269 (
		_w34918_,
		_w34925_,
		_w35096_
	);
	LUT4 #(
		.INIT('h0004)
	) name29270 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35097_
	);
	LUT4 #(
		.INIT('h0f04)
	) name29271 (
		_w34918_,
		_w35093_,
		_w35096_,
		_w35097_,
		_w35098_
	);
	LUT2 #(
		.INIT('h1)
	) name29272 (
		_w34918_,
		_w35091_,
		_w35099_
	);
	LUT2 #(
		.INIT('h2)
	) name29273 (
		_w34918_,
		_w34925_,
		_w35100_
	);
	LUT4 #(
		.INIT('h0100)
	) name29274 (
		_w35089_,
		_w35090_,
		_w35092_,
		_w35100_,
		_w35101_
	);
	LUT3 #(
		.INIT('h01)
	) name29275 (
		_w35099_,
		_w35098_,
		_w35101_,
		_w35102_
	);
	LUT3 #(
		.INIT('h65)
	) name29276 (
		\u0_L14_reg[7]/P0001 ,
		_w35095_,
		_w35102_,
		_w35103_
	);
	LUT4 #(
		.INIT('hfa6d)
	) name29277 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35104_
	);
	LUT4 #(
		.INIT('h4000)
	) name29278 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35105_
	);
	LUT4 #(
		.INIT('h9dba)
	) name29279 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35106_
	);
	LUT4 #(
		.INIT('h3120)
	) name29280 (
		_w34918_,
		_w35105_,
		_w35106_,
		_w35104_,
		_w35107_
	);
	LUT2 #(
		.INIT('h2)
	) name29281 (
		_w34925_,
		_w35107_,
		_w35108_
	);
	LUT3 #(
		.INIT('h10)
	) name29282 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w35109_
	);
	LUT4 #(
		.INIT('hef4f)
	) name29283 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35110_
	);
	LUT2 #(
		.INIT('h2)
	) name29284 (
		_w34918_,
		_w35110_,
		_w35111_
	);
	LUT4 #(
		.INIT('h6bff)
	) name29285 (
		_w34919_,
		_w34917_,
		_w34914_,
		_w34915_,
		_w35112_
	);
	LUT3 #(
		.INIT('hd0)
	) name29286 (
		_w34932_,
		_w35109_,
		_w35112_,
		_w35113_
	);
	LUT4 #(
		.INIT('h00e0)
	) name29287 (
		_w34919_,
		_w34917_,
		_w34915_,
		_w34918_,
		_w35114_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name29288 (
		_w34923_,
		_w35019_,
		_w35096_,
		_w35114_,
		_w35115_
	);
	LUT4 #(
		.INIT('hba00)
	) name29289 (
		_w34925_,
		_w35111_,
		_w35113_,
		_w35115_,
		_w35116_
	);
	LUT3 #(
		.INIT('h65)
	) name29290 (
		\u0_L14_reg[32]/P0001 ,
		_w35108_,
		_w35116_,
		_w35117_
	);
	LUT4 #(
		.INIT('h2022)
	) name29291 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35118_
	);
	LUT2 #(
		.INIT('h2)
	) name29292 (
		_w34750_,
		_w35118_,
		_w35119_
	);
	LUT3 #(
		.INIT('h02)
	) name29293 (
		_w24792_,
		_w24802_,
		_w34752_,
		_w35120_
	);
	LUT4 #(
		.INIT('hbecf)
	) name29294 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35121_
	);
	LUT4 #(
		.INIT('h0155)
	) name29295 (
		_w24791_,
		_w35119_,
		_w35120_,
		_w35121_,
		_w35122_
	);
	LUT4 #(
		.INIT('hf7f6)
	) name29296 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35123_
	);
	LUT3 #(
		.INIT('h02)
	) name29297 (
		_w24795_,
		_w24796_,
		_w24792_,
		_w35124_
	);
	LUT4 #(
		.INIT('h0031)
	) name29298 (
		_w24792_,
		_w35050_,
		_w35123_,
		_w35124_,
		_w35125_
	);
	LUT4 #(
		.INIT('haddf)
	) name29299 (
		_w24794_,
		_w24795_,
		_w24793_,
		_w24796_,
		_w35126_
	);
	LUT3 #(
		.INIT('hb1)
	) name29300 (
		_w24792_,
		_w24813_,
		_w35126_,
		_w35127_
	);
	LUT3 #(
		.INIT('hd0)
	) name29301 (
		_w24791_,
		_w35125_,
		_w35127_,
		_w35128_
	);
	LUT3 #(
		.INIT('h65)
	) name29302 (
		\u0_L14_reg[8]/P0001 ,
		_w35122_,
		_w35128_,
		_w35129_
	);
	LUT3 #(
		.INIT('h02)
	) name29303 (
		_w34765_,
		_w34773_,
		_w34910_,
		_w35130_
	);
	LUT3 #(
		.INIT('h02)
	) name29304 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w35131_
	);
	LUT4 #(
		.INIT('h00f7)
	) name29305 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w34765_,
		_w35132_
	);
	LUT2 #(
		.INIT('h4)
	) name29306 (
		_w35131_,
		_w35132_,
		_w35133_
	);
	LUT4 #(
		.INIT('h0600)
	) name29307 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w35134_
	);
	LUT3 #(
		.INIT('h01)
	) name29308 (
		_w34782_,
		_w34763_,
		_w35134_,
		_w35135_
	);
	LUT3 #(
		.INIT('he0)
	) name29309 (
		_w35130_,
		_w35133_,
		_w35135_,
		_w35136_
	);
	LUT3 #(
		.INIT('h40)
	) name29310 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w35137_
	);
	LUT4 #(
		.INIT('h0d00)
	) name29311 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w35138_
	);
	LUT3 #(
		.INIT('h01)
	) name29312 (
		_w34765_,
		_w35138_,
		_w35137_,
		_w35139_
	);
	LUT3 #(
		.INIT('hd0)
	) name29313 (
		_w34768_,
		_w34767_,
		_w34765_,
		_w35140_
	);
	LUT2 #(
		.INIT('h4)
	) name29314 (
		_w34905_,
		_w35140_,
		_w35141_
	);
	LUT4 #(
		.INIT('h2000)
	) name29315 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w35142_
	);
	LUT3 #(
		.INIT('h04)
	) name29316 (
		_w34783_,
		_w34763_,
		_w35142_,
		_w35143_
	);
	LUT3 #(
		.INIT('he0)
	) name29317 (
		_w35139_,
		_w35141_,
		_w35143_,
		_w35144_
	);
	LUT4 #(
		.INIT('hf7c4)
	) name29318 (
		_w34784_,
		_w34765_,
		_w34772_,
		_w35142_,
		_w35145_
	);
	LUT2 #(
		.INIT('h1)
	) name29319 (
		_w34904_,
		_w35145_,
		_w35146_
	);
	LUT4 #(
		.INIT('ha955)
	) name29320 (
		\u0_L14_reg[1]/P0001 ,
		_w35136_,
		_w35144_,
		_w35146_,
		_w35147_
	);
	LUT4 #(
		.INIT('h0100)
	) name29321 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w35148_
	);
	LUT4 #(
		.INIT('h0002)
	) name29322 (
		_w34763_,
		_w34895_,
		_w35142_,
		_w35148_,
		_w35149_
	);
	LUT4 #(
		.INIT('h7f7b)
	) name29323 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w35150_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name29324 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w34765_,
		_w35151_
	);
	LUT4 #(
		.INIT('hfc54)
	) name29325 (
		_w34766_,
		_w34765_,
		_w35150_,
		_w35151_,
		_w35152_
	);
	LUT2 #(
		.INIT('h8)
	) name29326 (
		_w35149_,
		_w35152_,
		_w35153_
	);
	LUT4 #(
		.INIT('hff8c)
	) name29327 (
		_w34764_,
		_w34768_,
		_w34766_,
		_w34767_,
		_w35154_
	);
	LUT2 #(
		.INIT('h1)
	) name29328 (
		_w34765_,
		_w35154_,
		_w35155_
	);
	LUT2 #(
		.INIT('h4)
	) name29329 (
		_w34777_,
		_w34794_,
		_w35156_
	);
	LUT4 #(
		.INIT('h00fd)
	) name29330 (
		_w34764_,
		_w34766_,
		_w34767_,
		_w34763_,
		_w35157_
	);
	LUT3 #(
		.INIT('h10)
	) name29331 (
		_w34786_,
		_w34796_,
		_w35157_,
		_w35158_
	);
	LUT3 #(
		.INIT('h10)
	) name29332 (
		_w35155_,
		_w35156_,
		_w35158_,
		_w35159_
	);
	LUT3 #(
		.INIT('h60)
	) name29333 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w35160_
	);
	LUT3 #(
		.INIT('h0d)
	) name29334 (
		_w34764_,
		_w34768_,
		_w34767_,
		_w35161_
	);
	LUT3 #(
		.INIT('h02)
	) name29335 (
		_w34769_,
		_w35161_,
		_w35160_,
		_w35162_
	);
	LUT2 #(
		.INIT('h8)
	) name29336 (
		_w34768_,
		_w34765_,
		_w35163_
	);
	LUT2 #(
		.INIT('h4)
	) name29337 (
		_w34906_,
		_w35163_,
		_w35164_
	);
	LUT2 #(
		.INIT('h1)
	) name29338 (
		_w35162_,
		_w35164_,
		_w35165_
	);
	LUT4 #(
		.INIT('ha955)
	) name29339 (
		\u0_L14_reg[26]/P0001 ,
		_w35153_,
		_w35159_,
		_w35165_,
		_w35166_
	);
	LUT4 #(
		.INIT('hc963)
	) name29340 (
		decrypt_pad,
		\u1_R14_reg[17]/NET0131 ,
		\u1_uk_K_r14_reg[31]/NET0131 ,
		\u1_uk_K_r14_reg[51]/NET0131 ,
		_w35167_
	);
	LUT4 #(
		.INIT('hc693)
	) name29341 (
		decrypt_pad,
		\u1_R14_reg[21]/NET0131 ,
		\u1_uk_K_r14_reg[45]/NET0131 ,
		\u1_uk_K_r14_reg[52]/NET0131 ,
		_w35168_
	);
	LUT4 #(
		.INIT('hc693)
	) name29342 (
		decrypt_pad,
		\u1_R14_reg[16]/NET0131 ,
		\u1_uk_K_r14_reg[29]/NET0131 ,
		\u1_uk_K_r14_reg[36]/NET0131 ,
		_w35169_
	);
	LUT3 #(
		.INIT('h20)
	) name29343 (
		_w35168_,
		_w35167_,
		_w35169_,
		_w35170_
	);
	LUT4 #(
		.INIT('hc693)
	) name29344 (
		decrypt_pad,
		\u1_R14_reg[19]/P0001 ,
		\u1_uk_K_r14_reg[1]/NET0131 ,
		\u1_uk_K_r14_reg[8]/P0001 ,
		_w35171_
	);
	LUT4 #(
		.INIT('hc693)
	) name29345 (
		decrypt_pad,
		\u1_R14_reg[18]/NET0131 ,
		\u1_uk_K_r14_reg[14]/NET0131 ,
		\u1_uk_K_r14_reg[21]/NET0131 ,
		_w35172_
	);
	LUT4 #(
		.INIT('h00fb)
	) name29346 (
		_w35172_,
		_w35167_,
		_w35169_,
		_w35171_,
		_w35173_
	);
	LUT3 #(
		.INIT('h80)
	) name29347 (
		_w35168_,
		_w35167_,
		_w35169_,
		_w35174_
	);
	LUT4 #(
		.INIT('h7c00)
	) name29348 (
		_w35168_,
		_w35167_,
		_w35169_,
		_w35171_,
		_w35175_
	);
	LUT4 #(
		.INIT('hfeba)
	) name29349 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35176_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name29350 (
		_w35170_,
		_w35173_,
		_w35175_,
		_w35176_,
		_w35177_
	);
	LUT2 #(
		.INIT('h4)
	) name29351 (
		_w35168_,
		_w35169_,
		_w35178_
	);
	LUT4 #(
		.INIT('h9fdf)
	) name29352 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35179_
	);
	LUT4 #(
		.INIT('hc693)
	) name29353 (
		decrypt_pad,
		\u1_R14_reg[20]/NET0131 ,
		\u1_uk_K_r14_reg[16]/NET0131 ,
		\u1_uk_K_r14_reg[23]/NET0131 ,
		_w35180_
	);
	LUT3 #(
		.INIT('hb0)
	) name29354 (
		_w35177_,
		_w35179_,
		_w35180_,
		_w35181_
	);
	LUT4 #(
		.INIT('hbff9)
	) name29355 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35182_
	);
	LUT2 #(
		.INIT('h2)
	) name29356 (
		_w35171_,
		_w35182_,
		_w35183_
	);
	LUT2 #(
		.INIT('h4)
	) name29357 (
		_w35168_,
		_w35171_,
		_w35184_
	);
	LUT4 #(
		.INIT('hfa3f)
	) name29358 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35185_
	);
	LUT3 #(
		.INIT('hb0)
	) name29359 (
		_w35168_,
		_w35167_,
		_w35171_,
		_w35186_
	);
	LUT4 #(
		.INIT('h5501)
	) name29360 (
		_w35172_,
		_w35167_,
		_w35169_,
		_w35171_,
		_w35187_
	);
	LUT4 #(
		.INIT('he0ee)
	) name29361 (
		_w35184_,
		_w35185_,
		_w35186_,
		_w35187_,
		_w35188_
	);
	LUT4 #(
		.INIT('h2000)
	) name29362 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35189_
	);
	LUT2 #(
		.INIT('h2)
	) name29363 (
		_w35172_,
		_w35171_,
		_w35190_
	);
	LUT4 #(
		.INIT('h0020)
	) name29364 (
		_w35172_,
		_w35167_,
		_w35169_,
		_w35171_,
		_w35191_
	);
	LUT2 #(
		.INIT('h1)
	) name29365 (
		_w35189_,
		_w35191_,
		_w35192_
	);
	LUT4 #(
		.INIT('h0e00)
	) name29366 (
		_w35180_,
		_w35188_,
		_w35183_,
		_w35192_,
		_w35193_
	);
	LUT3 #(
		.INIT('h65)
	) name29367 (
		\u1_L14_reg[25]/P0001 ,
		_w35181_,
		_w35193_,
		_w35194_
	);
	LUT4 #(
		.INIT('hc693)
	) name29368 (
		decrypt_pad,
		\u1_R14_reg[16]/NET0131 ,
		\u1_uk_K_r14_reg[33]/NET0131 ,
		\u1_uk_K_r14_reg[40]/NET0131 ,
		_w35195_
	);
	LUT4 #(
		.INIT('hc963)
	) name29369 (
		decrypt_pad,
		\u1_R14_reg[12]/NET0131 ,
		\u1_uk_K_r14_reg[4]/NET0131 ,
		\u1_uk_K_r14_reg[54]/NET0131 ,
		_w35196_
	);
	LUT4 #(
		.INIT('hc693)
	) name29370 (
		decrypt_pad,
		\u1_R14_reg[15]/NET0131 ,
		\u1_uk_K_r14_reg[25]/NET0131 ,
		\u1_uk_K_r14_reg[32]/NET0131 ,
		_w35197_
	);
	LUT4 #(
		.INIT('hc693)
	) name29371 (
		decrypt_pad,
		\u1_R14_reg[14]/NET0131 ,
		\u1_uk_K_r14_reg[17]/NET0131 ,
		\u1_uk_K_r14_reg[24]/NET0131 ,
		_w35198_
	);
	LUT4 #(
		.INIT('hc693)
	) name29372 (
		decrypt_pad,
		\u1_R14_reg[13]/NET0131 ,
		\u1_uk_K_r14_reg[48]/NET0131 ,
		\u1_uk_K_r14_reg[55]/NET0131 ,
		_w35199_
	);
	LUT4 #(
		.INIT('hc693)
	) name29373 (
		decrypt_pad,
		\u1_R14_reg[17]/NET0131 ,
		\u1_uk_K_r14_reg[13]/NET0131 ,
		\u1_uk_K_r14_reg[20]/NET0131 ,
		_w35200_
	);
	LUT4 #(
		.INIT('hc2cd)
	) name29374 (
		_w35200_,
		_w35198_,
		_w35199_,
		_w35197_,
		_w35201_
	);
	LUT2 #(
		.INIT('h2)
	) name29375 (
		_w35196_,
		_w35201_,
		_w35202_
	);
	LUT4 #(
		.INIT('h0001)
	) name29376 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35203_
	);
	LUT4 #(
		.INIT('heffe)
	) name29377 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35204_
	);
	LUT3 #(
		.INIT('h01)
	) name29378 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35205_
	);
	LUT4 #(
		.INIT('h0001)
	) name29379 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35197_,
		_w35206_
	);
	LUT2 #(
		.INIT('h2)
	) name29380 (
		_w35200_,
		_w35196_,
		_w35207_
	);
	LUT4 #(
		.INIT('h0200)
	) name29381 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35197_,
		_w35208_
	);
	LUT3 #(
		.INIT('h02)
	) name29382 (
		_w35204_,
		_w35206_,
		_w35208_,
		_w35209_
	);
	LUT3 #(
		.INIT('h45)
	) name29383 (
		_w35195_,
		_w35202_,
		_w35209_,
		_w35210_
	);
	LUT4 #(
		.INIT('h0008)
	) name29384 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35211_
	);
	LUT4 #(
		.INIT('heef7)
	) name29385 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35212_
	);
	LUT4 #(
		.INIT('h8000)
	) name29386 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35213_
	);
	LUT3 #(
		.INIT('h04)
	) name29387 (
		_w35196_,
		_w35198_,
		_w35199_,
		_w35214_
	);
	LUT4 #(
		.INIT('h7fdf)
	) name29388 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35215_
	);
	LUT4 #(
		.INIT('h0200)
	) name29389 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35216_
	);
	LUT4 #(
		.INIT('hbdbb)
	) name29390 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35217_
	);
	LUT4 #(
		.INIT('ha808)
	) name29391 (
		_w35215_,
		_w35217_,
		_w35197_,
		_w35212_,
		_w35218_
	);
	LUT4 #(
		.INIT('h7fde)
	) name29392 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35219_
	);
	LUT2 #(
		.INIT('h1)
	) name29393 (
		_w35197_,
		_w35219_,
		_w35220_
	);
	LUT3 #(
		.INIT('h80)
	) name29394 (
		_w35198_,
		_w35199_,
		_w35197_,
		_w35221_
	);
	LUT4 #(
		.INIT('h4000)
	) name29395 (
		_w35196_,
		_w35198_,
		_w35199_,
		_w35197_,
		_w35222_
	);
	LUT4 #(
		.INIT('h4000)
	) name29396 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35197_,
		_w35223_
	);
	LUT2 #(
		.INIT('h4)
	) name29397 (
		_w35198_,
		_w35223_,
		_w35224_
	);
	LUT3 #(
		.INIT('h23)
	) name29398 (
		_w35198_,
		_w35222_,
		_w35223_,
		_w35225_
	);
	LUT4 #(
		.INIT('h0d00)
	) name29399 (
		_w35195_,
		_w35218_,
		_w35220_,
		_w35225_,
		_w35226_
	);
	LUT3 #(
		.INIT('h65)
	) name29400 (
		\u1_L14_reg[10]/P0001 ,
		_w35210_,
		_w35226_,
		_w35227_
	);
	LUT3 #(
		.INIT('ha6)
	) name29401 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w35228_
	);
	LUT3 #(
		.INIT('h51)
	) name29402 (
		_w15393_,
		_w15388_,
		_w15392_,
		_w35229_
	);
	LUT2 #(
		.INIT('h8)
	) name29403 (
		_w35228_,
		_w35229_,
		_w35230_
	);
	LUT3 #(
		.INIT('h08)
	) name29404 (
		_w15393_,
		_w15389_,
		_w15391_,
		_w35231_
	);
	LUT3 #(
		.INIT('h15)
	) name29405 (
		_w15387_,
		_w15396_,
		_w35231_,
		_w35232_
	);
	LUT4 #(
		.INIT('h0034)
	) name29406 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35233_
	);
	LUT3 #(
		.INIT('h40)
	) name29407 (
		_w15388_,
		_w15389_,
		_w15392_,
		_w35234_
	);
	LUT4 #(
		.INIT('h4000)
	) name29408 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35235_
	);
	LUT4 #(
		.INIT('h0004)
	) name29409 (
		_w15393_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35236_
	);
	LUT3 #(
		.INIT('h01)
	) name29410 (
		_w35233_,
		_w35235_,
		_w35236_,
		_w35237_
	);
	LUT3 #(
		.INIT('h40)
	) name29411 (
		_w35230_,
		_w35232_,
		_w35237_,
		_w35238_
	);
	LUT2 #(
		.INIT('h6)
	) name29412 (
		_w15388_,
		_w15389_,
		_w35239_
	);
	LUT3 #(
		.INIT('h8c)
	) name29413 (
		_w15389_,
		_w15391_,
		_w15392_,
		_w35240_
	);
	LUT3 #(
		.INIT('h02)
	) name29414 (
		_w35229_,
		_w35240_,
		_w35239_,
		_w35241_
	);
	LUT3 #(
		.INIT('h82)
	) name29415 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w35242_
	);
	LUT4 #(
		.INIT('h0082)
	) name29416 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35243_
	);
	LUT4 #(
		.INIT('h80a0)
	) name29417 (
		_w15393_,
		_w15388_,
		_w15391_,
		_w15392_,
		_w35244_
	);
	LUT3 #(
		.INIT('h02)
	) name29418 (
		_w15387_,
		_w35243_,
		_w35244_,
		_w35245_
	);
	LUT2 #(
		.INIT('h4)
	) name29419 (
		_w35241_,
		_w35245_,
		_w35246_
	);
	LUT4 #(
		.INIT('h4004)
	) name29420 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35247_
	);
	LUT3 #(
		.INIT('h08)
	) name29421 (
		_w15388_,
		_w15391_,
		_w15392_,
		_w35248_
	);
	LUT4 #(
		.INIT('hfad8)
	) name29422 (
		_w15393_,
		_w15403_,
		_w35247_,
		_w35248_,
		_w35249_
	);
	LUT4 #(
		.INIT('h55a9)
	) name29423 (
		\u1_L14_reg[2]/P0001 ,
		_w35238_,
		_w35246_,
		_w35249_,
		_w35250_
	);
	LUT2 #(
		.INIT('h8)
	) name29424 (
		_w15293_,
		_w15295_,
		_w35251_
	);
	LUT3 #(
		.INIT('h28)
	) name29425 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w35252_
	);
	LUT4 #(
		.INIT('h8082)
	) name29426 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35253_
	);
	LUT4 #(
		.INIT('hfe54)
	) name29427 (
		_w15291_,
		_w15311_,
		_w35252_,
		_w35253_,
		_w35254_
	);
	LUT4 #(
		.INIT('h1000)
	) name29428 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35255_
	);
	LUT4 #(
		.INIT('hfb00)
	) name29429 (
		_w15292_,
		_w15293_,
		_w15294_,
		_w15299_,
		_w35256_
	);
	LUT3 #(
		.INIT('h10)
	) name29430 (
		_w15316_,
		_w35255_,
		_w35256_,
		_w35257_
	);
	LUT3 #(
		.INIT('h40)
	) name29431 (
		_w15291_,
		_w15293_,
		_w15295_,
		_w35258_
	);
	LUT4 #(
		.INIT('hafcf)
	) name29432 (
		_w15291_,
		_w15292_,
		_w15293_,
		_w15295_,
		_w35259_
	);
	LUT2 #(
		.INIT('h2)
	) name29433 (
		_w15294_,
		_w35259_,
		_w35260_
	);
	LUT4 #(
		.INIT('haaa2)
	) name29434 (
		_w15291_,
		_w15292_,
		_w15293_,
		_w15294_,
		_w35261_
	);
	LUT4 #(
		.INIT('h31bb)
	) name29435 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35262_
	);
	LUT4 #(
		.INIT('h0004)
	) name29436 (
		_w15291_,
		_w15292_,
		_w15293_,
		_w15295_,
		_w35263_
	);
	LUT4 #(
		.INIT('h0015)
	) name29437 (
		_w15299_,
		_w35261_,
		_w35262_,
		_w35263_,
		_w35264_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name29438 (
		_w35254_,
		_w35257_,
		_w35260_,
		_w35264_,
		_w35265_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name29439 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35266_
	);
	LUT4 #(
		.INIT('h0200)
	) name29440 (
		_w15291_,
		_w15292_,
		_w15293_,
		_w15294_,
		_w35267_
	);
	LUT4 #(
		.INIT('h0020)
	) name29441 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35268_
	);
	LUT4 #(
		.INIT('h2232)
	) name29442 (
		_w15291_,
		_w35267_,
		_w35266_,
		_w35268_,
		_w35269_
	);
	LUT3 #(
		.INIT('h65)
	) name29443 (
		\u1_L14_reg[27]/P0001 ,
		_w35265_,
		_w35269_,
		_w35270_
	);
	LUT4 #(
		.INIT('hc963)
	) name29444 (
		decrypt_pad,
		\u1_R14_reg[20]/NET0131 ,
		\u1_uk_K_r14_reg[14]/NET0131 ,
		\u1_uk_K_r14_reg[7]/NET0131 ,
		_w35271_
	);
	LUT4 #(
		.INIT('hc693)
	) name29445 (
		decrypt_pad,
		\u1_R14_reg[21]/NET0131 ,
		\u1_uk_K_r14_reg[22]/NET0131 ,
		\u1_uk_K_r14_reg[29]/NET0131 ,
		_w35272_
	);
	LUT4 #(
		.INIT('hc693)
	) name29446 (
		decrypt_pad,
		\u1_R14_reg[22]/P0001 ,
		\u1_uk_K_r14_reg[44]/NET0131 ,
		\u1_uk_K_r14_reg[51]/NET0131 ,
		_w35273_
	);
	LUT3 #(
		.INIT('h08)
	) name29447 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35274_
	);
	LUT4 #(
		.INIT('hc693)
	) name29448 (
		decrypt_pad,
		\u1_R14_reg[23]/P0001 ,
		\u1_uk_K_r14_reg[2]/NET0131 ,
		\u1_uk_K_r14_reg[9]/NET0131 ,
		_w35275_
	);
	LUT4 #(
		.INIT('hc693)
	) name29449 (
		decrypt_pad,
		\u1_R14_reg[25]/NET0131 ,
		\u1_uk_K_r14_reg[23]/NET0131 ,
		\u1_uk_K_r14_reg[30]/NET0131 ,
		_w35276_
	);
	LUT3 #(
		.INIT('h10)
	) name29450 (
		_w35271_,
		_w35272_,
		_w35276_,
		_w35277_
	);
	LUT4 #(
		.INIT('he0f0)
	) name29451 (
		_w35271_,
		_w35272_,
		_w35275_,
		_w35276_,
		_w35278_
	);
	LUT4 #(
		.INIT('h0200)
	) name29452 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35279_
	);
	LUT4 #(
		.INIT('hfda8)
	) name29453 (
		_w35275_,
		_w35274_,
		_w35277_,
		_w35279_,
		_w35280_
	);
	LUT4 #(
		.INIT('h0110)
	) name29454 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35281_
	);
	LUT4 #(
		.INIT('h4000)
	) name29455 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35282_
	);
	LUT3 #(
		.INIT('h02)
	) name29456 (
		_w35272_,
		_w35273_,
		_w35276_,
		_w35283_
	);
	LUT4 #(
		.INIT('hc693)
	) name29457 (
		decrypt_pad,
		\u1_R14_reg[24]/NET0131 ,
		\u1_uk_K_r14_reg[28]/NET0131 ,
		\u1_uk_K_r14_reg[35]/P0001 ,
		_w35284_
	);
	LUT4 #(
		.INIT('hfd00)
	) name29458 (
		_w35271_,
		_w35272_,
		_w35275_,
		_w35284_,
		_w35285_
	);
	LUT4 #(
		.INIT('h0100)
	) name29459 (
		_w35283_,
		_w35281_,
		_w35282_,
		_w35285_,
		_w35286_
	);
	LUT2 #(
		.INIT('h4)
	) name29460 (
		_w35280_,
		_w35286_,
		_w35287_
	);
	LUT3 #(
		.INIT('h01)
	) name29461 (
		_w35271_,
		_w35272_,
		_w35276_,
		_w35288_
	);
	LUT3 #(
		.INIT('hbe)
	) name29462 (
		_w35271_,
		_w35272_,
		_w35276_,
		_w35289_
	);
	LUT3 #(
		.INIT('h10)
	) name29463 (
		_w35275_,
		_w35279_,
		_w35289_,
		_w35290_
	);
	LUT3 #(
		.INIT('h04)
	) name29464 (
		_w35271_,
		_w35272_,
		_w35276_,
		_w35291_
	);
	LUT4 #(
		.INIT('h50d0)
	) name29465 (
		_w35271_,
		_w35272_,
		_w35275_,
		_w35273_,
		_w35292_
	);
	LUT2 #(
		.INIT('h4)
	) name29466 (
		_w35291_,
		_w35292_,
		_w35293_
	);
	LUT3 #(
		.INIT('h80)
	) name29467 (
		_w35271_,
		_w35272_,
		_w35276_,
		_w35294_
	);
	LUT4 #(
		.INIT('h8000)
	) name29468 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35295_
	);
	LUT2 #(
		.INIT('h1)
	) name29469 (
		_w35284_,
		_w35295_,
		_w35296_
	);
	LUT3 #(
		.INIT('he0)
	) name29470 (
		_w35290_,
		_w35293_,
		_w35296_,
		_w35297_
	);
	LUT2 #(
		.INIT('h1)
	) name29471 (
		_w35275_,
		_w35273_,
		_w35298_
	);
	LUT3 #(
		.INIT('h08)
	) name29472 (
		_w35271_,
		_w35272_,
		_w35276_,
		_w35299_
	);
	LUT4 #(
		.INIT('hcedf)
	) name29473 (
		_w35275_,
		_w35273_,
		_w35277_,
		_w35299_,
		_w35300_
	);
	LUT4 #(
		.INIT('ha955)
	) name29474 (
		\u1_L14_reg[19]/P0001 ,
		_w35287_,
		_w35297_,
		_w35300_,
		_w35301_
	);
	LUT4 #(
		.INIT('h14b0)
	) name29475 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35302_
	);
	LUT3 #(
		.INIT('h01)
	) name29476 (
		_w35275_,
		_w35279_,
		_w35302_,
		_w35303_
	);
	LUT4 #(
		.INIT('h0002)
	) name29477 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35304_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name29478 (
		_w35271_,
		_w35272_,
		_w35275_,
		_w35273_,
		_w35305_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name29479 (
		_w35284_,
		_w35294_,
		_w35304_,
		_w35305_,
		_w35306_
	);
	LUT2 #(
		.INIT('h4)
	) name29480 (
		_w35303_,
		_w35306_,
		_w35307_
	);
	LUT2 #(
		.INIT('h1)
	) name29481 (
		_w35271_,
		_w35273_,
		_w35308_
	);
	LUT4 #(
		.INIT('h0b07)
	) name29482 (
		_w35271_,
		_w35272_,
		_w35275_,
		_w35273_,
		_w35309_
	);
	LUT3 #(
		.INIT('h0d)
	) name29483 (
		_w35278_,
		_w35308_,
		_w35309_,
		_w35310_
	);
	LUT4 #(
		.INIT('h0002)
	) name29484 (
		_w35271_,
		_w35275_,
		_w35273_,
		_w35276_,
		_w35311_
	);
	LUT4 #(
		.INIT('h2000)
	) name29485 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35312_
	);
	LUT2 #(
		.INIT('h8)
	) name29486 (
		_w35275_,
		_w35273_,
		_w35313_
	);
	LUT4 #(
		.INIT('hbfb5)
	) name29487 (
		_w35272_,
		_w35275_,
		_w35273_,
		_w35276_,
		_w35314_
	);
	LUT4 #(
		.INIT('h0301)
	) name29488 (
		_w35271_,
		_w35311_,
		_w35312_,
		_w35314_,
		_w35315_
	);
	LUT3 #(
		.INIT('h45)
	) name29489 (
		_w35284_,
		_w35310_,
		_w35315_,
		_w35316_
	);
	LUT4 #(
		.INIT('h5ffb)
	) name29490 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35317_
	);
	LUT2 #(
		.INIT('h2)
	) name29491 (
		_w35275_,
		_w35317_,
		_w35318_
	);
	LUT2 #(
		.INIT('h8)
	) name29492 (
		_w35288_,
		_w35298_,
		_w35319_
	);
	LUT3 #(
		.INIT('h02)
	) name29493 (
		_w35300_,
		_w35319_,
		_w35318_,
		_w35320_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name29494 (
		\u1_L14_reg[11]/P0001 ,
		_w35316_,
		_w35307_,
		_w35320_,
		_w35321_
	);
	LUT4 #(
		.INIT('h0008)
	) name29495 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35322_
	);
	LUT4 #(
		.INIT('h0100)
	) name29496 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35323_
	);
	LUT3 #(
		.INIT('h02)
	) name29497 (
		_w35171_,
		_w35322_,
		_w35323_,
		_w35324_
	);
	LUT4 #(
		.INIT('h0001)
	) name29498 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35325_
	);
	LUT4 #(
		.INIT('h1000)
	) name29499 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35326_
	);
	LUT4 #(
		.INIT('h0800)
	) name29500 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35327_
	);
	LUT4 #(
		.INIT('he7ff)
	) name29501 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35328_
	);
	LUT3 #(
		.INIT('h10)
	) name29502 (
		_w35171_,
		_w35325_,
		_w35328_,
		_w35329_
	);
	LUT2 #(
		.INIT('h1)
	) name29503 (
		_w35324_,
		_w35329_,
		_w35330_
	);
	LUT2 #(
		.INIT('h2)
	) name29504 (
		_w35172_,
		_w35167_,
		_w35331_
	);
	LUT4 #(
		.INIT('h2022)
	) name29505 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35332_
	);
	LUT4 #(
		.INIT('h5051)
	) name29506 (
		_w35178_,
		_w35171_,
		_w35331_,
		_w35332_,
		_w35333_
	);
	LUT4 #(
		.INIT('hafdd)
	) name29507 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35334_
	);
	LUT3 #(
		.INIT('h31)
	) name29508 (
		_w35171_,
		_w35180_,
		_w35334_,
		_w35335_
	);
	LUT4 #(
		.INIT('hddaf)
	) name29509 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35336_
	);
	LUT2 #(
		.INIT('h2)
	) name29510 (
		_w35171_,
		_w35336_,
		_w35337_
	);
	LUT4 #(
		.INIT('h0008)
	) name29511 (
		_w35168_,
		_w35167_,
		_w35169_,
		_w35171_,
		_w35338_
	);
	LUT4 #(
		.INIT('h0400)
	) name29512 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35339_
	);
	LUT4 #(
		.INIT('h0002)
	) name29513 (
		_w35180_,
		_w35189_,
		_w35339_,
		_w35338_,
		_w35340_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name29514 (
		_w35333_,
		_w35335_,
		_w35337_,
		_w35340_,
		_w35341_
	);
	LUT3 #(
		.INIT('h56)
	) name29515 (
		\u1_L14_reg[3]/P0001 ,
		_w35330_,
		_w35341_,
		_w35342_
	);
	LUT4 #(
		.INIT('h0400)
	) name29516 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35343_
	);
	LUT4 #(
		.INIT('hfb55)
	) name29517 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35344_
	);
	LUT4 #(
		.INIT('h1000)
	) name29518 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35345_
	);
	LUT4 #(
		.INIT('h0020)
	) name29519 (
		_w15393_,
		_w35242_,
		_w35344_,
		_w35345_,
		_w35346_
	);
	LUT4 #(
		.INIT('h0408)
	) name29520 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35347_
	);
	LUT3 #(
		.INIT('h10)
	) name29521 (
		_w15388_,
		_w15391_,
		_w15392_,
		_w35348_
	);
	LUT4 #(
		.INIT('h4051)
	) name29522 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35349_
	);
	LUT4 #(
		.INIT('h0001)
	) name29523 (
		_w15393_,
		_w15397_,
		_w35348_,
		_w35349_,
		_w35350_
	);
	LUT4 #(
		.INIT('h8a88)
	) name29524 (
		_w15387_,
		_w35346_,
		_w35347_,
		_w35350_,
		_w35351_
	);
	LUT2 #(
		.INIT('h2)
	) name29525 (
		_w15393_,
		_w35349_,
		_w35352_
	);
	LUT3 #(
		.INIT('h10)
	) name29526 (
		_w15389_,
		_w15391_,
		_w15392_,
		_w35353_
	);
	LUT4 #(
		.INIT('ha4a6)
	) name29527 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35354_
	);
	LUT4 #(
		.INIT('h0001)
	) name29528 (
		_w15393_,
		_w15397_,
		_w35348_,
		_w35354_,
		_w35355_
	);
	LUT3 #(
		.INIT('h09)
	) name29529 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w35356_
	);
	LUT4 #(
		.INIT('h2900)
	) name29530 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35357_
	);
	LUT2 #(
		.INIT('h1)
	) name29531 (
		_w15387_,
		_w35357_,
		_w35358_
	);
	LUT3 #(
		.INIT('he0)
	) name29532 (
		_w35352_,
		_w35355_,
		_w35358_,
		_w35359_
	);
	LUT3 #(
		.INIT('ha9)
	) name29533 (
		\u1_L14_reg[28]/P0001 ,
		_w35351_,
		_w35359_,
		_w35360_
	);
	LUT4 #(
		.INIT('h0200)
	) name29534 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35197_,
		_w35361_
	);
	LUT4 #(
		.INIT('h0012)
	) name29535 (
		_w35196_,
		_w35198_,
		_w35199_,
		_w35197_,
		_w35362_
	);
	LUT4 #(
		.INIT('h0001)
	) name29536 (
		_w35216_,
		_w35223_,
		_w35362_,
		_w35361_,
		_w35363_
	);
	LUT4 #(
		.INIT('h020a)
	) name29537 (
		_w35195_,
		_w35198_,
		_w35213_,
		_w35206_,
		_w35364_
	);
	LUT3 #(
		.INIT('hd0)
	) name29538 (
		_w35200_,
		_w35199_,
		_w35197_,
		_w35365_
	);
	LUT4 #(
		.INIT('h8100)
	) name29539 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35197_,
		_w35366_
	);
	LUT4 #(
		.INIT('h0001)
	) name29540 (
		_w35195_,
		_w35211_,
		_w35222_,
		_w35366_,
		_w35367_
	);
	LUT4 #(
		.INIT('hbf15)
	) name29541 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35368_
	);
	LUT3 #(
		.INIT('hc8)
	) name29542 (
		_w35197_,
		_w35204_,
		_w35368_,
		_w35369_
	);
	LUT4 #(
		.INIT('h0777)
	) name29543 (
		_w35363_,
		_w35364_,
		_w35367_,
		_w35369_,
		_w35370_
	);
	LUT4 #(
		.INIT('h0040)
	) name29544 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35371_
	);
	LUT4 #(
		.INIT('heee2)
	) name29545 (
		_w35216_,
		_w35197_,
		_w35203_,
		_w35371_,
		_w35372_
	);
	LUT2 #(
		.INIT('h1)
	) name29546 (
		_w35224_,
		_w35372_,
		_w35373_
	);
	LUT3 #(
		.INIT('h65)
	) name29547 (
		\u1_L14_reg[20]/P0001 ,
		_w35370_,
		_w35373_,
		_w35374_
	);
	LUT4 #(
		.INIT('hc693)
	) name29548 (
		decrypt_pad,
		\u1_R14_reg[26]/NET0131 ,
		\u1_uk_K_r14_reg[15]/NET0131 ,
		\u1_uk_K_r14_reg[22]/NET0131 ,
		_w35375_
	);
	LUT4 #(
		.INIT('hc963)
	) name29549 (
		decrypt_pad,
		\u1_R14_reg[24]/NET0131 ,
		\u1_uk_K_r14_reg[2]/NET0131 ,
		\u1_uk_K_r14_reg[50]/NET0131 ,
		_w35376_
	);
	LUT4 #(
		.INIT('hc693)
	) name29550 (
		decrypt_pad,
		\u1_R14_reg[25]/NET0131 ,
		\u1_uk_K_r14_reg[30]/NET0131 ,
		\u1_uk_K_r14_reg[37]/NET0131 ,
		_w35377_
	);
	LUT4 #(
		.INIT('hc693)
	) name29551 (
		decrypt_pad,
		\u1_R14_reg[29]/NET0131 ,
		\u1_uk_K_r14_reg[31]/NET0131 ,
		\u1_uk_K_r14_reg[38]/NET0131 ,
		_w35378_
	);
	LUT3 #(
		.INIT('h40)
	) name29552 (
		_w35377_,
		_w35378_,
		_w35376_,
		_w35379_
	);
	LUT4 #(
		.INIT('h1428)
	) name29553 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35380_
	);
	LUT3 #(
		.INIT('h54)
	) name29554 (
		_w35377_,
		_w35375_,
		_w35376_,
		_w35381_
	);
	LUT4 #(
		.INIT('hc963)
	) name29555 (
		decrypt_pad,
		\u1_R14_reg[27]/P0001 ,
		\u1_uk_K_r14_reg[0]/P0001 ,
		\u1_uk_K_r14_reg[52]/NET0131 ,
		_w35382_
	);
	LUT4 #(
		.INIT('hf100)
	) name29556 (
		_w35377_,
		_w35378_,
		_w35376_,
		_w35382_,
		_w35383_
	);
	LUT2 #(
		.INIT('h4)
	) name29557 (
		_w35381_,
		_w35383_,
		_w35384_
	);
	LUT4 #(
		.INIT('h0040)
	) name29558 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35385_
	);
	LUT4 #(
		.INIT('hc693)
	) name29559 (
		decrypt_pad,
		\u1_R14_reg[28]/NET0131 ,
		\u1_uk_K_r14_reg[35]/P0001 ,
		\u1_uk_K_r14_reg[42]/P0001 ,
		_w35386_
	);
	LUT3 #(
		.INIT('hd0)
	) name29560 (
		_w35385_,
		_w35382_,
		_w35386_,
		_w35387_
	);
	LUT3 #(
		.INIT('h10)
	) name29561 (
		_w35380_,
		_w35384_,
		_w35387_,
		_w35388_
	);
	LUT4 #(
		.INIT('h0102)
	) name29562 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35389_
	);
	LUT3 #(
		.INIT('h08)
	) name29563 (
		_w35375_,
		_w35376_,
		_w35382_,
		_w35390_
	);
	LUT2 #(
		.INIT('h4)
	) name29564 (
		_w35377_,
		_w35382_,
		_w35391_
	);
	LUT4 #(
		.INIT('h0400)
	) name29565 (
		_w35377_,
		_w35378_,
		_w35376_,
		_w35382_,
		_w35392_
	);
	LUT3 #(
		.INIT('h01)
	) name29566 (
		_w35386_,
		_w35392_,
		_w35390_,
		_w35393_
	);
	LUT4 #(
		.INIT('h4000)
	) name29567 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35394_
	);
	LUT2 #(
		.INIT('h6)
	) name29568 (
		_w35377_,
		_w35378_,
		_w35395_
	);
	LUT3 #(
		.INIT('hd0)
	) name29569 (
		_w35375_,
		_w35376_,
		_w35382_,
		_w35396_
	);
	LUT3 #(
		.INIT('h54)
	) name29570 (
		_w35394_,
		_w35395_,
		_w35396_,
		_w35397_
	);
	LUT3 #(
		.INIT('h40)
	) name29571 (
		_w35389_,
		_w35393_,
		_w35397_,
		_w35398_
	);
	LUT3 #(
		.INIT('ha9)
	) name29572 (
		\u1_L14_reg[12]/P0001 ,
		_w35388_,
		_w35398_,
		_w35399_
	);
	LUT4 #(
		.INIT('hfb05)
	) name29573 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35400_
	);
	LUT2 #(
		.INIT('h2)
	) name29574 (
		_w15321_,
		_w35400_,
		_w35401_
	);
	LUT4 #(
		.INIT('hbf00)
	) name29575 (
		_w15321_,
		_w15322_,
		_w15323_,
		_w15331_,
		_w35402_
	);
	LUT4 #(
		.INIT('h0001)
	) name29576 (
		_w15321_,
		_w15322_,
		_w15325_,
		_w15323_,
		_w35403_
	);
	LUT4 #(
		.INIT('h0100)
	) name29577 (
		_w15332_,
		_w15338_,
		_w35403_,
		_w35402_,
		_w35404_
	);
	LUT2 #(
		.INIT('h4)
	) name29578 (
		_w35401_,
		_w35404_,
		_w35405_
	);
	LUT3 #(
		.INIT('h6f)
	) name29579 (
		_w15324_,
		_w15325_,
		_w15323_,
		_w35406_
	);
	LUT4 #(
		.INIT('h0040)
	) name29580 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35407_
	);
	LUT4 #(
		.INIT('h0020)
	) name29581 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35408_
	);
	LUT4 #(
		.INIT('h0200)
	) name29582 (
		_w15321_,
		_w35408_,
		_w35407_,
		_w35406_,
		_w35409_
	);
	LUT3 #(
		.INIT('h21)
	) name29583 (
		_w15324_,
		_w15325_,
		_w15323_,
		_w35410_
	);
	LUT4 #(
		.INIT('h5554)
	) name29584 (
		_w15321_,
		_w15322_,
		_w15324_,
		_w15323_,
		_w35411_
	);
	LUT2 #(
		.INIT('h4)
	) name29585 (
		_w35410_,
		_w35411_,
		_w35412_
	);
	LUT4 #(
		.INIT('h0008)
	) name29586 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35413_
	);
	LUT3 #(
		.INIT('h01)
	) name29587 (
		_w15331_,
		_w15343_,
		_w35413_,
		_w35414_
	);
	LUT3 #(
		.INIT('he0)
	) name29588 (
		_w35409_,
		_w35412_,
		_w35414_,
		_w35415_
	);
	LUT3 #(
		.INIT('ha9)
	) name29589 (
		\u1_L14_reg[17]/P0001 ,
		_w35405_,
		_w35415_,
		_w35416_
	);
	LUT4 #(
		.INIT('h1000)
	) name29590 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35417_
	);
	LUT3 #(
		.INIT('h20)
	) name29591 (
		_w35271_,
		_w35273_,
		_w35276_,
		_w35418_
	);
	LUT4 #(
		.INIT('he5bb)
	) name29592 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35419_
	);
	LUT4 #(
		.INIT('hda77)
	) name29593 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35420_
	);
	LUT4 #(
		.INIT('h3120)
	) name29594 (
		_w35275_,
		_w35304_,
		_w35420_,
		_w35419_,
		_w35421_
	);
	LUT4 #(
		.INIT('hfaf2)
	) name29595 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35422_
	);
	LUT4 #(
		.INIT('h3ffb)
	) name29596 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35423_
	);
	LUT4 #(
		.INIT('h7200)
	) name29597 (
		_w35275_,
		_w35418_,
		_w35422_,
		_w35423_,
		_w35424_
	);
	LUT3 #(
		.INIT('hb6)
	) name29598 (
		_w35271_,
		_w35272_,
		_w35276_,
		_w35425_
	);
	LUT4 #(
		.INIT('h70d0)
	) name29599 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35426_
	);
	LUT4 #(
		.INIT('h3031)
	) name29600 (
		_w35271_,
		_w35275_,
		_w35273_,
		_w35276_,
		_w35427_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name29601 (
		_w35313_,
		_w35425_,
		_w35426_,
		_w35427_,
		_w35428_
	);
	LUT4 #(
		.INIT('hd800)
	) name29602 (
		_w35284_,
		_w35424_,
		_w35421_,
		_w35428_,
		_w35429_
	);
	LUT2 #(
		.INIT('h9)
	) name29603 (
		\u1_L14_reg[4]/P0001 ,
		_w35429_,
		_w35430_
	);
	LUT4 #(
		.INIT('hbb7b)
	) name29604 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35431_
	);
	LUT2 #(
		.INIT('h2)
	) name29605 (
		_w35275_,
		_w35431_,
		_w35432_
	);
	LUT4 #(
		.INIT('h5fae)
	) name29606 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35433_
	);
	LUT2 #(
		.INIT('h1)
	) name29607 (
		_w35275_,
		_w35433_,
		_w35434_
	);
	LUT3 #(
		.INIT('h01)
	) name29608 (
		_w35281_,
		_w35311_,
		_w35312_,
		_w35435_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name29609 (
		_w35284_,
		_w35432_,
		_w35434_,
		_w35435_,
		_w35436_
	);
	LUT4 #(
		.INIT('h779c)
	) name29610 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35437_
	);
	LUT4 #(
		.INIT('h3032)
	) name29611 (
		_w35275_,
		_w35284_,
		_w35417_,
		_w35437_,
		_w35438_
	);
	LUT4 #(
		.INIT('hf17b)
	) name29612 (
		_w35271_,
		_w35272_,
		_w35273_,
		_w35276_,
		_w35439_
	);
	LUT2 #(
		.INIT('h1)
	) name29613 (
		_w35275_,
		_w35284_,
		_w35440_
	);
	LUT4 #(
		.INIT('h0800)
	) name29614 (
		_w35272_,
		_w35275_,
		_w35273_,
		_w35276_,
		_w35441_
	);
	LUT4 #(
		.INIT('h1011)
	) name29615 (
		_w35304_,
		_w35441_,
		_w35439_,
		_w35440_,
		_w35442_
	);
	LUT2 #(
		.INIT('h4)
	) name29616 (
		_w35438_,
		_w35442_,
		_w35443_
	);
	LUT3 #(
		.INIT('h9a)
	) name29617 (
		\u1_L14_reg[29]/P0001 ,
		_w35436_,
		_w35443_,
		_w35444_
	);
	LUT3 #(
		.INIT('h0d)
	) name29618 (
		_w15291_,
		_w15292_,
		_w15294_,
		_w35445_
	);
	LUT2 #(
		.INIT('h8)
	) name29619 (
		_w35251_,
		_w35445_,
		_w35446_
	);
	LUT3 #(
		.INIT('h01)
	) name29620 (
		_w15299_,
		_w15312_,
		_w35263_,
		_w35447_
	);
	LUT4 #(
		.INIT('h8fdf)
	) name29621 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35448_
	);
	LUT4 #(
		.INIT('h0400)
	) name29622 (
		_w15291_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35449_
	);
	LUT4 #(
		.INIT('he5ff)
	) name29623 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35450_
	);
	LUT4 #(
		.INIT('h3100)
	) name29624 (
		_w15291_,
		_w35449_,
		_w35448_,
		_w35450_,
		_w35451_
	);
	LUT3 #(
		.INIT('h40)
	) name29625 (
		_w35446_,
		_w35447_,
		_w35451_,
		_w35452_
	);
	LUT4 #(
		.INIT('h5545)
	) name29626 (
		_w15291_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35453_
	);
	LUT4 #(
		.INIT('haa2a)
	) name29627 (
		_w15291_,
		_w15292_,
		_w15293_,
		_w15295_,
		_w35454_
	);
	LUT4 #(
		.INIT('h5fbb)
	) name29628 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35455_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name29629 (
		_w15306_,
		_w35453_,
		_w35454_,
		_w35455_,
		_w35456_
	);
	LUT4 #(
		.INIT('h2100)
	) name29630 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35457_
	);
	LUT3 #(
		.INIT('h02)
	) name29631 (
		_w15299_,
		_w15315_,
		_w35457_,
		_w35458_
	);
	LUT2 #(
		.INIT('h4)
	) name29632 (
		_w35456_,
		_w35458_,
		_w35459_
	);
	LUT4 #(
		.INIT('h0002)
	) name29633 (
		_w15291_,
		_w15292_,
		_w15295_,
		_w15294_,
		_w35460_
	);
	LUT3 #(
		.INIT('h07)
	) name29634 (
		_w15301_,
		_w35258_,
		_w35460_,
		_w35461_
	);
	LUT4 #(
		.INIT('ha955)
	) name29635 (
		\u1_L14_reg[21]/P0001 ,
		_w35452_,
		_w35459_,
		_w35461_,
		_w35462_
	);
	LUT2 #(
		.INIT('h1)
	) name29636 (
		_w15387_,
		_w15393_,
		_w35463_
	);
	LUT4 #(
		.INIT('hefad)
	) name29637 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35464_
	);
	LUT3 #(
		.INIT('h40)
	) name29638 (
		_w35343_,
		_w35463_,
		_w35464_,
		_w35465_
	);
	LUT4 #(
		.INIT('haaa8)
	) name29639 (
		_w15393_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35466_
	);
	LUT4 #(
		.INIT('h5515)
	) name29640 (
		_w15393_,
		_w15388_,
		_w15389_,
		_w15391_,
		_w35467_
	);
	LUT4 #(
		.INIT('h8caf)
	) name29641 (
		_w35234_,
		_w35353_,
		_w35466_,
		_w35467_,
		_w35468_
	);
	LUT4 #(
		.INIT('h0002)
	) name29642 (
		_w15387_,
		_w15405_,
		_w35235_,
		_w35236_,
		_w35469_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name29643 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35470_
	);
	LUT4 #(
		.INIT('hba00)
	) name29644 (
		_w35465_,
		_w35468_,
		_w35469_,
		_w35470_,
		_w35471_
	);
	LUT4 #(
		.INIT('h0064)
	) name29645 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35472_
	);
	LUT4 #(
		.INIT('h8a00)
	) name29646 (
		_w15388_,
		_w15389_,
		_w15391_,
		_w15392_,
		_w35473_
	);
	LUT2 #(
		.INIT('h4)
	) name29647 (
		_w15387_,
		_w15393_,
		_w35474_
	);
	LUT4 #(
		.INIT('h0100)
	) name29648 (
		_w35356_,
		_w35472_,
		_w35473_,
		_w35474_,
		_w35475_
	);
	LUT3 #(
		.INIT('h56)
	) name29649 (
		\u1_L14_reg[13]/P0001 ,
		_w35471_,
		_w35475_,
		_w35476_
	);
	LUT3 #(
		.INIT('h23)
	) name29650 (
		_w15291_,
		_w15299_,
		_w35268_,
		_w35477_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name29651 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35478_
	);
	LUT4 #(
		.INIT('h4554)
	) name29652 (
		_w15291_,
		_w15292_,
		_w15295_,
		_w15294_,
		_w35479_
	);
	LUT4 #(
		.INIT('h4457)
	) name29653 (
		_w15291_,
		_w35268_,
		_w35478_,
		_w35479_,
		_w35480_
	);
	LUT3 #(
		.INIT('h32)
	) name29654 (
		_w15316_,
		_w35477_,
		_w35480_,
		_w35481_
	);
	LUT4 #(
		.INIT('hebfb)
	) name29655 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35482_
	);
	LUT2 #(
		.INIT('h2)
	) name29656 (
		_w15291_,
		_w35482_,
		_w35483_
	);
	LUT3 #(
		.INIT('h45)
	) name29657 (
		_w15293_,
		_w15295_,
		_w15294_,
		_w35484_
	);
	LUT3 #(
		.INIT('h45)
	) name29658 (
		_w15291_,
		_w15292_,
		_w15293_,
		_w35485_
	);
	LUT2 #(
		.INIT('h4)
	) name29659 (
		_w35484_,
		_w35485_,
		_w35486_
	);
	LUT4 #(
		.INIT('h8000)
	) name29660 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35487_
	);
	LUT3 #(
		.INIT('ha2)
	) name29661 (
		_w15291_,
		_w15292_,
		_w15293_,
		_w35488_
	);
	LUT3 #(
		.INIT('h31)
	) name29662 (
		_w15297_,
		_w35487_,
		_w35488_,
		_w35489_
	);
	LUT4 #(
		.INIT('h5455)
	) name29663 (
		_w15299_,
		_w35483_,
		_w35486_,
		_w35489_,
		_w35490_
	);
	LUT4 #(
		.INIT('hf9be)
	) name29664 (
		_w15292_,
		_w15293_,
		_w15295_,
		_w15294_,
		_w35491_
	);
	LUT2 #(
		.INIT('h2)
	) name29665 (
		_w15291_,
		_w35491_,
		_w35492_
	);
	LUT4 #(
		.INIT('haaa9)
	) name29666 (
		\u1_L14_reg[5]/P0001 ,
		_w35490_,
		_w35481_,
		_w35492_,
		_w35493_
	);
	LUT4 #(
		.INIT('h00ef)
	) name29667 (
		_w35377_,
		_w35378_,
		_w35376_,
		_w35382_,
		_w35494_
	);
	LUT4 #(
		.INIT('hf310)
	) name29668 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35495_
	);
	LUT2 #(
		.INIT('h8)
	) name29669 (
		_w35494_,
		_w35495_,
		_w35496_
	);
	LUT3 #(
		.INIT('h02)
	) name29670 (
		_w35378_,
		_w35375_,
		_w35376_,
		_w35497_
	);
	LUT2 #(
		.INIT('h4)
	) name29671 (
		_w35391_,
		_w35497_,
		_w35498_
	);
	LUT2 #(
		.INIT('h1)
	) name29672 (
		_w35377_,
		_w35375_,
		_w35499_
	);
	LUT2 #(
		.INIT('h8)
	) name29673 (
		_w35376_,
		_w35382_,
		_w35500_
	);
	LUT3 #(
		.INIT('h3b)
	) name29674 (
		_w35378_,
		_w35376_,
		_w35382_,
		_w35501_
	);
	LUT4 #(
		.INIT('h8000)
	) name29675 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35502_
	);
	LUT3 #(
		.INIT('h0d)
	) name29676 (
		_w35499_,
		_w35501_,
		_w35502_,
		_w35503_
	);
	LUT4 #(
		.INIT('h5455)
	) name29677 (
		_w35386_,
		_w35496_,
		_w35498_,
		_w35503_,
		_w35504_
	);
	LUT4 #(
		.INIT('hf070)
	) name29678 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35505_
	);
	LUT4 #(
		.INIT('h0048)
	) name29679 (
		_w35377_,
		_w35378_,
		_w35376_,
		_w35382_,
		_w35506_
	);
	LUT2 #(
		.INIT('h4)
	) name29680 (
		_w35505_,
		_w35506_,
		_w35507_
	);
	LUT2 #(
		.INIT('h6)
	) name29681 (
		_w35377_,
		_w35375_,
		_w35508_
	);
	LUT4 #(
		.INIT('he000)
	) name29682 (
		_w35378_,
		_w35375_,
		_w35376_,
		_w35382_,
		_w35509_
	);
	LUT4 #(
		.INIT('hffbe)
	) name29683 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35510_
	);
	LUT3 #(
		.INIT('h70)
	) name29684 (
		_w35508_,
		_w35509_,
		_w35510_,
		_w35511_
	);
	LUT4 #(
		.INIT('h0060)
	) name29685 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35512_
	);
	LUT4 #(
		.INIT('hee9f)
	) name29686 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35513_
	);
	LUT4 #(
		.INIT('h0100)
	) name29687 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35382_,
		_w35514_
	);
	LUT2 #(
		.INIT('h6)
	) name29688 (
		_w35375_,
		_w35376_,
		_w35515_
	);
	LUT4 #(
		.INIT('h0082)
	) name29689 (
		_w35377_,
		_w35375_,
		_w35376_,
		_w35382_,
		_w35516_
	);
	LUT4 #(
		.INIT('h0031)
	) name29690 (
		_w35382_,
		_w35514_,
		_w35513_,
		_w35516_,
		_w35517_
	);
	LUT4 #(
		.INIT('h7500)
	) name29691 (
		_w35386_,
		_w35507_,
		_w35511_,
		_w35517_,
		_w35518_
	);
	LUT3 #(
		.INIT('h65)
	) name29692 (
		\u1_L14_reg[22]/P0001 ,
		_w35504_,
		_w35518_,
		_w35519_
	);
	LUT3 #(
		.INIT('h01)
	) name29693 (
		_w35168_,
		_w35167_,
		_w35169_,
		_w35520_
	);
	LUT3 #(
		.INIT('h80)
	) name29694 (
		_w35168_,
		_w35172_,
		_w35169_,
		_w35521_
	);
	LUT4 #(
		.INIT('hfb00)
	) name29695 (
		_w35172_,
		_w35167_,
		_w35169_,
		_w35171_,
		_w35522_
	);
	LUT3 #(
		.INIT('h10)
	) name29696 (
		_w35520_,
		_w35521_,
		_w35522_,
		_w35523_
	);
	LUT3 #(
		.INIT('h40)
	) name29697 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35524_
	);
	LUT4 #(
		.INIT('h00fd)
	) name29698 (
		_w35168_,
		_w35167_,
		_w35169_,
		_w35171_,
		_w35525_
	);
	LUT4 #(
		.INIT('hdeff)
	) name29699 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35526_
	);
	LUT3 #(
		.INIT('h40)
	) name29700 (
		_w35524_,
		_w35525_,
		_w35526_,
		_w35527_
	);
	LUT4 #(
		.INIT('h0010)
	) name29701 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35528_
	);
	LUT3 #(
		.INIT('h01)
	) name29702 (
		_w35180_,
		_w35327_,
		_w35528_,
		_w35529_
	);
	LUT3 #(
		.INIT('he0)
	) name29703 (
		_w35523_,
		_w35527_,
		_w35529_,
		_w35530_
	);
	LUT3 #(
		.INIT('hea)
	) name29704 (
		_w35168_,
		_w35167_,
		_w35169_,
		_w35531_
	);
	LUT3 #(
		.INIT('h40)
	) name29705 (
		_w35521_,
		_w35522_,
		_w35531_,
		_w35532_
	);
	LUT3 #(
		.INIT('hf6)
	) name29706 (
		_w35168_,
		_w35167_,
		_w35169_,
		_w35533_
	);
	LUT2 #(
		.INIT('h1)
	) name29707 (
		_w35172_,
		_w35171_,
		_w35534_
	);
	LUT2 #(
		.INIT('h4)
	) name29708 (
		_w35533_,
		_w35534_,
		_w35535_
	);
	LUT3 #(
		.INIT('h02)
	) name29709 (
		_w35180_,
		_w35326_,
		_w35339_,
		_w35536_
	);
	LUT4 #(
		.INIT('h0200)
	) name29710 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35537_
	);
	LUT3 #(
		.INIT('h07)
	) name29711 (
		_w35174_,
		_w35190_,
		_w35537_,
		_w35538_
	);
	LUT4 #(
		.INIT('h1000)
	) name29712 (
		_w35535_,
		_w35532_,
		_w35536_,
		_w35538_,
		_w35539_
	);
	LUT4 #(
		.INIT('h0048)
	) name29713 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35540_
	);
	LUT4 #(
		.INIT('heffb)
	) name29714 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35541_
	);
	LUT3 #(
		.INIT('hb1)
	) name29715 (
		_w35171_,
		_w35540_,
		_w35541_,
		_w35542_
	);
	LUT4 #(
		.INIT('ha955)
	) name29716 (
		\u1_L14_reg[14]/P0001 ,
		_w35530_,
		_w35539_,
		_w35542_,
		_w35543_
	);
	LUT4 #(
		.INIT('h0800)
	) name29717 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35544_
	);
	LUT4 #(
		.INIT('h0200)
	) name29718 (
		_w15358_,
		_w15355_,
		_w15354_,
		_w15360_,
		_w35545_
	);
	LUT3 #(
		.INIT('h01)
	) name29719 (
		_w15353_,
		_w35545_,
		_w35544_,
		_w35546_
	);
	LUT2 #(
		.INIT('h8)
	) name29720 (
		_w15369_,
		_w15380_,
		_w35547_
	);
	LUT4 #(
		.INIT('h4182)
	) name29721 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35548_
	);
	LUT4 #(
		.INIT('h0405)
	) name29722 (
		_w15358_,
		_w15355_,
		_w15354_,
		_w15360_,
		_w35549_
	);
	LUT3 #(
		.INIT('h13)
	) name29723 (
		_w15372_,
		_w35548_,
		_w35549_,
		_w35550_
	);
	LUT3 #(
		.INIT('h31)
	) name29724 (
		_w15358_,
		_w15355_,
		_w15354_,
		_w35551_
	);
	LUT3 #(
		.INIT('h09)
	) name29725 (
		_w15358_,
		_w15356_,
		_w15360_,
		_w35552_
	);
	LUT4 #(
		.INIT('h0200)
	) name29726 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35553_
	);
	LUT4 #(
		.INIT('h2022)
	) name29727 (
		_w15353_,
		_w35553_,
		_w35551_,
		_w35552_,
		_w35554_
	);
	LUT4 #(
		.INIT('h00bf)
	) name29728 (
		_w35547_,
		_w35546_,
		_w35550_,
		_w35554_,
		_w35555_
	);
	LUT4 #(
		.INIT('h87a7)
	) name29729 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35556_
	);
	LUT4 #(
		.INIT('h0001)
	) name29730 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35557_
	);
	LUT4 #(
		.INIT('haffe)
	) name29731 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35558_
	);
	LUT4 #(
		.INIT('h08cc)
	) name29732 (
		_w15353_,
		_w15360_,
		_w35556_,
		_w35558_,
		_w35559_
	);
	LUT3 #(
		.INIT('h56)
	) name29733 (
		\u1_L14_reg[6]/P0001 ,
		_w35555_,
		_w35559_,
		_w35560_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name29734 (
		_w15321_,
		_w15322_,
		_w15324_,
		_w15323_,
		_w35561_
	);
	LUT2 #(
		.INIT('h4)
	) name29735 (
		_w15343_,
		_w35561_,
		_w35562_
	);
	LUT4 #(
		.INIT('h0051)
	) name29736 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35563_
	);
	LUT3 #(
		.INIT('h01)
	) name29737 (
		_w15321_,
		_w15327_,
		_w35563_,
		_w35564_
	);
	LUT4 #(
		.INIT('hff7c)
	) name29738 (
		_w15321_,
		_w15322_,
		_w15324_,
		_w15323_,
		_w35565_
	);
	LUT3 #(
		.INIT('h31)
	) name29739 (
		_w15325_,
		_w15346_,
		_w35565_,
		_w35566_
	);
	LUT4 #(
		.INIT('h0155)
	) name29740 (
		_w15331_,
		_w35562_,
		_w35564_,
		_w35566_,
		_w35567_
	);
	LUT4 #(
		.INIT('hf3d1)
	) name29741 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35568_
	);
	LUT2 #(
		.INIT('h2)
	) name29742 (
		_w15321_,
		_w35568_,
		_w35569_
	);
	LUT4 #(
		.INIT('hfe00)
	) name29743 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35570_
	);
	LUT3 #(
		.INIT('hd0)
	) name29744 (
		_w15321_,
		_w15322_,
		_w15325_,
		_w35571_
	);
	LUT4 #(
		.INIT('haff3)
	) name29745 (
		_w15321_,
		_w15322_,
		_w15325_,
		_w15323_,
		_w35572_
	);
	LUT4 #(
		.INIT('hfe00)
	) name29746 (
		_w15328_,
		_w35571_,
		_w35570_,
		_w35572_,
		_w35573_
	);
	LUT3 #(
		.INIT('h8a)
	) name29747 (
		_w15331_,
		_w35569_,
		_w35573_,
		_w35574_
	);
	LUT4 #(
		.INIT('h6fe7)
	) name29748 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35575_
	);
	LUT2 #(
		.INIT('h1)
	) name29749 (
		_w15321_,
		_w35575_,
		_w35576_
	);
	LUT3 #(
		.INIT('h07)
	) name29750 (
		_w15326_,
		_w15335_,
		_w15349_,
		_w35577_
	);
	LUT2 #(
		.INIT('h4)
	) name29751 (
		_w35576_,
		_w35577_,
		_w35578_
	);
	LUT4 #(
		.INIT('h5655)
	) name29752 (
		\u1_L14_reg[31]/P0001 ,
		_w35574_,
		_w35567_,
		_w35578_,
		_w35579_
	);
	LUT4 #(
		.INIT('hd3c3)
	) name29753 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35580_
	);
	LUT4 #(
		.INIT('h1555)
	) name29754 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35581_
	);
	LUT4 #(
		.INIT('h4802)
	) name29755 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35582_
	);
	LUT3 #(
		.INIT('he6)
	) name29756 (
		_w15324_,
		_w15325_,
		_w15323_,
		_w35583_
	);
	LUT4 #(
		.INIT('h0e04)
	) name29757 (
		_w15321_,
		_w35583_,
		_w35582_,
		_w35580_,
		_w35584_
	);
	LUT4 #(
		.INIT('h8228)
	) name29758 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35585_
	);
	LUT4 #(
		.INIT('h0501)
	) name29759 (
		_w15332_,
		_w15350_,
		_w35585_,
		_w35583_,
		_w35586_
	);
	LUT4 #(
		.INIT('haa2a)
	) name29760 (
		_w15322_,
		_w15324_,
		_w15325_,
		_w15323_,
		_w35587_
	);
	LUT3 #(
		.INIT('h01)
	) name29761 (
		_w15321_,
		_w35581_,
		_w35587_,
		_w35588_
	);
	LUT4 #(
		.INIT('h00d8)
	) name29762 (
		_w15331_,
		_w35586_,
		_w35584_,
		_w35588_,
		_w35589_
	);
	LUT2 #(
		.INIT('h9)
	) name29763 (
		\u1_L14_reg[9]/P0001 ,
		_w35589_,
		_w35590_
	);
	LUT4 #(
		.INIT('h134c)
	) name29764 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35591_
	);
	LUT4 #(
		.INIT('h2c82)
	) name29765 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35592_
	);
	LUT2 #(
		.INIT('h4)
	) name29766 (
		_w35382_,
		_w35386_,
		_w35593_
	);
	LUT2 #(
		.INIT('h9)
	) name29767 (
		_w35382_,
		_w35386_,
		_w35594_
	);
	LUT3 #(
		.INIT('h10)
	) name29768 (
		_w35379_,
		_w35592_,
		_w35594_,
		_w35595_
	);
	LUT4 #(
		.INIT('hfb00)
	) name29769 (
		_w35378_,
		_w35375_,
		_w35376_,
		_w35382_,
		_w35596_
	);
	LUT4 #(
		.INIT('h0100)
	) name29770 (
		_w35386_,
		_w35502_,
		_w35591_,
		_w35596_,
		_w35597_
	);
	LUT4 #(
		.INIT('h0010)
	) name29771 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35598_
	);
	LUT3 #(
		.INIT('h09)
	) name29772 (
		_w35377_,
		_w35375_,
		_w35376_,
		_w35599_
	);
	LUT3 #(
		.INIT('h28)
	) name29773 (
		_w35377_,
		_w35378_,
		_w35376_,
		_w35600_
	);
	LUT4 #(
		.INIT('h7000)
	) name29774 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35601_
	);
	LUT4 #(
		.INIT('h0002)
	) name29775 (
		_w35593_,
		_w35601_,
		_w35600_,
		_w35599_,
		_w35602_
	);
	LUT4 #(
		.INIT('h00f1)
	) name29776 (
		_w35595_,
		_w35597_,
		_w35598_,
		_w35602_,
		_w35603_
	);
	LUT2 #(
		.INIT('h6)
	) name29777 (
		\u1_L14_reg[7]/P0001 ,
		_w35603_,
		_w35604_
	);
	LUT4 #(
		.INIT('h0104)
	) name29778 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35605_
	);
	LUT4 #(
		.INIT('h00fd)
	) name29779 (
		_w35377_,
		_w35378_,
		_w35376_,
		_w35382_,
		_w35606_
	);
	LUT3 #(
		.INIT('h10)
	) name29780 (
		_w35394_,
		_w35605_,
		_w35606_,
		_w35607_
	);
	LUT3 #(
		.INIT('hb8)
	) name29781 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35608_
	);
	LUT4 #(
		.INIT('h3808)
	) name29782 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35609_
	);
	LUT4 #(
		.INIT('hfe00)
	) name29783 (
		_w35377_,
		_w35378_,
		_w35376_,
		_w35382_,
		_w35610_
	);
	LUT2 #(
		.INIT('h4)
	) name29784 (
		_w35609_,
		_w35610_,
		_w35611_
	);
	LUT4 #(
		.INIT('h2000)
	) name29785 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35612_
	);
	LUT2 #(
		.INIT('h2)
	) name29786 (
		_w35386_,
		_w35612_,
		_w35613_
	);
	LUT3 #(
		.INIT('he0)
	) name29787 (
		_w35607_,
		_w35611_,
		_w35613_,
		_w35614_
	);
	LUT3 #(
		.INIT('h10)
	) name29788 (
		_w35378_,
		_w35375_,
		_w35376_,
		_w35615_
	);
	LUT3 #(
		.INIT('h09)
	) name29789 (
		_w35377_,
		_w35378_,
		_w35382_,
		_w35616_
	);
	LUT2 #(
		.INIT('h4)
	) name29790 (
		_w35615_,
		_w35616_,
		_w35617_
	);
	LUT3 #(
		.INIT('h01)
	) name29791 (
		_w35386_,
		_w35502_,
		_w35512_,
		_w35618_
	);
	LUT4 #(
		.INIT('h0200)
	) name29792 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35376_,
		_w35619_
	);
	LUT3 #(
		.INIT('h0d)
	) name29793 (
		_w35500_,
		_w35608_,
		_w35619_,
		_w35620_
	);
	LUT3 #(
		.INIT('h40)
	) name29794 (
		_w35617_,
		_w35618_,
		_w35620_,
		_w35621_
	);
	LUT4 #(
		.INIT('h00a8)
	) name29795 (
		_w35377_,
		_w35378_,
		_w35375_,
		_w35382_,
		_w35622_
	);
	LUT4 #(
		.INIT('h0777)
	) name29796 (
		_w35385_,
		_w35382_,
		_w35515_,
		_w35622_,
		_w35623_
	);
	LUT4 #(
		.INIT('ha955)
	) name29797 (
		\u1_L14_reg[32]/P0001 ,
		_w35614_,
		_w35621_,
		_w35623_,
		_w35624_
	);
	LUT4 #(
		.INIT('hb8cd)
	) name29798 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35625_
	);
	LUT4 #(
		.INIT('h0400)
	) name29799 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35626_
	);
	LUT4 #(
		.INIT('h5504)
	) name29800 (
		_w15353_,
		_w15360_,
		_w35625_,
		_w35626_,
		_w35627_
	);
	LUT4 #(
		.INIT('hc7b6)
	) name29801 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35628_
	);
	LUT3 #(
		.INIT('h54)
	) name29802 (
		_w15353_,
		_w15360_,
		_w35628_,
		_w35629_
	);
	LUT3 #(
		.INIT('h2a)
	) name29803 (
		_w15353_,
		_w15372_,
		_w35549_,
		_w35630_
	);
	LUT3 #(
		.INIT('h0e)
	) name29804 (
		_w15358_,
		_w15354_,
		_w15360_,
		_w35631_
	);
	LUT2 #(
		.INIT('h4)
	) name29805 (
		_w15372_,
		_w35631_,
		_w35632_
	);
	LUT2 #(
		.INIT('h4)
	) name29806 (
		_w15354_,
		_w15360_,
		_w35633_
	);
	LUT3 #(
		.INIT('h45)
	) name29807 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w35634_
	);
	LUT3 #(
		.INIT('he0)
	) name29808 (
		_w15355_,
		_w15356_,
		_w15360_,
		_w35635_
	);
	LUT3 #(
		.INIT('hb0)
	) name29809 (
		_w15358_,
		_w15355_,
		_w15354_,
		_w35636_
	);
	LUT4 #(
		.INIT('h0777)
	) name29810 (
		_w35633_,
		_w35634_,
		_w35635_,
		_w35636_,
		_w35637_
	);
	LUT4 #(
		.INIT('h4555)
	) name29811 (
		_w35629_,
		_w35632_,
		_w35630_,
		_w35637_,
		_w35638_
	);
	LUT3 #(
		.INIT('h80)
	) name29812 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w35639_
	);
	LUT3 #(
		.INIT('hdb)
	) name29813 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w35640_
	);
	LUT4 #(
		.INIT('hdf9b)
	) name29814 (
		_w15354_,
		_w15360_,
		_w35639_,
		_w35640_,
		_w35641_
	);
	LUT4 #(
		.INIT('h5655)
	) name29815 (
		\u1_L14_reg[24]/P0001 ,
		_w35638_,
		_w35627_,
		_w35641_,
		_w35642_
	);
	LUT4 #(
		.INIT('hdf00)
	) name29816 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35643_
	);
	LUT3 #(
		.INIT('h90)
	) name29817 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w35644_
	);
	LUT4 #(
		.INIT('h0200)
	) name29818 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15360_,
		_w35645_
	);
	LUT4 #(
		.INIT('h00fb)
	) name29819 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35646_
	);
	LUT4 #(
		.INIT('h5455)
	) name29820 (
		_w35643_,
		_w35644_,
		_w35645_,
		_w35646_,
		_w35647_
	);
	LUT4 #(
		.INIT('h0012)
	) name29821 (
		_w15355_,
		_w15356_,
		_w15354_,
		_w15360_,
		_w35648_
	);
	LUT3 #(
		.INIT('ha8)
	) name29822 (
		_w15353_,
		_w35647_,
		_w35648_,
		_w35649_
	);
	LUT4 #(
		.INIT('h6f6c)
	) name29823 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35650_
	);
	LUT4 #(
		.INIT('h6800)
	) name29824 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15360_,
		_w35651_
	);
	LUT4 #(
		.INIT('h0032)
	) name29825 (
		_w15360_,
		_w35557_,
		_w35650_,
		_w35651_,
		_w35652_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name29826 (
		_w15358_,
		_w15355_,
		_w15356_,
		_w15354_,
		_w35653_
	);
	LUT4 #(
		.INIT('h0040)
	) name29827 (
		_w15358_,
		_w15355_,
		_w15354_,
		_w15360_,
		_w35654_
	);
	LUT3 #(
		.INIT('h0d)
	) name29828 (
		_w15360_,
		_w35653_,
		_w35654_,
		_w35655_
	);
	LUT3 #(
		.INIT('he0)
	) name29829 (
		_w15353_,
		_w35652_,
		_w35655_,
		_w35656_
	);
	LUT3 #(
		.INIT('h65)
	) name29830 (
		\u1_L14_reg[16]/P0001 ,
		_w35649_,
		_w35656_,
		_w35657_
	);
	LUT4 #(
		.INIT('hf55d)
	) name29831 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35658_
	);
	LUT4 #(
		.INIT('h5eff)
	) name29832 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35659_
	);
	LUT4 #(
		.INIT('hbfcb)
	) name29833 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35660_
	);
	LUT4 #(
		.INIT('hd800)
	) name29834 (
		_w35171_,
		_w35659_,
		_w35658_,
		_w35660_,
		_w35661_
	);
	LUT4 #(
		.INIT('hf5fe)
	) name29835 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35662_
	);
	LUT3 #(
		.INIT('h04)
	) name29836 (
		_w35172_,
		_w35169_,
		_w35171_,
		_w35663_
	);
	LUT4 #(
		.INIT('h0031)
	) name29837 (
		_w35171_,
		_w35540_,
		_w35662_,
		_w35663_,
		_w35664_
	);
	LUT4 #(
		.INIT('hbf9f)
	) name29838 (
		_w35168_,
		_w35172_,
		_w35167_,
		_w35169_,
		_w35665_
	);
	LUT4 #(
		.INIT('hd8fa)
	) name29839 (
		_w35171_,
		_w35322_,
		_w35339_,
		_w35665_,
		_w35666_
	);
	LUT4 #(
		.INIT('h0d08)
	) name29840 (
		_w35180_,
		_w35664_,
		_w35666_,
		_w35661_,
		_w35667_
	);
	LUT2 #(
		.INIT('h9)
	) name29841 (
		\u1_L14_reg[8]/P0001 ,
		_w35667_,
		_w35668_
	);
	LUT3 #(
		.INIT('h01)
	) name29842 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35669_
	);
	LUT3 #(
		.INIT('h02)
	) name29843 (
		_w35197_,
		_w35371_,
		_w35669_,
		_w35670_
	);
	LUT3 #(
		.INIT('h04)
	) name29844 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35671_
	);
	LUT4 #(
		.INIT('h00f7)
	) name29845 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35197_,
		_w35672_
	);
	LUT2 #(
		.INIT('h4)
	) name29846 (
		_w35671_,
		_w35672_,
		_w35673_
	);
	LUT4 #(
		.INIT('h0400)
	) name29847 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35674_
	);
	LUT4 #(
		.INIT('h0001)
	) name29848 (
		_w35195_,
		_w35213_,
		_w35216_,
		_w35674_,
		_w35675_
	);
	LUT3 #(
		.INIT('he0)
	) name29849 (
		_w35670_,
		_w35673_,
		_w35675_,
		_w35676_
	);
	LUT3 #(
		.INIT('h02)
	) name29850 (
		_w35196_,
		_w35198_,
		_w35199_,
		_w35677_
	);
	LUT2 #(
		.INIT('h2)
	) name29851 (
		_w35365_,
		_w35677_,
		_w35678_
	);
	LUT3 #(
		.INIT('h20)
	) name29852 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35679_
	);
	LUT4 #(
		.INIT('h0b00)
	) name29853 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35680_
	);
	LUT3 #(
		.INIT('h01)
	) name29854 (
		_w35197_,
		_w35680_,
		_w35679_,
		_w35681_
	);
	LUT4 #(
		.INIT('h4000)
	) name29855 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35682_
	);
	LUT3 #(
		.INIT('h02)
	) name29856 (
		_w35195_,
		_w35214_,
		_w35682_,
		_w35683_
	);
	LUT3 #(
		.INIT('he0)
	) name29857 (
		_w35678_,
		_w35681_,
		_w35683_,
		_w35684_
	);
	LUT4 #(
		.INIT('h6fdf)
	) name29858 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35685_
	);
	LUT2 #(
		.INIT('h2)
	) name29859 (
		_w35197_,
		_w35685_,
		_w35686_
	);
	LUT4 #(
		.INIT('hccdf)
	) name29860 (
		_w35198_,
		_w35197_,
		_w35205_,
		_w35682_,
		_w35687_
	);
	LUT2 #(
		.INIT('h4)
	) name29861 (
		_w35686_,
		_w35687_,
		_w35688_
	);
	LUT4 #(
		.INIT('ha955)
	) name29862 (
		\u1_L14_reg[1]/P0001 ,
		_w35676_,
		_w35684_,
		_w35688_,
		_w35689_
	);
	LUT4 #(
		.INIT('h006b)
	) name29863 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35197_,
		_w35690_
	);
	LUT4 #(
		.INIT('hd700)
	) name29864 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35197_,
		_w35691_
	);
	LUT3 #(
		.INIT('h01)
	) name29865 (
		_w35198_,
		_w35691_,
		_w35690_,
		_w35692_
	);
	LUT4 #(
		.INIT('h0100)
	) name29866 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35693_
	);
	LUT4 #(
		.INIT('h0100)
	) name29867 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35197_,
		_w35694_
	);
	LUT4 #(
		.INIT('h0002)
	) name29868 (
		_w35195_,
		_w35682_,
		_w35693_,
		_w35694_,
		_w35695_
	);
	LUT4 #(
		.INIT('h7f7d)
	) name29869 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35696_
	);
	LUT4 #(
		.INIT('hdddf)
	) name29870 (
		_w35200_,
		_w35196_,
		_w35199_,
		_w35197_,
		_w35697_
	);
	LUT4 #(
		.INIT('hfc54)
	) name29871 (
		_w35198_,
		_w35197_,
		_w35696_,
		_w35697_,
		_w35698_
	);
	LUT2 #(
		.INIT('h8)
	) name29872 (
		_w35695_,
		_w35698_,
		_w35699_
	);
	LUT4 #(
		.INIT('hff8a)
	) name29873 (
		_w35200_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35700_
	);
	LUT2 #(
		.INIT('h1)
	) name29874 (
		_w35197_,
		_w35700_,
		_w35701_
	);
	LUT2 #(
		.INIT('h4)
	) name29875 (
		_w35207_,
		_w35221_,
		_w35702_
	);
	LUT4 #(
		.INIT('h5551)
	) name29876 (
		_w35195_,
		_w35196_,
		_w35198_,
		_w35199_,
		_w35703_
	);
	LUT3 #(
		.INIT('h10)
	) name29877 (
		_w35216_,
		_w35223_,
		_w35703_,
		_w35704_
	);
	LUT3 #(
		.INIT('h10)
	) name29878 (
		_w35701_,
		_w35702_,
		_w35704_,
		_w35705_
	);
	LUT4 #(
		.INIT('h6665)
	) name29879 (
		\u1_L14_reg[26]/P0001 ,
		_w35692_,
		_w35699_,
		_w35705_,
		_w35706_
	);
	LUT4 #(
		.INIT('hc963)
	) name29880 (
		decrypt_pad,
		\u2_R14_reg[20]/NET0131 ,
		\u2_uk_K_r14_reg[16]/NET0131 ,
		\u2_uk_K_r14_reg[23]/NET0131 ,
		_w35707_
	);
	LUT4 #(
		.INIT('hc963)
	) name29881 (
		decrypt_pad,
		\u2_R14_reg[19]/P0001 ,
		\u2_uk_K_r14_reg[1]/NET0131 ,
		\u2_uk_K_r14_reg[8]/NET0131 ,
		_w35708_
	);
	LUT4 #(
		.INIT('hc693)
	) name29882 (
		decrypt_pad,
		\u2_R14_reg[17]/NET0131 ,
		\u2_uk_K_r14_reg[31]/NET0131 ,
		\u2_uk_K_r14_reg[51]/NET0131 ,
		_w35709_
	);
	LUT4 #(
		.INIT('hc963)
	) name29883 (
		decrypt_pad,
		\u2_R14_reg[16]/NET0131 ,
		\u2_uk_K_r14_reg[29]/NET0131 ,
		\u2_uk_K_r14_reg[36]/NET0131 ,
		_w35710_
	);
	LUT4 #(
		.INIT('hc963)
	) name29884 (
		decrypt_pad,
		\u2_R14_reg[21]/NET0131 ,
		\u2_uk_K_r14_reg[45]/NET0131 ,
		\u2_uk_K_r14_reg[52]/NET0131 ,
		_w35711_
	);
	LUT4 #(
		.INIT('h00bf)
	) name29885 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35708_,
		_w35712_
	);
	LUT4 #(
		.INIT('hc963)
	) name29886 (
		decrypt_pad,
		\u2_R14_reg[18]/NET0131 ,
		\u2_uk_K_r14_reg[14]/NET0131 ,
		\u2_uk_K_r14_reg[21]/NET0131 ,
		_w35713_
	);
	LUT3 #(
		.INIT('h02)
	) name29887 (
		_w35709_,
		_w35710_,
		_w35713_,
		_w35714_
	);
	LUT4 #(
		.INIT('h0305)
	) name29888 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35715_
	);
	LUT4 #(
		.INIT('h7f00)
	) name29889 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35708_,
		_w35716_
	);
	LUT4 #(
		.INIT('h6e00)
	) name29890 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35708_,
		_w35717_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name29891 (
		_w35712_,
		_w35714_,
		_w35715_,
		_w35717_,
		_w35718_
	);
	LUT4 #(
		.INIT('h08a0)
	) name29892 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35719_
	);
	LUT3 #(
		.INIT('ha8)
	) name29893 (
		_w35707_,
		_w35718_,
		_w35719_,
		_w35720_
	);
	LUT4 #(
		.INIT('hbcaf)
	) name29894 (
		_w35710_,
		_w35711_,
		_w35713_,
		_w35708_,
		_w35721_
	);
	LUT3 #(
		.INIT('h08)
	) name29895 (
		_w35710_,
		_w35711_,
		_w35713_,
		_w35722_
	);
	LUT4 #(
		.INIT('haa02)
	) name29896 (
		_w35709_,
		_w35707_,
		_w35721_,
		_w35722_,
		_w35723_
	);
	LUT3 #(
		.INIT('h08)
	) name29897 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35724_
	);
	LUT4 #(
		.INIT('h0900)
	) name29898 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35725_
	);
	LUT2 #(
		.INIT('h8)
	) name29899 (
		_w35725_,
		_w35708_,
		_w35726_
	);
	LUT4 #(
		.INIT('h0007)
	) name29900 (
		_w35710_,
		_w35711_,
		_w35713_,
		_w35707_,
		_w35727_
	);
	LUT3 #(
		.INIT('h07)
	) name29901 (
		_w35710_,
		_w35713_,
		_w35708_,
		_w35728_
	);
	LUT4 #(
		.INIT('hfb00)
	) name29902 (
		_w35710_,
		_w35711_,
		_w35713_,
		_w35708_,
		_w35729_
	);
	LUT4 #(
		.INIT('h1011)
	) name29903 (
		_w35709_,
		_w35729_,
		_w35727_,
		_w35728_,
		_w35730_
	);
	LUT3 #(
		.INIT('h01)
	) name29904 (
		_w35726_,
		_w35723_,
		_w35730_,
		_w35731_
	);
	LUT3 #(
		.INIT('h65)
	) name29905 (
		\u2_L14_reg[25]/P0001 ,
		_w35720_,
		_w35731_,
		_w35732_
	);
	LUT4 #(
		.INIT('hc963)
	) name29906 (
		decrypt_pad,
		\u2_R14_reg[8]/NET0131 ,
		\u2_uk_K_r14_reg[32]/NET0131 ,
		\u2_uk_K_r14_reg[39]/P0001 ,
		_w35733_
	);
	LUT4 #(
		.INIT('hc963)
	) name29907 (
		decrypt_pad,
		\u2_R14_reg[7]/P0001 ,
		\u2_uk_K_r14_reg[41]/NET0131 ,
		\u2_uk_K_r14_reg[48]/NET0131 ,
		_w35734_
	);
	LUT4 #(
		.INIT('hc963)
	) name29908 (
		decrypt_pad,
		\u2_R14_reg[5]/NET0131 ,
		\u2_uk_K_r14_reg[24]/NET0131 ,
		\u2_uk_K_r14_reg[6]/NET0131 ,
		_w35735_
	);
	LUT4 #(
		.INIT('hc963)
	) name29909 (
		decrypt_pad,
		\u2_R14_reg[9]/NET0131 ,
		\u2_uk_K_r14_reg[12]/NET0131 ,
		\u2_uk_K_r14_reg[19]/NET0131 ,
		_w35736_
	);
	LUT4 #(
		.INIT('hc963)
	) name29910 (
		decrypt_pad,
		\u2_R14_reg[4]/NET0131 ,
		\u2_uk_K_r14_reg[20]/NET0131 ,
		\u2_uk_K_r14_reg[27]/NET0131 ,
		_w35737_
	);
	LUT4 #(
		.INIT('hc963)
	) name29911 (
		decrypt_pad,
		\u2_R14_reg[6]/NET0131 ,
		\u2_uk_K_r14_reg[47]/NET0131 ,
		\u2_uk_K_r14_reg[54]/NET0131 ,
		_w35738_
	);
	LUT4 #(
		.INIT('hfb73)
	) name29912 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35739_
	);
	LUT2 #(
		.INIT('h4)
	) name29913 (
		_w35736_,
		_w35735_,
		_w35740_
	);
	LUT3 #(
		.INIT('had)
	) name29914 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35741_
	);
	LUT3 #(
		.INIT('h10)
	) name29915 (
		_w35737_,
		_w35735_,
		_w35738_,
		_w35742_
	);
	LUT4 #(
		.INIT('h0100)
	) name29916 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35743_
	);
	LUT4 #(
		.INIT('h00d8)
	) name29917 (
		_w35734_,
		_w35741_,
		_w35739_,
		_w35743_,
		_w35744_
	);
	LUT4 #(
		.INIT('h1005)
	) name29918 (
		_w35737_,
		_w35734_,
		_w35735_,
		_w35738_,
		_w35745_
	);
	LUT2 #(
		.INIT('h1)
	) name29919 (
		_w35735_,
		_w35738_,
		_w35746_
	);
	LUT4 #(
		.INIT('h8088)
	) name29920 (
		_w35736_,
		_w35737_,
		_w35734_,
		_w35735_,
		_w35747_
	);
	LUT4 #(
		.INIT('h4000)
	) name29921 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35748_
	);
	LUT4 #(
		.INIT('hbffa)
	) name29922 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35749_
	);
	LUT4 #(
		.INIT('h0b00)
	) name29923 (
		_w35746_,
		_w35747_,
		_w35745_,
		_w35749_,
		_w35750_
	);
	LUT4 #(
		.INIT('h0200)
	) name29924 (
		_w35736_,
		_w35737_,
		_w35734_,
		_w35735_,
		_w35751_
	);
	LUT4 #(
		.INIT('h0010)
	) name29925 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35752_
	);
	LUT4 #(
		.INIT('h77ef)
	) name29926 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35753_
	);
	LUT3 #(
		.INIT('h31)
	) name29927 (
		_w35734_,
		_w35751_,
		_w35753_,
		_w35754_
	);
	LUT4 #(
		.INIT('hd800)
	) name29928 (
		_w35733_,
		_w35744_,
		_w35750_,
		_w35754_,
		_w35755_
	);
	LUT2 #(
		.INIT('h9)
	) name29929 (
		\u2_L14_reg[18]/P0001 ,
		_w35755_,
		_w35756_
	);
	LUT4 #(
		.INIT('hc963)
	) name29930 (
		decrypt_pad,
		\u2_R14_reg[16]/NET0131 ,
		\u2_uk_K_r14_reg[33]/NET0131 ,
		\u2_uk_K_r14_reg[40]/NET0131 ,
		_w35757_
	);
	LUT4 #(
		.INIT('hc963)
	) name29931 (
		decrypt_pad,
		\u2_R14_reg[15]/NET0131 ,
		\u2_uk_K_r14_reg[25]/NET0131 ,
		\u2_uk_K_r14_reg[32]/NET0131 ,
		_w35758_
	);
	LUT4 #(
		.INIT('hc963)
	) name29932 (
		decrypt_pad,
		\u2_R14_reg[14]/NET0131 ,
		\u2_uk_K_r14_reg[17]/NET0131 ,
		\u2_uk_K_r14_reg[24]/NET0131 ,
		_w35759_
	);
	LUT4 #(
		.INIT('hc963)
	) name29933 (
		decrypt_pad,
		\u2_R14_reg[13]/NET0131 ,
		\u2_uk_K_r14_reg[48]/NET0131 ,
		\u2_uk_K_r14_reg[55]/NET0131 ,
		_w35760_
	);
	LUT4 #(
		.INIT('hc693)
	) name29934 (
		decrypt_pad,
		\u2_R14_reg[12]/NET0131 ,
		\u2_uk_K_r14_reg[4]/NET0131 ,
		\u2_uk_K_r14_reg[54]/NET0131 ,
		_w35761_
	);
	LUT4 #(
		.INIT('hc963)
	) name29935 (
		decrypt_pad,
		\u2_R14_reg[17]/NET0131 ,
		\u2_uk_K_r14_reg[13]/NET0131 ,
		\u2_uk_K_r14_reg[20]/NET0131 ,
		_w35762_
	);
	LUT2 #(
		.INIT('h4)
	) name29936 (
		_w35761_,
		_w35762_,
		_w35763_
	);
	LUT4 #(
		.INIT('h0400)
	) name29937 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35764_
	);
	LUT4 #(
		.INIT('hfb4f)
	) name29938 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35765_
	);
	LUT4 #(
		.INIT('h7dff)
	) name29939 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35766_
	);
	LUT2 #(
		.INIT('h2)
	) name29940 (
		_w35760_,
		_w35761_,
		_w35767_
	);
	LUT3 #(
		.INIT('h10)
	) name29941 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35768_
	);
	LUT4 #(
		.INIT('h1000)
	) name29942 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35769_
	);
	LUT4 #(
		.INIT('heff3)
	) name29943 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35770_
	);
	LUT4 #(
		.INIT('hc480)
	) name29944 (
		_w35758_,
		_w35766_,
		_w35770_,
		_w35765_,
		_w35771_
	);
	LUT2 #(
		.INIT('h2)
	) name29945 (
		_w35757_,
		_w35771_,
		_w35772_
	);
	LUT3 #(
		.INIT('h10)
	) name29946 (
		_w35758_,
		_w35759_,
		_w35762_,
		_w35773_
	);
	LUT4 #(
		.INIT('hc6c5)
	) name29947 (
		_w35758_,
		_w35759_,
		_w35760_,
		_w35762_,
		_w35774_
	);
	LUT2 #(
		.INIT('h2)
	) name29948 (
		_w35761_,
		_w35774_,
		_w35775_
	);
	LUT4 #(
		.INIT('h0008)
	) name29949 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35776_
	);
	LUT2 #(
		.INIT('h8)
	) name29950 (
		_w35758_,
		_w35759_,
		_w35777_
	);
	LUT3 #(
		.INIT('h01)
	) name29951 (
		_w35760_,
		_w35761_,
		_w35762_,
		_w35778_
	);
	LUT4 #(
		.INIT('hf5fc)
	) name29952 (
		_w35758_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35779_
	);
	LUT3 #(
		.INIT('h32)
	) name29953 (
		_w35777_,
		_w35776_,
		_w35779_,
		_w35780_
	);
	LUT3 #(
		.INIT('h45)
	) name29954 (
		_w35757_,
		_w35775_,
		_w35780_,
		_w35781_
	);
	LUT4 #(
		.INIT('h0001)
	) name29955 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35782_
	);
	LUT4 #(
		.INIT('h7dfe)
	) name29956 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35783_
	);
	LUT2 #(
		.INIT('h1)
	) name29957 (
		_w35758_,
		_w35783_,
		_w35784_
	);
	LUT3 #(
		.INIT('h80)
	) name29958 (
		_w35758_,
		_w35759_,
		_w35760_,
		_w35785_
	);
	LUT4 #(
		.INIT('h0080)
	) name29959 (
		_w35758_,
		_w35759_,
		_w35760_,
		_w35761_,
		_w35786_
	);
	LUT4 #(
		.INIT('h0080)
	) name29960 (
		_w35758_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35787_
	);
	LUT3 #(
		.INIT('h23)
	) name29961 (
		_w35759_,
		_w35786_,
		_w35787_,
		_w35788_
	);
	LUT2 #(
		.INIT('h4)
	) name29962 (
		_w35784_,
		_w35788_,
		_w35789_
	);
	LUT4 #(
		.INIT('h5655)
	) name29963 (
		\u2_L14_reg[10]/P0001 ,
		_w35772_,
		_w35781_,
		_w35789_,
		_w35790_
	);
	LUT4 #(
		.INIT('h2000)
	) name29964 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35791_
	);
	LUT4 #(
		.INIT('h0002)
	) name29965 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35792_
	);
	LUT3 #(
		.INIT('h01)
	) name29966 (
		_w35734_,
		_w35792_,
		_w35791_,
		_w35793_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name29967 (
		_w35737_,
		_w35734_,
		_w35735_,
		_w35738_,
		_w35794_
	);
	LUT2 #(
		.INIT('h4)
	) name29968 (
		_w35743_,
		_w35794_,
		_w35795_
	);
	LUT2 #(
		.INIT('h1)
	) name29969 (
		_w35793_,
		_w35795_,
		_w35796_
	);
	LUT4 #(
		.INIT('h39fd)
	) name29970 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35797_
	);
	LUT2 #(
		.INIT('h1)
	) name29971 (
		_w35734_,
		_w35797_,
		_w35798_
	);
	LUT2 #(
		.INIT('h8)
	) name29972 (
		_w35737_,
		_w35734_,
		_w35799_
	);
	LUT3 #(
		.INIT('h20)
	) name29973 (
		_w35736_,
		_w35735_,
		_w35738_,
		_w35800_
	);
	LUT3 #(
		.INIT('h15)
	) name29974 (
		_w35733_,
		_w35799_,
		_w35800_,
		_w35801_
	);
	LUT4 #(
		.INIT('h0052)
	) name29975 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35802_
	);
	LUT4 #(
		.INIT('h0002)
	) name29976 (
		_w35736_,
		_w35734_,
		_w35735_,
		_w35738_,
		_w35803_
	);
	LUT3 #(
		.INIT('h01)
	) name29977 (
		_w35791_,
		_w35802_,
		_w35803_,
		_w35804_
	);
	LUT3 #(
		.INIT('h40)
	) name29978 (
		_w35798_,
		_w35801_,
		_w35804_,
		_w35805_
	);
	LUT2 #(
		.INIT('h1)
	) name29979 (
		_w35734_,
		_w35735_,
		_w35806_
	);
	LUT4 #(
		.INIT('h0001)
	) name29980 (
		_w35736_,
		_w35737_,
		_w35734_,
		_w35735_,
		_w35807_
	);
	LUT4 #(
		.INIT('h80c0)
	) name29981 (
		_w35737_,
		_w35734_,
		_w35735_,
		_w35738_,
		_w35808_
	);
	LUT3 #(
		.INIT('h02)
	) name29982 (
		_w35733_,
		_w35808_,
		_w35807_,
		_w35809_
	);
	LUT2 #(
		.INIT('h9)
	) name29983 (
		_w35736_,
		_w35737_,
		_w35810_
	);
	LUT4 #(
		.INIT('h1300)
	) name29984 (
		_w35737_,
		_w35734_,
		_w35735_,
		_w35738_,
		_w35811_
	);
	LUT4 #(
		.INIT('hff7b)
	) name29985 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35812_
	);
	LUT3 #(
		.INIT('h70)
	) name29986 (
		_w35810_,
		_w35811_,
		_w35812_,
		_w35813_
	);
	LUT2 #(
		.INIT('h8)
	) name29987 (
		_w35809_,
		_w35813_,
		_w35814_
	);
	LUT4 #(
		.INIT('h6665)
	) name29988 (
		\u2_L14_reg[2]/P0001 ,
		_w35796_,
		_w35805_,
		_w35814_,
		_w35815_
	);
	LUT4 #(
		.INIT('hc963)
	) name29989 (
		decrypt_pad,
		\u2_R14_reg[32]/NET0131 ,
		\u2_uk_K_r14_reg[0]/NET0131 ,
		\u2_uk_K_r14_reg[7]/NET0131 ,
		_w35816_
	);
	LUT4 #(
		.INIT('hc693)
	) name29990 (
		decrypt_pad,
		\u2_R14_reg[31]/P0001 ,
		\u2_uk_K_r14_reg[1]/NET0131 ,
		\u2_uk_K_r14_reg[49]/P0001 ,
		_w35817_
	);
	LUT4 #(
		.INIT('hc693)
	) name29991 (
		decrypt_pad,
		\u2_R14_reg[28]/NET0131 ,
		\u2_uk_K_r14_reg[16]/NET0131 ,
		\u2_uk_K_r14_reg[9]/NET0131 ,
		_w35818_
	);
	LUT4 #(
		.INIT('hc963)
	) name29992 (
		decrypt_pad,
		\u2_R14_reg[30]/NET0131 ,
		\u2_uk_K_r14_reg[37]/NET0131 ,
		\u2_uk_K_r14_reg[44]/NET0131 ,
		_w35819_
	);
	LUT4 #(
		.INIT('hc963)
	) name29993 (
		decrypt_pad,
		\u2_R14_reg[29]/NET0131 ,
		\u2_uk_K_r14_reg[36]/NET0131 ,
		\u2_uk_K_r14_reg[43]/NET0131 ,
		_w35820_
	);
	LUT4 #(
		.INIT('hc963)
	) name29994 (
		decrypt_pad,
		\u2_R14_reg[1]/NET0131 ,
		\u2_uk_K_r14_reg[21]/NET0131 ,
		\u2_uk_K_r14_reg[28]/NET0131 ,
		_w35821_
	);
	LUT2 #(
		.INIT('h4)
	) name29995 (
		_w35821_,
		_w35820_,
		_w35822_
	);
	LUT4 #(
		.INIT('haf5c)
	) name29996 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w35823_
	);
	LUT2 #(
		.INIT('h1)
	) name29997 (
		_w35817_,
		_w35823_,
		_w35824_
	);
	LUT4 #(
		.INIT('hf010)
	) name29998 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w35825_
	);
	LUT2 #(
		.INIT('h4)
	) name29999 (
		_w35821_,
		_w35818_,
		_w35826_
	);
	LUT3 #(
		.INIT('hb0)
	) name30000 (
		_w35821_,
		_w35818_,
		_w35817_,
		_w35827_
	);
	LUT4 #(
		.INIT('h0400)
	) name30001 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w35828_
	);
	LUT4 #(
		.INIT('h0080)
	) name30002 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w35829_
	);
	LUT4 #(
		.INIT('hf97d)
	) name30003 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w35830_
	);
	LUT3 #(
		.INIT('h70)
	) name30004 (
		_w35825_,
		_w35827_,
		_w35830_,
		_w35831_
	);
	LUT3 #(
		.INIT('h8a)
	) name30005 (
		_w35816_,
		_w35824_,
		_w35831_,
		_w35832_
	);
	LUT4 #(
		.INIT('hef00)
	) name30006 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35817_,
		_w35833_
	);
	LUT4 #(
		.INIT('h7535)
	) name30007 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w35834_
	);
	LUT2 #(
		.INIT('h8)
	) name30008 (
		_w35833_,
		_w35834_,
		_w35835_
	);
	LUT4 #(
		.INIT('h0008)
	) name30009 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w35836_
	);
	LUT4 #(
		.INIT('h0004)
	) name30010 (
		_w35821_,
		_w35820_,
		_w35818_,
		_w35817_,
		_w35837_
	);
	LUT4 #(
		.INIT('h0080)
	) name30011 (
		_w35821_,
		_w35819_,
		_w35818_,
		_w35817_,
		_w35838_
	);
	LUT3 #(
		.INIT('h01)
	) name30012 (
		_w35836_,
		_w35837_,
		_w35838_,
		_w35839_
	);
	LUT3 #(
		.INIT('h45)
	) name30013 (
		_w35816_,
		_w35835_,
		_w35839_,
		_w35840_
	);
	LUT4 #(
		.INIT('hfdbf)
	) name30014 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w35841_
	);
	LUT2 #(
		.INIT('h1)
	) name30015 (
		_w35817_,
		_w35841_,
		_w35842_
	);
	LUT4 #(
		.INIT('h0400)
	) name30016 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35817_,
		_w35843_
	);
	LUT3 #(
		.INIT('h04)
	) name30017 (
		_w35819_,
		_w35818_,
		_w35817_,
		_w35844_
	);
	LUT3 #(
		.INIT('h13)
	) name30018 (
		_w35822_,
		_w35843_,
		_w35844_,
		_w35845_
	);
	LUT2 #(
		.INIT('h4)
	) name30019 (
		_w35842_,
		_w35845_,
		_w35846_
	);
	LUT4 #(
		.INIT('h5655)
	) name30020 (
		\u2_L14_reg[27]/P0001 ,
		_w35840_,
		_w35832_,
		_w35846_,
		_w35847_
	);
	LUT4 #(
		.INIT('hc963)
	) name30021 (
		decrypt_pad,
		\u2_R14_reg[23]/P0001 ,
		\u2_uk_K_r14_reg[2]/NET0131 ,
		\u2_uk_K_r14_reg[9]/NET0131 ,
		_w35848_
	);
	LUT4 #(
		.INIT('hc693)
	) name30022 (
		decrypt_pad,
		\u2_R14_reg[20]/NET0131 ,
		\u2_uk_K_r14_reg[14]/NET0131 ,
		\u2_uk_K_r14_reg[7]/NET0131 ,
		_w35849_
	);
	LUT4 #(
		.INIT('hc963)
	) name30023 (
		decrypt_pad,
		\u2_R14_reg[22]/P0001 ,
		\u2_uk_K_r14_reg[44]/NET0131 ,
		\u2_uk_K_r14_reg[51]/NET0131 ,
		_w35850_
	);
	LUT4 #(
		.INIT('hc963)
	) name30024 (
		decrypt_pad,
		\u2_R14_reg[21]/NET0131 ,
		\u2_uk_K_r14_reg[22]/NET0131 ,
		\u2_uk_K_r14_reg[29]/NET0131 ,
		_w35851_
	);
	LUT3 #(
		.INIT('h40)
	) name30025 (
		_w35850_,
		_w35849_,
		_w35851_,
		_w35852_
	);
	LUT4 #(
		.INIT('hc963)
	) name30026 (
		decrypt_pad,
		\u2_R14_reg[25]/NET0131 ,
		\u2_uk_K_r14_reg[23]/NET0131 ,
		\u2_uk_K_r14_reg[30]/NET0131 ,
		_w35853_
	);
	LUT4 #(
		.INIT('haff3)
	) name30027 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w35854_
	);
	LUT2 #(
		.INIT('h2)
	) name30028 (
		_w35848_,
		_w35854_,
		_w35855_
	);
	LUT3 #(
		.INIT('h0b)
	) name30029 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35856_
	);
	LUT2 #(
		.INIT('h1)
	) name30030 (
		_w35848_,
		_w35851_,
		_w35857_
	);
	LUT4 #(
		.INIT('hc963)
	) name30031 (
		decrypt_pad,
		\u2_R14_reg[24]/NET0131 ,
		\u2_uk_K_r14_reg[28]/NET0131 ,
		\u2_uk_K_r14_reg[35]/P0001 ,
		_w35858_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name30032 (
		_w35858_,
		_w35850_,
		_w35853_,
		_w35851_,
		_w35859_
	);
	LUT3 #(
		.INIT('hb0)
	) name30033 (
		_w35856_,
		_w35857_,
		_w35859_,
		_w35860_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name30034 (
		_w35853_,
		_w35849_,
		_w35848_,
		_w35851_,
		_w35861_
	);
	LUT4 #(
		.INIT('h8000)
	) name30035 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w35862_
	);
	LUT4 #(
		.INIT('h0405)
	) name30036 (
		_w35858_,
		_w35852_,
		_w35862_,
		_w35861_,
		_w35863_
	);
	LUT3 #(
		.INIT('h0b)
	) name30037 (
		_w35855_,
		_w35860_,
		_w35863_,
		_w35864_
	);
	LUT2 #(
		.INIT('h4)
	) name30038 (
		_w35853_,
		_w35849_,
		_w35865_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name30039 (
		_w35853_,
		_w35849_,
		_w35848_,
		_w35851_,
		_w35866_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name30040 (
		_w35853_,
		_w35849_,
		_w35848_,
		_w35851_,
		_w35867_
	);
	LUT3 #(
		.INIT('h01)
	) name30041 (
		_w35850_,
		_w35867_,
		_w35866_,
		_w35868_
	);
	LUT3 #(
		.INIT('h01)
	) name30042 (
		_w35853_,
		_w35849_,
		_w35851_,
		_w35869_
	);
	LUT3 #(
		.INIT('hde)
	) name30043 (
		_w35853_,
		_w35849_,
		_w35851_,
		_w35870_
	);
	LUT2 #(
		.INIT('h1)
	) name30044 (
		_w35858_,
		_w35848_,
		_w35871_
	);
	LUT3 #(
		.INIT('h72)
	) name30045 (
		_w35858_,
		_w35850_,
		_w35848_,
		_w35872_
	);
	LUT2 #(
		.INIT('h1)
	) name30046 (
		_w35850_,
		_w35848_,
		_w35873_
	);
	LUT4 #(
		.INIT('h0040)
	) name30047 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35848_,
		_w35874_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name30048 (
		_w35851_,
		_w35870_,
		_w35872_,
		_w35874_,
		_w35875_
	);
	LUT2 #(
		.INIT('h4)
	) name30049 (
		_w35868_,
		_w35875_,
		_w35876_
	);
	LUT3 #(
		.INIT('h65)
	) name30050 (
		\u2_L14_reg[19]/P0001 ,
		_w35864_,
		_w35876_,
		_w35877_
	);
	LUT4 #(
		.INIT('h202a)
	) name30051 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w35878_
	);
	LUT4 #(
		.INIT('h0440)
	) name30052 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w35879_
	);
	LUT3 #(
		.INIT('h01)
	) name30053 (
		_w35848_,
		_w35879_,
		_w35878_,
		_w35880_
	);
	LUT4 #(
		.INIT('h70f0)
	) name30054 (
		_w35853_,
		_w35849_,
		_w35848_,
		_w35851_,
		_w35881_
	);
	LUT4 #(
		.INIT('h0010)
	) name30055 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w35882_
	);
	LUT4 #(
		.INIT('hf5ef)
	) name30056 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w35883_
	);
	LUT2 #(
		.INIT('h8)
	) name30057 (
		_w35881_,
		_w35883_,
		_w35884_
	);
	LUT3 #(
		.INIT('ha8)
	) name30058 (
		_w35858_,
		_w35880_,
		_w35884_,
		_w35885_
	);
	LUT3 #(
		.INIT('he6)
	) name30059 (
		_w35850_,
		_w35849_,
		_w35851_,
		_w35886_
	);
	LUT4 #(
		.INIT('h090f)
	) name30060 (
		_w35850_,
		_w35849_,
		_w35848_,
		_w35851_,
		_w35887_
	);
	LUT3 #(
		.INIT('h07)
	) name30061 (
		_w35867_,
		_w35886_,
		_w35887_,
		_w35888_
	);
	LUT3 #(
		.INIT('hae)
	) name30062 (
		_w35850_,
		_w35848_,
		_w35851_,
		_w35889_
	);
	LUT4 #(
		.INIT('h0080)
	) name30063 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w35890_
	);
	LUT4 #(
		.INIT('h0501)
	) name30064 (
		_w35858_,
		_w35865_,
		_w35890_,
		_w35889_,
		_w35891_
	);
	LUT2 #(
		.INIT('h4)
	) name30065 (
		_w35888_,
		_w35891_,
		_w35892_
	);
	LUT4 #(
		.INIT('h0100)
	) name30066 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w35893_
	);
	LUT4 #(
		.INIT('h7e7f)
	) name30067 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w35894_
	);
	LUT2 #(
		.INIT('h2)
	) name30068 (
		_w35848_,
		_w35894_,
		_w35895_
	);
	LUT2 #(
		.INIT('h8)
	) name30069 (
		_w35869_,
		_w35873_,
		_w35896_
	);
	LUT3 #(
		.INIT('h01)
	) name30070 (
		_w35868_,
		_w35895_,
		_w35896_,
		_w35897_
	);
	LUT4 #(
		.INIT('h56aa)
	) name30071 (
		\u2_L14_reg[11]/P0001 ,
		_w35885_,
		_w35892_,
		_w35897_,
		_w35898_
	);
	LUT3 #(
		.INIT('h20)
	) name30072 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35899_
	);
	LUT4 #(
		.INIT('h0009)
	) name30073 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35900_
	);
	LUT4 #(
		.INIT('h4000)
	) name30074 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35901_
	);
	LUT4 #(
		.INIT('h0001)
	) name30075 (
		_w35708_,
		_w35899_,
		_w35900_,
		_w35901_,
		_w35902_
	);
	LUT4 #(
		.INIT('h0004)
	) name30076 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35903_
	);
	LUT4 #(
		.INIT('heffb)
	) name30077 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35904_
	);
	LUT3 #(
		.INIT('h02)
	) name30078 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35905_
	);
	LUT4 #(
		.INIT('hf700)
	) name30079 (
		_w35710_,
		_w35711_,
		_w35713_,
		_w35708_,
		_w35906_
	);
	LUT3 #(
		.INIT('h20)
	) name30080 (
		_w35904_,
		_w35905_,
		_w35906_,
		_w35907_
	);
	LUT4 #(
		.INIT('h0080)
	) name30081 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35908_
	);
	LUT4 #(
		.INIT('h0400)
	) name30082 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35909_
	);
	LUT4 #(
		.INIT('hfb7f)
	) name30083 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35910_
	);
	LUT4 #(
		.INIT('h02aa)
	) name30084 (
		_w35707_,
		_w35902_,
		_w35907_,
		_w35910_,
		_w35911_
	);
	LUT4 #(
		.INIT('h5100)
	) name30085 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35912_
	);
	LUT4 #(
		.INIT('h0cbc)
	) name30086 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w35913_
	);
	LUT4 #(
		.INIT('h0100)
	) name30087 (
		_w35708_,
		_w35900_,
		_w35901_,
		_w35913_,
		_w35914_
	);
	LUT3 #(
		.INIT('h40)
	) name30088 (
		_w35724_,
		_w35729_,
		_w35904_,
		_w35915_
	);
	LUT4 #(
		.INIT('h4445)
	) name30089 (
		_w35707_,
		_w35912_,
		_w35914_,
		_w35915_,
		_w35916_
	);
	LUT3 #(
		.INIT('h56)
	) name30090 (
		\u2_L14_reg[3]/P0001 ,
		_w35911_,
		_w35916_,
		_w35917_
	);
	LUT4 #(
		.INIT('h9080)
	) name30091 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35918_
	);
	LUT4 #(
		.INIT('hf0b0)
	) name30092 (
		_w35736_,
		_w35737_,
		_w35734_,
		_w35735_,
		_w35919_
	);
	LUT2 #(
		.INIT('h4)
	) name30093 (
		_w35918_,
		_w35919_,
		_w35920_
	);
	LUT4 #(
		.INIT('h2031)
	) name30094 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35921_
	);
	LUT4 #(
		.INIT('h3233)
	) name30095 (
		_w35737_,
		_w35734_,
		_w35735_,
		_w35738_,
		_w35922_
	);
	LUT3 #(
		.INIT('h04)
	) name30096 (
		_w35748_,
		_w35922_,
		_w35921_,
		_w35923_
	);
	LUT4 #(
		.INIT('h0008)
	) name30097 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35924_
	);
	LUT3 #(
		.INIT('h08)
	) name30098 (
		_w35737_,
		_w35734_,
		_w35738_,
		_w35925_
	);
	LUT4 #(
		.INIT('h0200)
	) name30099 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35926_
	);
	LUT4 #(
		.INIT('h0002)
	) name30100 (
		_w35733_,
		_w35924_,
		_w35925_,
		_w35926_,
		_w35927_
	);
	LUT3 #(
		.INIT('he0)
	) name30101 (
		_w35920_,
		_w35923_,
		_w35927_,
		_w35928_
	);
	LUT4 #(
		.INIT('h3d39)
	) name30102 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35929_
	);
	LUT4 #(
		.INIT('he4f5)
	) name30103 (
		_w35734_,
		_w35742_,
		_w35921_,
		_w35929_,
		_w35930_
	);
	LUT4 #(
		.INIT('h0900)
	) name30104 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w35931_
	);
	LUT3 #(
		.INIT('h01)
	) name30105 (
		_w35733_,
		_w35748_,
		_w35931_,
		_w35932_
	);
	LUT2 #(
		.INIT('h4)
	) name30106 (
		_w35930_,
		_w35932_,
		_w35933_
	);
	LUT3 #(
		.INIT('ha9)
	) name30107 (
		\u2_L14_reg[28]/P0001 ,
		_w35928_,
		_w35933_,
		_w35934_
	);
	LUT4 #(
		.INIT('h7bff)
	) name30108 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35935_
	);
	LUT4 #(
		.INIT('h0110)
	) name30109 (
		_w35758_,
		_w35759_,
		_w35760_,
		_w35761_,
		_w35936_
	);
	LUT3 #(
		.INIT('h02)
	) name30110 (
		_w35757_,
		_w35787_,
		_w35936_,
		_w35937_
	);
	LUT4 #(
		.INIT('h0200)
	) name30111 (
		_w35758_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35938_
	);
	LUT2 #(
		.INIT('h4)
	) name30112 (
		_w35758_,
		_w35759_,
		_w35939_
	);
	LUT3 #(
		.INIT('h13)
	) name30113 (
		_w35778_,
		_w35938_,
		_w35939_,
		_w35940_
	);
	LUT3 #(
		.INIT('h80)
	) name30114 (
		_w35935_,
		_w35937_,
		_w35940_,
		_w35941_
	);
	LUT4 #(
		.INIT('heff7)
	) name30115 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35942_
	);
	LUT3 #(
		.INIT('h8a)
	) name30116 (
		_w35758_,
		_w35760_,
		_w35762_,
		_w35943_
	);
	LUT4 #(
		.INIT('h8002)
	) name30117 (
		_w35758_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35944_
	);
	LUT3 #(
		.INIT('h10)
	) name30118 (
		_w35782_,
		_w35944_,
		_w35942_,
		_w35945_
	);
	LUT4 #(
		.INIT('hcc5f)
	) name30119 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35946_
	);
	LUT4 #(
		.INIT('h0302)
	) name30120 (
		_w35758_,
		_w35786_,
		_w35757_,
		_w35946_,
		_w35947_
	);
	LUT2 #(
		.INIT('h8)
	) name30121 (
		_w35945_,
		_w35947_,
		_w35948_
	);
	LUT4 #(
		.INIT('h0040)
	) name30122 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35949_
	);
	LUT4 #(
		.INIT('h0020)
	) name30123 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35950_
	);
	LUT4 #(
		.INIT('hff9e)
	) name30124 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w35951_
	);
	LUT4 #(
		.INIT('h3f15)
	) name30125 (
		_w35758_,
		_w35767_,
		_w35773_,
		_w35951_,
		_w35952_
	);
	LUT4 #(
		.INIT('ha955)
	) name30126 (
		\u2_L14_reg[20]/P0001 ,
		_w35941_,
		_w35948_,
		_w35952_,
		_w35953_
	);
	LUT4 #(
		.INIT('hc693)
	) name30127 (
		decrypt_pad,
		\u2_R14_reg[24]/NET0131 ,
		\u2_uk_K_r14_reg[2]/NET0131 ,
		\u2_uk_K_r14_reg[50]/NET0131 ,
		_w35954_
	);
	LUT4 #(
		.INIT('hc963)
	) name30128 (
		decrypt_pad,
		\u2_R14_reg[25]/NET0131 ,
		\u2_uk_K_r14_reg[30]/NET0131 ,
		\u2_uk_K_r14_reg[37]/NET0131 ,
		_w35955_
	);
	LUT4 #(
		.INIT('hc963)
	) name30129 (
		decrypt_pad,
		\u2_R14_reg[26]/P0001 ,
		\u2_uk_K_r14_reg[15]/NET0131 ,
		\u2_uk_K_r14_reg[22]/NET0131 ,
		_w35956_
	);
	LUT4 #(
		.INIT('hc963)
	) name30130 (
		decrypt_pad,
		\u2_R14_reg[29]/NET0131 ,
		\u2_uk_K_r14_reg[31]/NET0131 ,
		\u2_uk_K_r14_reg[38]/NET0131 ,
		_w35957_
	);
	LUT4 #(
		.INIT('h7776)
	) name30131 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w35958_
	);
	LUT4 #(
		.INIT('hc693)
	) name30132 (
		decrypt_pad,
		\u2_R14_reg[27]/P0001 ,
		\u2_uk_K_r14_reg[0]/NET0131 ,
		\u2_uk_K_r14_reg[52]/NET0131 ,
		_w35959_
	);
	LUT2 #(
		.INIT('h4)
	) name30133 (
		_w35958_,
		_w35959_,
		_w35960_
	);
	LUT4 #(
		.INIT('h0060)
	) name30134 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w35961_
	);
	LUT4 #(
		.INIT('hc963)
	) name30135 (
		decrypt_pad,
		\u2_R14_reg[28]/NET0131 ,
		\u2_uk_K_r14_reg[35]/P0001 ,
		\u2_uk_K_r14_reg[42]/P0001 ,
		_w35962_
	);
	LUT4 #(
		.INIT('h0200)
	) name30136 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w35963_
	);
	LUT3 #(
		.INIT('h04)
	) name30137 (
		_w35961_,
		_w35962_,
		_w35963_,
		_w35964_
	);
	LUT4 #(
		.INIT('h0400)
	) name30138 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w35965_
	);
	LUT4 #(
		.INIT('h1000)
	) name30139 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w35966_
	);
	LUT3 #(
		.INIT('h45)
	) name30140 (
		_w35965_,
		_w35959_,
		_w35966_,
		_w35967_
	);
	LUT3 #(
		.INIT('h40)
	) name30141 (
		_w35960_,
		_w35964_,
		_w35967_,
		_w35968_
	);
	LUT4 #(
		.INIT('h6000)
	) name30142 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w35969_
	);
	LUT4 #(
		.INIT('h0014)
	) name30143 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w35970_
	);
	LUT3 #(
		.INIT('h01)
	) name30144 (
		_w35962_,
		_w35970_,
		_w35969_,
		_w35971_
	);
	LUT2 #(
		.INIT('h6)
	) name30145 (
		_w35955_,
		_w35957_,
		_w35972_
	);
	LUT4 #(
		.INIT('h134c)
	) name30146 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w35973_
	);
	LUT3 #(
		.INIT('h02)
	) name30147 (
		_w35954_,
		_w35956_,
		_w35957_,
		_w35974_
	);
	LUT4 #(
		.INIT('h1102)
	) name30148 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w35975_
	);
	LUT4 #(
		.INIT('h04ee)
	) name30149 (
		_w35959_,
		_w35973_,
		_w35974_,
		_w35975_,
		_w35976_
	);
	LUT2 #(
		.INIT('h8)
	) name30150 (
		_w35971_,
		_w35976_,
		_w35977_
	);
	LUT3 #(
		.INIT('ha9)
	) name30151 (
		\u2_L14_reg[12]/P0001 ,
		_w35968_,
		_w35977_,
		_w35978_
	);
	LUT4 #(
		.INIT('hc693)
	) name30152 (
		decrypt_pad,
		\u2_R14_reg[1]/NET0131 ,
		\u2_uk_K_r14_reg[11]/NET0131 ,
		\u2_uk_K_r14_reg[4]/NET0131 ,
		_w35979_
	);
	LUT4 #(
		.INIT('hc963)
	) name30153 (
		decrypt_pad,
		\u2_R14_reg[5]/NET0131 ,
		\u2_uk_K_r14_reg[34]/NET0131 ,
		\u2_uk_K_r14_reg[41]/NET0131 ,
		_w35980_
	);
	LUT4 #(
		.INIT('hc963)
	) name30154 (
		decrypt_pad,
		\u2_R14_reg[32]/NET0131 ,
		\u2_uk_K_r14_reg[40]/NET0131 ,
		\u2_uk_K_r14_reg[47]/NET0131 ,
		_w35981_
	);
	LUT4 #(
		.INIT('hc963)
	) name30155 (
		decrypt_pad,
		\u2_R14_reg[2]/NET0131 ,
		\u2_uk_K_r14_reg[19]/NET0131 ,
		\u2_uk_K_r14_reg[26]/NET0131 ,
		_w35982_
	);
	LUT4 #(
		.INIT('h1020)
	) name30156 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w35983_
	);
	LUT4 #(
		.INIT('hc693)
	) name30157 (
		decrypt_pad,
		\u2_R14_reg[3]/NET0131 ,
		\u2_uk_K_r14_reg[3]/NET0131 ,
		\u2_uk_K_r14_reg[53]/NET0131 ,
		_w35984_
	);
	LUT4 #(
		.INIT('h7b00)
	) name30158 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35984_,
		_w35985_
	);
	LUT2 #(
		.INIT('h8)
	) name30159 (
		_w35980_,
		_w35981_,
		_w35986_
	);
	LUT3 #(
		.INIT('h09)
	) name30160 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35987_
	);
	LUT4 #(
		.INIT('h00fe)
	) name30161 (
		_w35980_,
		_w35981_,
		_w35982_,
		_w35984_,
		_w35988_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name30162 (
		_w35983_,
		_w35985_,
		_w35987_,
		_w35988_,
		_w35989_
	);
	LUT4 #(
		.INIT('hc693)
	) name30163 (
		decrypt_pad,
		\u2_R14_reg[4]/NET0131 ,
		\u2_uk_K_r14_reg[13]/NET0131 ,
		\u2_uk_K_r14_reg[6]/NET0131 ,
		_w35990_
	);
	LUT4 #(
		.INIT('h4200)
	) name30164 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w35991_
	);
	LUT2 #(
		.INIT('h1)
	) name30165 (
		_w35990_,
		_w35991_,
		_w35992_
	);
	LUT4 #(
		.INIT('h005e)
	) name30166 (
		_w35981_,
		_w35979_,
		_w35982_,
		_w35984_,
		_w35993_
	);
	LUT3 #(
		.INIT('h02)
	) name30167 (
		_w35981_,
		_w35979_,
		_w35982_,
		_w35994_
	);
	LUT4 #(
		.INIT('h0008)
	) name30168 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w35995_
	);
	LUT4 #(
		.INIT('hab00)
	) name30169 (
		_w35981_,
		_w35979_,
		_w35982_,
		_w35984_,
		_w35996_
	);
	LUT3 #(
		.INIT('h45)
	) name30170 (
		_w35993_,
		_w35995_,
		_w35996_,
		_w35997_
	);
	LUT3 #(
		.INIT('h40)
	) name30171 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35998_
	);
	LUT4 #(
		.INIT('h0040)
	) name30172 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w35999_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name30173 (
		_w35990_,
		_w35980_,
		_w35979_,
		_w35982_,
		_w36000_
	);
	LUT2 #(
		.INIT('h4)
	) name30174 (
		_w35999_,
		_w36000_,
		_w36001_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name30175 (
		_w35989_,
		_w35992_,
		_w35997_,
		_w36001_,
		_w36002_
	);
	LUT2 #(
		.INIT('h6)
	) name30176 (
		\u2_L14_reg[17]/P0001 ,
		_w36002_,
		_w36003_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name30177 (
		_w35853_,
		_w35849_,
		_w35848_,
		_w35851_,
		_w36004_
	);
	LUT4 #(
		.INIT('h0484)
	) name30178 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w36005_
	);
	LUT4 #(
		.INIT('h0008)
	) name30179 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w36006_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name30180 (
		_w35853_,
		_w35849_,
		_w35848_,
		_w35851_,
		_w36007_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name30181 (
		_w36004_,
		_w36005_,
		_w36006_,
		_w36007_,
		_w36008_
	);
	LUT2 #(
		.INIT('h1)
	) name30182 (
		_w35874_,
		_w35882_,
		_w36009_
	);
	LUT3 #(
		.INIT('h45)
	) name30183 (
		_w35858_,
		_w36008_,
		_w36009_,
		_w36010_
	);
	LUT4 #(
		.INIT('heafa)
	) name30184 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w36011_
	);
	LUT2 #(
		.INIT('h1)
	) name30185 (
		_w35848_,
		_w36011_,
		_w36012_
	);
	LUT3 #(
		.INIT('h80)
	) name30186 (
		_w35850_,
		_w35853_,
		_w35851_,
		_w36013_
	);
	LUT4 #(
		.INIT('h4000)
	) name30187 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35848_,
		_w36014_
	);
	LUT3 #(
		.INIT('h01)
	) name30188 (
		_w35893_,
		_w36013_,
		_w36014_,
		_w36015_
	);
	LUT4 #(
		.INIT('h90e0)
	) name30189 (
		_w35853_,
		_w35849_,
		_w35848_,
		_w35851_,
		_w36016_
	);
	LUT4 #(
		.INIT('h070b)
	) name30190 (
		_w35853_,
		_w35849_,
		_w35848_,
		_w35851_,
		_w36017_
	);
	LUT4 #(
		.INIT('h0001)
	) name30191 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35848_,
		_w36018_
	);
	LUT4 #(
		.INIT('h00fd)
	) name30192 (
		_w35850_,
		_w36017_,
		_w36016_,
		_w36018_,
		_w36019_
	);
	LUT4 #(
		.INIT('h7500)
	) name30193 (
		_w35858_,
		_w36012_,
		_w36015_,
		_w36019_,
		_w36020_
	);
	LUT3 #(
		.INIT('h65)
	) name30194 (
		\u2_L14_reg[4]/P0001 ,
		_w36010_,
		_w36020_,
		_w36021_
	);
	LUT4 #(
		.INIT('hf010)
	) name30195 (
		_w35850_,
		_w35853_,
		_w35848_,
		_w35851_,
		_w36022_
	);
	LUT4 #(
		.INIT('h9297)
	) name30196 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w36023_
	);
	LUT2 #(
		.INIT('h4)
	) name30197 (
		_w36022_,
		_w36023_,
		_w36024_
	);
	LUT4 #(
		.INIT('hd2ff)
	) name30198 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w36025_
	);
	LUT3 #(
		.INIT('ha2)
	) name30199 (
		_w35858_,
		_w35848_,
		_w36025_,
		_w36026_
	);
	LUT4 #(
		.INIT('h3dce)
	) name30200 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w36027_
	);
	LUT4 #(
		.INIT('h0501)
	) name30201 (
		_w35858_,
		_w35848_,
		_w36006_,
		_w36027_,
		_w36028_
	);
	LUT4 #(
		.INIT('h9abf)
	) name30202 (
		_w35850_,
		_w35853_,
		_w35849_,
		_w35851_,
		_w36029_
	);
	LUT4 #(
		.INIT('h4000)
	) name30203 (
		_w35850_,
		_w35853_,
		_w35848_,
		_w35851_,
		_w36030_
	);
	LUT4 #(
		.INIT('h0031)
	) name30204 (
		_w35871_,
		_w35882_,
		_w36029_,
		_w36030_,
		_w36031_
	);
	LUT4 #(
		.INIT('hf400)
	) name30205 (
		_w36024_,
		_w36026_,
		_w36028_,
		_w36031_,
		_w36032_
	);
	LUT2 #(
		.INIT('h6)
	) name30206 (
		\u2_L14_reg[29]/P0001 ,
		_w36032_,
		_w36033_
	);
	LUT4 #(
		.INIT('h0800)
	) name30207 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36034_
	);
	LUT4 #(
		.INIT('hff10)
	) name30208 (
		_w35821_,
		_w35819_,
		_w35818_,
		_w35817_,
		_w36035_
	);
	LUT4 #(
		.INIT('hf700)
	) name30209 (
		_w35821_,
		_w35820_,
		_w35818_,
		_w35817_,
		_w36036_
	);
	LUT3 #(
		.INIT('h80)
	) name30210 (
		_w35819_,
		_w35820_,
		_w35818_,
		_w36037_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name30211 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36038_
	);
	LUT4 #(
		.INIT('h0eee)
	) name30212 (
		_w36034_,
		_w36035_,
		_w36036_,
		_w36038_,
		_w36039_
	);
	LUT4 #(
		.INIT('h4004)
	) name30213 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36040_
	);
	LUT4 #(
		.INIT('h0002)
	) name30214 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36041_
	);
	LUT3 #(
		.INIT('h02)
	) name30215 (
		_w35816_,
		_w36041_,
		_w36040_,
		_w36042_
	);
	LUT2 #(
		.INIT('h4)
	) name30216 (
		_w36039_,
		_w36042_,
		_w36043_
	);
	LUT4 #(
		.INIT('h5515)
	) name30217 (
		_w35816_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36044_
	);
	LUT4 #(
		.INIT('h0020)
	) name30218 (
		_w35821_,
		_w35819_,
		_w35818_,
		_w35817_,
		_w36045_
	);
	LUT4 #(
		.INIT('h0001)
	) name30219 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36046_
	);
	LUT4 #(
		.INIT('h0100)
	) name30220 (
		_w35828_,
		_w36045_,
		_w36046_,
		_w36044_,
		_w36047_
	);
	LUT4 #(
		.INIT('ha3ff)
	) name30221 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36048_
	);
	LUT2 #(
		.INIT('h2)
	) name30222 (
		_w35817_,
		_w36048_,
		_w36049_
	);
	LUT4 #(
		.INIT('h2000)
	) name30223 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36050_
	);
	LUT4 #(
		.INIT('h0008)
	) name30224 (
		_w35821_,
		_w35819_,
		_w35818_,
		_w35817_,
		_w36051_
	);
	LUT3 #(
		.INIT('h01)
	) name30225 (
		_w35837_,
		_w36051_,
		_w36050_,
		_w36052_
	);
	LUT3 #(
		.INIT('h40)
	) name30226 (
		_w36049_,
		_w36052_,
		_w36047_,
		_w36053_
	);
	LUT4 #(
		.INIT('h0100)
	) name30227 (
		_w35819_,
		_w35820_,
		_w35818_,
		_w35817_,
		_w36054_
	);
	LUT3 #(
		.INIT('h07)
	) name30228 (
		_w35820_,
		_w36045_,
		_w36054_,
		_w36055_
	);
	LUT4 #(
		.INIT('ha955)
	) name30229 (
		\u2_L14_reg[21]/P0001 ,
		_w36043_,
		_w36053_,
		_w36055_,
		_w36056_
	);
	LUT4 #(
		.INIT('hbf7f)
	) name30230 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w36057_
	);
	LUT4 #(
		.INIT('hedeb)
	) name30231 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w36058_
	);
	LUT4 #(
		.INIT('h0515)
	) name30232 (
		_w35734_,
		_w35733_,
		_w36057_,
		_w36058_,
		_w36059_
	);
	LUT4 #(
		.INIT('h72f6)
	) name30233 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w36060_
	);
	LUT2 #(
		.INIT('h2)
	) name30234 (
		_w35734_,
		_w36060_,
		_w36061_
	);
	LUT3 #(
		.INIT('h02)
	) name30235 (
		_w35736_,
		_w35737_,
		_w35738_,
		_w36062_
	);
	LUT2 #(
		.INIT('h4)
	) name30236 (
		_w35806_,
		_w36062_,
		_w36063_
	);
	LUT3 #(
		.INIT('h15)
	) name30237 (
		_w35733_,
		_w35740_,
		_w35925_,
		_w36064_
	);
	LUT3 #(
		.INIT('h10)
	) name30238 (
		_w36061_,
		_w36063_,
		_w36064_,
		_w36065_
	);
	LUT3 #(
		.INIT('h27)
	) name30239 (
		_w35736_,
		_w35737_,
		_w35738_,
		_w36066_
	);
	LUT4 #(
		.INIT('h2202)
	) name30240 (
		_w35733_,
		_w35752_,
		_w35806_,
		_w36066_,
		_w36067_
	);
	LUT4 #(
		.INIT('hddfa)
	) name30241 (
		_w35736_,
		_w35737_,
		_w35735_,
		_w35738_,
		_w36068_
	);
	LUT2 #(
		.INIT('h2)
	) name30242 (
		_w35734_,
		_w36068_,
		_w36069_
	);
	LUT3 #(
		.INIT('h10)
	) name30243 (
		_w35791_,
		_w35803_,
		_w36057_,
		_w36070_
	);
	LUT3 #(
		.INIT('h40)
	) name30244 (
		_w36069_,
		_w36067_,
		_w36070_,
		_w36071_
	);
	LUT4 #(
		.INIT('h999a)
	) name30245 (
		\u2_L14_reg[13]/P0001 ,
		_w36059_,
		_w36065_,
		_w36071_,
		_w36072_
	);
	LUT4 #(
		.INIT('hfbf5)
	) name30246 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36073_
	);
	LUT2 #(
		.INIT('h2)
	) name30247 (
		_w35817_,
		_w36073_,
		_w36074_
	);
	LUT4 #(
		.INIT('h00e4)
	) name30248 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35817_,
		_w36075_
	);
	LUT3 #(
		.INIT('h54)
	) name30249 (
		_w35826_,
		_w36037_,
		_w36075_,
		_w36076_
	);
	LUT4 #(
		.INIT('h1000)
	) name30250 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36077_
	);
	LUT2 #(
		.INIT('h1)
	) name30251 (
		_w35844_,
		_w36077_,
		_w36078_
	);
	LUT4 #(
		.INIT('h5455)
	) name30252 (
		_w35816_,
		_w36076_,
		_w36074_,
		_w36078_,
		_w36079_
	);
	LUT4 #(
		.INIT('h6350)
	) name30253 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36080_
	);
	LUT4 #(
		.INIT('h00df)
	) name30254 (
		_w35819_,
		_w35820_,
		_w35818_,
		_w35817_,
		_w36081_
	);
	LUT4 #(
		.INIT('h00de)
	) name30255 (
		_w35819_,
		_w35820_,
		_w35818_,
		_w35817_,
		_w36082_
	);
	LUT4 #(
		.INIT('h3302)
	) name30256 (
		_w35817_,
		_w35829_,
		_w36080_,
		_w36082_,
		_w36083_
	);
	LUT4 #(
		.INIT('hffbe)
	) name30257 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36084_
	);
	LUT4 #(
		.INIT('hfdb6)
	) name30258 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36085_
	);
	LUT4 #(
		.INIT('h3f15)
	) name30259 (
		_w35817_,
		_w35822_,
		_w35844_,
		_w36085_,
		_w36086_
	);
	LUT3 #(
		.INIT('hd0)
	) name30260 (
		_w35816_,
		_w36083_,
		_w36086_,
		_w36087_
	);
	LUT3 #(
		.INIT('h9a)
	) name30261 (
		\u2_L14_reg[5]/P0001 ,
		_w36079_,
		_w36087_,
		_w36088_
	);
	LUT4 #(
		.INIT('hc963)
	) name30262 (
		decrypt_pad,
		\u2_R14_reg[12]/NET0131 ,
		\u2_uk_K_r14_reg[10]/P0001 ,
		\u2_uk_K_r14_reg[17]/NET0131 ,
		_w36089_
	);
	LUT4 #(
		.INIT('hc963)
	) name30263 (
		decrypt_pad,
		\u2_R14_reg[8]/NET0131 ,
		\u2_uk_K_r14_reg[46]/NET0131 ,
		\u2_uk_K_r14_reg[53]/NET0131 ,
		_w36090_
	);
	LUT4 #(
		.INIT('hc963)
	) name30264 (
		decrypt_pad,
		\u2_R14_reg[10]/P0001 ,
		\u2_uk_K_r14_reg[26]/NET0131 ,
		\u2_uk_K_r14_reg[33]/NET0131 ,
		_w36091_
	);
	LUT2 #(
		.INIT('h8)
	) name30265 (
		_w36090_,
		_w36091_,
		_w36092_
	);
	LUT4 #(
		.INIT('hc963)
	) name30266 (
		decrypt_pad,
		\u2_R14_reg[13]/NET0131 ,
		\u2_uk_K_r14_reg[55]/NET0131 ,
		\u2_uk_K_r14_reg[5]/NET0131 ,
		_w36093_
	);
	LUT4 #(
		.INIT('hc963)
	) name30267 (
		decrypt_pad,
		\u2_R14_reg[9]/NET0131 ,
		\u2_uk_K_r14_reg[18]/NET0131 ,
		\u2_uk_K_r14_reg[25]/NET0131 ,
		_w36094_
	);
	LUT3 #(
		.INIT('h08)
	) name30268 (
		_w36093_,
		_w36091_,
		_w36094_,
		_w36095_
	);
	LUT4 #(
		.INIT('hc963)
	) name30269 (
		decrypt_pad,
		\u2_R14_reg[11]/P0001 ,
		\u2_uk_K_r14_reg[27]/NET0131 ,
		\u2_uk_K_r14_reg[34]/NET0131 ,
		_w36096_
	);
	LUT3 #(
		.INIT('hca)
	) name30270 (
		_w36090_,
		_w36093_,
		_w36094_,
		_w36097_
	);
	LUT4 #(
		.INIT('h5044)
	) name30271 (
		_w36096_,
		_w36090_,
		_w36093_,
		_w36094_,
		_w36098_
	);
	LUT3 #(
		.INIT('h54)
	) name30272 (
		_w36092_,
		_w36095_,
		_w36098_,
		_w36099_
	);
	LUT4 #(
		.INIT('h000b)
	) name30273 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36100_
	);
	LUT4 #(
		.INIT('h0009)
	) name30274 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36101_
	);
	LUT4 #(
		.INIT('h7c5f)
	) name30275 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36102_
	);
	LUT3 #(
		.INIT('h31)
	) name30276 (
		_w36096_,
		_w36101_,
		_w36102_,
		_w36103_
	);
	LUT3 #(
		.INIT('h45)
	) name30277 (
		_w36089_,
		_w36099_,
		_w36103_,
		_w36104_
	);
	LUT2 #(
		.INIT('h8)
	) name30278 (
		_w36089_,
		_w36096_,
		_w36105_
	);
	LUT2 #(
		.INIT('h1)
	) name30279 (
		_w36090_,
		_w36093_,
		_w36106_
	);
	LUT4 #(
		.INIT('hebe9)
	) name30280 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36107_
	);
	LUT2 #(
		.INIT('h2)
	) name30281 (
		_w36105_,
		_w36107_,
		_w36108_
	);
	LUT4 #(
		.INIT('h4e5f)
	) name30282 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36109_
	);
	LUT2 #(
		.INIT('h2)
	) name30283 (
		_w36089_,
		_w36096_,
		_w36110_
	);
	LUT2 #(
		.INIT('h4)
	) name30284 (
		_w36109_,
		_w36110_,
		_w36111_
	);
	LUT2 #(
		.INIT('h8)
	) name30285 (
		_w36096_,
		_w36090_,
		_w36112_
	);
	LUT2 #(
		.INIT('h8)
	) name30286 (
		_w36095_,
		_w36112_,
		_w36113_
	);
	LUT2 #(
		.INIT('h8)
	) name30287 (
		_w36090_,
		_w36093_,
		_w36114_
	);
	LUT3 #(
		.INIT('h80)
	) name30288 (
		_w36089_,
		_w36091_,
		_w36094_,
		_w36115_
	);
	LUT2 #(
		.INIT('h4)
	) name30289 (
		_w36096_,
		_w36091_,
		_w36116_
	);
	LUT4 #(
		.INIT('h1000)
	) name30290 (
		_w36096_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36117_
	);
	LUT3 #(
		.INIT('h0b)
	) name30291 (
		_w36114_,
		_w36115_,
		_w36117_,
		_w36118_
	);
	LUT4 #(
		.INIT('h0100)
	) name30292 (
		_w36108_,
		_w36111_,
		_w36113_,
		_w36118_,
		_w36119_
	);
	LUT3 #(
		.INIT('h9a)
	) name30293 (
		\u2_L14_reg[30]/P0001 ,
		_w36104_,
		_w36119_,
		_w36120_
	);
	LUT4 #(
		.INIT('h0010)
	) name30294 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36121_
	);
	LUT4 #(
		.INIT('h5a65)
	) name30295 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36122_
	);
	LUT2 #(
		.INIT('h1)
	) name30296 (
		_w35959_,
		_w36122_,
		_w36123_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name30297 (
		_w35954_,
		_w35955_,
		_w35957_,
		_w35959_,
		_w36124_
	);
	LUT4 #(
		.INIT('h8000)
	) name30298 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36125_
	);
	LUT3 #(
		.INIT('h0e)
	) name30299 (
		_w35956_,
		_w36124_,
		_w36125_,
		_w36126_
	);
	LUT3 #(
		.INIT('h45)
	) name30300 (
		_w35962_,
		_w36123_,
		_w36126_,
		_w36127_
	);
	LUT4 #(
		.INIT('hd7df)
	) name30301 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36128_
	);
	LUT4 #(
		.INIT('hb9ff)
	) name30302 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36129_
	);
	LUT4 #(
		.INIT('heffe)
	) name30303 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36130_
	);
	LUT4 #(
		.INIT('he400)
	) name30304 (
		_w35959_,
		_w36129_,
		_w36128_,
		_w36130_,
		_w36131_
	);
	LUT4 #(
		.INIT('hef9d)
	) name30305 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36132_
	);
	LUT4 #(
		.INIT('h0100)
	) name30306 (
		_w35955_,
		_w35956_,
		_w35957_,
		_w35959_,
		_w36133_
	);
	LUT4 #(
		.INIT('h0084)
	) name30307 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35959_,
		_w36134_
	);
	LUT4 #(
		.INIT('h000d)
	) name30308 (
		_w35959_,
		_w36132_,
		_w36133_,
		_w36134_,
		_w36135_
	);
	LUT3 #(
		.INIT('hd0)
	) name30309 (
		_w35962_,
		_w36131_,
		_w36135_,
		_w36136_
	);
	LUT3 #(
		.INIT('h65)
	) name30310 (
		\u2_L14_reg[22]/P0001 ,
		_w36127_,
		_w36136_,
		_w36137_
	);
	LUT4 #(
		.INIT('hfe00)
	) name30311 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35708_,
		_w36138_
	);
	LUT4 #(
		.INIT('h3fdd)
	) name30312 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36139_
	);
	LUT2 #(
		.INIT('h8)
	) name30313 (
		_w36138_,
		_w36139_,
		_w36140_
	);
	LUT4 #(
		.INIT('he5ef)
	) name30314 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36141_
	);
	LUT4 #(
		.INIT('h0100)
	) name30315 (
		_w35708_,
		_w35908_,
		_w35903_,
		_w36141_,
		_w36142_
	);
	LUT4 #(
		.INIT('hbffd)
	) name30316 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36143_
	);
	LUT4 #(
		.INIT('h0155)
	) name30317 (
		_w35707_,
		_w36140_,
		_w36142_,
		_w36143_,
		_w36144_
	);
	LUT4 #(
		.INIT('h0021)
	) name30318 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35708_,
		_w36145_
	);
	LUT4 #(
		.INIT('h00b7)
	) name30319 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36146_
	);
	LUT4 #(
		.INIT('h0080)
	) name30320 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35708_,
		_w36147_
	);
	LUT4 #(
		.INIT('hfb00)
	) name30321 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36148_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name30322 (
		_w36145_,
		_w36146_,
		_w36147_,
		_w36148_,
		_w36149_
	);
	LUT4 #(
		.INIT('hc727)
	) name30323 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36150_
	);
	LUT2 #(
		.INIT('h2)
	) name30324 (
		_w35708_,
		_w36150_,
		_w36151_
	);
	LUT4 #(
		.INIT('h0108)
	) name30325 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36152_
	);
	LUT4 #(
		.INIT('h1200)
	) name30326 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36153_
	);
	LUT3 #(
		.INIT('hd8)
	) name30327 (
		_w35708_,
		_w36152_,
		_w36153_,
		_w36154_
	);
	LUT4 #(
		.INIT('h0057)
	) name30328 (
		_w35707_,
		_w36149_,
		_w36151_,
		_w36154_,
		_w36155_
	);
	LUT3 #(
		.INIT('h65)
	) name30329 (
		\u2_L14_reg[14]/P0001 ,
		_w36144_,
		_w36155_,
		_w36156_
	);
	LUT2 #(
		.INIT('h9)
	) name30330 (
		_w36090_,
		_w36093_,
		_w36157_
	);
	LUT4 #(
		.INIT('h9990)
	) name30331 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36158_
	);
	LUT4 #(
		.INIT('h0990)
	) name30332 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36159_
	);
	LUT4 #(
		.INIT('h4000)
	) name30333 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36160_
	);
	LUT2 #(
		.INIT('h4)
	) name30334 (
		_w36096_,
		_w36160_,
		_w36161_
	);
	LUT4 #(
		.INIT('h000d)
	) name30335 (
		_w36096_,
		_w36090_,
		_w36091_,
		_w36094_,
		_w36162_
	);
	LUT4 #(
		.INIT('h0200)
	) name30336 (
		_w36096_,
		_w36090_,
		_w36091_,
		_w36094_,
		_w36163_
	);
	LUT4 #(
		.INIT('h2000)
	) name30337 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36164_
	);
	LUT4 #(
		.INIT('h000b)
	) name30338 (
		_w36157_,
		_w36162_,
		_w36163_,
		_w36164_,
		_w36165_
	);
	LUT4 #(
		.INIT('h5455)
	) name30339 (
		_w36089_,
		_w36161_,
		_w36159_,
		_w36165_,
		_w36166_
	);
	LUT4 #(
		.INIT('h0001)
	) name30340 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36167_
	);
	LUT4 #(
		.INIT('hff3e)
	) name30341 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36168_
	);
	LUT2 #(
		.INIT('h2)
	) name30342 (
		_w36096_,
		_w36168_,
		_w36169_
	);
	LUT4 #(
		.INIT('h9d33)
	) name30343 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36170_
	);
	LUT2 #(
		.INIT('h2)
	) name30344 (
		_w36105_,
		_w36170_,
		_w36171_
	);
	LUT3 #(
		.INIT('h45)
	) name30345 (
		_w36090_,
		_w36091_,
		_w36094_,
		_w36172_
	);
	LUT4 #(
		.INIT('h2002)
	) name30346 (
		_w36089_,
		_w36096_,
		_w36093_,
		_w36094_,
		_w36173_
	);
	LUT4 #(
		.INIT('h7077)
	) name30347 (
		_w36106_,
		_w36115_,
		_w36172_,
		_w36173_,
		_w36174_
	);
	LUT3 #(
		.INIT('h10)
	) name30348 (
		_w36171_,
		_w36169_,
		_w36174_,
		_w36175_
	);
	LUT3 #(
		.INIT('h65)
	) name30349 (
		\u2_L14_reg[6]/P0001 ,
		_w36166_,
		_w36175_,
		_w36176_
	);
	LUT2 #(
		.INIT('h4)
	) name30350 (
		_w35982_,
		_w35984_,
		_w36177_
	);
	LUT4 #(
		.INIT('h2a22)
	) name30351 (
		_w35980_,
		_w35979_,
		_w35982_,
		_w35984_,
		_w36178_
	);
	LUT3 #(
		.INIT('h54)
	) name30352 (
		_w35986_,
		_w35994_,
		_w36178_,
		_w36179_
	);
	LUT4 #(
		.INIT('he4f5)
	) name30353 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36180_
	);
	LUT3 #(
		.INIT('h08)
	) name30354 (
		_w35981_,
		_w35979_,
		_w35984_,
		_w36181_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name30355 (
		_w35990_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36182_
	);
	LUT4 #(
		.INIT('h0d00)
	) name30356 (
		_w35984_,
		_w36180_,
		_w36181_,
		_w36182_,
		_w36183_
	);
	LUT2 #(
		.INIT('h4)
	) name30357 (
		_w36179_,
		_w36183_,
		_w36184_
	);
	LUT3 #(
		.INIT('hce)
	) name30358 (
		_w35979_,
		_w35982_,
		_w35984_,
		_w36185_
	);
	LUT2 #(
		.INIT('h2)
	) name30359 (
		_w35986_,
		_w36185_,
		_w36186_
	);
	LUT2 #(
		.INIT('h8)
	) name30360 (
		_w35982_,
		_w35984_,
		_w36187_
	);
	LUT3 #(
		.INIT('h15)
	) name30361 (
		_w35990_,
		_w35998_,
		_w36187_,
		_w36188_
	);
	LUT4 #(
		.INIT('hfbce)
	) name30362 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36189_
	);
	LUT4 #(
		.INIT('h2000)
	) name30363 (
		_w35980_,
		_w35981_,
		_w35982_,
		_w35984_,
		_w36190_
	);
	LUT4 #(
		.INIT('hdefe)
	) name30364 (
		_w35980_,
		_w35981_,
		_w35982_,
		_w35984_,
		_w36191_
	);
	LUT4 #(
		.INIT('hfc54)
	) name30365 (
		_w35979_,
		_w35984_,
		_w36189_,
		_w36191_,
		_w36192_
	);
	LUT3 #(
		.INIT('h40)
	) name30366 (
		_w36186_,
		_w36188_,
		_w36192_,
		_w36193_
	);
	LUT4 #(
		.INIT('hfd00)
	) name30367 (
		_w35981_,
		_w35979_,
		_w35982_,
		_w35984_,
		_w36194_
	);
	LUT4 #(
		.INIT('h0250)
	) name30368 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36195_
	);
	LUT4 #(
		.INIT('h8000)
	) name30369 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36196_
	);
	LUT4 #(
		.INIT('h3332)
	) name30370 (
		_w35984_,
		_w36194_,
		_w36195_,
		_w36196_,
		_w36197_
	);
	LUT3 #(
		.INIT('h01)
	) name30371 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w36198_
	);
	LUT2 #(
		.INIT('h8)
	) name30372 (
		_w36187_,
		_w36198_,
		_w36199_
	);
	LUT2 #(
		.INIT('h1)
	) name30373 (
		_w36197_,
		_w36199_,
		_w36200_
	);
	LUT4 #(
		.INIT('ha955)
	) name30374 (
		\u2_L14_reg[31]/P0001 ,
		_w36184_,
		_w36193_,
		_w36200_,
		_w36201_
	);
	LUT4 #(
		.INIT('h9600)
	) name30375 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36202_
	);
	LUT3 #(
		.INIT('hda)
	) name30376 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w36203_
	);
	LUT4 #(
		.INIT('h0051)
	) name30377 (
		_w35999_,
		_w36177_,
		_w36203_,
		_w36202_,
		_w36204_
	);
	LUT2 #(
		.INIT('h2)
	) name30378 (
		_w35990_,
		_w36204_,
		_w36205_
	);
	LUT4 #(
		.INIT('h0080)
	) name30379 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36206_
	);
	LUT4 #(
		.INIT('hdf7f)
	) name30380 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36207_
	);
	LUT2 #(
		.INIT('h1)
	) name30381 (
		_w35984_,
		_w36207_,
		_w36208_
	);
	LUT4 #(
		.INIT('ha5e5)
	) name30382 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36209_
	);
	LUT2 #(
		.INIT('h2)
	) name30383 (
		_w35984_,
		_w36209_,
		_w36210_
	);
	LUT4 #(
		.INIT('h0900)
	) name30384 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36211_
	);
	LUT4 #(
		.INIT('h0025)
	) name30385 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35984_,
		_w36212_
	);
	LUT3 #(
		.INIT('h01)
	) name30386 (
		_w36206_,
		_w36212_,
		_w36211_,
		_w36213_
	);
	LUT4 #(
		.INIT('h2322)
	) name30387 (
		_w35990_,
		_w36208_,
		_w36210_,
		_w36213_,
		_w36214_
	);
	LUT3 #(
		.INIT('h65)
	) name30388 (
		\u2_L14_reg[9]/P0001 ,
		_w36205_,
		_w36214_,
		_w36215_
	);
	LUT4 #(
		.INIT('h0010)
	) name30389 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36216_
	);
	LUT2 #(
		.INIT('h2)
	) name30390 (
		_w36194_,
		_w36216_,
		_w36217_
	);
	LUT4 #(
		.INIT('h0208)
	) name30391 (
		_w35990_,
		_w35980_,
		_w35981_,
		_w35979_,
		_w36218_
	);
	LUT4 #(
		.INIT('h1555)
	) name30392 (
		_w35990_,
		_w35980_,
		_w35981_,
		_w35979_,
		_w36219_
	);
	LUT4 #(
		.INIT('h8400)
	) name30393 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36220_
	);
	LUT2 #(
		.INIT('h4)
	) name30394 (
		_w36219_,
		_w36220_,
		_w36221_
	);
	LUT4 #(
		.INIT('h0002)
	) name30395 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35982_,
		_w36222_
	);
	LUT3 #(
		.INIT('h01)
	) name30396 (
		_w35984_,
		_w35999_,
		_w36222_,
		_w36223_
	);
	LUT4 #(
		.INIT('h5455)
	) name30397 (
		_w36217_,
		_w36221_,
		_w36218_,
		_w36223_,
		_w36224_
	);
	LUT4 #(
		.INIT('h3f1f)
	) name30398 (
		_w35981_,
		_w35979_,
		_w35982_,
		_w35984_,
		_w36225_
	);
	LUT2 #(
		.INIT('h2)
	) name30399 (
		_w35980_,
		_w36225_,
		_w36226_
	);
	LUT4 #(
		.INIT('h1000)
	) name30400 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35984_,
		_w36227_
	);
	LUT4 #(
		.INIT('h5515)
	) name30401 (
		_w35990_,
		_w35981_,
		_w35979_,
		_w35984_,
		_w36228_
	);
	LUT3 #(
		.INIT('h01)
	) name30402 (
		_w35980_,
		_w35979_,
		_w35982_,
		_w36229_
	);
	LUT4 #(
		.INIT('h0100)
	) name30403 (
		_w36190_,
		_w36229_,
		_w36227_,
		_w36228_,
		_w36230_
	);
	LUT2 #(
		.INIT('h2)
	) name30404 (
		_w35990_,
		_w35995_,
		_w36231_
	);
	LUT4 #(
		.INIT('h2000)
	) name30405 (
		_w35980_,
		_w35981_,
		_w35979_,
		_w35984_,
		_w36232_
	);
	LUT4 #(
		.INIT('h0037)
	) name30406 (
		_w35998_,
		_w36187_,
		_w36198_,
		_w36232_,
		_w36233_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name30407 (
		_w36226_,
		_w36230_,
		_w36231_,
		_w36233_,
		_w36234_
	);
	LUT3 #(
		.INIT('ha9)
	) name30408 (
		\u2_L14_reg[23]/P0001 ,
		_w36224_,
		_w36234_,
		_w36235_
	);
	LUT4 #(
		.INIT('h0fe5)
	) name30409 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36236_
	);
	LUT4 #(
		.INIT('h0100)
	) name30410 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36237_
	);
	LUT4 #(
		.INIT('h0501)
	) name30411 (
		_w35816_,
		_w35817_,
		_w36237_,
		_w36236_,
		_w36238_
	);
	LUT4 #(
		.INIT('h0008)
	) name30412 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35817_,
		_w36239_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name30413 (
		_w35816_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36240_
	);
	LUT4 #(
		.INIT('h0100)
	) name30414 (
		_w35821_,
		_w35820_,
		_w35818_,
		_w35817_,
		_w36241_
	);
	LUT4 #(
		.INIT('hf7bf)
	) name30415 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36242_
	);
	LUT4 #(
		.INIT('h1000)
	) name30416 (
		_w36241_,
		_w36239_,
		_w36240_,
		_w36242_,
		_w36243_
	);
	LUT4 #(
		.INIT('h0020)
	) name30417 (
		_w35821_,
		_w35819_,
		_w35820_,
		_w35818_,
		_w36244_
	);
	LUT3 #(
		.INIT('h10)
	) name30418 (
		_w35816_,
		_w35820_,
		_w35818_,
		_w36245_
	);
	LUT4 #(
		.INIT('h0008)
	) name30419 (
		_w36084_,
		_w36081_,
		_w36244_,
		_w36245_,
		_w36246_
	);
	LUT3 #(
		.INIT('h02)
	) name30420 (
		_w35817_,
		_w35829_,
		_w36041_,
		_w36247_
	);
	LUT4 #(
		.INIT('heee0)
	) name30421 (
		_w36238_,
		_w36243_,
		_w36246_,
		_w36247_,
		_w36248_
	);
	LUT2 #(
		.INIT('h9)
	) name30422 (
		\u2_L14_reg[15]/P0001 ,
		_w36248_,
		_w36249_
	);
	LUT4 #(
		.INIT('h0a04)
	) name30423 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36250_
	);
	LUT4 #(
		.INIT('h4080)
	) name30424 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36251_
	);
	LUT2 #(
		.INIT('h2)
	) name30425 (
		_w35962_,
		_w35959_,
		_w36252_
	);
	LUT2 #(
		.INIT('h4)
	) name30426 (
		_w35962_,
		_w35959_,
		_w36253_
	);
	LUT2 #(
		.INIT('h9)
	) name30427 (
		_w35962_,
		_w35959_,
		_w36254_
	);
	LUT4 #(
		.INIT('h0100)
	) name30428 (
		_w36121_,
		_w36250_,
		_w36251_,
		_w36254_,
		_w36255_
	);
	LUT4 #(
		.INIT('h44a8)
	) name30429 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36256_
	);
	LUT3 #(
		.INIT('h41)
	) name30430 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w36257_
	);
	LUT3 #(
		.INIT('h02)
	) name30431 (
		_w36252_,
		_w36257_,
		_w36256_,
		_w36258_
	);
	LUT4 #(
		.INIT('h2000)
	) name30432 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36259_
	);
	LUT3 #(
		.INIT('h20)
	) name30433 (
		_w35954_,
		_w35955_,
		_w35957_,
		_w36260_
	);
	LUT4 #(
		.INIT('h957a)
	) name30434 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36261_
	);
	LUT3 #(
		.INIT('h04)
	) name30435 (
		_w36121_,
		_w36253_,
		_w36261_,
		_w36262_
	);
	LUT4 #(
		.INIT('h00f1)
	) name30436 (
		_w36255_,
		_w36258_,
		_w36259_,
		_w36262_,
		_w36263_
	);
	LUT2 #(
		.INIT('h6)
	) name30437 (
		\u2_L14_reg[7]/P0001 ,
		_w36263_,
		_w36264_
	);
	LUT4 #(
		.INIT('hdeb9)
	) name30438 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36265_
	);
	LUT2 #(
		.INIT('h1)
	) name30439 (
		_w35959_,
		_w36265_,
		_w36266_
	);
	LUT4 #(
		.INIT('h0080)
	) name30440 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36267_
	);
	LUT4 #(
		.INIT('h134e)
	) name30441 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36268_
	);
	LUT3 #(
		.INIT('h70)
	) name30442 (
		_w35956_,
		_w35957_,
		_w35959_,
		_w36269_
	);
	LUT3 #(
		.INIT('h45)
	) name30443 (
		_w36267_,
		_w36268_,
		_w36269_,
		_w36270_
	);
	LUT3 #(
		.INIT('h8a)
	) name30444 (
		_w35962_,
		_w36266_,
		_w36270_,
		_w36271_
	);
	LUT4 #(
		.INIT('h6fb7)
	) name30445 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36272_
	);
	LUT4 #(
		.INIT('h545e)
	) name30446 (
		_w35959_,
		_w35972_,
		_w35974_,
		_w36260_,
		_w36273_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name30447 (
		_w35954_,
		_w35955_,
		_w35956_,
		_w35957_,
		_w36274_
	);
	LUT3 #(
		.INIT('h72)
	) name30448 (
		_w35959_,
		_w35966_,
		_w36274_,
		_w36275_
	);
	LUT4 #(
		.INIT('hea00)
	) name30449 (
		_w35962_,
		_w36272_,
		_w36273_,
		_w36275_,
		_w36276_
	);
	LUT3 #(
		.INIT('h65)
	) name30450 (
		\u2_L14_reg[32]/P0001 ,
		_w36271_,
		_w36276_,
		_w36277_
	);
	LUT4 #(
		.INIT('h6260)
	) name30451 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36278_
	);
	LUT3 #(
		.INIT('h01)
	) name30452 (
		_w36096_,
		_w36101_,
		_w36278_,
		_w36279_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name30453 (
		_w36096_,
		_w36090_,
		_w36093_,
		_w36094_,
		_w36280_
	);
	LUT4 #(
		.INIT('heb4b)
	) name30454 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36281_
	);
	LUT2 #(
		.INIT('h8)
	) name30455 (
		_w36280_,
		_w36281_,
		_w36282_
	);
	LUT3 #(
		.INIT('h54)
	) name30456 (
		_w36089_,
		_w36279_,
		_w36282_,
		_w36283_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name30457 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36284_
	);
	LUT4 #(
		.INIT('hd8fa)
	) name30458 (
		_w36096_,
		_w36100_,
		_w36158_,
		_w36284_,
		_w36285_
	);
	LUT3 #(
		.INIT('h8a)
	) name30459 (
		_w36089_,
		_w36157_,
		_w36162_,
		_w36286_
	);
	LUT2 #(
		.INIT('h4)
	) name30460 (
		_w36285_,
		_w36286_,
		_w36287_
	);
	LUT3 #(
		.INIT('h80)
	) name30461 (
		_w36090_,
		_w36093_,
		_w36094_,
		_w36288_
	);
	LUT4 #(
		.INIT('h002a)
	) name30462 (
		_w36096_,
		_w36090_,
		_w36093_,
		_w36091_,
		_w36289_
	);
	LUT4 #(
		.INIT('h135f)
	) name30463 (
		_w36116_,
		_w36097_,
		_w36288_,
		_w36289_,
		_w36290_
	);
	LUT4 #(
		.INIT('ha955)
	) name30464 (
		\u2_L14_reg[24]/P0001 ,
		_w36283_,
		_w36287_,
		_w36290_,
		_w36291_
	);
	LUT4 #(
		.INIT('h3dc3)
	) name30465 (
		_w36096_,
		_w36090_,
		_w36093_,
		_w36094_,
		_w36292_
	);
	LUT4 #(
		.INIT('h0104)
	) name30466 (
		_w36096_,
		_w36090_,
		_w36093_,
		_w36091_,
		_w36293_
	);
	LUT4 #(
		.INIT('h0302)
	) name30467 (
		_w36091_,
		_w36160_,
		_w36293_,
		_w36292_,
		_w36294_
	);
	LUT4 #(
		.INIT('h2880)
	) name30468 (
		_w36096_,
		_w36090_,
		_w36093_,
		_w36094_,
		_w36295_
	);
	LUT4 #(
		.INIT('h76ba)
	) name30469 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36296_
	);
	LUT4 #(
		.INIT('h0f02)
	) name30470 (
		_w36096_,
		_w36167_,
		_w36295_,
		_w36296_,
		_w36297_
	);
	LUT4 #(
		.INIT('hdfef)
	) name30471 (
		_w36090_,
		_w36093_,
		_w36091_,
		_w36094_,
		_w36298_
	);
	LUT4 #(
		.INIT('h0040)
	) name30472 (
		_w36096_,
		_w36090_,
		_w36091_,
		_w36094_,
		_w36299_
	);
	LUT3 #(
		.INIT('h0d)
	) name30473 (
		_w36096_,
		_w36298_,
		_w36299_,
		_w36300_
	);
	LUT4 #(
		.INIT('hd800)
	) name30474 (
		_w36089_,
		_w36294_,
		_w36297_,
		_w36300_,
		_w36301_
	);
	LUT2 #(
		.INIT('h9)
	) name30475 (
		\u2_L14_reg[16]/P0001 ,
		_w36301_,
		_w36302_
	);
	LUT4 #(
		.INIT('hbfbe)
	) name30476 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36303_
	);
	LUT3 #(
		.INIT('h02)
	) name30477 (
		_w35710_,
		_w35713_,
		_w35708_,
		_w36304_
	);
	LUT4 #(
		.INIT('h0031)
	) name30478 (
		_w35708_,
		_w36153_,
		_w36303_,
		_w36304_,
		_w36305_
	);
	LUT2 #(
		.INIT('h2)
	) name30479 (
		_w35707_,
		_w36305_,
		_w36306_
	);
	LUT4 #(
		.INIT('h2030)
	) name30480 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36307_
	);
	LUT4 #(
		.INIT('hf351)
	) name30481 (
		_w35712_,
		_w35716_,
		_w35903_,
		_w36307_,
		_w36308_
	);
	LUT4 #(
		.INIT('hf6dd)
	) name30482 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36309_
	);
	LUT4 #(
		.INIT('he5df)
	) name30483 (
		_w35709_,
		_w35710_,
		_w35711_,
		_w35713_,
		_w36310_
	);
	LUT3 #(
		.INIT('hb1)
	) name30484 (
		_w35708_,
		_w35909_,
		_w36310_,
		_w36311_
	);
	LUT4 #(
		.INIT('hba00)
	) name30485 (
		_w35707_,
		_w36308_,
		_w36309_,
		_w36311_,
		_w36312_
	);
	LUT3 #(
		.INIT('h65)
	) name30486 (
		\u2_L14_reg[8]/P0001 ,
		_w36306_,
		_w36312_,
		_w36313_
	);
	LUT4 #(
		.INIT('h3050)
	) name30487 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36314_
	);
	LUT3 #(
		.INIT('h01)
	) name30488 (
		_w35759_,
		_w35761_,
		_w35762_,
		_w36315_
	);
	LUT4 #(
		.INIT('hfad8)
	) name30489 (
		_w35758_,
		_w35950_,
		_w36314_,
		_w36315_,
		_w36316_
	);
	LUT3 #(
		.INIT('h10)
	) name30490 (
		_w35757_,
		_w35949_,
		_w35935_,
		_w36317_
	);
	LUT4 #(
		.INIT('h4404)
	) name30491 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36318_
	);
	LUT4 #(
		.INIT('h5155)
	) name30492 (
		_w35758_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36319_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name30493 (
		_w35768_,
		_w35943_,
		_w36318_,
		_w36319_,
		_w36320_
	);
	LUT4 #(
		.INIT('h0080)
	) name30494 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36321_
	);
	LUT4 #(
		.INIT('hfd00)
	) name30495 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35757_,
		_w36322_
	);
	LUT2 #(
		.INIT('h4)
	) name30496 (
		_w36321_,
		_w36322_,
		_w36323_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name30497 (
		_w36316_,
		_w36317_,
		_w36320_,
		_w36323_,
		_w36324_
	);
	LUT4 #(
		.INIT('h7df7)
	) name30498 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36325_
	);
	LUT2 #(
		.INIT('h2)
	) name30499 (
		_w35758_,
		_w36325_,
		_w36326_
	);
	LUT4 #(
		.INIT('haabf)
	) name30500 (
		_w35758_,
		_w35759_,
		_w35778_,
		_w36321_,
		_w36327_
	);
	LUT2 #(
		.INIT('h4)
	) name30501 (
		_w36326_,
		_w36327_,
		_w36328_
	);
	LUT3 #(
		.INIT('h65)
	) name30502 (
		\u2_L14_reg[1]/P0001 ,
		_w36324_,
		_w36328_,
		_w36329_
	);
	LUT4 #(
		.INIT('h0eff)
	) name30503 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36330_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name30504 (
		_w35758_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36331_
	);
	LUT4 #(
		.INIT('h04cc)
	) name30505 (
		_w35758_,
		_w35759_,
		_w36330_,
		_w36331_,
		_w36332_
	);
	LUT3 #(
		.INIT('h01)
	) name30506 (
		_w35758_,
		_w35761_,
		_w36330_,
		_w36333_
	);
	LUT4 #(
		.INIT('h0002)
	) name30507 (
		_w35758_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36334_
	);
	LUT4 #(
		.INIT('hff7b)
	) name30508 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36335_
	);
	LUT2 #(
		.INIT('h4)
	) name30509 (
		_w36334_,
		_w36335_,
		_w36336_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name30510 (
		_w35757_,
		_w36332_,
		_w36333_,
		_w36336_,
		_w36337_
	);
	LUT2 #(
		.INIT('h2)
	) name30511 (
		_w35785_,
		_w35763_,
		_w36338_
	);
	LUT3 #(
		.INIT('h01)
	) name30512 (
		_w35768_,
		_w35764_,
		_w35787_,
		_w36339_
	);
	LUT3 #(
		.INIT('h45)
	) name30513 (
		_w35757_,
		_w36338_,
		_w36339_,
		_w36340_
	);
	LUT4 #(
		.INIT('h4014)
	) name30514 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36341_
	);
	LUT4 #(
		.INIT('hfdcc)
	) name30515 (
		_w35759_,
		_w35760_,
		_w35761_,
		_w35762_,
		_w36342_
	);
	LUT4 #(
		.INIT('h0504)
	) name30516 (
		_w35758_,
		_w35757_,
		_w36341_,
		_w36342_,
		_w36343_
	);
	LUT3 #(
		.INIT('h02)
	) name30517 (
		_w35758_,
		_w35769_,
		_w35764_,
		_w36344_
	);
	LUT2 #(
		.INIT('h1)
	) name30518 (
		_w36343_,
		_w36344_,
		_w36345_
	);
	LUT4 #(
		.INIT('h5556)
	) name30519 (
		\u2_L14_reg[26]/P0001 ,
		_w36337_,
		_w36340_,
		_w36345_,
		_w36346_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g16/_0_  = _w5855_ ;
	assign \g191647/_3_  = _w5883_ ;
	assign \g191648/_3_  = _w5916_ ;
	assign \g191819/_3_  = _w5949_ ;
	assign \g191821/_0_  = _w5981_ ;
	assign \g191940/_3_  = _w6010_ ;
	assign \g191941/_0_  = _w6024_ ;
	assign \g191942/_0_  = _w6058_ ;
	assign \g191944/_0_  = _w6073_ ;
	assign \g191945/_0_  = _w6091_ ;
	assign \g191946/_0_  = _w6111_ ;
	assign \g191947/_3_  = _w6129_ ;
	assign \g191948/_0_  = _w6146_ ;
	assign \g191949/_0_  = _w6160_ ;
	assign \g191950/_0_  = _w6186_ ;
	assign \g191951/_3_  = _w6205_ ;
	assign \g191952/_0_  = _w6222_ ;
	assign \g192015/_3_  = _w6239_ ;
	assign \g192016/_3_  = _w6253_ ;
	assign \g192017/_3_  = _w6272_ ;
	assign \g192018/_3_  = _w6287_ ;
	assign \g192019/_3_  = _w6306_ ;
	assign \g192020/_0_  = _w6340_ ;
	assign \g192021/_3_  = _w6353_ ;
	assign \g192022/_0_  = _w6365_ ;
	assign \g192047/_0_  = _w6381_ ;
	assign \g192048/_0_  = _w6397_ ;
	assign \g192049/_0_  = _w6412_ ;
	assign \g192050/_0_  = _w6427_ ;
	assign \g192051/_0_  = _w6439_ ;
	assign \g192081/_0_  = _w6452_ ;
	assign \g193428/_3_  = _w6484_ ;
	assign \g193720/_0_  = _w6517_ ;
	assign \g193721/_0_  = _w6549_ ;
	assign \g193877/_0_  = _w6585_ ;
	assign \g193878/_0_  = _w6599_ ;
	assign \g193879/_0_  = _w6613_ ;
	assign \g193880/_3_  = _w6648_ ;
	assign \g193881/_0_  = _w6678_ ;
	assign \g193882/_0_  = _w6695_ ;
	assign \g193998/_0_  = _w6714_ ;
	assign \g193999/_0_  = _w6732_ ;
	assign \g194000/_3_  = _w6748_ ;
	assign \g194001/_0_  = _w6766_ ;
	assign \g194002/_0_  = _w6801_ ;
	assign \g194003/_0_  = _w6815_ ;
	assign \g194004/_0_  = _w6834_ ;
	assign \g194005/_0_  = _w6854_ ;
	assign \g194006/_0_  = _w6871_ ;
	assign \g194007/_0_  = _w6888_ ;
	assign \g194008/_0_  = _w6904_ ;
	assign \g194009/_0_  = _w6921_ ;
	assign \g194010/_0_  = _w6938_ ;
	assign \g194055/_3_  = _w6953_ ;
	assign \g194056/_3_  = _w6969_ ;
	assign \g194057/_0_  = _w6981_ ;
	assign \g194058/_0_  = _w7012_ ;
	assign \g194059/_0_  = _w7025_ ;
	assign \g194060/_0_  = _w7038_ ;
	assign \g194090/_0_  = _w7055_ ;
	assign \g194091/_0_  = _w7067_ ;
	assign \g194092/_0_  = _w7085_ ;
	assign \g194093/_0_  = _w7101_ ;
	assign \g195671/_0_  = _w7137_ ;
	assign \g195672/_3_  = _w7169_ ;
	assign \g195868/_0_  = _w7198_ ;
	assign \g195869/_0_  = _w7236_ ;
	assign \g195870/_0_  = _w7267_ ;
	assign \g196010/_0_  = _w7282_ ;
	assign \g196011/_0_  = _w7297_ ;
	assign \g196012/_0_  = _w7328_ ;
	assign \g196013/_0_  = _w7344_ ;
	assign \g196014/_0_  = _w7360_ ;
	assign \g196015/_0_  = _w7378_ ;
	assign \g196016/_0_  = _w7399_ ;
	assign \g196017/_0_  = _w7425_ ;
	assign \g196018/_0_  = _w7440_ ;
	assign \g196019/_3_  = _w7459_ ;
	assign \g196020/_0_  = _w7476_ ;
	assign \g196021/_0_  = _w7494_ ;
	assign \g196022/_0_  = _w7511_ ;
	assign \g196096/_3_  = _w7528_ ;
	assign \g196097/_0_  = _w7544_ ;
	assign \g196098/_0_  = _w7560_ ;
	assign \g196099/_0_  = _w7577_ ;
	assign \g196100/_3_  = _w7599_ ;
	assign \g196101/_0_  = _w7630_ ;
	assign \g196102/_0_  = _w7641_ ;
	assign \g196103/_0_  = _w7653_ ;
	assign \g196136/_0_  = _w7670_ ;
	assign \g196137/_0_  = _w7688_ ;
	assign \g196138/_0_  = _w7704_ ;
	assign \g196139/_0_  = _w7717_ ;
	assign \g196140/_0_  = _w7727_ ;
	assign \g196170/_0_  = _w7740_ ;
	assign \g197520/_3_  = _w7772_ ;
	assign \g197821/_0_  = _w7806_ ;
	assign \g197923/_0_  = _w7834_ ;
	assign \g197996/_0_  = _w7870_ ;
	assign \g197997/_3_  = _w7899_ ;
	assign \g197998/_0_  = _w7914_ ;
	assign \g197999/_0_  = _w7947_ ;
	assign \g198000/_0_  = _w7966_ ;
	assign \g198071/_0_  = _w7980_ ;
	assign \g198123/_0_  = _w7992_ ;
	assign \g198124/_0_  = _w8012_ ;
	assign \g198125/_0_  = _w8034_ ;
	assign \g198126/_0_  = _w8051_ ;
	assign \g198127/_0_  = _w8079_ ;
	assign \g198128/_0_  = _w8096_ ;
	assign \g198129/_0_  = _w8113_ ;
	assign \g198130/_0_  = _w8136_ ;
	assign \g198131/_0_  = _w8150_ ;
	assign \g198132/_0_  = _w8167_ ;
	assign \g198133/_0_  = _w8184_ ;
	assign \g198134/_3_  = _w8202_ ;
	assign \g198135/_0_  = _w8220_ ;
	assign \g198182/_0_  = _w8236_ ;
	assign \g198183/_3_  = _w8255_ ;
	assign \g198184/_0_  = _w8269_ ;
	assign \g198185/_0_  = _w8299_ ;
	assign \g198186/_0_  = _w8308_ ;
	assign \g198187/_0_  = _w8321_ ;
	assign \g198219/_0_  = _w8334_ ;
	assign \g198220/_0_  = _w8354_ ;
	assign \g198221/_0_  = _w8369_ ;
	assign \g198222/_0_  = _w8382_ ;
	assign \g199794/_0_  = _w8413_ ;
	assign \g199795/_3_  = _w8445_ ;
	assign \g200006/_0_  = _w8476_ ;
	assign \g200007/_0_  = _w8513_ ;
	assign \g200008/_0_  = _w8543_ ;
	assign \g200139/_0_  = _w8558_ ;
	assign \g200140/_0_  = _w8573_ ;
	assign \g200141/_0_  = _w8603_ ;
	assign \g200142/_0_  = _w8622_ ;
	assign \g200143/_0_  = _w8638_ ;
	assign \g200144/_0_  = _w8659_ ;
	assign \g200145/_0_  = _w8677_ ;
	assign \g200146/_0_  = _w8691_ ;
	assign \g200147/_0_  = _w8717_ ;
	assign \g200148/_0_  = _w8729_ ;
	assign \g200149/_0_  = _w8744_ ;
	assign \g200150/_3_  = _w8763_ ;
	assign \g200151/_0_  = _w8781_ ;
	assign \g200228/_3_  = _w8798_ ;
	assign \g200229/_0_  = _w8813_ ;
	assign \g200230/_0_  = _w8829_ ;
	assign \g200231/_0_  = _w8847_ ;
	assign \g200232/_3_  = _w8863_ ;
	assign \g200233/_0_  = _w8894_ ;
	assign \g200234/_0_  = _w8907_ ;
	assign \g200235/_0_  = _w8919_ ;
	assign \g200268/_0_  = _w8936_ ;
	assign \g200269/_0_  = _w8954_ ;
	assign \g200270/_0_  = _w8970_ ;
	assign \g200271/_0_  = _w8986_ ;
	assign \g200272/_0_  = _w8996_ ;
	assign \g200299/_0_  = _w9009_ ;
	assign \g201655/_3_  = _w9039_ ;
	assign \g201960/_0_  = _w9070_ ;
	assign \g201961/_0_  = _w9098_ ;
	assign \g202131/_0_  = _w9113_ ;
	assign \g202132/_0_  = _w9149_ ;
	assign \g202133/_3_  = _w9181_ ;
	assign \g202134/_0_  = _w9193_ ;
	assign \g202135/_0_  = _w9211_ ;
	assign \g202136/_0_  = _w9239_ ;
	assign \g202257/_0_  = _w9257_ ;
	assign \g202258/_0_  = _w9275_ ;
	assign \g202259/_3_  = _w9293_ ;
	assign \g202260/_0_  = _w9322_ ;
	assign \g202261/_0_  = _w9339_ ;
	assign \g202262/_0_  = _w9354_ ;
	assign \g202263/_0_  = _w9369_ ;
	assign \g202264/_0_  = _w9387_ ;
	assign \g202265/_0_  = _w9403_ ;
	assign \g202266/_0_  = _w9419_ ;
	assign \g202267/_0_  = _w9435_ ;
	assign \g202268/_0_  = _w9450_ ;
	assign \g202269/_0_  = _w9463_ ;
	assign \g202317/_0_  = _w9478_ ;
	assign \g202318/_3_  = _w9494_ ;
	assign \g202319/_0_  = _w9509_ ;
	assign \g202320/_0_  = _w9534_ ;
	assign \g202321/_0_  = _w9545_ ;
	assign \g202322/_0_  = _w9557_ ;
	assign \g202354/_0_  = _w9572_ ;
	assign \g202355/_0_  = _w9584_ ;
	assign \g202356/_0_  = _w9603_ ;
	assign \g202357/_0_  = _w9620_ ;
	assign \g203927/_0_  = _w9647_ ;
	assign \g203928/_3_  = _w9676_ ;
	assign \g204142/_0_  = _w9705_ ;
	assign \g204143/_0_  = _w9740_ ;
	assign \g204144/_0_  = _w9774_ ;
	assign \g204275/_0_  = _w9794_ ;
	assign \g204276/_0_  = _w9808_ ;
	assign \g204277/_0_  = _w9826_ ;
	assign \g204278/_0_  = _w9842_ ;
	assign \g204279/_0_  = _w9872_ ;
	assign \g204280/_0_  = _w9888_ ;
	assign \g204281/_0_  = _w9910_ ;
	assign \g204282/_0_  = _w9928_ ;
	assign \g204283/_0_  = _w9948_ ;
	assign \g204284/_0_  = _w9971_ ;
	assign \g204285/_0_  = _w9985_ ;
	assign \g204286/_3_  = _w10005_ ;
	assign \g204287/_0_  = _w10023_ ;
	assign \g204363/_3_  = _w10039_ ;
	assign \g204364/_0_  = _w10051_ ;
	assign \g204365/_0_  = _w10067_ ;
	assign \g204366/_0_  = _w10082_ ;
	assign \g204367/_3_  = _w10097_ ;
	assign \g204368/_0_  = _w10131_ ;
	assign \g204369/_0_  = _w10145_ ;
	assign \g204370/_0_  = _w10157_ ;
	assign \g204403/_0_  = _w10173_ ;
	assign \g204404/_0_  = _w10189_ ;
	assign \g204405/_0_  = _w10204_ ;
	assign \g204406/_0_  = _w10221_ ;
	assign \g204407/_0_  = _w10236_ ;
	assign \g204434/_0_  = _w10248_ ;
	assign \g205833/_3_  = _w10277_ ;
	assign \g206103/_0_  = _w10310_ ;
	assign \g206104/_0_  = _w10340_ ;
	assign \g206266/_0_  = _w10354_ ;
	assign \g206267/_0_  = _w10386_ ;
	assign \g206268/_0_  = _w10400_ ;
	assign \g206269/_3_  = _w10431_ ;
	assign \g206270/_0_  = _w10448_ ;
	assign \g206271/_0_  = _w10473_ ;
	assign \g206387/_0_  = _w10493_ ;
	assign \g206388/_0_  = _w10509_ ;
	assign \g206389/_3_  = _w10529_ ;
	assign \g206390/_0_  = _w10558_ ;
	assign \g206391/_0_  = _w10576_ ;
	assign \g206392/_0_  = _w10590_ ;
	assign \g206393/_0_  = _w10607_ ;
	assign \g206394/_0_  = _w10625_ ;
	assign \g206395/_0_  = _w10641_ ;
	assign \g206396/_0_  = _w10657_ ;
	assign \g206397/_0_  = _w10677_ ;
	assign \g206398/_0_  = _w10694_ ;
	assign \g206399/_0_  = _w10707_ ;
	assign \g206446/_0_  = _w10723_ ;
	assign \g206447/_3_  = _w10739_ ;
	assign \g206448/_0_  = _w10754_ ;
	assign \g206449/_0_  = _w10779_ ;
	assign \g206450/_0_  = _w10791_ ;
	assign \g206451/_0_  = _w10801_ ;
	assign \g206483/_0_  = _w10816_ ;
	assign \g206484/_0_  = _w10828_ ;
	assign \g206485/_0_  = _w10847_ ;
	assign \g206486/_0_  = _w10864_ ;
	assign \g208069/_0_  = _w10892_ ;
	assign \g208070/_3_  = _w10924_ ;
	assign \g208253/_0_  = _w10955_ ;
	assign \g208254/_0_  = _w10989_ ;
	assign \g208255/_0_  = _w11013_ ;
	assign \g208406/_0_  = _w11029_ ;
	assign \g208407/_0_  = _w11046_ ;
	assign \g208408/_0_  = _w11076_ ;
	assign \g208409/_0_  = _w11094_ ;
	assign \g208410/_0_  = _w11110_ ;
	assign \g208411/_0_  = _w11127_ ;
	assign \g208412/_0_  = _w11149_ ;
	assign \g208413/_0_  = _w11167_ ;
	assign \g208414/_0_  = _w11182_ ;
	assign \g208415/_3_  = _w11217_ ;
	assign \g208416/_0_  = _w11229_ ;
	assign \g208417/_0_  = _w11247_ ;
	assign \g208418/_0_  = _w11265_ ;
	assign \g208493/_3_  = _w11281_ ;
	assign \g208494/_0_  = _w11296_ ;
	assign \g208495/_0_  = _w11313_ ;
	assign \g208496/_0_  = _w11329_ ;
	assign \g208497/_3_  = _w11343_ ;
	assign \g208498/_0_  = _w11374_ ;
	assign \g208499/_0_  = _w11388_ ;
	assign \g208500/_0_  = _w11400_ ;
	assign \g208533/_0_  = _w11417_ ;
	assign \g208534/_0_  = _w11435_ ;
	assign \g208535/_0_  = _w11451_ ;
	assign \g208536/_0_  = _w11468_ ;
	assign \g208537/_0_  = _w11479_ ;
	assign \g208564/_0_  = _w11492_ ;
	assign \g209938/_3_  = _w11527_ ;
	assign \g210205/_0_  = _w11558_ ;
	assign \g210206/_0_  = _w11589_ ;
	assign \g210380/_0_  = _w11607_ ;
	assign \g210381/_0_  = _w11638_ ;
	assign \g210382/_0_  = _w11650_ ;
	assign \g210383/_3_  = _w11681_ ;
	assign \g210384/_0_  = _w11699_ ;
	assign \g210385/_0_  = _w11727_ ;
	assign \g210499/_0_  = _w11747_ ;
	assign \g210500/_0_  = _w11761_ ;
	assign \g210501/_3_  = _w11781_ ;
	assign \g210502/_0_  = _w11799_ ;
	assign \g210503/_0_  = _w11832_ ;
	assign \g210504/_0_  = _w11847_ ;
	assign \g210505/_0_  = _w11862_ ;
	assign \g210506/_0_  = _w11882_ ;
	assign \g210507/_0_  = _w11899_ ;
	assign \g210508/_0_  = _w11916_ ;
	assign \g210509/_0_  = _w11934_ ;
	assign \g210510/_0_  = _w11951_ ;
	assign \g210511/_0_  = _w11963_ ;
	assign \g210558/_0_  = _w11979_ ;
	assign \g210559/_3_  = _w11996_ ;
	assign \g210560/_0_  = _w12012_ ;
	assign \g210561/_0_  = _w12041_ ;
	assign \g210562/_0_  = _w12053_ ;
	assign \g210563/_0_  = _w12064_ ;
	assign \g210595/_0_  = _w12081_ ;
	assign \g210596/_0_  = _w12093_ ;
	assign \g210597/_0_  = _w12108_ ;
	assign \g210598/_0_  = _w12124_ ;
	assign \g212159/_0_  = _w12154_ ;
	assign \g212160/_3_  = _w12187_ ;
	assign \g212384/_0_  = _w12218_ ;
	assign \g212385/_0_  = _w12255_ ;
	assign \g212386/_0_  = _w12287_ ;
	assign \g212536/_0_  = _w12301_ ;
	assign \g212537/_0_  = _w12318_ ;
	assign \g212538/_0_  = _w12348_ ;
	assign \g212539/_0_  = _w12363_ ;
	assign \g212540/_0_  = _w12378_ ;
	assign \g212541/_0_  = _w12395_ ;
	assign \g212542/_0_  = _w12413_ ;
	assign \g212543/_0_  = _w12427_ ;
	assign \g212544/_0_  = _w12439_ ;
	assign \g212545/_0_  = _w12457_ ;
	assign \g212546/_3_  = _w12488_ ;
	assign \g212547/_0_  = _w12506_ ;
	assign \g212623/_3_  = _w12526_ ;
	assign \g212624/_0_  = _w12541_ ;
	assign \g212625/_0_  = _w12559_ ;
	assign \g212626/_0_  = _w12577_ ;
	assign \g212627/_0_  = _w12594_ ;
	assign \g212628/_3_  = _w12610_ ;
	assign \g212629/_0_  = _w12641_ ;
	assign \g212630/_0_  = _w12654_ ;
	assign \g212631/_0_  = _w12666_ ;
	assign \g212667/_0_  = _w12683_ ;
	assign \g212668/_0_  = _w12701_ ;
	assign \g212669/_0_  = _w12717_ ;
	assign \g212670/_0_  = _w12734_ ;
	assign \g212671/_0_  = _w12745_ ;
	assign \g212699/_0_  = _w12757_ ;
	assign \g214033/_3_  = _w12787_ ;
	assign \g214309/_3_  = _w12818_ ;
	assign \g214310/_0_  = _w12849_ ;
	assign \g214494/_0_  = _w12865_ ;
	assign \g214495/_0_  = _w12901_ ;
	assign \g214496/_0_  = _w12913_ ;
	assign \g214497/_3_  = _w12944_ ;
	assign \g214632/_0_  = _w12962_ ;
	assign \g214633/_0_  = _w12980_ ;
	assign \g214634/_3_  = _w13000_ ;
	assign \g214635/_0_  = _w13034_ ;
	assign \g214636/_0_  = _w13061_ ;
	assign \g214637/_0_  = _w13076_ ;
	assign \g214638/_0_  = _w13100_ ;
	assign \g214639/_0_  = _w13117_ ;
	assign \g214640/_0_  = _w13133_ ;
	assign \g214641/_0_  = _w13150_ ;
	assign \g214642/_0_  = _w13167_ ;
	assign \g214643/_0_  = _w13185_ ;
	assign \g214691/_0_  = _w13200_ ;
	assign \g214692/_0_  = _w13222_ ;
	assign \g214693/_3_  = _w13238_ ;
	assign \g214694/_0_  = _w13263_ ;
	assign \g214695/_0_  = _w13278_ ;
	assign \g214696/_0_  = _w13292_ ;
	assign \g214697/_0_  = _w13303_ ;
	assign \g214729/_0_  = _w13318_ ;
	assign \g214730/_0_  = _w13330_ ;
	assign \g214731/_0_  = _w13349_ ;
	assign \g214732/_0_  = _w13366_ ;
	assign \g214733/_0_  = _w13382_ ;
	assign \g216157/_0_  = _w13409_ ;
	assign \g216158/_3_  = _w13442_ ;
	assign \g216492/_0_  = _w13473_ ;
	assign \g216493/_0_  = _w13501_ ;
	assign \g216671/_0_  = _w13515_ ;
	assign \g216672/_0_  = _w13529_ ;
	assign \g216673/_0_  = _w13565_ ;
	assign \g216674/_0_  = _w13590_ ;
	assign \g216675/_0_  = _w13605_ ;
	assign \g216676/_3_  = _w13626_ ;
	assign \g216677/_0_  = _w13641_ ;
	assign \g216735/_0_  = _w13658_ ;
	assign \g216736/_3_  = _w13677_ ;
	assign \g216737/_0_  = _w13695_ ;
	assign \g216738/_0_  = _w13729_ ;
	assign \g216739/_0_  = _w13744_ ;
	assign \g216740/_0_  = _w13764_ ;
	assign \g216741/_0_  = _w13782_ ;
	assign \g216742/_0_  = _w13800_ ;
	assign \g216743/_0_  = _w13816_ ;
	assign \g216744/_0_  = _w13831_ ;
	assign \g216745/_0_  = _w13847_ ;
	assign \g216746/_3_  = _w13862_ ;
	assign \g216747/_0_  = _w13893_ ;
	assign \g216748/_0_  = _w13907_ ;
	assign \g216749/_0_  = _w13921_ ;
	assign \g216788/_0_  = _w13938_ ;
	assign \g216789/_0_  = _w13956_ ;
	assign \g216790/_0_  = _w13972_ ;
	assign \g216791/_0_  = _w13987_ ;
	assign \g216792/_0_  = _w14001_ ;
	assign \g216829/_0_  = _w14013_ ;
	assign \g218407/_3_  = _w14045_ ;
	assign \g218408/_0_  = _w14072_ ;
	assign \g218423/_3_  = _w14105_ ;
	assign \g218601/_0_  = _w14140_ ;
	assign \g218602/_0_  = _w14154_ ;
	assign \g218603/_0_  = _w14171_ ;
	assign \g218604/_0_  = _w14199_ ;
	assign \g218724/_0_  = _w14213_ ;
	assign \g218725/_0_  = _w14231_ ;
	assign \g218726/_0_  = _w14263_ ;
	assign \g218727/_0_  = _w14278_ ;
	assign \g218728/_0_  = _w14292_ ;
	assign \g218729/_0_  = _w14312_ ;
	assign \g218730/_0_  = _w14330_ ;
	assign \g218731/_0_  = _w14350_ ;
	assign \g218732/_0_  = _w14368_ ;
	assign \g218733/_0_  = _w14385_ ;
	assign \g218734/_0_  = _w14408_ ;
	assign \g218735/_3_  = _w14428_ ;
	assign \g218736/_0_  = _w14441_ ;
	assign \g218808/_3_  = _w14457_ ;
	assign \g218809/_0_  = _w14475_ ;
	assign \g218810/_0_  = _w14491_ ;
	assign \g218811/_3_  = _w14504_ ;
	assign \g218812/_0_  = _w14519_ ;
	assign \g218813/_0_  = _w14548_ ;
	assign \g218814/_0_  = _w14562_ ;
	assign \g218846/_0_  = _w14580_ ;
	assign \g218847/_0_  = _w14594_ ;
	assign \g218848/_0_  = _w14609_ ;
	assign \g218849/_0_  = _w14620_ ;
	assign \g218877/_0_  = _w14632_ ;
	assign \g22/_0_  = _w14655_ ;
	assign \g220545/_0_  = _w14684_ ;
	assign \g220546/_3_  = _w14723_ ;
	assign \g220725/_3_  = _w14754_ ;
	assign \g220726/_0_  = _w14790_ ;
	assign \g220793/_0_  = _w14807_ ;
	assign \g220794/_0_  = _w14824_ ;
	assign \g220795/_0_  = _w14857_ ;
	assign \g220796/_0_  = _w14884_ ;
	assign \g220797/_0_  = _w14898_ ;
	assign \g220798/_0_  = _w14912_ ;
	assign \g220799/_0_  = _w14930_ ;
	assign \g220800/_0_  = _w14953_ ;
	assign \g220801/_0_  = _w14968_ ;
	assign \g220802/_0_  = _w14991_ ;
	assign \g220803/_0_  = _w15006_ ;
	assign \g220804/_3_  = _w15026_ ;
	assign \g220805/_0_  = _w15042_ ;
	assign \g220806/_0_  = _w15058_ ;
	assign \g220807/_0_  = _w15075_ ;
	assign \g220872/_3_  = _w15091_ ;
	assign \g220873/_0_  = _w15110_ ;
	assign \g220874/_3_  = _w15127_ ;
	assign \g220875/_0_  = _w15158_ ;
	assign \g220876/_0_  = _w15173_ ;
	assign \g220877/_0_  = _w15185_ ;
	assign \g220921/_0_  = _w15202_ ;
	assign \g220922/_0_  = _w15220_ ;
	assign \g220923/_0_  = _w15234_ ;
	assign \g220924/_0_  = _w15250_ ;
	assign \g220925/_0_  = _w15265_ ;
	assign \g220926/_0_  = _w15278_ ;
	assign \g220969/_0_  = _w15290_ ;
	assign \g221011/_3_  = _w15320_ ;
	assign \g221039/_3_  = _w15352_ ;
	assign \g221086/_3_  = _w15386_ ;
	assign \g221131/_0_  = _w15410_ ;
	assign \g224010/_3_  = _w15444_ ;
	assign \g224368/_3_  = _w15472_ ;
	assign \g224369/_3_  = _w15500_ ;
	assign \g224532/_0_  = _w15521_ ;
	assign \g224533/_0_  = _w15535_ ;
	assign \g224534/_0_  = _w15570_ ;
	assign \g224535/_3_  = _w15601_ ;
	assign \g224536/_0_  = _w15616_ ;
	assign \g224537/_0_  = _w15651_ ;
	assign \g224640/_3_  = _w15671_ ;
	assign \g224641/_0_  = _w15701_ ;
	assign \g224642/_0_  = _w15720_ ;
	assign \g224643/_3_  = _w15736_ ;
	assign \g224644/_0_  = _w15754_ ;
	assign \g224645/_0_  = _w15771_ ;
	assign \g224646/_3_  = _w15782_ ;
	assign \g224647/_0_  = _w15799_ ;
	assign \g224648/_3_  = _w15818_ ;
	assign \g224649/_0_  = _w15836_ ;
	assign \g224650/_0_  = _w15851_ ;
	assign \g224651/_0_  = _w15868_ ;
	assign \g224652/_0_  = _w15882_ ;
	assign \g224690/_0_  = _w15892_ ;
	assign \g224691/_3_  = _w15907_ ;
	assign \g224692/_3_  = _w15923_ ;
	assign \g224693/_0_  = _w15939_ ;
	assign \g224694/_0_  = _w15964_ ;
	assign \g224695/_3_  = _w15980_ ;
	assign \g224723/_0_  = _w16001_ ;
	assign \g224724/_0_  = _w16017_ ;
	assign \g224725/_0_  = _w16031_ ;
	assign \g224726/_0_  = _w16049_ ;
	assign \g226372/_0_  = _w16079_ ;
	assign \g226373/_3_  = _w16113_ ;
	assign \g226549/_3_  = _w16147_ ;
	assign \g226550/_0_  = _w16185_ ;
	assign \g226616/_0_  = _w16201_ ;
	assign \g226635/_0_  = _w16215_ ;
	assign \g226636/_0_  = _w16248_ ;
	assign \g226637/_0_  = _w16266_ ;
	assign \g226638/_0_  = _w16283_ ;
	assign \g226639/_0_  = _w16299_ ;
	assign \g226640/_0_  = _w16316_ ;
	assign \g226641/_3_  = _w16347_ ;
	assign \g226642/_0_  = _w16366_ ;
	assign \g226643/_0_  = _w16384_ ;
	assign \g226644/_0_  = _w16401_ ;
	assign \g226645/_0_  = _w16432_ ;
	assign \g226646/_0_  = _w16448_ ;
	assign \g226692/_3_  = _w16467_ ;
	assign \g226693/_0_  = _w16480_ ;
	assign \g226694/_3_  = _w16498_ ;
	assign \g226695/_3_  = _w16517_ ;
	assign \g226696/_3_  = _w16534_ ;
	assign \g226697/_0_  = _w16565_ ;
	assign \g226698/_0_  = _w16578_ ;
	assign \g226699/_0_  = _w16592_ ;
	assign \g226728/_0_  = _w16611_ ;
	assign \g226729/_0_  = _w16628_ ;
	assign \g226730/_0_  = _w16643_ ;
	assign \g226731/_0_  = _w16653_ ;
	assign \g226732/_0_  = _w16668_ ;
	assign \g226759/_0_  = _w16680_ ;
	assign \g228250/_0_  = _w16718_ ;
	assign \g228396/_0_  = _w16752_ ;
	assign \g228397/_0_  = _w16782_ ;
	assign \g228566/_0_  = _w16818_ ;
	assign \g228567/_0_  = _w16834_ ;
	assign \g228568/_0_  = _w16863_ ;
	assign \g228609/_0_  = _w16878_ ;
	assign \g228610/_3_  = _w16912_ ;
	assign \g228688/_0_  = _w16929_ ;
	assign \g228689/_0_  = _w16943_ ;
	assign \g228690/_3_  = _w16963_ ;
	assign \g228691/_0_  = _w16980_ ;
	assign \g228692/_0_  = _w16992_ ;
	assign \g228693/_0_  = _w17013_ ;
	assign \g228694/_0_  = _w17028_ ;
	assign \g228695/_0_  = _w17045_ ;
	assign \g228696/_0_  = _w17073_ ;
	assign \g228697/_0_  = _w17090_ ;
	assign \g228698/_0_  = _w17117_ ;
	assign \g228699/_0_  = _w17134_ ;
	assign \g228700/_0_  = _w17149_ ;
	assign \g228748/_0_  = _w17167_ ;
	assign \g228749/_3_  = _w17185_ ;
	assign \g228750/_0_  = _w17200_ ;
	assign \g228751/_0_  = _w17227_ ;
	assign \g228752/_0_  = _w17243_ ;
	assign \g228753/_0_  = _w17256_ ;
	assign \g228784/_0_  = _w17272_ ;
	assign \g228785/_0_  = _w17290_ ;
	assign \g228786/_0_  = _w17306_ ;
	assign \g228787/_3_  = _w17318_ ;
	assign \g230339/_0_  = _w17349_ ;
	assign \g230340/_0_  = _w17378_ ;
	assign \g230546/_0_  = _w17415_ ;
	assign \g230580/_0_  = _w17452_ ;
	assign \g230679/_0_  = _w17468_ ;
	assign \g230680/_0_  = _w17484_ ;
	assign \g230681/_0_  = _w17520_ ;
	assign \g230682/_0_  = _w17533_ ;
	assign \g230683/_0_  = _w17562_ ;
	assign \g230684/_0_  = _w17577_ ;
	assign \g230685/_0_  = _w17599_ ;
	assign \g230686/_0_  = _w17615_ ;
	assign \g230687/_0_  = _w17642_ ;
	assign \g230688/_0_  = _w17657_ ;
	assign \g230689/_3_  = _w17680_ ;
	assign \g230690/_0_  = _w17698_ ;
	assign \g230710/_0_  = _w17715_ ;
	assign \g230766/_0_  = _w17727_ ;
	assign \g230767/_0_  = _w17747_ ;
	assign \g230768/_0_  = _w17763_ ;
	assign \g230769/_3_  = _w17778_ ;
	assign \g230770/_0_  = _w17804_ ;
	assign \g230771/_0_  = _w17817_ ;
	assign \g230772/_0_  = _w17831_ ;
	assign \g230773/_3_  = _w17848_ ;
	assign \g230810/_0_  = _w17864_ ;
	assign \g230811/_0_  = _w17882_ ;
	assign \g230812/_0_  = _w17898_ ;
	assign \g230813/_0_  = _w17912_ ;
	assign \g230814/_0_  = _w17924_ ;
	assign \g230840/_3_  = _w17936_ ;
	assign \g232196/_3_  = _w17972_ ;
	assign \g232469/_0_  = _w17998_ ;
	assign \g232470/_0_  = _w18029_ ;
	assign \g232633/_0_  = _w18068_ ;
	assign \g232635/_3_  = _w18104_ ;
	assign \g232636/_0_  = _w18119_ ;
	assign \g232637/_0_  = _w18132_ ;
	assign \g232691/_0_  = _w18164_ ;
	assign \g232747/_0_  = _w18182_ ;
	assign \g232748/_0_  = _w18198_ ;
	assign \g232749/_3_  = _w18219_ ;
	assign \g232750/_0_  = _w18251_ ;
	assign \g232751/_0_  = _w18268_ ;
	assign \g232752/_0_  = _w18284_ ;
	assign \g232753/_0_  = _w18298_ ;
	assign \g232754/_0_  = _w18318_ ;
	assign \g232755/_0_  = _w18340_ ;
	assign \g232756/_0_  = _w18356_ ;
	assign \g232757/_0_  = _w18374_ ;
	assign \g232758/_0_  = _w18387_ ;
	assign \g232759/_0_  = _w18400_ ;
	assign \g232804/_0_  = _w18417_ ;
	assign \g232805/_0_  = _w18432_ ;
	assign \g232806/_0_  = _w18458_ ;
	assign \g232807/_0_  = _w18473_ ;
	assign \g232808/_3_  = _w18488_ ;
	assign \g232809/_0_  = _w18501_ ;
	assign \g232841/_0_  = _w18520_ ;
	assign \g232842/_3_  = _w18533_ ;
	assign \g232843/_0_  = _w18549_ ;
	assign \g232844/_0_  = _w18565_ ;
	assign \g234520/_0_  = _w18590_ ;
	assign \g234687/_0_  = _w18622_ ;
	assign \g234688/_0_  = _w18654_ ;
	assign \g234689/_0_  = _w18687_ ;
	assign \g234764/_0_  = _w18707_ ;
	assign \g234765/_0_  = _w18726_ ;
	assign \g234766/_0_  = _w18756_ ;
	assign \g234767/_3_  = _w18771_ ;
	assign \g234768/_0_  = _w18788_ ;
	assign \g234769/_0_  = _w18811_ ;
	assign \g234770/_0_  = _w18831_ ;
	assign \g234771/_0_  = _w18855_ ;
	assign \g234772/_0_  = _w18868_ ;
	assign \g234773/_0_  = _w18884_ ;
	assign \g234774/_3_  = _w18914_ ;
	assign \g234775/_0_  = _w18931_ ;
	assign \g234776/_0_  = _w18947_ ;
	assign \g234824/_3_  = _w18966_ ;
	assign \g234825/_0_  = _w18979_ ;
	assign \g234826/_0_  = _w18999_ ;
	assign \g234827/_0_  = _w19014_ ;
	assign \g234828/_3_  = _w19029_ ;
	assign \g234829/_0_  = _w19057_ ;
	assign \g234830/_0_  = _w19073_ ;
	assign \g234831/_0_  = _w19086_ ;
	assign \g234867/_0_  = _w19107_ ;
	assign \g234868/_0_  = _w19123_ ;
	assign \g234869/_0_  = _w19137_ ;
	assign \g234870/_0_  = _w19153_ ;
	assign \g234896/_0_  = _w19165_ ;
	assign \g236294/_3_  = _w19199_ ;
	assign \g236541/_0_  = _w19232_ ;
	assign \g236542/_0_  = _w19263_ ;
	assign \g236724/_0_  = _w19280_ ;
	assign \g236725/_0_  = _w19316_ ;
	assign \g236726/_0_  = _w19331_ ;
	assign \g236727/_3_  = _w19359_ ;
	assign \g236728/_0_  = _w19373_ ;
	assign \g236729/_0_  = _w19398_ ;
	assign \g236821/_0_  = _w19414_ ;
	assign \g236822/_3_  = _w19441_ ;
	assign \g236823/_0_  = _w19473_ ;
	assign \g236824/_3_  = _w19489_ ;
	assign \g236825/_0_  = _w19503_ ;
	assign \g236826/_0_  = _w19518_ ;
	assign \g236827/_0_  = _w19538_ ;
	assign \g236828/_0_  = _w19555_ ;
	assign \g236829/_0_  = _w19576_ ;
	assign \g236830/_0_  = _w19596_ ;
	assign \g236831/_0_  = _w19610_ ;
	assign \g236832/_0_  = _w19623_ ;
	assign \g236877/_0_  = _w19638_ ;
	assign \g236878/_3_  = _w19653_ ;
	assign \g236879/_0_  = _w19667_ ;
	assign \g236880/_0_  = _w19694_ ;
	assign \g236881/_0_  = _w19707_ ;
	assign \g236882/_0_  = _w19719_ ;
	assign \g236914/_0_  = _w19737_ ;
	assign \g236915/_0_  = _w19751_ ;
	assign \g236916/_0_  = _w19771_ ;
	assign \g236917/_0_  = _w19788_ ;
	assign \g238530/_0_  = _w19819_ ;
	assign \g238531/_3_  = _w19850_ ;
	assign \g238723/_0_  = _w19884_ ;
	assign \g238724/_0_  = _w19923_ ;
	assign \g238725/_0_  = _w19949_ ;
	assign \g238840/_0_  = _w19967_ ;
	assign \g238841/_0_  = _w19983_ ;
	assign \g238842/_0_  = _w20012_ ;
	assign \g238843/_3_  = _w20030_ ;
	assign \g238844/_0_  = _w20045_ ;
	assign \g238845/_0_  = _w20061_ ;
	assign \g238846/_0_  = _w20083_ ;
	assign \g238847/_0_  = _w20104_ ;
	assign \g238848/_0_  = _w20122_ ;
	assign \g238849/_0_  = _w20144_ ;
	assign \g238850/_0_  = _w20160_ ;
	assign \g238851/_3_  = _w20181_ ;
	assign \g238852/_0_  = _w20196_ ;
	assign \g238924/_0_  = _w20208_ ;
	assign \g238925/_0_  = _w20220_ ;
	assign \g238926/_0_  = _w20235_ ;
	assign \g238927/_3_  = _w20250_ ;
	assign \g238928/_0_  = _w20273_ ;
	assign \g238929/_0_  = _w20286_ ;
	assign \g238930/_0_  = _w20299_ ;
	assign \g238965/_0_  = _w20313_ ;
	assign \g238966/_0_  = _w20331_ ;
	assign \g238967/_0_  = _w20347_ ;
	assign \g238968/_0_  = _w20363_ ;
	assign \g238969/_0_  = _w20377_ ;
	assign \g238996/_0_  = _w20391_ ;
	assign \g240353/_3_  = _w20419_ ;
	assign \g240640/_0_  = _w20453_ ;
	assign \g240641/_0_  = _w20484_ ;
	assign \g240813/_0_  = _w20501_ ;
	assign \g240814/_0_  = _w20537_ ;
	assign \g240815/_3_  = _w20572_ ;
	assign \g240816/_0_  = _w20588_ ;
	assign \g240817/_0_  = _w20618_ ;
	assign \g240818/_0_  = _w20632_ ;
	assign \g240925/_0_  = _w20655_ ;
	assign \g240926/_0_  = _w20671_ ;
	assign \g240927/_3_  = _w20687_ ;
	assign \g240928/_0_  = _w20718_ ;
	assign \g240929/_3_  = _w20736_ ;
	assign \g240930/_0_  = _w20752_ ;
	assign \g240931/_0_  = _w20770_ ;
	assign \g240932/_0_  = _w20788_ ;
	assign \g240933/_0_  = _w20804_ ;
	assign \g240934/_0_  = _w20824_ ;
	assign \g240935/_0_  = _w20842_ ;
	assign \g240936/_0_  = _w20859_ ;
	assign \g240937/_0_  = _w20872_ ;
	assign \g240984/_0_  = _w20890_ ;
	assign \g240985/_3_  = _w20905_ ;
	assign \g240986/_0_  = _w20920_ ;
	assign \g240987/_0_  = _w20948_ ;
	assign \g240988/_0_  = _w20961_ ;
	assign \g240989/_0_  = _w20975_ ;
	assign \g241021/_0_  = _w20989_ ;
	assign \g241022/_0_  = _w21001_ ;
	assign \g241023/_0_  = _w21017_ ;
	assign \g241024/_0_  = _w21034_ ;
	assign \g242616/_0_  = _w21062_ ;
	assign \g242617/_3_  = _w21094_ ;
	assign \g242815/_0_  = _w21127_ ;
	assign \g242816/_0_  = _w21163_ ;
	assign \g242817/_0_  = _w21195_ ;
	assign \g242955/_0_  = _w21213_ ;
	assign \g242956/_0_  = _w21230_ ;
	assign \g242957/_0_  = _w21263_ ;
	assign \g242958/_3_  = _w21280_ ;
	assign \g242959/_0_  = _w21296_ ;
	assign \g242960/_0_  = _w21311_ ;
	assign \g242961/_0_  = _w21331_ ;
	assign \g242962/_0_  = _w21348_ ;
	assign \g242963/_3_  = _w21376_ ;
	assign \g242964/_0_  = _w21392_ ;
	assign \g242965/_0_  = _w21410_ ;
	assign \g242966/_0_  = _w21425_ ;
	assign \g242967/_0_  = _w21443_ ;
	assign \g243037/_3_  = _w21464_ ;
	assign \g243038/_0_  = _w21477_ ;
	assign \g243039/_0_  = _w21497_ ;
	assign \g243040/_0_  = _w21515_ ;
	assign \g243041/_3_  = _w21529_ ;
	assign \g243042/_0_  = _w21558_ ;
	assign \g243043/_0_  = _w21575_ ;
	assign \g243044/_0_  = _w21587_ ;
	assign \g243078/_0_  = _w21598_ ;
	assign \g243079/_0_  = _w21616_ ;
	assign \g243080/_0_  = _w21632_ ;
	assign \g243081/_0_  = _w21645_ ;
	assign \g243082/_0_  = _w21656_ ;
	assign \g243109/_0_  = _w21669_ ;
	assign \g244465/_3_  = _w21694_ ;
	assign \g244753/_3_  = _w21729_ ;
	assign \g244754/_0_  = _w21760_ ;
	assign \g244924/_0_  = _w21797_ ;
	assign \g244925/_0_  = _w21813_ ;
	assign \g244926/_3_  = _w21841_ ;
	assign \g244927/_0_  = _w21858_ ;
	assign \g244928/_0_  = _w21890_ ;
	assign \g245035/_0_  = _w21906_ ;
	assign \g245036/_0_  = _w21922_ ;
	assign \g245037/_0_  = _w21958_ ;
	assign \g245038/_3_  = _w21975_ ;
	assign \g245039/_3_  = _w22002_ ;
	assign \g245040/_0_  = _w22014_ ;
	assign \g245041/_0_  = _w22030_ ;
	assign \g245043/_0_  = _w22048_ ;
	assign \g245045/_0_  = _w22062_ ;
	assign \g245046/_0_  = _w22078_ ;
	assign \g245047/_0_  = _w22089_ ;
	assign \g245092/_0_  = _w22109_ ;
	assign \g245093/_3_  = _w22124_ ;
	assign \g245094/_0_  = _w22137_ ;
	assign \g245095/_0_  = _w22150_ ;
	assign \g245096/_0_  = _w22175_ ;
	assign \g245097/_0_  = _w22185_ ;
	assign \g245129/_0_  = _w22202_ ;
	assign \g245130/_0_  = _w22216_ ;
	assign \g245131/_0_  = _w22234_ ;
	assign \g245132/_0_  = _w22252_ ;
	assign \g246715/_0_  = _w22283_ ;
	assign \g246716/_3_  = _w22314_ ;
	assign \g246911/_0_  = _w22348_ ;
	assign \g246912/_0_  = _w22384_ ;
	assign \g246913/_0_  = _w22415_ ;
	assign \g247057/_0_  = _w22432_ ;
	assign \g247058/_0_  = _w22448_ ;
	assign \g247059/_0_  = _w22481_ ;
	assign \g247060/_0_  = _w22497_ ;
	assign \g247061/_0_  = _w22512_ ;
	assign \g247062/_3_  = _w22532_ ;
	assign \g247063/_0_  = _w22550_ ;
	assign \g247064/_0_  = _w22567_ ;
	assign \g247065/_0_  = _w22584_ ;
	assign \g247066/_0_  = _w22600_ ;
	assign \g247067/_3_  = _w22628_ ;
	assign \g247068/_0_  = _w22646_ ;
	assign \g247069/_0_  = _w22661_ ;
	assign \g247137/_3_  = _w22682_ ;
	assign \g247138/_0_  = _w22694_ ;
	assign \g247139/_0_  = _w22708_ ;
	assign \g247140/_0_  = _w22723_ ;
	assign \g247141/_3_  = _w22738_ ;
	assign \g247142/_0_  = _w22765_ ;
	assign \g247143/_0_  = _w22778_ ;
	assign \g247144/_0_  = _w22790_ ;
	assign \g247179/_0_  = _w22804_ ;
	assign \g247180/_0_  = _w22823_ ;
	assign \g247181/_0_  = _w22837_ ;
	assign \g247182/_0_  = _w22850_ ;
	assign \g247183/_0_  = _w22864_ ;
	assign \g247210/_0_  = _w22877_ ;
	assign \g248581/_3_  = _w22908_ ;
	assign \g248828/_0_  = _w22939_ ;
	assign \g248829/_0_  = _w22967_ ;
	assign \g249033/_0_  = _w22983_ ;
	assign \g249035/_0_  = _w22998_ ;
	assign \g249036/_3_  = _w23025_ ;
	assign \g249037/_0_  = _w23038_ ;
	assign \g249038/_0_  = _w23067_ ;
	assign \g249147/_0_  = _w23099_ ;
	assign \g249148/_0_  = _w23116_ ;
	assign \g249149/_3_  = _w23142_ ;
	assign \g249150/_0_  = _w23164_ ;
	assign \g249152/_0_  = _w23187_ ;
	assign \g249153/_0_  = _w23201_ ;
	assign \g249155/_0_  = _w23217_ ;
	assign \g249156/_0_  = _w23231_ ;
	assign \g249157/_0_  = _w23243_ ;
	assign \g249200/_3_  = _w23261_ ;
	assign \g249201/_0_  = _w23283_ ;
	assign \g249202/_0_  = _w23300_ ;
	assign \g249203/_3_  = _w23314_ ;
	assign \g249204/_0_  = _w23329_ ;
	assign \g249205/_0_  = _w23358_ ;
	assign \g249206/_0_  = _w23375_ ;
	assign \g249207/_0_  = _w23389_ ;
	assign \g249239/_0_  = _w23400_ ;
	assign \g249240/_0_  = _w23412_ ;
	assign \g249241/_0_  = _w23430_ ;
	assign \g249242/_0_  = _w23446_ ;
	assign \g250815/_0_  = _w23473_ ;
	assign \g251006/_0_  = _w23506_ ;
	assign \g251007/_0_  = _w23539_ ;
	assign \g251008/_0_  = _w23570_ ;
	assign \g251009/_3_  = _w23598_ ;
	assign \g251160/_0_  = _w23611_ ;
	assign \g251161/_0_  = _w23628_ ;
	assign \g251162/_0_  = _w23663_ ;
	assign \g251163/_3_  = _w23683_ ;
	assign \g251164/_0_  = _w23707_ ;
	assign \g251165/_0_  = _w23723_ ;
	assign \g251166/_0_  = _w23741_ ;
	assign \g251167/_0_  = _w23756_ ;
	assign \g251168/_0_  = _w23784_ ;
	assign \g251169/_0_  = _w23799_ ;
	assign \g251170/_3_  = _w23823_ ;
	assign \g251171/_0_  = _w23837_ ;
	assign \g251245/_3_  = _w23850_ ;
	assign \g251246/_0_  = _w23865_ ;
	assign \g251247/_0_  = _w23879_ ;
	assign \g251248/_0_  = _w23894_ ;
	assign \g251249/_3_  = _w23905_ ;
	assign \g251250/_0_  = _w23932_ ;
	assign \g251251/_0_  = _w23947_ ;
	assign \g251252/_0_  = _w23959_ ;
	assign \g251286/_0_  = _w23972_ ;
	assign \g251287/_0_  = _w23989_ ;
	assign \g251288/_0_  = _w24006_ ;
	assign \g251289/_0_  = _w24025_ ;
	assign \g251290/_0_  = _w24039_ ;
	assign \g251291/_0_  = _w24049_ ;
	assign \g251318/_0_  = _w24061_ ;
	assign \g252698/_3_  = _w24092_ ;
	assign \g252942/_0_  = _w24121_ ;
	assign \g252943/_0_  = _w24149_ ;
	assign \g253118/_0_  = _w24165_ ;
	assign \g253119/_0_  = _w24181_ ;
	assign \g253120/_0_  = _w24221_ ;
	assign \g253121/_0_  = _w24238_ ;
	assign \g253122/_3_  = _w24266_ ;
	assign \g253123/_0_  = _w24283_ ;
	assign \g253236/_0_  = _w24301_ ;
	assign \g253237/_3_  = _w24328_ ;
	assign \g253238/_3_  = _w24352_ ;
	assign \g253239/_0_  = _w24384_ ;
	assign \g253240/_0_  = _w24404_ ;
	assign \g253241/_0_  = _w24424_ ;
	assign \g253242/_0_  = _w24438_ ;
	assign \g253243/_0_  = _w24457_ ;
	assign \g253244/_0_  = _w24471_ ;
	assign \g253245/_0_  = _w24486_ ;
	assign \g253246/_0_  = _w24500_ ;
	assign \g253247/_0_  = _w24512_ ;
	assign \g253248/_0_  = _w24526_ ;
	assign \g253306/_0_  = _w24543_ ;
	assign \g253307/_3_  = _w24556_ ;
	assign \g253308/_0_  = _w24568_ ;
	assign \g253309/_0_  = _w24601_ ;
	assign \g253310/_0_  = _w24618_ ;
	assign \g253311/_0_  = _w24632_ ;
	assign \g253356/_0_  = _w24649_ ;
	assign \g253357/_0_  = _w24663_ ;
	assign \g253358/_0_  = _w24681_ ;
	assign \g253359/_0_  = _w24696_ ;
	assign \g253436/_3_  = _w24724_ ;
	assign \g253437/_0_  = _w24759_ ;
	assign \g253438/_0_  = _w24774_ ;
	assign \g253469/_3_  = _w24790_ ;
	assign \g253470/_3_  = _w24818_ ;
	assign \g253471/_3_  = _w24830_ ;
	assign \g253521/_0_  = _w24853_ ;
	assign \g253522/_0_  = _w24886_ ;
	assign \g253523/_0_  = _w24907_ ;
	assign \g253524/_3_  = _w24921_ ;
	assign \g256730/_3_  = _w24949_ ;
	assign \g256731/_3_  = _w24977_ ;
	assign \g256927/_0_  = _w25008_ ;
	assign \g256928/_0_  = _w25040_ ;
	assign \g256929/_3_  = _w25074_ ;
	assign \g257049/_0_  = _w25089_ ;
	assign \g257050/_0_  = _w25105_ ;
	assign \g257051/_3_  = _w25121_ ;
	assign \g257052/_0_  = _w25137_ ;
	assign \g257053/_0_  = _w25148_ ;
	assign \g257054/_0_  = _w25172_ ;
	assign \g257055/_3_  = _w25189_ ;
	assign \g257056/_0_  = _w25212_ ;
	assign \g257057/_0_  = _w25227_ ;
	assign \g257058/_3_  = _w25245_ ;
	assign \g257059/_0_  = _w25266_ ;
	assign \g257060/_0_  = _w25282_ ;
	assign \g257082/_0_  = _w25300_ ;
	assign \g257125/_3_  = _w25319_ ;
	assign \g257126/_0_  = _w25334_ ;
	assign \g257127/_0_  = _w25351_ ;
	assign \g257128/_3_  = _w25368_ ;
	assign \g257129/_3_  = _w25388_ ;
	assign \g257130/_0_  = _w25416_ ;
	assign \g257131/_0_  = _w25428_ ;
	assign \g257132/_0_  = _w25443_ ;
	assign \g257163/_0_  = _w25463_ ;
	assign \g257164/_0_  = _w25476_ ;
	assign \g257165/_0_  = _w25489_ ;
	assign \g257166/_0_  = _w25499_ ;
	assign \g257167/_0_  = _w25512_ ;
	assign \g257194/_0_  = _w25525_ ;
	assign \g258552/_0_  = _w25557_ ;
	assign \g258850/_0_  = _w25585_ ;
	assign \g258851/_3_  = _w25613_ ;
	assign \g258993/_0_  = _w25629_ ;
	assign \g258994/_0_  = _w25666_ ;
	assign \g258995/_0_  = _w25681_ ;
	assign \g258996/_0_  = _w25712_ ;
	assign \g259026/_3_  = _w25740_ ;
	assign \g259027/_0_  = _w25753_ ;
	assign \g259105/_0_  = _w25771_ ;
	assign \g259106/_0_  = _w25789_ ;
	assign \g259107/_3_  = _w25816_ ;
	assign \g259108/_0_  = _w25848_ ;
	assign \g259109/_3_  = _w25864_ ;
	assign \g259110/_0_  = _w25881_ ;
	assign \g259111/_0_  = _w25897_ ;
	assign \g259112/_0_  = _w25914_ ;
	assign \g259113/_0_  = _w25928_ ;
	assign \g259114/_0_  = _w25943_ ;
	assign \g259115/_0_  = _w25957_ ;
	assign \g259116/_0_  = _w25970_ ;
	assign \g259117/_0_  = _w25984_ ;
	assign \g259163/_3_  = _w26001_ ;
	assign \g259164/_3_  = _w26016_ ;
	assign \g259165/_0_  = _w26031_ ;
	assign \g259166/_0_  = _w26061_ ;
	assign \g259167/_0_  = _w26074_ ;
	assign \g259168/_0_  = _w26088_ ;
	assign \g259197/_0_  = _w26104_ ;
	assign \g259198/_0_  = _w26121_ ;
	assign \g259199/_0_  = _w26136_ ;
	assign \g259200/_0_  = _w26150_ ;
	assign \g260774/_0_  = _w26181_ ;
	assign \g260792/_3_  = _w26211_ ;
	assign \g260991/_0_  = _w26244_ ;
	assign \g261013/_0_  = _w26275_ ;
	assign \g261070/_0_  = _w26312_ ;
	assign \g261125/_0_  = _w26332_ ;
	assign \g261126/_0_  = _w26350_ ;
	assign \g261128/_0_  = _w26376_ ;
	assign \g261129/_0_  = _w26398_ ;
	assign \g261130/_0_  = _w26412_ ;
	assign \g261131/_0_  = _w26426_ ;
	assign \g261132/_0_  = _w26450_ ;
	assign \g261133/_0_  = _w26465_ ;
	assign \g261134/_3_  = _w26488_ ;
	assign \g261135/_0_  = _w26509_ ;
	assign \g261136/_0_  = _w26526_ ;
	assign \g261158/_3_  = _w26540_ ;
	assign \g261206/_0_  = _w26556_ ;
	assign \g261207/_0_  = _w26571_ ;
	assign \g261208/_0_  = _w26584_ ;
	assign \g261209/_0_  = _w26602_ ;
	assign \g261210/_3_  = _w26621_ ;
	assign \g261211/_0_  = _w26647_ ;
	assign \g261212/_3_  = _w26665_ ;
	assign \g261213/_0_  = _w26677_ ;
	assign \g261248/_0_  = _w26695_ ;
	assign \g261249/_0_  = _w26711_ ;
	assign \g261250/_0_  = _w26724_ ;
	assign \g261251/_0_  = _w26738_ ;
	assign \g261252/_0_  = _w26753_ ;
	assign \g261279/_0_  = _w26765_ ;
	assign \g262658/_3_  = _w26797_ ;
	assign \g262949/_0_  = _w26829_ ;
	assign \g263008/_3_  = _w26861_ ;
	assign \g263092/_0_  = _w26876_ ;
	assign \g263093/_0_  = _w26910_ ;
	assign \g263099/_0_  = _w26925_ ;
	assign \g263100/_0_  = _w26955_ ;
	assign \g263101/_0_  = _w26974_ ;
	assign \g263159/_3_  = _w27006_ ;
	assign \g263204/_3_  = _w27024_ ;
	assign \g263205/_0_  = _w27042_ ;
	assign \g263206/_0_  = _w27066_ ;
	assign \g263208/_0_  = _w27080_ ;
	assign \g263209/_0_  = _w27100_ ;
	assign \g263210/_0_  = _w27114_ ;
	assign \g263211/_0_  = _w27134_ ;
	assign \g263212/_0_  = _w27151_ ;
	assign \g263213/_0_  = _w27167_ ;
	assign \g263214/_0_  = _w27181_ ;
	assign \g263215/_3_  = _w27200_ ;
	assign \g263216/_0_  = _w27221_ ;
	assign \g263260/_0_  = _w27237_ ;
	assign \g263261/_0_  = _w27255_ ;
	assign \g263262/_3_  = _w27270_ ;
	assign \g263263/_0_  = _w27299_ ;
	assign \g263264/_0_  = _w27314_ ;
	assign \g263265/_0_  = _w27328_ ;
	assign \g263297/_0_  = _w27342_ ;
	assign \g263298/_0_  = _w27353_ ;
	assign \g263299/_0_  = _w27371_ ;
	assign \g263300/_0_  = _w27387_ ;
	assign \g264930/_0_  = _w27414_ ;
	assign \g264946/_3_  = _w27442_ ;
	assign \g265143/_0_  = _w27475_ ;
	assign \g265144/_0_  = _w27513_ ;
	assign \g265152/_0_  = _w27545_ ;
	assign \g265222/_0_  = _w27564_ ;
	assign \g265223/_0_  = _w27592_ ;
	assign \g265224/_0_  = _w27608_ ;
	assign \g265225/_0_  = _w27626_ ;
	assign \g265226/_0_  = _w27662_ ;
	assign \g265227/_3_  = _w27679_ ;
	assign \g265228/_0_  = _w27696_ ;
	assign \g265229/_0_  = _w27708_ ;
	assign \g265230/_0_  = _w27728_ ;
	assign \g265231/_0_  = _w27744_ ;
	assign \g265232/_0_  = _w27759_ ;
	assign \g265233/_3_  = _w27779_ ;
	assign \g265234/_0_  = _w27793_ ;
	assign \g265306/_0_  = _w27810_ ;
	assign \g265307/_0_  = _w27828_ ;
	assign \g265308/_3_  = _w27843_ ;
	assign \g265309/_3_  = _w27858_ ;
	assign \g265310/_0_  = _w27887_ ;
	assign \g265311/_0_  = _w27900_ ;
	assign \g265312/_0_  = _w27914_ ;
	assign \g265313/_0_  = _w27926_ ;
	assign \g265348/_0_  = _w27939_ ;
	assign \g265349/_0_  = _w27955_ ;
	assign \g265350/_0_  = _w27971_ ;
	assign \g265351/_0_  = _w27985_ ;
	assign \g265379/_0_  = _w27997_ ;
	assign \g266965/_3_  = _w28029_ ;
	assign \g267049/_3_  = _w28061_ ;
	assign \g267050/_0_  = _w28091_ ;
	assign \g267215/_0_  = _w28106_ ;
	assign \g267216/_0_  = _w28142_ ;
	assign \g267263/_0_  = _w28157_ ;
	assign \g267264/_3_  = _w28185_ ;
	assign \g267265/_0_  = _w28203_ ;
	assign \g267266/_0_  = _w28233_ ;
	assign \g267314/_3_  = _w28253_ ;
	assign \g267315/_0_  = _w28289_ ;
	assign \g267316/_0_  = _w28307_ ;
	assign \g267317/_0_  = _w28321_ ;
	assign \g267318/_0_  = _w28336_ ;
	assign \g267319/_0_  = _w28360_ ;
	assign \g267320/_3_  = _w28374_ ;
	assign \g267321/_0_  = _w28387_ ;
	assign \g267322/_0_  = _w28401_ ;
	assign \g267324/_0_  = _w28415_ ;
	assign \g267325/_0_  = _w28429_ ;
	assign \g267326/_0_  = _w28444_ ;
	assign \g267372/_0_  = _w28458_ ;
	assign \g267373/_3_  = _w28477_ ;
	assign \g267374/_0_  = _w28491_ ;
	assign \g267375/_0_  = _w28520_ ;
	assign \g267376/_0_  = _w28534_ ;
	assign \g267377/_0_  = _w28550_ ;
	assign \g267409/_0_  = _w28561_ ;
	assign \g267410/_0_  = _w28579_ ;
	assign \g267411/_0_  = _w28595_ ;
	assign \g267412/_0_  = _w28607_ ;
	assign \g269004/_0_  = _w28634_ ;
	assign \g269099/_3_  = _w28665_ ;
	assign \g269202/_0_  = _w28704_ ;
	assign \g269226/_0_  = _w28731_ ;
	assign \g269333/_3_  = _w28751_ ;
	assign \g269334/_0_  = _w28783_ ;
	assign \g269335/_0_  = _w28800_ ;
	assign \g269355/_0_  = _w28823_ ;
	assign \g269356/_0_  = _w28839_ ;
	assign \g269357/_3_  = _w28871_ ;
	assign \g269358/_0_  = _w28891_ ;
	assign \g269359/_0_  = _w28906_ ;
	assign \g269360/_0_  = _w28942_ ;
	assign \g269361/_0_  = _w28962_ ;
	assign \g269362/_0_  = _w28977_ ;
	assign \g269363/_0_  = _w28995_ ;
	assign \g269364/_0_  = _w29011_ ;
	assign \g269414/_0_  = _w29024_ ;
	assign \g269415/_0_  = _w29038_ ;
	assign \g269416/_0_  = _w29053_ ;
	assign \g269417/_0_  = _w29067_ ;
	assign \g269418/_3_  = _w29085_ ;
	assign \g269419/_0_  = _w29103_ ;
	assign \g269420/_3_  = _w29122_ ;
	assign \g269421/_0_  = _w29147_ ;
	assign \g269456/_0_  = _w29170_ ;
	assign \g269457/_0_  = _w29182_ ;
	assign \g269458/_0_  = _w29202_ ;
	assign \g269459/_0_  = _w29216_ ;
	assign \g269460/_0_  = _w29227_ ;
	assign \g269487/_0_  = _w29241_ ;
	assign \g271006/_3_  = _w29270_ ;
	assign \g271186/_3_  = _w29300_ ;
	assign \g271187/_0_  = _w29330_ ;
	assign \g271299/_0_  = _w29368_ ;
	assign \g271300/_0_  = _w29395_ ;
	assign \g271301/_3_  = _w29427_ ;
	assign \g271302/_0_  = _w29442_ ;
	assign \g271303/_0_  = _w29459_ ;
	assign \g271352/_0_  = _w29480_ ;
	assign \g271410/_0_  = _w29496_ ;
	assign \g271411/_0_  = _w29509_ ;
	assign \g271412/_0_  = _w29535_ ;
	assign \g271413/_0_  = _w29557_ ;
	assign \g271414/_0_  = _w29576_ ;
	assign \g271415/_0_  = _w29596_ ;
	assign \g271416/_0_  = _w29613_ ;
	assign \g271417/_3_  = _w29628_ ;
	assign \g271418/_3_  = _w29647_ ;
	assign \g271419/_0_  = _w29663_ ;
	assign \g271420/_0_  = _w29681_ ;
	assign \g271421/_0_  = _w29695_ ;
	assign \g271422/_0_  = _w29711_ ;
	assign \g271468/_3_  = _w29727_ ;
	assign \g271469/_0_  = _w29744_ ;
	assign \g271470/_0_  = _w29773_ ;
	assign \g271471/_0_  = _w29789_ ;
	assign \g271472/_0_  = _w29802_ ;
	assign \g271473/_0_  = _w29813_ ;
	assign \g271505/_0_  = _w29827_ ;
	assign \g271506/_0_  = _w29839_ ;
	assign \g271507/_0_  = _w29861_ ;
	assign \g271508/_0_  = _w29876_ ;
	assign \g273135/_0_  = _w29906_ ;
	assign \g273136/_3_  = _w29937_ ;
	assign \g273362/_0_  = _w29970_ ;
	assign \g273373/_0_  = _w30005_ ;
	assign \g273374/_0_  = _w30037_ ;
	assign \g273431/_0_  = _w30055_ ;
	assign \g273432/_0_  = _w30070_ ;
	assign \g273433/_3_  = _w30100_ ;
	assign \g273434/_0_  = _w30118_ ;
	assign \g273435/_0_  = _w30130_ ;
	assign \g273436/_0_  = _w30161_ ;
	assign \g273437/_3_  = _w30178_ ;
	assign \g273438/_0_  = _w30196_ ;
	assign \g273439/_0_  = _w30216_ ;
	assign \g273441/_0_  = _w30235_ ;
	assign \g273442/_0_  = _w30252_ ;
	assign \g273443/_0_  = _w30268_ ;
	assign \g273515/_3_  = _w30287_ ;
	assign \g273516/_0_  = _w30305_ ;
	assign \g273517/_0_  = _w30325_ ;
	assign \g273518/_3_  = _w30345_ ;
	assign \g273519/_0_  = _w30358_ ;
	assign \g273520/_0_  = _w30371_ ;
	assign \g273521/_0_  = _w30385_ ;
	assign \g273522/_0_  = _w30410_ ;
	assign \g273557/_0_  = _w30429_ ;
	assign \g273558/_0_  = _w30445_ ;
	assign \g273559/_0_  = _w30460_ ;
	assign \g273560/_0_  = _w30474_ ;
	assign \g273561/_0_  = _w30485_ ;
	assign \g273588/_0_  = _w30497_ ;
	assign \g274960/_3_  = _w30528_ ;
	assign \g275266/_3_  = _w30563_ ;
	assign \g275327/_0_  = _w30593_ ;
	assign \g275396/_0_  = _w30612_ ;
	assign \g275397/_3_  = _w30642_ ;
	assign \g275398/_0_  = _w30659_ ;
	assign \g275455/_0_  = _w30689_ ;
	assign \g275456/_0_  = _w30704_ ;
	assign \g275463/_0_  = _w30740_ ;
	assign \g275510/_3_  = _w30761_ ;
	assign \g275511/_0_  = _w30781_ ;
	assign \g275512/_0_  = _w30792_ ;
	assign \g275513/_0_  = _w30809_ ;
	assign \g275514/_3_  = _w30828_ ;
	assign \g275515/_0_  = _w30844_ ;
	assign \g275516/_0_  = _w30871_ ;
	assign \g275517/_0_  = _w30887_ ;
	assign \g275518/_0_  = _w30909_ ;
	assign \g275519/_0_  = _w30924_ ;
	assign \g275520/_0_  = _w30942_ ;
	assign \g275521/_0_  = _w30958_ ;
	assign \g275522/_0_  = _w30974_ ;
	assign \g275568/_0_  = _w30988_ ;
	assign \g275569/_0_  = _w31002_ ;
	assign \g275570/_0_  = _w31017_ ;
	assign \g275571/_0_  = _w31043_ ;
	assign \g275572/_3_  = _w31061_ ;
	assign \g275573/_0_  = _w31074_ ;
	assign \g275605/_0_  = _w31093_ ;
	assign \g275606/_0_  = _w31105_ ;
	assign \g275607/_0_  = _w31118_ ;
	assign \g275608/_0_  = _w31135_ ;
	assign \g277189/_0_  = _w31163_ ;
	assign \g277294/_3_  = _w31200_ ;
	assign \g277367/_0_  = _w31232_ ;
	assign \g277456/_0_  = _w31262_ ;
	assign \g277457/_0_  = _w31294_ ;
	assign \g277512/_0_  = _w31316_ ;
	assign \g277513/_0_  = _w31348_ ;
	assign \g277514/_3_  = _w31380_ ;
	assign \g277515/_0_  = _w31396_ ;
	assign \g277516/_0_  = _w31415_ ;
	assign \g277517/_3_  = _w31429_ ;
	assign \g277518/_0_  = _w31446_ ;
	assign \g277519/_0_  = _w31466_ ;
	assign \g277520/_0_  = _w31480_ ;
	assign \g277521/_0_  = _w31494_ ;
	assign \g277594/_0_  = _w31511_ ;
	assign \g277595/_0_  = _w31527_ ;
	assign \g277596/_3_  = _w31544_ ;
	assign \g277597/_0_  = _w31556_ ;
	assign \g277598/_0_  = _w31574_ ;
	assign \g277599/_0_  = _w31600_ ;
	assign \g277600/_0_  = _w31615_ ;
	assign \g277601/_3_  = _w31634_ ;
	assign \g277635/_0_  = _w31648_ ;
	assign \g277636/_0_  = _w31670_ ;
	assign \g277637/_0_  = _w31689_ ;
	assign \g277638/_0_  = _w31701_ ;
	assign \g277639/_0_  = _w31714_ ;
	assign \g277666/_0_  = _w31728_ ;
	assign \g279090/_3_  = _w31758_ ;
	assign \g279330/_0_  = _w31792_ ;
	assign \g279331/_0_  = _w31820_ ;
	assign \g279493/_3_  = _w31849_ ;
	assign \g279494/_0_  = _w31868_ ;
	assign \g279495/_0_  = _w31883_ ;
	assign \g279502/_0_  = _w31899_ ;
	assign \g279503/_0_  = _w31932_ ;
	assign \g279504/_0_  = _w31968_ ;
	assign \g279590/_0_  = _w31985_ ;
	assign \g279591/_0_  = _w32005_ ;
	assign \g279592/_0_  = _w32020_ ;
	assign \g279593/_0_  = _w32050_ ;
	assign \g279594/_3_  = _w32069_ ;
	assign \g279595/_3_  = _w32084_ ;
	assign \g279596/_0_  = _w32104_ ;
	assign \g279597/_0_  = _w32121_ ;
	assign \g279598/_0_  = _w32135_ ;
	assign \g279599/_0_  = _w32154_ ;
	assign \g279600/_0_  = _w32168_ ;
	assign \g279601/_0_  = _w32180_ ;
	assign \g279602/_0_  = _w32198_ ;
	assign \g279649/_0_  = _w32228_ ;
	assign \g279650/_0_  = _w32243_ ;
	assign \g279651/_0_  = _w32256_ ;
	assign \g279652/_0_  = _w32268_ ;
	assign \g279653/_0_  = _w32287_ ;
	assign \g279654/_3_  = _w32300_ ;
	assign \g279686/_0_  = _w32319_ ;
	assign \g279687/_0_  = _w32333_ ;
	assign \g279688/_0_  = _w32350_ ;
	assign \g279689/_0_  = _w32363_ ;
	assign \g281329/_0_  = _w32390_ ;
	assign \g281394/_0_  = _w32432_ ;
	assign \g281483/_0_  = _w32456_ ;
	assign \g281498/_0_  = _w32492_ ;
	assign \g281532/_0_  = _w32528_ ;
	assign \g281616/_0_  = _w32560_ ;
	assign \g281617/_0_  = _w32581_ ;
	assign \g281618/_0_  = _w32600_ ;
	assign \g281619/_0_  = _w32619_ ;
	assign \g281620/_0_  = _w32633_ ;
	assign \g281621/_0_  = _w32651_ ;
	assign \g281622/_0_  = _w32678_ ;
	assign \g281623/_3_  = _w32696_ ;
	assign \g281624/_0_  = _w32713_ ;
	assign \g281642/_0_  = _w32735_ ;
	assign \g281643/_0_  = _w32749_ ;
	assign \g281644/_3_  = _w32773_ ;
	assign \g281645/_0_  = _w32789_ ;
	assign \g281696/_0_  = _w32801_ ;
	assign \g281697/_3_  = _w32819_ ;
	assign \g281698/_0_  = _w32830_ ;
	assign \g281699/_0_  = _w32854_ ;
	assign \g281700/_0_  = _w32869_ ;
	assign \g281701/_0_  = _w32886_ ;
	assign \g281702/_3_  = _w32902_ ;
	assign \g281703/_0_  = _w32915_ ;
	assign \g281799/_0_  = _w32936_ ;
	assign \g281800/_0_  = _w32953_ ;
	assign \g281801/_0_  = _w32969_ ;
	assign \g281802/_0_  = _w32982_ ;
	assign \g281803/_0_  = _w32994_ ;
	assign \g281965/_0_  = _w33008_ ;
	assign \g287377/_0_  = _w33046_ ;
	assign \g287867/_0_  = _w33082_ ;
	assign \g287899/_0_  = _w33110_ ;
	assign \g288304/_0_  = _w33123_ ;
	assign \g288334/_0_  = _w33140_ ;
	assign \g288350/_0_  = _w33175_ ;
	assign \g288351/_0_  = _w33189_ ;
	assign \g288352/_3_  = _w33221_ ;
	assign \g288353/_0_  = _w33242_ ;
	assign \g288668/_0_  = _w33261_ ;
	assign \g288669/_0_  = _w33278_ ;
	assign \g288670/_0_  = _w33297_ ;
	assign \g288671/_0_  = _w33316_ ;
	assign \g288673/_0_  = _w33336_ ;
	assign \g288674/_3_  = _w33352_ ;
	assign \g288675/_0_  = _w33385_ ;
	assign \g288676/_0_  = _w33412_ ;
	assign \g288677/_0_  = _w33424_ ;
	assign \g288678/_0_  = _w33441_ ;
	assign \g288679/_0_  = _w33457_ ;
	assign \g288680/_3_  = _w33475_ ;
	assign \g288889/_0_  = _w33489_ ;
	assign \g288890/_0_  = _w33504_ ;
	assign \g288891/_0_  = _w33519_ ;
	assign \g288892/_0_  = _w33532_ ;
	assign \g288893/_3_  = _w33548_ ;
	assign \g288894/_0_  = _w33563_ ;
	assign \g288895/_0_  = _w33579_ ;
	assign \g288984/_0_  = _w33593_ ;
	assign \g288985/_0_  = _w33608_ ;
	assign \g288986/_0_  = _w33622_ ;
	assign \g294974/_0_  = _w33651_ ;
	assign \g295054/_0_  = _w33683_ ;
	assign \g295601/_0_  = _w33717_ ;
	assign \g295607/_0_  = _w33746_ ;
	assign \g296036/_0_  = _w33779_ ;
	assign \g296037/_0_  = _w33806_ ;
	assign \g296038/_0_  = _w33837_ ;
	assign \g296039/_0_  = _w33856_ ;
	assign \g296040/_0_  = _w33875_ ;
	assign \g296041/_0_  = _w33889_ ;
	assign \g296042/_0_  = _w33907_ ;
	assign \g296043/_3_  = _w33943_ ;
	assign \g296044/_0_  = _w33961_ ;
	assign \g296045/_0_  = _w33977_ ;
	assign \g296046/_0_  = _w33995_ ;
	assign \g296047/_0_  = _w34009_ ;
	assign \g296048/_0_  = _w34024_ ;
	assign \g296049/_3_  = _w34040_ ;
	assign \g296522/_3_  = _w34058_ ;
	assign \g296523/_3_  = _w34070_ ;
	assign \g296524/_0_  = _w34087_ ;
	assign \g296525/_0_  = _w34108_ ;
	assign \g296526/_0_  = _w34122_ ;
	assign \g296527/_0_  = _w34140_ ;
	assign \g296528/_3_  = _w34154_ ;
	assign \g296529/_0_  = _w34167_ ;
	assign \g296530/_0_  = _w34185_ ;
	assign \g296531/_0_  = _w34198_ ;
	assign \g297026/_0_  = _w34211_ ;
	assign \g297027/_0_  = _w34229_ ;
	assign \g305620/_3_  = _w34230_ ;
	assign \g305621/_3_  = _w34231_ ;
	assign \g305622/_3_  = _w34232_ ;
	assign \g305623/_3_  = _w34233_ ;
	assign \g305624/_3_  = _w34234_ ;
	assign \g305625/_3_  = _w34235_ ;
	assign \g305626/_3_  = _w34236_ ;
	assign \g305627/_3_  = _w34237_ ;
	assign \g305628/_3_  = _w34238_ ;
	assign \g305629/_3_  = _w34239_ ;
	assign \g305630/_3_  = _w34240_ ;
	assign \g305631/_3_  = _w34241_ ;
	assign \g305632/_3_  = _w34242_ ;
	assign \g305633/_3_  = _w34243_ ;
	assign \g305634/_3_  = _w34244_ ;
	assign \g305635/_3_  = _w34245_ ;
	assign \g305636/_3_  = _w34246_ ;
	assign \g305637/_3_  = _w34247_ ;
	assign \g305638/_3_  = _w34248_ ;
	assign \g305639/_3_  = _w34249_ ;
	assign \g305640/_3_  = _w34250_ ;
	assign \g305641/_3_  = _w34251_ ;
	assign \g305642/_3_  = _w34252_ ;
	assign \g305643/_3_  = _w34253_ ;
	assign \g305644/_3_  = _w34254_ ;
	assign \g305645/_3_  = _w34255_ ;
	assign \g305646/_3_  = _w34256_ ;
	assign \g305647/_3_  = _w34257_ ;
	assign \g305648/_3_  = _w34258_ ;
	assign \g305649/_3_  = _w34259_ ;
	assign \g305650/_3_  = _w34260_ ;
	assign \g305651/_3_  = _w34261_ ;
	assign \g305652/_3_  = _w34262_ ;
	assign \g305653/_3_  = _w34263_ ;
	assign \g305654/_3_  = _w34264_ ;
	assign \g305655/_3_  = _w34265_ ;
	assign \g305656/_3_  = _w34266_ ;
	assign \g305657/_3_  = _w34267_ ;
	assign \g305658/_3_  = _w34268_ ;
	assign \g305659/_3_  = _w34269_ ;
	assign \g305660/_3_  = _w34270_ ;
	assign \g305661/_3_  = _w34271_ ;
	assign \g305662/_3_  = _w34272_ ;
	assign \g305663/_3_  = _w34273_ ;
	assign \g305664/_3_  = _w34274_ ;
	assign \g305665/_3_  = _w34275_ ;
	assign \g305666/_3_  = _w34276_ ;
	assign \g305667/_3_  = _w34277_ ;
	assign \g305668/_3_  = _w34278_ ;
	assign \g305669/_3_  = _w34279_ ;
	assign \g305670/_3_  = _w34280_ ;
	assign \g305671/_3_  = _w34281_ ;
	assign \g305672/_3_  = _w34282_ ;
	assign \g305673/_3_  = _w34283_ ;
	assign \g305674/_3_  = _w34284_ ;
	assign \g305675/_3_  = _w34285_ ;
	assign \g305676/_3_  = _w34286_ ;
	assign \g305677/_3_  = _w34287_ ;
	assign \g305678/_3_  = _w34288_ ;
	assign \g305679/_3_  = _w34289_ ;
	assign \g305680/_3_  = _w34290_ ;
	assign \g305681/_3_  = _w34291_ ;
	assign \g305682/_3_  = _w34292_ ;
	assign \g305683/_3_  = _w34293_ ;
	assign \g305684/_3_  = _w34294_ ;
	assign \g305685/_3_  = _w34295_ ;
	assign \g305686/_3_  = _w34296_ ;
	assign \g305687/_3_  = _w34297_ ;
	assign \g305688/_3_  = _w34298_ ;
	assign \g305689/_3_  = _w34299_ ;
	assign \g305690/_3_  = _w34300_ ;
	assign \g305691/_3_  = _w34301_ ;
	assign \g305692/_3_  = _w34302_ ;
	assign \g305693/_3_  = _w34303_ ;
	assign \g305694/_3_  = _w34304_ ;
	assign \g305695/_3_  = _w34305_ ;
	assign \g305696/_3_  = _w34306_ ;
	assign \g305697/_3_  = _w34307_ ;
	assign \g305698/_3_  = _w34308_ ;
	assign \g305699/_3_  = _w34309_ ;
	assign \g305700/_3_  = _w34310_ ;
	assign \g305701/_3_  = _w34311_ ;
	assign \g305702/_3_  = _w34312_ ;
	assign \g305703/_3_  = _w34313_ ;
	assign \g305704/_3_  = _w34314_ ;
	assign \g305705/_3_  = _w34315_ ;
	assign \g305706/_3_  = _w34316_ ;
	assign \g305707/_3_  = _w34317_ ;
	assign \g305708/_3_  = _w34318_ ;
	assign \g305709/_3_  = _w34319_ ;
	assign \g305710/_3_  = _w34320_ ;
	assign \g305711/_3_  = _w34321_ ;
	assign \g305712/_3_  = _w34322_ ;
	assign \g305713/_3_  = _w34323_ ;
	assign \g305714/_3_  = _w34324_ ;
	assign \g305715/_3_  = _w34325_ ;
	assign \g305716/_3_  = _w34326_ ;
	assign \g305717/_3_  = _w34327_ ;
	assign \g305718/_3_  = _w34328_ ;
	assign \g305719/_3_  = _w34329_ ;
	assign \g305720/_3_  = _w34330_ ;
	assign \g305721/_3_  = _w34331_ ;
	assign \g305722/_3_  = _w34332_ ;
	assign \g305723/_3_  = _w34333_ ;
	assign \g305724/_3_  = _w34334_ ;
	assign \g305725/_3_  = _w34335_ ;
	assign \g305726/_3_  = _w34336_ ;
	assign \g305727/_3_  = _w34337_ ;
	assign \g305728/_3_  = _w34338_ ;
	assign \g305729/_3_  = _w34339_ ;
	assign \g305730/_3_  = _w34340_ ;
	assign \g305731/_3_  = _w34341_ ;
	assign \g321371/_0_  = _w34356_ ;
	assign \g321424/_0_  = _w34366_ ;
	assign \g321474/_3_  = _w34383_ ;
	assign \g321637/_3_  = _w34398_ ;
	assign \g321688/_0_  = _w34414_ ;
	assign \g321712/_0_  = _w34432_ ;
	assign \g321772/_3_  = _w34448_ ;
	assign \g321832/_0_  = _w34465_ ;
	assign \g321999/_0_  = _w34480_ ;
	assign \g322013/_3_  = _w34494_ ;
	assign \g322109/_0_  = _w34514_ ;
	assign \g322184/_0_  = _w34526_ ;
	assign \g322250/_0_  = _w34544_ ;
	assign \g322274/_0_  = _w34556_ ;
	assign \g322293/_3_  = _w34567_ ;
	assign \g322437/_0_  = _w34580_ ;
	assign \g322537/_3_  = _w34592_ ;
	assign \g322584/_0_  = _w34608_ ;
	assign \g322830/_0_  = _w34619_ ;
	assign \g322871/_0_  = _w34635_ ;
	assign \g322882/_0_  = _w34653_ ;
	assign \g322933/_0_  = _w34666_ ;
	assign \g323004/_0_  = _w34681_ ;
	assign \g323104/_0_  = _w34693_ ;
	assign \g323125/_0_  = _w34713_ ;
	assign \g323138/_3_  = _w34726_ ;
	assign \g323273/_0_  = _w34742_ ;
	assign \u0_desOut_reg[0]/_05_  = _w34762_ ;
	assign \u0_desOut_reg[12]/_05_  = _w34800_ ;
	assign \u0_desOut_reg[14]/_05_  = _w34824_ ;
	assign \u0_desOut_reg[18]/_05_  = _w34853_ ;
	assign \u0_desOut_reg[20]/_05_  = _w34874_ ;
	assign \u0_desOut_reg[24]/_05_  = _w34893_ ;
	assign \u0_desOut_reg[26]/_05_  = _w34913_ ;
	assign \u0_desOut_reg[28]/_05_  = _w34936_ ;
	assign \u0_desOut_reg[2]/_05_  = _w34948_ ;
	assign \u0_desOut_reg[30]/_05_  = _w34965_ ;
	assign \u0_desOut_reg[32]/_05_  = _w34979_ ;
	assign \u0_desOut_reg[34]/_05_  = _w35000_ ;
	assign \u0_desOut_reg[36]/_05_  = _w35016_ ;
	assign \u0_desOut_reg[42]/_05_  = _w35037_ ;
	assign \u0_desOut_reg[44]/_05_  = _w35054_ ;
	assign \u0_desOut_reg[46]/_05_  = _w35066_ ;
	assign \u0_desOut_reg[48]/_05_  = _w35085_ ;
	assign \u0_desOut_reg[54]/_05_  = _w35103_ ;
	assign \u0_desOut_reg[56]/_05_  = _w35117_ ;
	assign \u0_desOut_reg[62]/_05_  = _w35129_ ;
	assign \u0_desOut_reg[6]/_05_  = _w35147_ ;
	assign \u0_desOut_reg[8]/_05_  = _w35166_ ;
	assign \u1_desOut_reg[0]/_05_  = _w35194_ ;
	assign \u1_desOut_reg[12]/_05_  = _w35227_ ;
	assign \u1_desOut_reg[14]/_05_  = _w35250_ ;
	assign \u1_desOut_reg[16]/_05_  = _w35270_ ;
	assign \u1_desOut_reg[18]/_05_  = _w35301_ ;
	assign \u1_desOut_reg[20]/_05_  = _w35321_ ;
	assign \u1_desOut_reg[22]/_05_  = _w35342_ ;
	assign \u1_desOut_reg[24]/_05_  = _w35360_ ;
	assign \u1_desOut_reg[26]/_05_  = _w35374_ ;
	assign \u1_desOut_reg[28]/_05_  = _w35399_ ;
	assign \u1_desOut_reg[2]/_05_  = _w35416_ ;
	assign \u1_desOut_reg[30]/_05_  = _w35430_ ;
	assign \u1_desOut_reg[32]/_05_  = _w35444_ ;
	assign \u1_desOut_reg[34]/_05_  = _w35462_ ;
	assign \u1_desOut_reg[36]/_05_  = _w35476_ ;
	assign \u1_desOut_reg[38]/_05_  = _w35493_ ;
	assign \u1_desOut_reg[42]/_05_  = _w35519_ ;
	assign \u1_desOut_reg[44]/_05_  = _w35543_ ;
	assign \u1_desOut_reg[46]/_05_  = _w35560_ ;
	assign \u1_desOut_reg[48]/_05_  = _w35579_ ;
	assign \u1_desOut_reg[4]/_05_  = _w35590_ ;
	assign \u1_desOut_reg[54]/_05_  = _w35604_ ;
	assign \u1_desOut_reg[56]/_05_  = _w35624_ ;
	assign \u1_desOut_reg[58]/_05_  = _w35642_ ;
	assign \u1_desOut_reg[60]/_05_  = _w35657_ ;
	assign \u1_desOut_reg[62]/_05_  = _w35668_ ;
	assign \u1_desOut_reg[6]/_05_  = _w35689_ ;
	assign \u1_desOut_reg[8]/_05_  = _w35706_ ;
	assign \u2_desOut_reg[0]/_05_  = _w35732_ ;
	assign \u2_desOut_reg[10]/_05_  = _w35756_ ;
	assign \u2_desOut_reg[12]/_05_  = _w35790_ ;
	assign \u2_desOut_reg[14]/_05_  = _w35815_ ;
	assign \u2_desOut_reg[16]/_05_  = _w35847_ ;
	assign \u2_desOut_reg[18]/_05_  = _w35877_ ;
	assign \u2_desOut_reg[20]/_05_  = _w35898_ ;
	assign \u2_desOut_reg[22]/_05_  = _w35917_ ;
	assign \u2_desOut_reg[24]/_05_  = _w35934_ ;
	assign \u2_desOut_reg[26]/_05_  = _w35953_ ;
	assign \u2_desOut_reg[28]/_05_  = _w35978_ ;
	assign \u2_desOut_reg[2]/_05_  = _w36003_ ;
	assign \u2_desOut_reg[30]/_05_  = _w36021_ ;
	assign \u2_desOut_reg[32]/_05_  = _w36033_ ;
	assign \u2_desOut_reg[34]/_05_  = _w36056_ ;
	assign \u2_desOut_reg[36]/_05_  = _w36072_ ;
	assign \u2_desOut_reg[38]/_05_  = _w36088_ ;
	assign \u2_desOut_reg[40]/_05_  = _w36120_ ;
	assign \u2_desOut_reg[42]/_05_  = _w36137_ ;
	assign \u2_desOut_reg[44]/_05_  = _w36156_ ;
	assign \u2_desOut_reg[46]/_05_  = _w36176_ ;
	assign \u2_desOut_reg[48]/_05_  = _w36201_ ;
	assign \u2_desOut_reg[4]/_05_  = _w36215_ ;
	assign \u2_desOut_reg[50]/_05_  = _w36235_ ;
	assign \u2_desOut_reg[52]/_05_  = _w36249_ ;
	assign \u2_desOut_reg[54]/_05_  = _w36264_ ;
	assign \u2_desOut_reg[56]/_05_  = _w36277_ ;
	assign \u2_desOut_reg[58]/_05_  = _w36291_ ;
	assign \u2_desOut_reg[60]/_05_  = _w36302_ ;
	assign \u2_desOut_reg[62]/_05_  = _w36313_ ;
	assign \u2_desOut_reg[6]/_05_  = _w36329_ ;
	assign \u2_desOut_reg[8]/_05_  = _w36346_ ;
endmodule;