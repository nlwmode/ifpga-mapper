module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	output q_pad ;
	output r_pad ;
	output s_pad ;
	output t_pad ;
	output u_pad ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		e_pad,
		f_pad,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		a_pad,
		_w17_,
		_w18_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		c_pad,
		d_pad,
		_w19_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		j_pad,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		j_pad,
		_w19_,
		_w21_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		e_pad,
		f_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		_w20_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w21_,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w18_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		b_pad,
		_w17_,
		_w26_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		l_pad,
		_w20_,
		_w27_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		l_pad,
		_w20_,
		_w28_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		_w22_,
		_w27_,
		_w29_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w28_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w26_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		g_pad,
		_w17_,
		_w32_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		m_pad,
		_w27_,
		_w33_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		l_pad,
		m_pad,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w20_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		_w22_,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w33_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w32_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		h_pad,
		_w17_,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		n_pad,
		_w35_,
		_w40_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		n_pad,
		_w35_,
		_w41_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		_w22_,
		_w40_,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w41_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w39_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		d_pad,
		i_pad,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		k_pad,
		o_pad,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		p_pad,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w45_,
		_w47_,
		_w48_
	);
	assign q_pad = _w25_ ;
	assign r_pad = _w31_ ;
	assign s_pad = _w38_ ;
	assign t_pad = _w44_ ;
	assign u_pad = _w48_ ;
endmodule;