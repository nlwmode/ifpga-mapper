module top (\a0_pad , a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, \h0_pad , h_pad, \i0_pad , i_pad, \j0_pad , j_pad, \k0_pad , k_pad, \l0_pad , l_pad, \m0_pad , m_pad, \n0_pad , n_pad, \o0_pad , o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \a1_pad , \b1_pad , \c1_pad , \d1_pad , \e1_pad , \f1_pad , \g1_pad , \h1_pad , \i1_pad , \j1_pad , \j4 , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , \u277_syn_3 , \v0_pad , \w0_pad , \y0_pad , \z0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \a1_pad  ;
	output \b1_pad  ;
	output \c1_pad  ;
	output \d1_pad  ;
	output \e1_pad  ;
	output \f1_pad  ;
	output \g1_pad  ;
	output \h1_pad  ;
	output \i1_pad  ;
	output \j1_pad  ;
	output \j4  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output \u277_syn_3  ;
	output \v0_pad  ;
	output \w0_pad  ;
	output \y0_pad  ;
	output \z0_pad  ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\c0_pad ,
		\j0_pad ,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\b0_pad ,
		i_pad,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\b0_pad ,
		e_pad,
		_w45_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\d0_pad ,
		i_pad,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\n0_pad ,
		\o0_pad ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\e0_pad ,
		j_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		_w46_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\k0_pad ,
		_w42_,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\b0_pad ,
		e_pad,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w53_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		e_pad,
		k_pad,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		_w48_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\c0_pad ,
		\j0_pad ,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\l0_pad ,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\b0_pad ,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w58_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		s_pad,
		t_pad,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		u_pad,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w61_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\e0_pad ,
		\g0_pad ,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\j0_pad ,
		\k0_pad ,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\c0_pad ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\b0_pad ,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		_w66_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		e_pad,
		n_pad,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w48_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w70_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w65_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\a0_pad ,
		\b0_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\i0_pad ,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		m_pad,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		b_pad,
		w_pad,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		x_pad,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		x_pad,
		y_pad,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w78_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\c0_pad ,
		i_pad,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\b0_pad ,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h2)
	) name42 (
		\j0_pad ,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		_w51_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\b0_pad ,
		\c0_pad ,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\l0_pad ,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		p_pad,
		_w62_,
		_w88_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		q_pad,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\b0_pad ,
		_w53_,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		_w66_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		e_pad,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		c_pad,
		_w47_,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		e_pad,
		_w44_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		_w48_,
		_w93_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		\b0_pad ,
		\l0_pad ,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		\j0_pad ,
		_w86_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w97_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		v_pad,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		v_pad,
		_w99_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		p_pad,
		r_pad,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\f0_pad ,
		\h0_pad ,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w102_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		o_pad,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		o_pad,
		z_pad,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		a_pad,
		z_pad,
		_w107_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\m0_pad ,
		_w106_,
		_w108_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		_w107_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		d_pad,
		_w105_,
		_w110_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w109_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		l_pad,
		_w76_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\b0_pad ,
		g_pad,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\l0_pad ,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		h_pad,
		_w48_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w55_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		e_pad,
		f_pad,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w48_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		_w91_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w114_,
		_w116_,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		_w119_,
		_w120_,
		_w121_
	);
	assign \a1_pad  = _w52_ ;
	assign \b1_pad  = _w62_ ;
	assign \c1_pad  = _w74_ ;
	assign \d1_pad  = _w74_ ;
	assign \e1_pad  = _w77_ ;
	assign \f1_pad  = _w79_ ;
	assign \g1_pad  = _w81_ ;
	assign \h1_pad  = _w52_ ;
	assign \i1_pad  = _w52_ ;
	assign \j1_pad  = _w85_ ;
	assign \j4  = _w87_ ;
	assign \p0_pad  = _w89_ ;
	assign \q0_pad  = _w92_ ;
	assign \r0_pad  = _w96_ ;
	assign \s0_pad  = _w100_ ;
	assign \t0_pad  = _w101_ ;
	assign \u277_syn_3  = _w48_ ;
	assign \v0_pad  = _w87_ ;
	assign \w0_pad  = _w111_ ;
	assign \y0_pad  = _w112_ ;
	assign \z0_pad  = _w121_ ;
endmodule;