module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  output q_pad ;
  output r_pad ;
  output s_pad ;
  output t_pad ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 ;
  assign n21 = c_pad & d_pad ;
  assign n22 = e_pad & j_pad ;
  assign n23 = n21 & n22 ;
  assign n17 = h_pad & i_pad ;
  assign n20 = a_pad & b_pad ;
  assign n24 = n17 & n20 ;
  assign n18 = k_pad & l_pad ;
  assign n19 = f_pad & g_pad ;
  assign n25 = n18 & n19 ;
  assign n26 = n24 & n25 ;
  assign n27 = n23 & n26 ;
  assign n28 = ~i_pad & ~j_pad ;
  assign n29 = ~n17 & ~n28 ;
  assign n35 = ~j_pad & k_pad ;
  assign n41 = ~n29 & ~n35 ;
  assign n30 = ~l_pad & ~m_pad ;
  assign n31 = ~n18 & ~n30 ;
  assign n32 = ~n_pad & ~o_pad ;
  assign n33 = m_pad & n_pad ;
  assign n34 = ~n32 & ~n33 ;
  assign n42 = ~n31 & ~n34 ;
  assign n36 = ~g_pad & ~h_pad ;
  assign n37 = ~n19 & ~n36 ;
  assign n38 = ~e_pad & ~f_pad ;
  assign n39 = e_pad & p_pad ;
  assign n40 = ~n38 & ~n39 ;
  assign n43 = ~n37 & ~n40 ;
  assign n44 = n42 & n43 ;
  assign n45 = n41 & n44 ;
  assign n46 = ~p_pad & n45 ;
  assign n47 = o_pad & n45 ;
  assign n48 = ~k_pad & ~p_pad ;
  assign n49 = n28 & n48 ;
  assign n50 = n30 & n32 ;
  assign n51 = n36 & n38 ;
  assign n52 = n50 & n51 ;
  assign n53 = n49 & n52 ;
  assign q_pad = n27 ;
  assign r_pad = ~n46 ;
  assign s_pad = ~n47 ;
  assign t_pad = n53 ;
endmodule
