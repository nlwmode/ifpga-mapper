module top( \G0_pad  , \G10_pad  , \G11_pad  , \G12_pad  , \G13_pad  , \G14_pad  , \G15_pad  , \G16_pad  , \G18_pad  , \G1_pad  , \G2_pad  , \G38_reg/NET0131  , \G39_reg/NET0131  , \G3_pad  , \G40_reg/NET0131  , \G41_reg/NET0131  , \G42_reg/NET0131  , \G4_pad  , \G5_pad  , \G6_pad  , \G7_pad  , \G8_pad  , \G9_pad  , \G288_pad  , \G290_pad  , \G296_pad  , \G302_pad  , \G315_pad  , \G325_pad  , \G327_pad  , \G45_pad  , \G47_pad  , \G49_pad  , \G53_pad  , \G55_pad  , \_al_n0  , \_al_n1  , \g1404/_0_  , \g1412/_0_  , \g1416/_0_  , \g1451/_2_  , \g1459/_3_  , \g1511/_3_  , \g1527/_3_  , \g1529/_3_  , \g31/_0_  , \g33/_1_  , \g56/_3_  );
  input \G0_pad  ;
  input \G10_pad  ;
  input \G11_pad  ;
  input \G12_pad  ;
  input \G13_pad  ;
  input \G14_pad  ;
  input \G15_pad  ;
  input \G16_pad  ;
  input \G18_pad  ;
  input \G1_pad  ;
  input \G2_pad  ;
  input \G38_reg/NET0131  ;
  input \G39_reg/NET0131  ;
  input \G3_pad  ;
  input \G40_reg/NET0131  ;
  input \G41_reg/NET0131  ;
  input \G42_reg/NET0131  ;
  input \G4_pad  ;
  input \G5_pad  ;
  input \G6_pad  ;
  input \G7_pad  ;
  input \G8_pad  ;
  input \G9_pad  ;
  output \G288_pad  ;
  output \G290_pad  ;
  output \G296_pad  ;
  output \G302_pad  ;
  output \G315_pad  ;
  output \G325_pad  ;
  output \G327_pad  ;
  output \G45_pad  ;
  output \G47_pad  ;
  output \G49_pad  ;
  output \G53_pad  ;
  output \G55_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1404/_0_  ;
  output \g1412/_0_  ;
  output \g1416/_0_  ;
  output \g1451/_2_  ;
  output \g1459/_3_  ;
  output \g1511/_3_  ;
  output \g1527/_3_  ;
  output \g1529/_3_  ;
  output \g31/_0_  ;
  output \g33/_1_  ;
  output \g56/_3_  ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 ;
  assign n24 = \G39_reg/NET0131  & \G40_reg/NET0131  ;
  assign n25 = ~\G38_reg/NET0131  & ~\G41_reg/NET0131  ;
  assign n26 = ~\G42_reg/NET0131  & n25 ;
  assign n27 = n24 & n26 ;
  assign n29 = \G15_pad  & \G39_reg/NET0131  ;
  assign n28 = ~\G40_reg/NET0131  & ~\G41_reg/NET0131  ;
  assign n30 = ~\G42_reg/NET0131  & n28 ;
  assign n31 = n29 & n30 ;
  assign n32 = \G40_reg/NET0131  & \G41_reg/NET0131  ;
  assign n33 = ~\G42_reg/NET0131  & n32 ;
  assign n34 = ~\G38_reg/NET0131  & n33 ;
  assign n35 = \G39_reg/NET0131  & n34 ;
  assign n44 = ~\G41_reg/NET0131  & ~\G42_reg/NET0131  ;
  assign n45 = \G38_reg/NET0131  & n44 ;
  assign n46 = \G40_reg/NET0131  & ~n45 ;
  assign n47 = \G4_pad  & ~n46 ;
  assign n37 = \G41_reg/NET0131  & \G42_reg/NET0131  ;
  assign n48 = ~\G16_pad  & ~n37 ;
  assign n49 = ~\G40_reg/NET0131  & n48 ;
  assign n50 = ~n47 & ~n49 ;
  assign n51 = \G39_reg/NET0131  & ~n50 ;
  assign n36 = \G16_pad  & ~\G4_pad  ;
  assign n38 = \G40_reg/NET0131  & n37 ;
  assign n39 = \G38_reg/NET0131  & ~n38 ;
  assign n40 = ~\G40_reg/NET0131  & ~n37 ;
  assign n41 = ~\G39_reg/NET0131  & ~n40 ;
  assign n42 = ~n39 & n41 ;
  assign n43 = ~n36 & n42 ;
  assign n53 = ~\G39_reg/NET0131  & ~\G40_reg/NET0131  ;
  assign n54 = n44 & n53 ;
  assign n52 = \G16_pad  & ~\G38_reg/NET0131  ;
  assign n55 = ~\G1_pad  & n52 ;
  assign n56 = n54 & n55 ;
  assign n57 = ~n43 & ~n56 ;
  assign n58 = ~n51 & n57 ;
  assign n59 = n24 & n37 ;
  assign n60 = ~n54 & ~n59 ;
  assign n61 = ~\G38_reg/NET0131  & ~n60 ;
  assign n62 = \G42_reg/NET0131  & n24 ;
  assign n63 = n25 & n62 ;
  assign n64 = \G42_reg/NET0131  & n29 ;
  assign n65 = n28 & n64 ;
  assign n70 = \G15_pad  & n52 ;
  assign n66 = ~\G10_pad  & ~\G11_pad  ;
  assign n69 = ~\G39_reg/NET0131  & ~\G4_pad  ;
  assign n71 = ~n66 & n69 ;
  assign n72 = n70 & n71 ;
  assign n67 = \G10_pad  & \G11_pad  ;
  assign n68 = ~\G12_pad  & ~n67 ;
  assign n73 = n33 & ~n68 ;
  assign n74 = n72 & n73 ;
  assign n75 = ~\G5_pad  & n27 ;
  assign n76 = \G39_reg/NET0131  & ~n46 ;
  assign n77 = ~n42 & ~n76 ;
  assign n78 = ~\G40_reg/NET0131  & \G41_reg/NET0131  ;
  assign n79 = ~\G42_reg/NET0131  & n78 ;
  assign n80 = ~\G38_reg/NET0131  & ~\G39_reg/NET0131  ;
  assign n81 = n79 & n80 ;
  assign n82 = \G5_pad  & n27 ;
  assign n92 = \G13_pad  & \G15_pad  ;
  assign n93 = \G42_reg/NET0131  & n92 ;
  assign n90 = \G38_reg/NET0131  & ~\G42_reg/NET0131  ;
  assign n91 = \G40_reg/NET0131  & ~n90 ;
  assign n94 = ~\G15_pad  & ~\G42_reg/NET0131  ;
  assign n95 = n91 & ~n94 ;
  assign n96 = ~n93 & n95 ;
  assign n97 = ~\G39_reg/NET0131  & ~n96 ;
  assign n83 = \G6_pad  & \G7_pad  ;
  assign n84 = \G8_pad  & \G9_pad  ;
  assign n85 = n83 & n84 ;
  assign n86 = ~\G40_reg/NET0131  & ~n85 ;
  assign n87 = \G38_reg/NET0131  & \G39_reg/NET0131  ;
  assign n88 = ~n86 & n87 ;
  assign n89 = ~\G15_pad  & ~\G40_reg/NET0131  ;
  assign n98 = \G41_reg/NET0131  & ~n89 ;
  assign n99 = ~n88 & n98 ;
  assign n100 = ~n97 & n99 ;
  assign n101 = ~\G1_pad  & n28 ;
  assign n104 = ~\G7_pad  & ~\G8_pad  ;
  assign n105 = \G9_pad  & n104 ;
  assign n102 = \G15_pad  & \G40_reg/NET0131  ;
  assign n103 = ~\G42_reg/NET0131  & \G6_pad  ;
  assign n106 = n102 & n103 ;
  assign n107 = n105 & n106 ;
  assign n108 = ~n101 & ~n107 ;
  assign n109 = n80 & ~n108 ;
  assign n110 = ~\G41_reg/NET0131  & \G42_reg/NET0131  ;
  assign n111 = ~\G39_reg/NET0131  & ~n110 ;
  assign n112 = ~\G40_reg/NET0131  & ~n94 ;
  assign n113 = ~n64 & n112 ;
  assign n114 = ~n111 & n113 ;
  assign n115 = ~\G15_pad  & ~\G38_reg/NET0131  ;
  assign n116 = ~\G39_reg/NET0131  & \G42_reg/NET0131  ;
  assign n117 = n115 & n116 ;
  assign n118 = ~n114 & ~n117 ;
  assign n119 = ~n109 & n118 ;
  assign n120 = ~n100 & n119 ;
  assign n121 = \G16_pad  & ~n120 ;
  assign n127 = ~\G41_reg/NET0131  & \G5_pad  ;
  assign n128 = ~\G42_reg/NET0131  & ~n127 ;
  assign n130 = ~\G1_pad  & ~\G3_pad  ;
  assign n131 = n110 & n130 ;
  assign n132 = ~n128 & ~n131 ;
  assign n129 = \G2_pad  & ~n128 ;
  assign n133 = n24 & ~n129 ;
  assign n134 = ~n132 & n133 ;
  assign n122 = \G15_pad  & ~\G39_reg/NET0131  ;
  assign n123 = \G14_pad  & n122 ;
  assign n124 = n79 & n123 ;
  assign n125 = \G4_pad  & ~n40 ;
  assign n126 = ~\G39_reg/NET0131  & n125 ;
  assign n135 = ~n124 & ~n126 ;
  assign n136 = ~n134 & n135 ;
  assign n137 = ~\G38_reg/NET0131  & ~n136 ;
  assign n138 = \G4_pad  & n76 ;
  assign n139 = \G0_pad  & \G39_reg/NET0131  ;
  assign n140 = \G38_reg/NET0131  & ~n69 ;
  assign n141 = ~n139 & n140 ;
  assign n142 = n38 & n141 ;
  assign n143 = ~n138 & ~n142 ;
  assign n144 = ~n137 & n143 ;
  assign n145 = ~n121 & n144 ;
  assign n146 = ~\G18_pad  & ~n145 ;
  assign n149 = ~\G4_pad  & n44 ;
  assign n148 = ~\G0_pad  & n37 ;
  assign n150 = \G38_reg/NET0131  & ~n148 ;
  assign n151 = ~n149 & n150 ;
  assign n147 = ~\G38_reg/NET0131  & n132 ;
  assign n152 = n24 & ~n147 ;
  assign n153 = ~n151 & n152 ;
  assign n173 = \G15_pad  & \G38_reg/NET0131  ;
  assign n174 = n85 & n173 ;
  assign n175 = \G16_pad  & ~n174 ;
  assign n171 = \G39_reg/NET0131  & ~\G4_pad  ;
  assign n172 = ~\G40_reg/NET0131  & n171 ;
  assign n176 = n37 & n172 ;
  assign n177 = ~n175 & n176 ;
  assign n157 = \G16_pad  & n69 ;
  assign n158 = ~n89 & n157 ;
  assign n159 = ~n40 & n158 ;
  assign n154 = ~\G42_reg/NET0131  & ~n66 ;
  assign n155 = \G15_pad  & n32 ;
  assign n156 = ~n154 & n155 ;
  assign n160 = ~n39 & ~n156 ;
  assign n161 = n159 & n160 ;
  assign n166 = \G2_pad  & n130 ;
  assign n167 = ~\G16_pad  & n166 ;
  assign n168 = ~\G41_reg/NET0131  & ~n167 ;
  assign n162 = ~\G40_reg/NET0131  & ~\G42_reg/NET0131  ;
  assign n163 = ~\G14_pad  & \G15_pad  ;
  assign n164 = \G41_reg/NET0131  & ~n163 ;
  assign n165 = n162 & ~n164 ;
  assign n169 = n80 & n165 ;
  assign n170 = ~n168 & n169 ;
  assign n178 = ~n161 & ~n170 ;
  assign n179 = ~n177 & n178 ;
  assign n180 = ~n153 & n179 ;
  assign n181 = ~\G18_pad  & ~n180 ;
  assign n183 = \G38_reg/NET0131  & ~n33 ;
  assign n182 = ~\G39_reg/NET0131  & ~n32 ;
  assign n184 = ~n62 & ~n182 ;
  assign n185 = n183 & n184 ;
  assign n186 = \G10_pad  & \G12_pad  ;
  assign n187 = ~\G11_pad  & ~n186 ;
  assign n188 = n122 & ~n187 ;
  assign n189 = n34 & n188 ;
  assign n190 = ~n185 & ~n189 ;
  assign n191 = n36 & ~n190 ;
  assign n193 = \G16_pad  & \G38_reg/NET0131  ;
  assign n194 = ~\G16_pad  & ~\G1_pad  ;
  assign n195 = ~\G38_reg/NET0131  & n194 ;
  assign n196 = ~\G42_reg/NET0131  & ~n195 ;
  assign n197 = ~n193 & ~n196 ;
  assign n192 = \G0_pad  & n90 ;
  assign n198 = ~\G39_reg/NET0131  & n28 ;
  assign n199 = ~n192 & n198 ;
  assign n200 = ~n197 & n199 ;
  assign n201 = ~\G0_pad  & n87 ;
  assign n202 = \G1_pad  & \G39_reg/NET0131  ;
  assign n203 = ~\G41_reg/NET0131  & n202 ;
  assign n204 = ~n201 & ~n203 ;
  assign n205 = \G38_reg/NET0131  & ~\G41_reg/NET0131  ;
  assign n206 = \G40_reg/NET0131  & \G42_reg/NET0131  ;
  assign n207 = ~n205 & n206 ;
  assign n208 = ~n204 & n207 ;
  assign n209 = ~n200 & ~n208 ;
  assign n210 = ~n191 & n209 ;
  assign n211 = ~\G18_pad  & ~n210 ;
  assign n212 = ~\G42_reg/NET0131  & n53 ;
  assign n213 = ~n62 & ~n212 ;
  assign n214 = \G1_pad  & n25 ;
  assign n215 = ~n213 & n214 ;
  assign n216 = \G3_pad  & n54 ;
  assign n217 = n195 & n216 ;
  assign n218 = n52 & n59 ;
  assign n219 = \G15_pad  & n81 ;
  assign n220 = ~\G38_reg/NET0131  & n124 ;
  assign n236 = ~\G39_reg/NET0131  & ~n125 ;
  assign n233 = n102 & n110 ;
  assign n234 = \G16_pad  & ~n162 ;
  assign n235 = ~n233 & n234 ;
  assign n237 = ~n165 & ~n235 ;
  assign n238 = n236 & n237 ;
  assign n223 = \G41_reg/NET0131  & ~\G4_pad  ;
  assign n224 = ~\G41_reg/NET0131  & ~\G5_pad  ;
  assign n225 = \G39_reg/NET0131  & ~n224 ;
  assign n226 = ~n223 & ~n225 ;
  assign n221 = ~\G16_pad  & \G41_reg/NET0131  ;
  assign n222 = \G42_reg/NET0131  & ~n221 ;
  assign n227 = \G40_reg/NET0131  & ~n222 ;
  assign n228 = ~n226 & n227 ;
  assign n229 = ~\G16_pad  & n53 ;
  assign n230 = ~n62 & ~n229 ;
  assign n231 = ~\G41_reg/NET0131  & n166 ;
  assign n232 = ~n230 & n231 ;
  assign n239 = ~n228 & ~n232 ;
  assign n240 = ~n238 & n239 ;
  assign n241 = ~\G38_reg/NET0131  & ~n240 ;
  assign n250 = ~\G39_reg/NET0131  & ~n115 ;
  assign n251 = ~\G40_reg/NET0131  & n223 ;
  assign n252 = ~n250 & n251 ;
  assign n253 = n175 & n252 ;
  assign n242 = \G16_pad  & n92 ;
  assign n243 = n69 & ~n242 ;
  assign n244 = ~n201 & ~n243 ;
  assign n245 = n38 & ~n244 ;
  assign n246 = \G15_pad  & ~n44 ;
  assign n247 = \G16_pad  & ~n246 ;
  assign n248 = n40 & n171 ;
  assign n249 = ~n247 & n248 ;
  assign n254 = ~n245 & ~n249 ;
  assign n255 = ~n253 & n254 ;
  assign n256 = ~n241 & n255 ;
  assign n257 = ~\G18_pad  & ~n256 ;
  assign n259 = n68 & n154 ;
  assign n260 = \G16_pad  & n122 ;
  assign n261 = n223 & n260 ;
  assign n262 = n91 & n261 ;
  assign n263 = ~n259 & n262 ;
  assign n258 = ~n48 & n172 ;
  assign n264 = n26 & n53 ;
  assign n265 = n167 & n264 ;
  assign n266 = ~n258 & ~n265 ;
  assign n267 = ~n263 & n266 ;
  assign n268 = ~n153 & n267 ;
  assign n269 = ~\G18_pad  & ~n268 ;
  assign \G288_pad  = n27 ;
  assign \G290_pad  = n31 ;
  assign \G296_pad  = n35 ;
  assign \G302_pad  = ~n58 ;
  assign \G315_pad  = n61 ;
  assign \G325_pad  = n63 ;
  assign \G327_pad  = n65 ;
  assign \G45_pad  = n74 ;
  assign \G47_pad  = n75 ;
  assign \G49_pad  = ~n77 ;
  assign \G53_pad  = n81 ;
  assign \G55_pad  = n82 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1404/_0_  = n146 ;
  assign \g1412/_0_  = n181 ;
  assign \g1416/_0_  = n211 ;
  assign \g1451/_2_  = n215 ;
  assign \g1459/_3_  = n217 ;
  assign \g1511/_3_  = n218 ;
  assign \g1527/_3_  = n219 ;
  assign \g1529/_3_  = n220 ;
  assign \g31/_0_  = n257 ;
  assign \g33/_1_  = n269 ;
  assign \g56/_3_  = n177 ;
endmodule
