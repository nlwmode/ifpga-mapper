module top( \priority[0]  , \priority[1]  , \priority[2]  , \priority[3]  , \priority[4]  , \priority[5]  , \priority[6]  , \priority[7]  , \priority[8]  , \priority[9]  , \priority[10]  , \priority[11]  , \priority[12]  , \priority[13]  , \priority[14]  , \priority[15]  , \priority[16]  , \priority[17]  , \priority[18]  , \priority[19]  , \priority[20]  , \priority[21]  , \priority[22]  , \priority[23]  , \priority[24]  , \priority[25]  , \priority[26]  , \priority[27]  , \priority[28]  , \priority[29]  , \priority[30]  , \priority[31]  , \priority[32]  , \priority[33]  , \priority[34]  , \priority[35]  , \priority[36]  , \priority[37]  , \priority[38]  , \priority[39]  , \priority[40]  , \priority[41]  , \priority[42]  , \priority[43]  , \priority[44]  , \priority[45]  , \priority[46]  , \priority[47]  , \priority[48]  , \priority[49]  , \priority[50]  , \priority[51]  , \priority[52]  , \priority[53]  , \priority[54]  , \priority[55]  , \priority[56]  , \priority[57]  , \priority[58]  , \priority[59]  , \priority[60]  , \priority[61]  , \priority[62]  , \priority[63]  , \priority[64]  , \priority[65]  , \priority[66]  , \priority[67]  , \priority[68]  , \priority[69]  , \priority[70]  , \priority[71]  , \priority[72]  , \priority[73]  , \priority[74]  , \priority[75]  , \priority[76]  , \priority[77]  , \priority[78]  , \priority[79]  , \priority[80]  , \priority[81]  , \priority[82]  , \priority[83]  , \priority[84]  , \priority[85]  , \priority[86]  , \priority[87]  , \priority[88]  , \priority[89]  , \priority[90]  , \priority[91]  , \priority[92]  , \priority[93]  , \priority[94]  , \priority[95]  , \priority[96]  , \priority[97]  , \priority[98]  , \priority[99]  , \priority[100]  , \priority[101]  , \priority[102]  , \priority[103]  , \priority[104]  , \priority[105]  , \priority[106]  , \priority[107]  , \priority[108]  , \priority[109]  , \priority[110]  , \priority[111]  , \priority[112]  , \priority[113]  , \priority[114]  , \priority[115]  , \priority[116]  , \priority[117]  , \priority[118]  , \priority[119]  , \priority[120]  , \priority[121]  , \priority[122]  , \priority[123]  , \priority[124]  , \priority[125]  , \priority[126]  , \priority[127]  , \req[0]  , \req[1]  , \req[2]  , \req[3]  , \req[4]  , \req[5]  , \req[6]  , \req[7]  , \req[8]  , \req[9]  , \req[10]  , \req[11]  , \req[12]  , \req[13]  , \req[14]  , \req[15]  , \req[16]  , \req[17]  , \req[18]  , \req[19]  , \req[20]  , \req[21]  , \req[22]  , \req[23]  , \req[24]  , \req[25]  , \req[26]  , \req[27]  , \req[28]  , \req[29]  , \req[30]  , \req[31]  , \req[32]  , \req[33]  , \req[34]  , \req[35]  , \req[36]  , \req[37]  , \req[38]  , \req[39]  , \req[40]  , \req[41]  , \req[42]  , \req[43]  , \req[44]  , \req[45]  , \req[46]  , \req[47]  , \req[48]  , \req[49]  , \req[50]  , \req[51]  , \req[52]  , \req[53]  , \req[54]  , \req[55]  , \req[56]  , \req[57]  , \req[58]  , \req[59]  , \req[60]  , \req[61]  , \req[62]  , \req[63]  , \req[64]  , \req[65]  , \req[66]  , \req[67]  , \req[68]  , \req[69]  , \req[70]  , \req[71]  , \req[72]  , \req[73]  , \req[74]  , \req[75]  , \req[76]  , \req[77]  , \req[78]  , \req[79]  , \req[80]  , \req[81]  , \req[82]  , \req[83]  , \req[84]  , \req[85]  , \req[86]  , \req[87]  , \req[88]  , \req[89]  , \req[90]  , \req[91]  , \req[92]  , \req[93]  , \req[94]  , \req[95]  , \req[96]  , \req[97]  , \req[98]  , \req[99]  , \req[100]  , \req[101]  , \req[102]  , \req[103]  , \req[104]  , \req[105]  , \req[106]  , \req[107]  , \req[108]  , \req[109]  , \req[110]  , \req[111]  , \req[112]  , \req[113]  , \req[114]  , \req[115]  , \req[116]  , \req[117]  , \req[118]  , \req[119]  , \req[120]  , \req[121]  , \req[122]  , \req[123]  , \req[124]  , \req[125]  , \req[126]  , \req[127]  , \grant[0]  , \grant[1]  , \grant[2]  , \grant[3]  , \grant[4]  , \grant[5]  , \grant[6]  , \grant[7]  , \grant[8]  , \grant[9]  , \grant[10]  , \grant[11]  , \grant[12]  , \grant[13]  , \grant[14]  , \grant[15]  , \grant[16]  , \grant[17]  , \grant[18]  , \grant[19]  , \grant[20]  , \grant[21]  , \grant[22]  , \grant[23]  , \grant[24]  , \grant[25]  , \grant[26]  , \grant[27]  , \grant[28]  , \grant[29]  , \grant[30]  , \grant[31]  , \grant[32]  , \grant[33]  , \grant[34]  , \grant[35]  , \grant[36]  , \grant[37]  , \grant[38]  , \grant[39]  , \grant[40]  , \grant[41]  , \grant[42]  , \grant[43]  , \grant[44]  , \grant[45]  , \grant[46]  , \grant[47]  , \grant[48]  , \grant[49]  , \grant[50]  , \grant[51]  , \grant[52]  , \grant[53]  , \grant[54]  , \grant[55]  , \grant[56]  , \grant[57]  , \grant[58]  , \grant[59]  , \grant[60]  , \grant[61]  , \grant[62]  , \grant[63]  , \grant[64]  , \grant[65]  , \grant[66]  , \grant[67]  , \grant[68]  , \grant[69]  , \grant[70]  , \grant[71]  , \grant[72]  , \grant[73]  , \grant[74]  , \grant[75]  , \grant[76]  , \grant[77]  , \grant[78]  , \grant[79]  , \grant[80]  , \grant[81]  , \grant[82]  , \grant[83]  , \grant[84]  , \grant[85]  , \grant[86]  , \grant[87]  , \grant[88]  , \grant[89]  , \grant[90]  , \grant[91]  , \grant[92]  , \grant[93]  , \grant[94]  , \grant[95]  , \grant[96]  , \grant[97]  , \grant[98]  , \grant[99]  , \grant[100]  , \grant[101]  , \grant[102]  , \grant[103]  , \grant[104]  , \grant[105]  , \grant[106]  , \grant[107]  , \grant[108]  , \grant[109]  , \grant[110]  , \grant[111]  , \grant[112]  , \grant[113]  , \grant[114]  , \grant[115]  , \grant[116]  , \grant[117]  , \grant[118]  , \grant[119]  , \grant[120]  , \grant[121]  , \grant[122]  , \grant[123]  , \grant[124]  , \grant[125]  , \grant[126]  , \grant[127]  , anyGrant );
  input \priority[0]  ;
  input \priority[1]  ;
  input \priority[2]  ;
  input \priority[3]  ;
  input \priority[4]  ;
  input \priority[5]  ;
  input \priority[6]  ;
  input \priority[7]  ;
  input \priority[8]  ;
  input \priority[9]  ;
  input \priority[10]  ;
  input \priority[11]  ;
  input \priority[12]  ;
  input \priority[13]  ;
  input \priority[14]  ;
  input \priority[15]  ;
  input \priority[16]  ;
  input \priority[17]  ;
  input \priority[18]  ;
  input \priority[19]  ;
  input \priority[20]  ;
  input \priority[21]  ;
  input \priority[22]  ;
  input \priority[23]  ;
  input \priority[24]  ;
  input \priority[25]  ;
  input \priority[26]  ;
  input \priority[27]  ;
  input \priority[28]  ;
  input \priority[29]  ;
  input \priority[30]  ;
  input \priority[31]  ;
  input \priority[32]  ;
  input \priority[33]  ;
  input \priority[34]  ;
  input \priority[35]  ;
  input \priority[36]  ;
  input \priority[37]  ;
  input \priority[38]  ;
  input \priority[39]  ;
  input \priority[40]  ;
  input \priority[41]  ;
  input \priority[42]  ;
  input \priority[43]  ;
  input \priority[44]  ;
  input \priority[45]  ;
  input \priority[46]  ;
  input \priority[47]  ;
  input \priority[48]  ;
  input \priority[49]  ;
  input \priority[50]  ;
  input \priority[51]  ;
  input \priority[52]  ;
  input \priority[53]  ;
  input \priority[54]  ;
  input \priority[55]  ;
  input \priority[56]  ;
  input \priority[57]  ;
  input \priority[58]  ;
  input \priority[59]  ;
  input \priority[60]  ;
  input \priority[61]  ;
  input \priority[62]  ;
  input \priority[63]  ;
  input \priority[64]  ;
  input \priority[65]  ;
  input \priority[66]  ;
  input \priority[67]  ;
  input \priority[68]  ;
  input \priority[69]  ;
  input \priority[70]  ;
  input \priority[71]  ;
  input \priority[72]  ;
  input \priority[73]  ;
  input \priority[74]  ;
  input \priority[75]  ;
  input \priority[76]  ;
  input \priority[77]  ;
  input \priority[78]  ;
  input \priority[79]  ;
  input \priority[80]  ;
  input \priority[81]  ;
  input \priority[82]  ;
  input \priority[83]  ;
  input \priority[84]  ;
  input \priority[85]  ;
  input \priority[86]  ;
  input \priority[87]  ;
  input \priority[88]  ;
  input \priority[89]  ;
  input \priority[90]  ;
  input \priority[91]  ;
  input \priority[92]  ;
  input \priority[93]  ;
  input \priority[94]  ;
  input \priority[95]  ;
  input \priority[96]  ;
  input \priority[97]  ;
  input \priority[98]  ;
  input \priority[99]  ;
  input \priority[100]  ;
  input \priority[101]  ;
  input \priority[102]  ;
  input \priority[103]  ;
  input \priority[104]  ;
  input \priority[105]  ;
  input \priority[106]  ;
  input \priority[107]  ;
  input \priority[108]  ;
  input \priority[109]  ;
  input \priority[110]  ;
  input \priority[111]  ;
  input \priority[112]  ;
  input \priority[113]  ;
  input \priority[114]  ;
  input \priority[115]  ;
  input \priority[116]  ;
  input \priority[117]  ;
  input \priority[118]  ;
  input \priority[119]  ;
  input \priority[120]  ;
  input \priority[121]  ;
  input \priority[122]  ;
  input \priority[123]  ;
  input \priority[124]  ;
  input \priority[125]  ;
  input \priority[126]  ;
  input \priority[127]  ;
  input \req[0]  ;
  input \req[1]  ;
  input \req[2]  ;
  input \req[3]  ;
  input \req[4]  ;
  input \req[5]  ;
  input \req[6]  ;
  input \req[7]  ;
  input \req[8]  ;
  input \req[9]  ;
  input \req[10]  ;
  input \req[11]  ;
  input \req[12]  ;
  input \req[13]  ;
  input \req[14]  ;
  input \req[15]  ;
  input \req[16]  ;
  input \req[17]  ;
  input \req[18]  ;
  input \req[19]  ;
  input \req[20]  ;
  input \req[21]  ;
  input \req[22]  ;
  input \req[23]  ;
  input \req[24]  ;
  input \req[25]  ;
  input \req[26]  ;
  input \req[27]  ;
  input \req[28]  ;
  input \req[29]  ;
  input \req[30]  ;
  input \req[31]  ;
  input \req[32]  ;
  input \req[33]  ;
  input \req[34]  ;
  input \req[35]  ;
  input \req[36]  ;
  input \req[37]  ;
  input \req[38]  ;
  input \req[39]  ;
  input \req[40]  ;
  input \req[41]  ;
  input \req[42]  ;
  input \req[43]  ;
  input \req[44]  ;
  input \req[45]  ;
  input \req[46]  ;
  input \req[47]  ;
  input \req[48]  ;
  input \req[49]  ;
  input \req[50]  ;
  input \req[51]  ;
  input \req[52]  ;
  input \req[53]  ;
  input \req[54]  ;
  input \req[55]  ;
  input \req[56]  ;
  input \req[57]  ;
  input \req[58]  ;
  input \req[59]  ;
  input \req[60]  ;
  input \req[61]  ;
  input \req[62]  ;
  input \req[63]  ;
  input \req[64]  ;
  input \req[65]  ;
  input \req[66]  ;
  input \req[67]  ;
  input \req[68]  ;
  input \req[69]  ;
  input \req[70]  ;
  input \req[71]  ;
  input \req[72]  ;
  input \req[73]  ;
  input \req[74]  ;
  input \req[75]  ;
  input \req[76]  ;
  input \req[77]  ;
  input \req[78]  ;
  input \req[79]  ;
  input \req[80]  ;
  input \req[81]  ;
  input \req[82]  ;
  input \req[83]  ;
  input \req[84]  ;
  input \req[85]  ;
  input \req[86]  ;
  input \req[87]  ;
  input \req[88]  ;
  input \req[89]  ;
  input \req[90]  ;
  input \req[91]  ;
  input \req[92]  ;
  input \req[93]  ;
  input \req[94]  ;
  input \req[95]  ;
  input \req[96]  ;
  input \req[97]  ;
  input \req[98]  ;
  input \req[99]  ;
  input \req[100]  ;
  input \req[101]  ;
  input \req[102]  ;
  input \req[103]  ;
  input \req[104]  ;
  input \req[105]  ;
  input \req[106]  ;
  input \req[107]  ;
  input \req[108]  ;
  input \req[109]  ;
  input \req[110]  ;
  input \req[111]  ;
  input \req[112]  ;
  input \req[113]  ;
  input \req[114]  ;
  input \req[115]  ;
  input \req[116]  ;
  input \req[117]  ;
  input \req[118]  ;
  input \req[119]  ;
  input \req[120]  ;
  input \req[121]  ;
  input \req[122]  ;
  input \req[123]  ;
  input \req[124]  ;
  input \req[125]  ;
  input \req[126]  ;
  input \req[127]  ;
  output \grant[0]  ;
  output \grant[1]  ;
  output \grant[2]  ;
  output \grant[3]  ;
  output \grant[4]  ;
  output \grant[5]  ;
  output \grant[6]  ;
  output \grant[7]  ;
  output \grant[8]  ;
  output \grant[9]  ;
  output \grant[10]  ;
  output \grant[11]  ;
  output \grant[12]  ;
  output \grant[13]  ;
  output \grant[14]  ;
  output \grant[15]  ;
  output \grant[16]  ;
  output \grant[17]  ;
  output \grant[18]  ;
  output \grant[19]  ;
  output \grant[20]  ;
  output \grant[21]  ;
  output \grant[22]  ;
  output \grant[23]  ;
  output \grant[24]  ;
  output \grant[25]  ;
  output \grant[26]  ;
  output \grant[27]  ;
  output \grant[28]  ;
  output \grant[29]  ;
  output \grant[30]  ;
  output \grant[31]  ;
  output \grant[32]  ;
  output \grant[33]  ;
  output \grant[34]  ;
  output \grant[35]  ;
  output \grant[36]  ;
  output \grant[37]  ;
  output \grant[38]  ;
  output \grant[39]  ;
  output \grant[40]  ;
  output \grant[41]  ;
  output \grant[42]  ;
  output \grant[43]  ;
  output \grant[44]  ;
  output \grant[45]  ;
  output \grant[46]  ;
  output \grant[47]  ;
  output \grant[48]  ;
  output \grant[49]  ;
  output \grant[50]  ;
  output \grant[51]  ;
  output \grant[52]  ;
  output \grant[53]  ;
  output \grant[54]  ;
  output \grant[55]  ;
  output \grant[56]  ;
  output \grant[57]  ;
  output \grant[58]  ;
  output \grant[59]  ;
  output \grant[60]  ;
  output \grant[61]  ;
  output \grant[62]  ;
  output \grant[63]  ;
  output \grant[64]  ;
  output \grant[65]  ;
  output \grant[66]  ;
  output \grant[67]  ;
  output \grant[68]  ;
  output \grant[69]  ;
  output \grant[70]  ;
  output \grant[71]  ;
  output \grant[72]  ;
  output \grant[73]  ;
  output \grant[74]  ;
  output \grant[75]  ;
  output \grant[76]  ;
  output \grant[77]  ;
  output \grant[78]  ;
  output \grant[79]  ;
  output \grant[80]  ;
  output \grant[81]  ;
  output \grant[82]  ;
  output \grant[83]  ;
  output \grant[84]  ;
  output \grant[85]  ;
  output \grant[86]  ;
  output \grant[87]  ;
  output \grant[88]  ;
  output \grant[89]  ;
  output \grant[90]  ;
  output \grant[91]  ;
  output \grant[92]  ;
  output \grant[93]  ;
  output \grant[94]  ;
  output \grant[95]  ;
  output \grant[96]  ;
  output \grant[97]  ;
  output \grant[98]  ;
  output \grant[99]  ;
  output \grant[100]  ;
  output \grant[101]  ;
  output \grant[102]  ;
  output \grant[103]  ;
  output \grant[104]  ;
  output \grant[105]  ;
  output \grant[106]  ;
  output \grant[107]  ;
  output \grant[108]  ;
  output \grant[109]  ;
  output \grant[110]  ;
  output \grant[111]  ;
  output \grant[112]  ;
  output \grant[113]  ;
  output \grant[114]  ;
  output \grant[115]  ;
  output \grant[116]  ;
  output \grant[117]  ;
  output \grant[118]  ;
  output \grant[119]  ;
  output \grant[120]  ;
  output \grant[121]  ;
  output \grant[122]  ;
  output \grant[123]  ;
  output \grant[124]  ;
  output \grant[125]  ;
  output \grant[126]  ;
  output \grant[127]  ;
  output anyGrant ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 ;
  assign n257 = \priority[126]  & ~\req[126]  ;
  assign n258 = ~\priority[0]  & ~\priority[127]  ;
  assign n259 = ~n257 & n258 ;
  assign n260 = ~\priority[0]  & \req[127]  ;
  assign n261 = \req[0]  & ~n260 ;
  assign n262 = ~n259 & n261 ;
  assign n263 = \priority[1]  & ~\req[1]  ;
  assign n264 = ~\priority[2]  & ~n263 ;
  assign n265 = ~\req[2]  & ~\req[3]  ;
  assign n266 = ~n264 & n265 ;
  assign n267 = \priority[6]  & ~\req[6]  ;
  assign n268 = ~\priority[7]  & ~\priority[8]  ;
  assign n269 = ~n267 & n268 ;
  assign n270 = \priority[3]  & ~\req[3]  ;
  assign n271 = ~\priority[4]  & ~\priority[5]  ;
  assign n272 = ~n270 & n271 ;
  assign n273 = n269 & n272 ;
  assign n274 = ~n266 & n273 ;
  assign n275 = ~\priority[5]  & \req[4]  ;
  assign n276 = ~\req[5]  & ~\req[6]  ;
  assign n277 = ~n275 & n276 ;
  assign n278 = n269 & ~n277 ;
  assign n279 = ~\priority[11]  & \req[10]  ;
  assign n280 = ~\req[11]  & ~\req[12]  ;
  assign n281 = ~n279 & n280 ;
  assign n282 = ~\priority[8]  & \req[7]  ;
  assign n283 = ~\req[8]  & ~\req[9]  ;
  assign n284 = ~n282 & n283 ;
  assign n285 = n281 & n284 ;
  assign n286 = ~n278 & n285 ;
  assign n287 = ~n274 & n286 ;
  assign n288 = \priority[9]  & ~\req[9]  ;
  assign n289 = ~\priority[10]  & ~\priority[11]  ;
  assign n290 = ~n288 & n289 ;
  assign n291 = n281 & ~n290 ;
  assign n292 = \priority[15]  & ~\req[15]  ;
  assign n293 = ~\priority[16]  & ~\priority[17]  ;
  assign n294 = ~n292 & n293 ;
  assign n295 = \priority[12]  & ~\req[12]  ;
  assign n296 = ~\priority[13]  & ~\priority[14]  ;
  assign n297 = ~n295 & n296 ;
  assign n298 = n294 & n297 ;
  assign n299 = ~n291 & n298 ;
  assign n300 = ~n287 & n299 ;
  assign n301 = ~\priority[14]  & \req[13]  ;
  assign n302 = ~\req[14]  & ~\req[15]  ;
  assign n303 = ~n301 & n302 ;
  assign n304 = n294 & ~n303 ;
  assign n305 = ~\priority[20]  & \req[19]  ;
  assign n306 = ~\req[20]  & ~\req[21]  ;
  assign n307 = ~n305 & n306 ;
  assign n308 = ~\priority[17]  & \req[16]  ;
  assign n309 = ~\req[17]  & ~\req[18]  ;
  assign n310 = ~n308 & n309 ;
  assign n311 = n307 & n310 ;
  assign n312 = ~n304 & n311 ;
  assign n313 = ~n300 & n312 ;
  assign n314 = \priority[18]  & ~\req[18]  ;
  assign n315 = ~\priority[19]  & ~\priority[20]  ;
  assign n316 = ~n314 & n315 ;
  assign n317 = n307 & ~n316 ;
  assign n318 = \priority[24]  & ~\req[24]  ;
  assign n319 = ~\priority[25]  & ~\priority[26]  ;
  assign n320 = ~n318 & n319 ;
  assign n321 = \priority[21]  & ~\req[21]  ;
  assign n322 = ~\priority[22]  & ~\priority[23]  ;
  assign n323 = ~n321 & n322 ;
  assign n324 = n320 & n323 ;
  assign n325 = ~n317 & n324 ;
  assign n326 = ~n313 & n325 ;
  assign n327 = ~\priority[23]  & \req[22]  ;
  assign n328 = ~\req[23]  & ~\req[24]  ;
  assign n329 = ~n327 & n328 ;
  assign n330 = n320 & ~n329 ;
  assign n331 = ~\priority[29]  & \req[28]  ;
  assign n332 = ~\req[29]  & ~\req[30]  ;
  assign n333 = ~n331 & n332 ;
  assign n334 = ~\priority[26]  & \req[25]  ;
  assign n335 = ~\req[26]  & ~\req[27]  ;
  assign n336 = ~n334 & n335 ;
  assign n337 = n333 & n336 ;
  assign n338 = ~n330 & n337 ;
  assign n339 = ~n326 & n338 ;
  assign n340 = \priority[27]  & ~\req[27]  ;
  assign n341 = ~\priority[28]  & ~\priority[29]  ;
  assign n342 = ~n340 & n341 ;
  assign n343 = n333 & ~n342 ;
  assign n344 = \priority[33]  & ~\req[33]  ;
  assign n345 = ~\priority[34]  & ~\priority[35]  ;
  assign n346 = ~n344 & n345 ;
  assign n347 = \priority[30]  & ~\req[30]  ;
  assign n348 = ~\priority[31]  & ~\priority[32]  ;
  assign n349 = ~n347 & n348 ;
  assign n350 = n346 & n349 ;
  assign n351 = ~n343 & n350 ;
  assign n352 = ~n339 & n351 ;
  assign n353 = ~\priority[32]  & \req[31]  ;
  assign n354 = ~\req[32]  & ~\req[33]  ;
  assign n355 = ~n353 & n354 ;
  assign n356 = n346 & ~n355 ;
  assign n357 = ~\priority[38]  & \req[37]  ;
  assign n358 = ~\req[38]  & ~\req[39]  ;
  assign n359 = ~n357 & n358 ;
  assign n360 = ~\priority[35]  & \req[34]  ;
  assign n361 = ~\req[35]  & ~\req[36]  ;
  assign n362 = ~n360 & n361 ;
  assign n363 = n359 & n362 ;
  assign n364 = ~n356 & n363 ;
  assign n365 = ~n352 & n364 ;
  assign n366 = \priority[36]  & ~\req[36]  ;
  assign n367 = ~\priority[37]  & ~\priority[38]  ;
  assign n368 = ~n366 & n367 ;
  assign n369 = n359 & ~n368 ;
  assign n370 = \priority[42]  & ~\req[42]  ;
  assign n371 = ~\priority[43]  & ~\priority[44]  ;
  assign n372 = ~n370 & n371 ;
  assign n373 = \priority[39]  & ~\req[39]  ;
  assign n374 = ~\priority[40]  & ~\priority[41]  ;
  assign n375 = ~n373 & n374 ;
  assign n376 = n372 & n375 ;
  assign n377 = ~n369 & n376 ;
  assign n378 = ~n365 & n377 ;
  assign n379 = ~\priority[41]  & \req[40]  ;
  assign n380 = ~\req[41]  & ~\req[42]  ;
  assign n381 = ~n379 & n380 ;
  assign n382 = n372 & ~n381 ;
  assign n383 = ~\priority[47]  & \req[46]  ;
  assign n384 = ~\req[47]  & ~\req[48]  ;
  assign n385 = ~n383 & n384 ;
  assign n386 = ~\priority[44]  & \req[43]  ;
  assign n387 = ~\req[44]  & ~\req[45]  ;
  assign n388 = ~n386 & n387 ;
  assign n389 = n385 & n388 ;
  assign n390 = ~n382 & n389 ;
  assign n391 = ~n378 & n390 ;
  assign n392 = \priority[45]  & ~\req[45]  ;
  assign n393 = ~\priority[46]  & ~\priority[47]  ;
  assign n394 = ~n392 & n393 ;
  assign n395 = n385 & ~n394 ;
  assign n396 = \priority[51]  & ~\req[51]  ;
  assign n397 = ~\priority[52]  & ~\priority[53]  ;
  assign n398 = ~n396 & n397 ;
  assign n399 = \priority[48]  & ~\req[48]  ;
  assign n400 = ~\priority[49]  & ~\priority[50]  ;
  assign n401 = ~n399 & n400 ;
  assign n402 = n398 & n401 ;
  assign n403 = ~n395 & n402 ;
  assign n404 = ~n391 & n403 ;
  assign n405 = ~\priority[50]  & \req[49]  ;
  assign n406 = ~\req[50]  & ~\req[51]  ;
  assign n407 = ~n405 & n406 ;
  assign n408 = n398 & ~n407 ;
  assign n409 = ~\priority[56]  & \req[55]  ;
  assign n410 = ~\req[56]  & ~\req[57]  ;
  assign n411 = ~n409 & n410 ;
  assign n412 = ~\priority[53]  & \req[52]  ;
  assign n413 = ~\req[53]  & ~\req[54]  ;
  assign n414 = ~n412 & n413 ;
  assign n415 = n411 & n414 ;
  assign n416 = ~n408 & n415 ;
  assign n417 = ~n404 & n416 ;
  assign n418 = \priority[54]  & ~\req[54]  ;
  assign n419 = ~\priority[55]  & ~\priority[56]  ;
  assign n420 = ~n418 & n419 ;
  assign n421 = n411 & ~n420 ;
  assign n422 = \priority[60]  & ~\req[60]  ;
  assign n423 = ~\priority[61]  & ~\priority[62]  ;
  assign n424 = ~n422 & n423 ;
  assign n425 = \priority[57]  & ~\req[57]  ;
  assign n426 = ~\priority[58]  & ~\priority[59]  ;
  assign n427 = ~n425 & n426 ;
  assign n428 = n424 & n427 ;
  assign n429 = ~n421 & n428 ;
  assign n430 = ~n417 & n429 ;
  assign n431 = ~\priority[59]  & \req[58]  ;
  assign n432 = ~\req[59]  & ~\req[60]  ;
  assign n433 = ~n431 & n432 ;
  assign n434 = n424 & ~n433 ;
  assign n435 = ~\priority[65]  & \req[64]  ;
  assign n436 = ~\req[65]  & ~\req[66]  ;
  assign n437 = ~n435 & n436 ;
  assign n438 = ~\priority[62]  & \req[61]  ;
  assign n439 = ~\req[62]  & ~\req[63]  ;
  assign n440 = ~n438 & n439 ;
  assign n441 = n437 & n440 ;
  assign n442 = ~n434 & n441 ;
  assign n443 = ~n430 & n442 ;
  assign n444 = \priority[63]  & ~\req[63]  ;
  assign n445 = ~\priority[64]  & ~\priority[65]  ;
  assign n446 = ~n444 & n445 ;
  assign n447 = n437 & ~n446 ;
  assign n448 = \priority[69]  & ~\req[69]  ;
  assign n449 = ~\priority[70]  & ~\priority[71]  ;
  assign n450 = ~n448 & n449 ;
  assign n451 = \priority[66]  & ~\req[66]  ;
  assign n452 = ~\priority[67]  & ~\priority[68]  ;
  assign n453 = ~n451 & n452 ;
  assign n454 = n450 & n453 ;
  assign n455 = ~n447 & n454 ;
  assign n456 = ~n443 & n455 ;
  assign n457 = ~\priority[68]  & \req[67]  ;
  assign n458 = ~\req[68]  & ~\req[69]  ;
  assign n459 = ~n457 & n458 ;
  assign n460 = n450 & ~n459 ;
  assign n461 = ~\priority[74]  & \req[73]  ;
  assign n462 = ~\req[74]  & ~\req[75]  ;
  assign n463 = ~n461 & n462 ;
  assign n464 = ~\priority[71]  & \req[70]  ;
  assign n465 = ~\req[71]  & ~\req[72]  ;
  assign n466 = ~n464 & n465 ;
  assign n467 = n463 & n466 ;
  assign n468 = ~n460 & n467 ;
  assign n469 = ~n456 & n468 ;
  assign n470 = \priority[72]  & ~\req[72]  ;
  assign n471 = ~\priority[73]  & ~\priority[74]  ;
  assign n472 = ~n470 & n471 ;
  assign n473 = n463 & ~n472 ;
  assign n474 = \priority[78]  & ~\req[78]  ;
  assign n475 = ~\priority[79]  & ~\priority[80]  ;
  assign n476 = ~n474 & n475 ;
  assign n477 = \priority[75]  & ~\req[75]  ;
  assign n478 = ~\priority[76]  & ~\priority[77]  ;
  assign n479 = ~n477 & n478 ;
  assign n480 = n476 & n479 ;
  assign n481 = ~n473 & n480 ;
  assign n482 = ~n469 & n481 ;
  assign n483 = ~\priority[77]  & \req[76]  ;
  assign n484 = ~\req[77]  & ~\req[78]  ;
  assign n485 = ~n483 & n484 ;
  assign n486 = n476 & ~n485 ;
  assign n487 = ~\priority[83]  & \req[82]  ;
  assign n488 = ~\req[83]  & ~\req[84]  ;
  assign n489 = ~n487 & n488 ;
  assign n490 = ~\priority[80]  & \req[79]  ;
  assign n491 = ~\req[80]  & ~\req[81]  ;
  assign n492 = ~n490 & n491 ;
  assign n493 = n489 & n492 ;
  assign n494 = ~n486 & n493 ;
  assign n495 = ~n482 & n494 ;
  assign n496 = \priority[81]  & ~\req[81]  ;
  assign n497 = ~\priority[82]  & ~\priority[83]  ;
  assign n498 = ~n496 & n497 ;
  assign n499 = n489 & ~n498 ;
  assign n500 = \priority[87]  & ~\req[87]  ;
  assign n501 = ~\priority[88]  & ~\priority[89]  ;
  assign n502 = ~n500 & n501 ;
  assign n503 = \priority[84]  & ~\req[84]  ;
  assign n504 = ~\priority[85]  & ~\priority[86]  ;
  assign n505 = ~n503 & n504 ;
  assign n506 = n502 & n505 ;
  assign n507 = ~n499 & n506 ;
  assign n508 = ~n495 & n507 ;
  assign n509 = ~\priority[86]  & \req[85]  ;
  assign n510 = ~\req[86]  & ~\req[87]  ;
  assign n511 = ~n509 & n510 ;
  assign n512 = n502 & ~n511 ;
  assign n513 = ~\priority[92]  & \req[91]  ;
  assign n514 = ~\req[92]  & ~\req[93]  ;
  assign n515 = ~n513 & n514 ;
  assign n516 = ~\priority[89]  & \req[88]  ;
  assign n517 = ~\req[89]  & ~\req[90]  ;
  assign n518 = ~n516 & n517 ;
  assign n519 = n515 & n518 ;
  assign n520 = ~n512 & n519 ;
  assign n521 = ~n508 & n520 ;
  assign n522 = \priority[90]  & ~\req[90]  ;
  assign n523 = ~\priority[91]  & ~\priority[92]  ;
  assign n524 = ~n522 & n523 ;
  assign n525 = n515 & ~n524 ;
  assign n526 = \priority[96]  & ~\req[96]  ;
  assign n527 = ~\priority[97]  & ~\priority[98]  ;
  assign n528 = ~n526 & n527 ;
  assign n529 = \priority[93]  & ~\req[93]  ;
  assign n530 = ~\priority[94]  & ~\priority[95]  ;
  assign n531 = ~n529 & n530 ;
  assign n532 = n528 & n531 ;
  assign n533 = ~n525 & n532 ;
  assign n534 = ~n521 & n533 ;
  assign n535 = ~\priority[95]  & \req[94]  ;
  assign n536 = ~\req[95]  & ~\req[96]  ;
  assign n537 = ~n535 & n536 ;
  assign n538 = n528 & ~n537 ;
  assign n539 = ~\priority[101]  & \req[100]  ;
  assign n540 = ~\req[101]  & ~\req[102]  ;
  assign n541 = ~n539 & n540 ;
  assign n542 = ~\priority[98]  & \req[97]  ;
  assign n543 = ~\req[98]  & ~\req[99]  ;
  assign n544 = ~n542 & n543 ;
  assign n545 = n541 & n544 ;
  assign n546 = ~n538 & n545 ;
  assign n547 = ~n534 & n546 ;
  assign n548 = \priority[99]  & ~\req[99]  ;
  assign n549 = ~\priority[100]  & ~\priority[101]  ;
  assign n550 = ~n548 & n549 ;
  assign n551 = n541 & ~n550 ;
  assign n552 = \priority[105]  & ~\req[105]  ;
  assign n553 = ~\priority[106]  & ~\priority[107]  ;
  assign n554 = ~n552 & n553 ;
  assign n555 = \priority[102]  & ~\req[102]  ;
  assign n556 = ~\priority[103]  & ~\priority[104]  ;
  assign n557 = ~n555 & n556 ;
  assign n558 = n554 & n557 ;
  assign n559 = ~n551 & n558 ;
  assign n560 = ~n547 & n559 ;
  assign n561 = ~\priority[104]  & \req[103]  ;
  assign n562 = ~\req[104]  & ~\req[105]  ;
  assign n563 = ~n561 & n562 ;
  assign n564 = n554 & ~n563 ;
  assign n565 = ~\priority[110]  & \req[109]  ;
  assign n566 = ~\req[110]  & ~\req[111]  ;
  assign n567 = ~n565 & n566 ;
  assign n568 = ~\priority[107]  & \req[106]  ;
  assign n569 = ~\req[107]  & ~\req[108]  ;
  assign n570 = ~n568 & n569 ;
  assign n571 = n567 & n570 ;
  assign n572 = ~n564 & n571 ;
  assign n573 = ~n560 & n572 ;
  assign n574 = \priority[108]  & ~\req[108]  ;
  assign n575 = ~\priority[109]  & ~\priority[110]  ;
  assign n576 = ~n574 & n575 ;
  assign n577 = n567 & ~n576 ;
  assign n578 = \priority[114]  & ~\req[114]  ;
  assign n579 = ~\priority[115]  & ~\priority[116]  ;
  assign n580 = ~n578 & n579 ;
  assign n581 = \priority[111]  & ~\req[111]  ;
  assign n582 = ~\priority[112]  & ~\priority[113]  ;
  assign n583 = ~n581 & n582 ;
  assign n584 = n580 & n583 ;
  assign n585 = ~n577 & n584 ;
  assign n586 = ~n573 & n585 ;
  assign n587 = ~\priority[113]  & \req[112]  ;
  assign n588 = ~\req[113]  & ~\req[114]  ;
  assign n589 = ~n587 & n588 ;
  assign n590 = n580 & ~n589 ;
  assign n591 = ~\priority[119]  & \req[118]  ;
  assign n592 = ~\req[119]  & ~\req[120]  ;
  assign n593 = ~n591 & n592 ;
  assign n594 = ~\priority[116]  & \req[115]  ;
  assign n595 = ~\req[116]  & ~\req[117]  ;
  assign n596 = ~n594 & n595 ;
  assign n597 = n593 & n596 ;
  assign n598 = ~n590 & n597 ;
  assign n599 = ~n586 & n598 ;
  assign n600 = \priority[117]  & ~\req[117]  ;
  assign n601 = ~\priority[118]  & ~\priority[119]  ;
  assign n602 = ~n600 & n601 ;
  assign n603 = n593 & ~n602 ;
  assign n604 = \priority[123]  & ~\req[123]  ;
  assign n605 = ~\priority[124]  & ~\priority[125]  ;
  assign n606 = ~n604 & n605 ;
  assign n607 = \priority[120]  & ~\req[120]  ;
  assign n608 = ~\priority[121]  & ~\priority[122]  ;
  assign n609 = ~n607 & n608 ;
  assign n610 = n606 & n609 ;
  assign n611 = ~n603 & n610 ;
  assign n612 = ~n599 & n611 ;
  assign n613 = ~\priority[122]  & \req[121]  ;
  assign n614 = ~\req[122]  & ~\req[123]  ;
  assign n615 = ~n613 & n614 ;
  assign n616 = n606 & ~n615 ;
  assign n617 = ~\priority[125]  & \req[124]  ;
  assign n618 = ~\req[125]  & ~\req[126]  ;
  assign n619 = ~n617 & n618 ;
  assign n620 = n261 & n619 ;
  assign n621 = ~n616 & n620 ;
  assign n622 = ~n612 & n621 ;
  assign n623 = ~n262 & ~n622 ;
  assign n624 = \priority[127]  & ~\req[127]  ;
  assign n625 = ~\priority[0]  & ~\priority[1]  ;
  assign n626 = ~n624 & n625 ;
  assign n627 = ~\priority[1]  & \req[0]  ;
  assign n628 = \req[1]  & ~n627 ;
  assign n629 = ~n626 & n628 ;
  assign n630 = \priority[2]  & ~\req[2]  ;
  assign n631 = ~\priority[3]  & ~n630 ;
  assign n632 = ~\req[3]  & ~\req[4]  ;
  assign n633 = ~n631 & n632 ;
  assign n634 = \priority[7]  & ~\req[7]  ;
  assign n635 = ~\priority[8]  & ~\priority[9]  ;
  assign n636 = ~n634 & n635 ;
  assign n637 = \priority[4]  & ~\req[4]  ;
  assign n638 = ~\priority[5]  & ~\priority[6]  ;
  assign n639 = ~n637 & n638 ;
  assign n640 = n636 & n639 ;
  assign n641 = ~n633 & n640 ;
  assign n642 = ~\priority[6]  & \req[5]  ;
  assign n643 = ~\req[6]  & ~\req[7]  ;
  assign n644 = ~n642 & n643 ;
  assign n645 = n636 & ~n644 ;
  assign n646 = ~\priority[12]  & \req[11]  ;
  assign n647 = ~\req[12]  & ~\req[13]  ;
  assign n648 = ~n646 & n647 ;
  assign n649 = ~\priority[9]  & \req[8]  ;
  assign n650 = ~\req[9]  & ~\req[10]  ;
  assign n651 = ~n649 & n650 ;
  assign n652 = n648 & n651 ;
  assign n653 = ~n645 & n652 ;
  assign n654 = ~n641 & n653 ;
  assign n655 = \priority[10]  & ~\req[10]  ;
  assign n656 = ~\priority[11]  & ~\priority[12]  ;
  assign n657 = ~n655 & n656 ;
  assign n658 = n648 & ~n657 ;
  assign n659 = \priority[16]  & ~\req[16]  ;
  assign n660 = ~\priority[17]  & ~\priority[18]  ;
  assign n661 = ~n659 & n660 ;
  assign n662 = \priority[13]  & ~\req[13]  ;
  assign n663 = ~\priority[14]  & ~\priority[15]  ;
  assign n664 = ~n662 & n663 ;
  assign n665 = n661 & n664 ;
  assign n666 = ~n658 & n665 ;
  assign n667 = ~n654 & n666 ;
  assign n668 = ~\priority[15]  & \req[14]  ;
  assign n669 = ~\req[15]  & ~\req[16]  ;
  assign n670 = ~n668 & n669 ;
  assign n671 = n661 & ~n670 ;
  assign n672 = ~\priority[21]  & \req[20]  ;
  assign n673 = ~\req[21]  & ~\req[22]  ;
  assign n674 = ~n672 & n673 ;
  assign n675 = ~\priority[18]  & \req[17]  ;
  assign n676 = ~\req[18]  & ~\req[19]  ;
  assign n677 = ~n675 & n676 ;
  assign n678 = n674 & n677 ;
  assign n679 = ~n671 & n678 ;
  assign n680 = ~n667 & n679 ;
  assign n681 = \priority[19]  & ~\req[19]  ;
  assign n682 = ~\priority[20]  & ~\priority[21]  ;
  assign n683 = ~n681 & n682 ;
  assign n684 = n674 & ~n683 ;
  assign n685 = \priority[25]  & ~\req[25]  ;
  assign n686 = ~\priority[26]  & ~\priority[27]  ;
  assign n687 = ~n685 & n686 ;
  assign n688 = \priority[22]  & ~\req[22]  ;
  assign n689 = ~\priority[23]  & ~\priority[24]  ;
  assign n690 = ~n688 & n689 ;
  assign n691 = n687 & n690 ;
  assign n692 = ~n684 & n691 ;
  assign n693 = ~n680 & n692 ;
  assign n694 = ~\priority[24]  & \req[23]  ;
  assign n695 = ~\req[24]  & ~\req[25]  ;
  assign n696 = ~n694 & n695 ;
  assign n697 = n687 & ~n696 ;
  assign n698 = ~\priority[30]  & \req[29]  ;
  assign n699 = ~\req[30]  & ~\req[31]  ;
  assign n700 = ~n698 & n699 ;
  assign n701 = ~\priority[27]  & \req[26]  ;
  assign n702 = ~\req[27]  & ~\req[28]  ;
  assign n703 = ~n701 & n702 ;
  assign n704 = n700 & n703 ;
  assign n705 = ~n697 & n704 ;
  assign n706 = ~n693 & n705 ;
  assign n707 = \priority[28]  & ~\req[28]  ;
  assign n708 = ~\priority[29]  & ~\priority[30]  ;
  assign n709 = ~n707 & n708 ;
  assign n710 = n700 & ~n709 ;
  assign n711 = \priority[34]  & ~\req[34]  ;
  assign n712 = ~\priority[35]  & ~\priority[36]  ;
  assign n713 = ~n711 & n712 ;
  assign n714 = \priority[31]  & ~\req[31]  ;
  assign n715 = ~\priority[32]  & ~\priority[33]  ;
  assign n716 = ~n714 & n715 ;
  assign n717 = n713 & n716 ;
  assign n718 = ~n710 & n717 ;
  assign n719 = ~n706 & n718 ;
  assign n720 = ~\priority[33]  & \req[32]  ;
  assign n721 = ~\req[33]  & ~\req[34]  ;
  assign n722 = ~n720 & n721 ;
  assign n723 = n713 & ~n722 ;
  assign n724 = ~\priority[39]  & \req[38]  ;
  assign n725 = ~\req[39]  & ~\req[40]  ;
  assign n726 = ~n724 & n725 ;
  assign n727 = ~\priority[36]  & \req[35]  ;
  assign n728 = ~\req[36]  & ~\req[37]  ;
  assign n729 = ~n727 & n728 ;
  assign n730 = n726 & n729 ;
  assign n731 = ~n723 & n730 ;
  assign n732 = ~n719 & n731 ;
  assign n733 = \priority[37]  & ~\req[37]  ;
  assign n734 = ~\priority[38]  & ~\priority[39]  ;
  assign n735 = ~n733 & n734 ;
  assign n736 = n726 & ~n735 ;
  assign n737 = \priority[43]  & ~\req[43]  ;
  assign n738 = ~\priority[44]  & ~\priority[45]  ;
  assign n739 = ~n737 & n738 ;
  assign n740 = \priority[40]  & ~\req[40]  ;
  assign n741 = ~\priority[41]  & ~\priority[42]  ;
  assign n742 = ~n740 & n741 ;
  assign n743 = n739 & n742 ;
  assign n744 = ~n736 & n743 ;
  assign n745 = ~n732 & n744 ;
  assign n746 = ~\priority[42]  & \req[41]  ;
  assign n747 = ~\req[42]  & ~\req[43]  ;
  assign n748 = ~n746 & n747 ;
  assign n749 = n739 & ~n748 ;
  assign n750 = ~\priority[48]  & \req[47]  ;
  assign n751 = ~\req[48]  & ~\req[49]  ;
  assign n752 = ~n750 & n751 ;
  assign n753 = ~\priority[45]  & \req[44]  ;
  assign n754 = ~\req[45]  & ~\req[46]  ;
  assign n755 = ~n753 & n754 ;
  assign n756 = n752 & n755 ;
  assign n757 = ~n749 & n756 ;
  assign n758 = ~n745 & n757 ;
  assign n759 = \priority[46]  & ~\req[46]  ;
  assign n760 = ~\priority[47]  & ~\priority[48]  ;
  assign n761 = ~n759 & n760 ;
  assign n762 = n752 & ~n761 ;
  assign n763 = \priority[52]  & ~\req[52]  ;
  assign n764 = ~\priority[53]  & ~\priority[54]  ;
  assign n765 = ~n763 & n764 ;
  assign n766 = \priority[49]  & ~\req[49]  ;
  assign n767 = ~\priority[50]  & ~\priority[51]  ;
  assign n768 = ~n766 & n767 ;
  assign n769 = n765 & n768 ;
  assign n770 = ~n762 & n769 ;
  assign n771 = ~n758 & n770 ;
  assign n772 = ~\priority[51]  & \req[50]  ;
  assign n773 = ~\req[51]  & ~\req[52]  ;
  assign n774 = ~n772 & n773 ;
  assign n775 = n765 & ~n774 ;
  assign n776 = ~\priority[57]  & \req[56]  ;
  assign n777 = ~\req[57]  & ~\req[58]  ;
  assign n778 = ~n776 & n777 ;
  assign n779 = ~\priority[54]  & \req[53]  ;
  assign n780 = ~\req[54]  & ~\req[55]  ;
  assign n781 = ~n779 & n780 ;
  assign n782 = n778 & n781 ;
  assign n783 = ~n775 & n782 ;
  assign n784 = ~n771 & n783 ;
  assign n785 = \priority[55]  & ~\req[55]  ;
  assign n786 = ~\priority[56]  & ~\priority[57]  ;
  assign n787 = ~n785 & n786 ;
  assign n788 = n778 & ~n787 ;
  assign n789 = \priority[61]  & ~\req[61]  ;
  assign n790 = ~\priority[62]  & ~\priority[63]  ;
  assign n791 = ~n789 & n790 ;
  assign n792 = \priority[58]  & ~\req[58]  ;
  assign n793 = ~\priority[59]  & ~\priority[60]  ;
  assign n794 = ~n792 & n793 ;
  assign n795 = n791 & n794 ;
  assign n796 = ~n788 & n795 ;
  assign n797 = ~n784 & n796 ;
  assign n798 = ~\priority[60]  & \req[59]  ;
  assign n799 = ~\req[60]  & ~\req[61]  ;
  assign n800 = ~n798 & n799 ;
  assign n801 = n791 & ~n800 ;
  assign n802 = ~\priority[66]  & \req[65]  ;
  assign n803 = ~\req[66]  & ~\req[67]  ;
  assign n804 = ~n802 & n803 ;
  assign n805 = ~\priority[63]  & \req[62]  ;
  assign n806 = ~\req[63]  & ~\req[64]  ;
  assign n807 = ~n805 & n806 ;
  assign n808 = n804 & n807 ;
  assign n809 = ~n801 & n808 ;
  assign n810 = ~n797 & n809 ;
  assign n811 = \priority[64]  & ~\req[64]  ;
  assign n812 = ~\priority[65]  & ~\priority[66]  ;
  assign n813 = ~n811 & n812 ;
  assign n814 = n804 & ~n813 ;
  assign n815 = \priority[70]  & ~\req[70]  ;
  assign n816 = ~\priority[71]  & ~\priority[72]  ;
  assign n817 = ~n815 & n816 ;
  assign n818 = \priority[67]  & ~\req[67]  ;
  assign n819 = ~\priority[68]  & ~\priority[69]  ;
  assign n820 = ~n818 & n819 ;
  assign n821 = n817 & n820 ;
  assign n822 = ~n814 & n821 ;
  assign n823 = ~n810 & n822 ;
  assign n824 = ~\priority[69]  & \req[68]  ;
  assign n825 = ~\req[69]  & ~\req[70]  ;
  assign n826 = ~n824 & n825 ;
  assign n827 = n817 & ~n826 ;
  assign n828 = ~\priority[75]  & \req[74]  ;
  assign n829 = ~\req[75]  & ~\req[76]  ;
  assign n830 = ~n828 & n829 ;
  assign n831 = ~\priority[72]  & \req[71]  ;
  assign n832 = ~\req[72]  & ~\req[73]  ;
  assign n833 = ~n831 & n832 ;
  assign n834 = n830 & n833 ;
  assign n835 = ~n827 & n834 ;
  assign n836 = ~n823 & n835 ;
  assign n837 = \priority[73]  & ~\req[73]  ;
  assign n838 = ~\priority[74]  & ~\priority[75]  ;
  assign n839 = ~n837 & n838 ;
  assign n840 = n830 & ~n839 ;
  assign n841 = \priority[79]  & ~\req[79]  ;
  assign n842 = ~\priority[80]  & ~\priority[81]  ;
  assign n843 = ~n841 & n842 ;
  assign n844 = \priority[76]  & ~\req[76]  ;
  assign n845 = ~\priority[77]  & ~\priority[78]  ;
  assign n846 = ~n844 & n845 ;
  assign n847 = n843 & n846 ;
  assign n848 = ~n840 & n847 ;
  assign n849 = ~n836 & n848 ;
  assign n850 = ~\priority[78]  & \req[77]  ;
  assign n851 = ~\req[78]  & ~\req[79]  ;
  assign n852 = ~n850 & n851 ;
  assign n853 = n843 & ~n852 ;
  assign n854 = ~\priority[84]  & \req[83]  ;
  assign n855 = ~\req[84]  & ~\req[85]  ;
  assign n856 = ~n854 & n855 ;
  assign n857 = ~\priority[81]  & \req[80]  ;
  assign n858 = ~\req[81]  & ~\req[82]  ;
  assign n859 = ~n857 & n858 ;
  assign n860 = n856 & n859 ;
  assign n861 = ~n853 & n860 ;
  assign n862 = ~n849 & n861 ;
  assign n863 = \priority[82]  & ~\req[82]  ;
  assign n864 = ~\priority[83]  & ~\priority[84]  ;
  assign n865 = ~n863 & n864 ;
  assign n866 = n856 & ~n865 ;
  assign n867 = \priority[88]  & ~\req[88]  ;
  assign n868 = ~\priority[89]  & ~\priority[90]  ;
  assign n869 = ~n867 & n868 ;
  assign n870 = \priority[85]  & ~\req[85]  ;
  assign n871 = ~\priority[86]  & ~\priority[87]  ;
  assign n872 = ~n870 & n871 ;
  assign n873 = n869 & n872 ;
  assign n874 = ~n866 & n873 ;
  assign n875 = ~n862 & n874 ;
  assign n876 = ~\priority[87]  & \req[86]  ;
  assign n877 = ~\req[87]  & ~\req[88]  ;
  assign n878 = ~n876 & n877 ;
  assign n879 = n869 & ~n878 ;
  assign n880 = ~\priority[93]  & \req[92]  ;
  assign n881 = ~\req[93]  & ~\req[94]  ;
  assign n882 = ~n880 & n881 ;
  assign n883 = ~\priority[90]  & \req[89]  ;
  assign n884 = ~\req[90]  & ~\req[91]  ;
  assign n885 = ~n883 & n884 ;
  assign n886 = n882 & n885 ;
  assign n887 = ~n879 & n886 ;
  assign n888 = ~n875 & n887 ;
  assign n889 = \priority[91]  & ~\req[91]  ;
  assign n890 = ~\priority[92]  & ~\priority[93]  ;
  assign n891 = ~n889 & n890 ;
  assign n892 = n882 & ~n891 ;
  assign n893 = \priority[97]  & ~\req[97]  ;
  assign n894 = ~\priority[98]  & ~\priority[99]  ;
  assign n895 = ~n893 & n894 ;
  assign n896 = \priority[94]  & ~\req[94]  ;
  assign n897 = ~\priority[95]  & ~\priority[96]  ;
  assign n898 = ~n896 & n897 ;
  assign n899 = n895 & n898 ;
  assign n900 = ~n892 & n899 ;
  assign n901 = ~n888 & n900 ;
  assign n902 = ~\priority[96]  & \req[95]  ;
  assign n903 = ~\req[96]  & ~\req[97]  ;
  assign n904 = ~n902 & n903 ;
  assign n905 = n895 & ~n904 ;
  assign n906 = ~\priority[102]  & \req[101]  ;
  assign n907 = ~\req[102]  & ~\req[103]  ;
  assign n908 = ~n906 & n907 ;
  assign n909 = ~\priority[99]  & \req[98]  ;
  assign n910 = ~\req[99]  & ~\req[100]  ;
  assign n911 = ~n909 & n910 ;
  assign n912 = n908 & n911 ;
  assign n913 = ~n905 & n912 ;
  assign n914 = ~n901 & n913 ;
  assign n915 = \priority[100]  & ~\req[100]  ;
  assign n916 = ~\priority[101]  & ~\priority[102]  ;
  assign n917 = ~n915 & n916 ;
  assign n918 = n908 & ~n917 ;
  assign n919 = \priority[106]  & ~\req[106]  ;
  assign n920 = ~\priority[107]  & ~\priority[108]  ;
  assign n921 = ~n919 & n920 ;
  assign n922 = \priority[103]  & ~\req[103]  ;
  assign n923 = ~\priority[104]  & ~\priority[105]  ;
  assign n924 = ~n922 & n923 ;
  assign n925 = n921 & n924 ;
  assign n926 = ~n918 & n925 ;
  assign n927 = ~n914 & n926 ;
  assign n928 = ~\priority[105]  & \req[104]  ;
  assign n929 = ~\req[105]  & ~\req[106]  ;
  assign n930 = ~n928 & n929 ;
  assign n931 = n921 & ~n930 ;
  assign n932 = ~\priority[111]  & \req[110]  ;
  assign n933 = ~\req[111]  & ~\req[112]  ;
  assign n934 = ~n932 & n933 ;
  assign n935 = ~\priority[108]  & \req[107]  ;
  assign n936 = ~\req[108]  & ~\req[109]  ;
  assign n937 = ~n935 & n936 ;
  assign n938 = n934 & n937 ;
  assign n939 = ~n931 & n938 ;
  assign n940 = ~n927 & n939 ;
  assign n941 = \priority[109]  & ~\req[109]  ;
  assign n942 = ~\priority[110]  & ~\priority[111]  ;
  assign n943 = ~n941 & n942 ;
  assign n944 = n934 & ~n943 ;
  assign n945 = \priority[115]  & ~\req[115]  ;
  assign n946 = ~\priority[116]  & ~\priority[117]  ;
  assign n947 = ~n945 & n946 ;
  assign n948 = \priority[112]  & ~\req[112]  ;
  assign n949 = ~\priority[113]  & ~\priority[114]  ;
  assign n950 = ~n948 & n949 ;
  assign n951 = n947 & n950 ;
  assign n952 = ~n944 & n951 ;
  assign n953 = ~n940 & n952 ;
  assign n954 = ~\priority[114]  & \req[113]  ;
  assign n955 = ~\req[114]  & ~\req[115]  ;
  assign n956 = ~n954 & n955 ;
  assign n957 = n947 & ~n956 ;
  assign n958 = ~\priority[120]  & \req[119]  ;
  assign n959 = ~\req[120]  & ~\req[121]  ;
  assign n960 = ~n958 & n959 ;
  assign n961 = ~\priority[117]  & \req[116]  ;
  assign n962 = ~\req[117]  & ~\req[118]  ;
  assign n963 = ~n961 & n962 ;
  assign n964 = n960 & n963 ;
  assign n965 = ~n957 & n964 ;
  assign n966 = ~n953 & n965 ;
  assign n967 = \priority[118]  & ~\req[118]  ;
  assign n968 = ~\priority[119]  & ~\priority[120]  ;
  assign n969 = ~n967 & n968 ;
  assign n970 = n960 & ~n969 ;
  assign n971 = \priority[124]  & ~\req[124]  ;
  assign n972 = ~\priority[125]  & ~\priority[126]  ;
  assign n973 = ~n971 & n972 ;
  assign n974 = \priority[121]  & ~\req[121]  ;
  assign n975 = ~\priority[122]  & ~\priority[123]  ;
  assign n976 = ~n974 & n975 ;
  assign n977 = n973 & n976 ;
  assign n978 = ~n970 & n977 ;
  assign n979 = ~n966 & n978 ;
  assign n980 = ~\priority[123]  & \req[122]  ;
  assign n981 = ~\req[123]  & ~\req[124]  ;
  assign n982 = ~n980 & n981 ;
  assign n983 = n973 & ~n982 ;
  assign n984 = ~\priority[126]  & \req[125]  ;
  assign n985 = ~\req[126]  & ~\req[127]  ;
  assign n986 = ~n984 & n985 ;
  assign n987 = n628 & n986 ;
  assign n988 = ~n983 & n987 ;
  assign n989 = ~n979 & n988 ;
  assign n990 = ~n629 & ~n989 ;
  assign n991 = \priority[0]  & ~\req[0]  ;
  assign n992 = ~\priority[1]  & ~\priority[2]  ;
  assign n993 = ~n991 & n992 ;
  assign n994 = ~\priority[2]  & \req[1]  ;
  assign n995 = \req[2]  & ~n994 ;
  assign n996 = ~n993 & n995 ;
  assign n997 = ~\priority[4]  & ~n270 ;
  assign n998 = ~\req[4]  & ~\req[5]  ;
  assign n999 = ~n997 & n998 ;
  assign n1000 = \priority[8]  & ~\req[8]  ;
  assign n1001 = ~\priority[9]  & ~\priority[10]  ;
  assign n1002 = ~n1000 & n1001 ;
  assign n1003 = \priority[5]  & ~\req[5]  ;
  assign n1004 = ~\priority[6]  & ~\priority[7]  ;
  assign n1005 = ~n1003 & n1004 ;
  assign n1006 = n1002 & n1005 ;
  assign n1007 = ~n999 & n1006 ;
  assign n1008 = ~\priority[7]  & \req[6]  ;
  assign n1009 = ~\req[7]  & ~\req[8]  ;
  assign n1010 = ~n1008 & n1009 ;
  assign n1011 = n1002 & ~n1010 ;
  assign n1012 = ~\priority[13]  & \req[12]  ;
  assign n1013 = ~\req[13]  & ~\req[14]  ;
  assign n1014 = ~n1012 & n1013 ;
  assign n1015 = ~\priority[10]  & \req[9]  ;
  assign n1016 = ~\req[10]  & ~\req[11]  ;
  assign n1017 = ~n1015 & n1016 ;
  assign n1018 = n1014 & n1017 ;
  assign n1019 = ~n1011 & n1018 ;
  assign n1020 = ~n1007 & n1019 ;
  assign n1021 = \priority[11]  & ~\req[11]  ;
  assign n1022 = ~\priority[12]  & ~\priority[13]  ;
  assign n1023 = ~n1021 & n1022 ;
  assign n1024 = n1014 & ~n1023 ;
  assign n1025 = \priority[17]  & ~\req[17]  ;
  assign n1026 = ~\priority[18]  & ~\priority[19]  ;
  assign n1027 = ~n1025 & n1026 ;
  assign n1028 = \priority[14]  & ~\req[14]  ;
  assign n1029 = ~\priority[15]  & ~\priority[16]  ;
  assign n1030 = ~n1028 & n1029 ;
  assign n1031 = n1027 & n1030 ;
  assign n1032 = ~n1024 & n1031 ;
  assign n1033 = ~n1020 & n1032 ;
  assign n1034 = ~\priority[16]  & \req[15]  ;
  assign n1035 = ~\req[16]  & ~\req[17]  ;
  assign n1036 = ~n1034 & n1035 ;
  assign n1037 = n1027 & ~n1036 ;
  assign n1038 = ~\priority[22]  & \req[21]  ;
  assign n1039 = ~\req[22]  & ~\req[23]  ;
  assign n1040 = ~n1038 & n1039 ;
  assign n1041 = ~\priority[19]  & \req[18]  ;
  assign n1042 = ~\req[19]  & ~\req[20]  ;
  assign n1043 = ~n1041 & n1042 ;
  assign n1044 = n1040 & n1043 ;
  assign n1045 = ~n1037 & n1044 ;
  assign n1046 = ~n1033 & n1045 ;
  assign n1047 = \priority[20]  & ~\req[20]  ;
  assign n1048 = ~\priority[21]  & ~\priority[22]  ;
  assign n1049 = ~n1047 & n1048 ;
  assign n1050 = n1040 & ~n1049 ;
  assign n1051 = \priority[26]  & ~\req[26]  ;
  assign n1052 = ~\priority[27]  & ~\priority[28]  ;
  assign n1053 = ~n1051 & n1052 ;
  assign n1054 = \priority[23]  & ~\req[23]  ;
  assign n1055 = ~\priority[24]  & ~\priority[25]  ;
  assign n1056 = ~n1054 & n1055 ;
  assign n1057 = n1053 & n1056 ;
  assign n1058 = ~n1050 & n1057 ;
  assign n1059 = ~n1046 & n1058 ;
  assign n1060 = ~\priority[25]  & \req[24]  ;
  assign n1061 = ~\req[25]  & ~\req[26]  ;
  assign n1062 = ~n1060 & n1061 ;
  assign n1063 = n1053 & ~n1062 ;
  assign n1064 = ~\priority[31]  & \req[30]  ;
  assign n1065 = ~\req[31]  & ~\req[32]  ;
  assign n1066 = ~n1064 & n1065 ;
  assign n1067 = ~\priority[28]  & \req[27]  ;
  assign n1068 = ~\req[28]  & ~\req[29]  ;
  assign n1069 = ~n1067 & n1068 ;
  assign n1070 = n1066 & n1069 ;
  assign n1071 = ~n1063 & n1070 ;
  assign n1072 = ~n1059 & n1071 ;
  assign n1073 = \priority[29]  & ~\req[29]  ;
  assign n1074 = ~\priority[30]  & ~\priority[31]  ;
  assign n1075 = ~n1073 & n1074 ;
  assign n1076 = n1066 & ~n1075 ;
  assign n1077 = \priority[35]  & ~\req[35]  ;
  assign n1078 = ~\priority[36]  & ~\priority[37]  ;
  assign n1079 = ~n1077 & n1078 ;
  assign n1080 = \priority[32]  & ~\req[32]  ;
  assign n1081 = ~\priority[33]  & ~\priority[34]  ;
  assign n1082 = ~n1080 & n1081 ;
  assign n1083 = n1079 & n1082 ;
  assign n1084 = ~n1076 & n1083 ;
  assign n1085 = ~n1072 & n1084 ;
  assign n1086 = ~\priority[34]  & \req[33]  ;
  assign n1087 = ~\req[34]  & ~\req[35]  ;
  assign n1088 = ~n1086 & n1087 ;
  assign n1089 = n1079 & ~n1088 ;
  assign n1090 = ~\priority[40]  & \req[39]  ;
  assign n1091 = ~\req[40]  & ~\req[41]  ;
  assign n1092 = ~n1090 & n1091 ;
  assign n1093 = ~\priority[37]  & \req[36]  ;
  assign n1094 = ~\req[37]  & ~\req[38]  ;
  assign n1095 = ~n1093 & n1094 ;
  assign n1096 = n1092 & n1095 ;
  assign n1097 = ~n1089 & n1096 ;
  assign n1098 = ~n1085 & n1097 ;
  assign n1099 = \priority[38]  & ~\req[38]  ;
  assign n1100 = ~\priority[39]  & ~\priority[40]  ;
  assign n1101 = ~n1099 & n1100 ;
  assign n1102 = n1092 & ~n1101 ;
  assign n1103 = \priority[44]  & ~\req[44]  ;
  assign n1104 = ~\priority[45]  & ~\priority[46]  ;
  assign n1105 = ~n1103 & n1104 ;
  assign n1106 = \priority[41]  & ~\req[41]  ;
  assign n1107 = ~\priority[42]  & ~\priority[43]  ;
  assign n1108 = ~n1106 & n1107 ;
  assign n1109 = n1105 & n1108 ;
  assign n1110 = ~n1102 & n1109 ;
  assign n1111 = ~n1098 & n1110 ;
  assign n1112 = ~\priority[43]  & \req[42]  ;
  assign n1113 = ~\req[43]  & ~\req[44]  ;
  assign n1114 = ~n1112 & n1113 ;
  assign n1115 = n1105 & ~n1114 ;
  assign n1116 = ~\priority[49]  & \req[48]  ;
  assign n1117 = ~\req[49]  & ~\req[50]  ;
  assign n1118 = ~n1116 & n1117 ;
  assign n1119 = ~\priority[46]  & \req[45]  ;
  assign n1120 = ~\req[46]  & ~\req[47]  ;
  assign n1121 = ~n1119 & n1120 ;
  assign n1122 = n1118 & n1121 ;
  assign n1123 = ~n1115 & n1122 ;
  assign n1124 = ~n1111 & n1123 ;
  assign n1125 = \priority[47]  & ~\req[47]  ;
  assign n1126 = ~\priority[48]  & ~\priority[49]  ;
  assign n1127 = ~n1125 & n1126 ;
  assign n1128 = n1118 & ~n1127 ;
  assign n1129 = \priority[53]  & ~\req[53]  ;
  assign n1130 = ~\priority[54]  & ~\priority[55]  ;
  assign n1131 = ~n1129 & n1130 ;
  assign n1132 = \priority[50]  & ~\req[50]  ;
  assign n1133 = ~\priority[51]  & ~\priority[52]  ;
  assign n1134 = ~n1132 & n1133 ;
  assign n1135 = n1131 & n1134 ;
  assign n1136 = ~n1128 & n1135 ;
  assign n1137 = ~n1124 & n1136 ;
  assign n1138 = ~\priority[52]  & \req[51]  ;
  assign n1139 = ~\req[52]  & ~\req[53]  ;
  assign n1140 = ~n1138 & n1139 ;
  assign n1141 = n1131 & ~n1140 ;
  assign n1142 = ~\priority[58]  & \req[57]  ;
  assign n1143 = ~\req[58]  & ~\req[59]  ;
  assign n1144 = ~n1142 & n1143 ;
  assign n1145 = ~\priority[55]  & \req[54]  ;
  assign n1146 = ~\req[55]  & ~\req[56]  ;
  assign n1147 = ~n1145 & n1146 ;
  assign n1148 = n1144 & n1147 ;
  assign n1149 = ~n1141 & n1148 ;
  assign n1150 = ~n1137 & n1149 ;
  assign n1151 = \priority[56]  & ~\req[56]  ;
  assign n1152 = ~\priority[57]  & ~\priority[58]  ;
  assign n1153 = ~n1151 & n1152 ;
  assign n1154 = n1144 & ~n1153 ;
  assign n1155 = \priority[62]  & ~\req[62]  ;
  assign n1156 = ~\priority[63]  & ~\priority[64]  ;
  assign n1157 = ~n1155 & n1156 ;
  assign n1158 = \priority[59]  & ~\req[59]  ;
  assign n1159 = ~\priority[60]  & ~\priority[61]  ;
  assign n1160 = ~n1158 & n1159 ;
  assign n1161 = n1157 & n1160 ;
  assign n1162 = ~n1154 & n1161 ;
  assign n1163 = ~n1150 & n1162 ;
  assign n1164 = ~\priority[61]  & \req[60]  ;
  assign n1165 = ~\req[61]  & ~\req[62]  ;
  assign n1166 = ~n1164 & n1165 ;
  assign n1167 = n1157 & ~n1166 ;
  assign n1168 = ~\priority[67]  & \req[66]  ;
  assign n1169 = ~\req[67]  & ~\req[68]  ;
  assign n1170 = ~n1168 & n1169 ;
  assign n1171 = ~\priority[64]  & \req[63]  ;
  assign n1172 = ~\req[64]  & ~\req[65]  ;
  assign n1173 = ~n1171 & n1172 ;
  assign n1174 = n1170 & n1173 ;
  assign n1175 = ~n1167 & n1174 ;
  assign n1176 = ~n1163 & n1175 ;
  assign n1177 = \priority[65]  & ~\req[65]  ;
  assign n1178 = ~\priority[66]  & ~\priority[67]  ;
  assign n1179 = ~n1177 & n1178 ;
  assign n1180 = n1170 & ~n1179 ;
  assign n1181 = \priority[71]  & ~\req[71]  ;
  assign n1182 = ~\priority[72]  & ~\priority[73]  ;
  assign n1183 = ~n1181 & n1182 ;
  assign n1184 = \priority[68]  & ~\req[68]  ;
  assign n1185 = ~\priority[69]  & ~\priority[70]  ;
  assign n1186 = ~n1184 & n1185 ;
  assign n1187 = n1183 & n1186 ;
  assign n1188 = ~n1180 & n1187 ;
  assign n1189 = ~n1176 & n1188 ;
  assign n1190 = ~\priority[70]  & \req[69]  ;
  assign n1191 = ~\req[70]  & ~\req[71]  ;
  assign n1192 = ~n1190 & n1191 ;
  assign n1193 = n1183 & ~n1192 ;
  assign n1194 = ~\priority[76]  & \req[75]  ;
  assign n1195 = ~\req[76]  & ~\req[77]  ;
  assign n1196 = ~n1194 & n1195 ;
  assign n1197 = ~\priority[73]  & \req[72]  ;
  assign n1198 = ~\req[73]  & ~\req[74]  ;
  assign n1199 = ~n1197 & n1198 ;
  assign n1200 = n1196 & n1199 ;
  assign n1201 = ~n1193 & n1200 ;
  assign n1202 = ~n1189 & n1201 ;
  assign n1203 = \priority[74]  & ~\req[74]  ;
  assign n1204 = ~\priority[75]  & ~\priority[76]  ;
  assign n1205 = ~n1203 & n1204 ;
  assign n1206 = n1196 & ~n1205 ;
  assign n1207 = \priority[80]  & ~\req[80]  ;
  assign n1208 = ~\priority[81]  & ~\priority[82]  ;
  assign n1209 = ~n1207 & n1208 ;
  assign n1210 = \priority[77]  & ~\req[77]  ;
  assign n1211 = ~\priority[78]  & ~\priority[79]  ;
  assign n1212 = ~n1210 & n1211 ;
  assign n1213 = n1209 & n1212 ;
  assign n1214 = ~n1206 & n1213 ;
  assign n1215 = ~n1202 & n1214 ;
  assign n1216 = ~\priority[79]  & \req[78]  ;
  assign n1217 = ~\req[79]  & ~\req[80]  ;
  assign n1218 = ~n1216 & n1217 ;
  assign n1219 = n1209 & ~n1218 ;
  assign n1220 = ~\priority[85]  & \req[84]  ;
  assign n1221 = ~\req[85]  & ~\req[86]  ;
  assign n1222 = ~n1220 & n1221 ;
  assign n1223 = ~\priority[82]  & \req[81]  ;
  assign n1224 = ~\req[82]  & ~\req[83]  ;
  assign n1225 = ~n1223 & n1224 ;
  assign n1226 = n1222 & n1225 ;
  assign n1227 = ~n1219 & n1226 ;
  assign n1228 = ~n1215 & n1227 ;
  assign n1229 = \priority[83]  & ~\req[83]  ;
  assign n1230 = ~\priority[84]  & ~\priority[85]  ;
  assign n1231 = ~n1229 & n1230 ;
  assign n1232 = n1222 & ~n1231 ;
  assign n1233 = \priority[89]  & ~\req[89]  ;
  assign n1234 = ~\priority[90]  & ~\priority[91]  ;
  assign n1235 = ~n1233 & n1234 ;
  assign n1236 = \priority[86]  & ~\req[86]  ;
  assign n1237 = ~\priority[87]  & ~\priority[88]  ;
  assign n1238 = ~n1236 & n1237 ;
  assign n1239 = n1235 & n1238 ;
  assign n1240 = ~n1232 & n1239 ;
  assign n1241 = ~n1228 & n1240 ;
  assign n1242 = ~\priority[88]  & \req[87]  ;
  assign n1243 = ~\req[88]  & ~\req[89]  ;
  assign n1244 = ~n1242 & n1243 ;
  assign n1245 = n1235 & ~n1244 ;
  assign n1246 = ~\priority[94]  & \req[93]  ;
  assign n1247 = ~\req[94]  & ~\req[95]  ;
  assign n1248 = ~n1246 & n1247 ;
  assign n1249 = ~\priority[91]  & \req[90]  ;
  assign n1250 = ~\req[91]  & ~\req[92]  ;
  assign n1251 = ~n1249 & n1250 ;
  assign n1252 = n1248 & n1251 ;
  assign n1253 = ~n1245 & n1252 ;
  assign n1254 = ~n1241 & n1253 ;
  assign n1255 = \priority[92]  & ~\req[92]  ;
  assign n1256 = ~\priority[93]  & ~\priority[94]  ;
  assign n1257 = ~n1255 & n1256 ;
  assign n1258 = n1248 & ~n1257 ;
  assign n1259 = \priority[98]  & ~\req[98]  ;
  assign n1260 = ~\priority[99]  & ~\priority[100]  ;
  assign n1261 = ~n1259 & n1260 ;
  assign n1262 = \priority[95]  & ~\req[95]  ;
  assign n1263 = ~\priority[96]  & ~\priority[97]  ;
  assign n1264 = ~n1262 & n1263 ;
  assign n1265 = n1261 & n1264 ;
  assign n1266 = ~n1258 & n1265 ;
  assign n1267 = ~n1254 & n1266 ;
  assign n1268 = ~\priority[97]  & \req[96]  ;
  assign n1269 = ~\req[97]  & ~\req[98]  ;
  assign n1270 = ~n1268 & n1269 ;
  assign n1271 = n1261 & ~n1270 ;
  assign n1272 = ~\priority[103]  & \req[102]  ;
  assign n1273 = ~\req[103]  & ~\req[104]  ;
  assign n1274 = ~n1272 & n1273 ;
  assign n1275 = ~\priority[100]  & \req[99]  ;
  assign n1276 = ~\req[100]  & ~\req[101]  ;
  assign n1277 = ~n1275 & n1276 ;
  assign n1278 = n1274 & n1277 ;
  assign n1279 = ~n1271 & n1278 ;
  assign n1280 = ~n1267 & n1279 ;
  assign n1281 = \priority[101]  & ~\req[101]  ;
  assign n1282 = ~\priority[102]  & ~\priority[103]  ;
  assign n1283 = ~n1281 & n1282 ;
  assign n1284 = n1274 & ~n1283 ;
  assign n1285 = \priority[107]  & ~\req[107]  ;
  assign n1286 = ~\priority[108]  & ~\priority[109]  ;
  assign n1287 = ~n1285 & n1286 ;
  assign n1288 = \priority[104]  & ~\req[104]  ;
  assign n1289 = ~\priority[105]  & ~\priority[106]  ;
  assign n1290 = ~n1288 & n1289 ;
  assign n1291 = n1287 & n1290 ;
  assign n1292 = ~n1284 & n1291 ;
  assign n1293 = ~n1280 & n1292 ;
  assign n1294 = ~\priority[106]  & \req[105]  ;
  assign n1295 = ~\req[106]  & ~\req[107]  ;
  assign n1296 = ~n1294 & n1295 ;
  assign n1297 = n1287 & ~n1296 ;
  assign n1298 = ~\priority[112]  & \req[111]  ;
  assign n1299 = ~\req[112]  & ~\req[113]  ;
  assign n1300 = ~n1298 & n1299 ;
  assign n1301 = ~\priority[109]  & \req[108]  ;
  assign n1302 = ~\req[109]  & ~\req[110]  ;
  assign n1303 = ~n1301 & n1302 ;
  assign n1304 = n1300 & n1303 ;
  assign n1305 = ~n1297 & n1304 ;
  assign n1306 = ~n1293 & n1305 ;
  assign n1307 = \priority[110]  & ~\req[110]  ;
  assign n1308 = ~\priority[111]  & ~\priority[112]  ;
  assign n1309 = ~n1307 & n1308 ;
  assign n1310 = n1300 & ~n1309 ;
  assign n1311 = \priority[116]  & ~\req[116]  ;
  assign n1312 = ~\priority[117]  & ~\priority[118]  ;
  assign n1313 = ~n1311 & n1312 ;
  assign n1314 = \priority[113]  & ~\req[113]  ;
  assign n1315 = ~\priority[114]  & ~\priority[115]  ;
  assign n1316 = ~n1314 & n1315 ;
  assign n1317 = n1313 & n1316 ;
  assign n1318 = ~n1310 & n1317 ;
  assign n1319 = ~n1306 & n1318 ;
  assign n1320 = ~\priority[115]  & \req[114]  ;
  assign n1321 = ~\req[115]  & ~\req[116]  ;
  assign n1322 = ~n1320 & n1321 ;
  assign n1323 = n1313 & ~n1322 ;
  assign n1324 = ~\priority[121]  & \req[120]  ;
  assign n1325 = ~\req[121]  & ~\req[122]  ;
  assign n1326 = ~n1324 & n1325 ;
  assign n1327 = ~\priority[118]  & \req[117]  ;
  assign n1328 = ~\req[118]  & ~\req[119]  ;
  assign n1329 = ~n1327 & n1328 ;
  assign n1330 = n1326 & n1329 ;
  assign n1331 = ~n1323 & n1330 ;
  assign n1332 = ~n1319 & n1331 ;
  assign n1333 = \priority[119]  & ~\req[119]  ;
  assign n1334 = ~\priority[120]  & ~\priority[121]  ;
  assign n1335 = ~n1333 & n1334 ;
  assign n1336 = n1326 & ~n1335 ;
  assign n1337 = \priority[125]  & ~\req[125]  ;
  assign n1338 = ~\priority[126]  & ~\priority[127]  ;
  assign n1339 = ~n1337 & n1338 ;
  assign n1340 = \priority[122]  & ~\req[122]  ;
  assign n1341 = ~\priority[123]  & ~\priority[124]  ;
  assign n1342 = ~n1340 & n1341 ;
  assign n1343 = n1339 & n1342 ;
  assign n1344 = ~n1336 & n1343 ;
  assign n1345 = ~n1332 & n1344 ;
  assign n1346 = ~\priority[124]  & \req[123]  ;
  assign n1347 = ~\req[124]  & ~\req[125]  ;
  assign n1348 = ~n1346 & n1347 ;
  assign n1349 = n1339 & ~n1348 ;
  assign n1350 = ~\priority[127]  & \req[126]  ;
  assign n1351 = ~\req[0]  & ~\req[127]  ;
  assign n1352 = ~n1350 & n1351 ;
  assign n1353 = n995 & n1352 ;
  assign n1354 = ~n1349 & n1353 ;
  assign n1355 = ~n1345 & n1354 ;
  assign n1356 = ~n996 & ~n1355 ;
  assign n1357 = ~\priority[2]  & ~\priority[3]  ;
  assign n1358 = ~n263 & n1357 ;
  assign n1359 = ~\priority[3]  & \req[2]  ;
  assign n1360 = \req[3]  & ~n1359 ;
  assign n1361 = ~n1358 & n1360 ;
  assign n1362 = ~\priority[5]  & ~n637 ;
  assign n1363 = n276 & ~n1362 ;
  assign n1364 = n269 & n290 ;
  assign n1365 = ~n1363 & n1364 ;
  assign n1366 = ~n284 & n290 ;
  assign n1367 = n281 & n303 ;
  assign n1368 = ~n1366 & n1367 ;
  assign n1369 = ~n1365 & n1368 ;
  assign n1370 = ~n297 & n303 ;
  assign n1371 = n294 & n316 ;
  assign n1372 = ~n1370 & n1371 ;
  assign n1373 = ~n1369 & n1372 ;
  assign n1374 = ~n310 & n316 ;
  assign n1375 = n307 & n329 ;
  assign n1376 = ~n1374 & n1375 ;
  assign n1377 = ~n1373 & n1376 ;
  assign n1378 = ~n323 & n329 ;
  assign n1379 = n320 & n342 ;
  assign n1380 = ~n1378 & n1379 ;
  assign n1381 = ~n1377 & n1380 ;
  assign n1382 = ~n336 & n342 ;
  assign n1383 = n333 & n355 ;
  assign n1384 = ~n1382 & n1383 ;
  assign n1385 = ~n1381 & n1384 ;
  assign n1386 = ~n349 & n355 ;
  assign n1387 = n346 & n368 ;
  assign n1388 = ~n1386 & n1387 ;
  assign n1389 = ~n1385 & n1388 ;
  assign n1390 = ~n362 & n368 ;
  assign n1391 = n359 & n381 ;
  assign n1392 = ~n1390 & n1391 ;
  assign n1393 = ~n1389 & n1392 ;
  assign n1394 = ~n375 & n381 ;
  assign n1395 = n372 & n394 ;
  assign n1396 = ~n1394 & n1395 ;
  assign n1397 = ~n1393 & n1396 ;
  assign n1398 = ~n388 & n394 ;
  assign n1399 = n385 & n407 ;
  assign n1400 = ~n1398 & n1399 ;
  assign n1401 = ~n1397 & n1400 ;
  assign n1402 = ~n401 & n407 ;
  assign n1403 = n398 & n420 ;
  assign n1404 = ~n1402 & n1403 ;
  assign n1405 = ~n1401 & n1404 ;
  assign n1406 = ~n414 & n420 ;
  assign n1407 = n411 & n433 ;
  assign n1408 = ~n1406 & n1407 ;
  assign n1409 = ~n1405 & n1408 ;
  assign n1410 = ~n427 & n433 ;
  assign n1411 = n424 & n446 ;
  assign n1412 = ~n1410 & n1411 ;
  assign n1413 = ~n1409 & n1412 ;
  assign n1414 = ~n440 & n446 ;
  assign n1415 = n437 & n459 ;
  assign n1416 = ~n1414 & n1415 ;
  assign n1417 = ~n1413 & n1416 ;
  assign n1418 = ~n453 & n459 ;
  assign n1419 = n450 & n472 ;
  assign n1420 = ~n1418 & n1419 ;
  assign n1421 = ~n1417 & n1420 ;
  assign n1422 = ~n466 & n472 ;
  assign n1423 = n463 & n485 ;
  assign n1424 = ~n1422 & n1423 ;
  assign n1425 = ~n1421 & n1424 ;
  assign n1426 = ~n479 & n485 ;
  assign n1427 = n476 & n498 ;
  assign n1428 = ~n1426 & n1427 ;
  assign n1429 = ~n1425 & n1428 ;
  assign n1430 = ~n492 & n498 ;
  assign n1431 = n489 & n511 ;
  assign n1432 = ~n1430 & n1431 ;
  assign n1433 = ~n1429 & n1432 ;
  assign n1434 = ~n505 & n511 ;
  assign n1435 = n502 & n524 ;
  assign n1436 = ~n1434 & n1435 ;
  assign n1437 = ~n1433 & n1436 ;
  assign n1438 = ~n518 & n524 ;
  assign n1439 = n515 & n537 ;
  assign n1440 = ~n1438 & n1439 ;
  assign n1441 = ~n1437 & n1440 ;
  assign n1442 = ~n531 & n537 ;
  assign n1443 = n528 & n550 ;
  assign n1444 = ~n1442 & n1443 ;
  assign n1445 = ~n1441 & n1444 ;
  assign n1446 = ~n544 & n550 ;
  assign n1447 = n541 & n563 ;
  assign n1448 = ~n1446 & n1447 ;
  assign n1449 = ~n1445 & n1448 ;
  assign n1450 = ~n557 & n563 ;
  assign n1451 = n554 & n576 ;
  assign n1452 = ~n1450 & n1451 ;
  assign n1453 = ~n1449 & n1452 ;
  assign n1454 = ~n570 & n576 ;
  assign n1455 = n567 & n589 ;
  assign n1456 = ~n1454 & n1455 ;
  assign n1457 = ~n1453 & n1456 ;
  assign n1458 = ~n583 & n589 ;
  assign n1459 = n580 & n602 ;
  assign n1460 = ~n1458 & n1459 ;
  assign n1461 = ~n1457 & n1460 ;
  assign n1462 = ~n596 & n602 ;
  assign n1463 = n593 & n615 ;
  assign n1464 = ~n1462 & n1463 ;
  assign n1465 = ~n1461 & n1464 ;
  assign n1466 = ~n609 & n615 ;
  assign n1467 = n259 & n606 ;
  assign n1468 = ~n1466 & n1467 ;
  assign n1469 = ~n1465 & n1468 ;
  assign n1470 = n259 & ~n619 ;
  assign n1471 = ~\req[0]  & ~\req[1]  ;
  assign n1472 = ~n260 & n1471 ;
  assign n1473 = n1360 & n1472 ;
  assign n1474 = ~n1470 & n1473 ;
  assign n1475 = ~n1469 & n1474 ;
  assign n1476 = ~n1361 & ~n1475 ;
  assign n1477 = ~\priority[3]  & ~\priority[4]  ;
  assign n1478 = ~n630 & n1477 ;
  assign n1479 = ~\priority[4]  & \req[3]  ;
  assign n1480 = \req[4]  & ~n1479 ;
  assign n1481 = ~n1478 & n1480 ;
  assign n1482 = ~\priority[6]  & ~n1003 ;
  assign n1483 = n643 & ~n1482 ;
  assign n1484 = n636 & n657 ;
  assign n1485 = ~n1483 & n1484 ;
  assign n1486 = ~n651 & n657 ;
  assign n1487 = n648 & n670 ;
  assign n1488 = ~n1486 & n1487 ;
  assign n1489 = ~n1485 & n1488 ;
  assign n1490 = ~n664 & n670 ;
  assign n1491 = n661 & n683 ;
  assign n1492 = ~n1490 & n1491 ;
  assign n1493 = ~n1489 & n1492 ;
  assign n1494 = ~n677 & n683 ;
  assign n1495 = n674 & n696 ;
  assign n1496 = ~n1494 & n1495 ;
  assign n1497 = ~n1493 & n1496 ;
  assign n1498 = ~n690 & n696 ;
  assign n1499 = n687 & n709 ;
  assign n1500 = ~n1498 & n1499 ;
  assign n1501 = ~n1497 & n1500 ;
  assign n1502 = ~n703 & n709 ;
  assign n1503 = n700 & n722 ;
  assign n1504 = ~n1502 & n1503 ;
  assign n1505 = ~n1501 & n1504 ;
  assign n1506 = ~n716 & n722 ;
  assign n1507 = n713 & n735 ;
  assign n1508 = ~n1506 & n1507 ;
  assign n1509 = ~n1505 & n1508 ;
  assign n1510 = ~n729 & n735 ;
  assign n1511 = n726 & n748 ;
  assign n1512 = ~n1510 & n1511 ;
  assign n1513 = ~n1509 & n1512 ;
  assign n1514 = ~n742 & n748 ;
  assign n1515 = n739 & n761 ;
  assign n1516 = ~n1514 & n1515 ;
  assign n1517 = ~n1513 & n1516 ;
  assign n1518 = ~n755 & n761 ;
  assign n1519 = n752 & n774 ;
  assign n1520 = ~n1518 & n1519 ;
  assign n1521 = ~n1517 & n1520 ;
  assign n1522 = ~n768 & n774 ;
  assign n1523 = n765 & n787 ;
  assign n1524 = ~n1522 & n1523 ;
  assign n1525 = ~n1521 & n1524 ;
  assign n1526 = ~n781 & n787 ;
  assign n1527 = n778 & n800 ;
  assign n1528 = ~n1526 & n1527 ;
  assign n1529 = ~n1525 & n1528 ;
  assign n1530 = ~n794 & n800 ;
  assign n1531 = n791 & n813 ;
  assign n1532 = ~n1530 & n1531 ;
  assign n1533 = ~n1529 & n1532 ;
  assign n1534 = ~n807 & n813 ;
  assign n1535 = n804 & n826 ;
  assign n1536 = ~n1534 & n1535 ;
  assign n1537 = ~n1533 & n1536 ;
  assign n1538 = ~n820 & n826 ;
  assign n1539 = n817 & n839 ;
  assign n1540 = ~n1538 & n1539 ;
  assign n1541 = ~n1537 & n1540 ;
  assign n1542 = ~n833 & n839 ;
  assign n1543 = n830 & n852 ;
  assign n1544 = ~n1542 & n1543 ;
  assign n1545 = ~n1541 & n1544 ;
  assign n1546 = ~n846 & n852 ;
  assign n1547 = n843 & n865 ;
  assign n1548 = ~n1546 & n1547 ;
  assign n1549 = ~n1545 & n1548 ;
  assign n1550 = ~n859 & n865 ;
  assign n1551 = n856 & n878 ;
  assign n1552 = ~n1550 & n1551 ;
  assign n1553 = ~n1549 & n1552 ;
  assign n1554 = ~n872 & n878 ;
  assign n1555 = n869 & n891 ;
  assign n1556 = ~n1554 & n1555 ;
  assign n1557 = ~n1553 & n1556 ;
  assign n1558 = ~n885 & n891 ;
  assign n1559 = n882 & n904 ;
  assign n1560 = ~n1558 & n1559 ;
  assign n1561 = ~n1557 & n1560 ;
  assign n1562 = ~n898 & n904 ;
  assign n1563 = n895 & n917 ;
  assign n1564 = ~n1562 & n1563 ;
  assign n1565 = ~n1561 & n1564 ;
  assign n1566 = ~n911 & n917 ;
  assign n1567 = n908 & n930 ;
  assign n1568 = ~n1566 & n1567 ;
  assign n1569 = ~n1565 & n1568 ;
  assign n1570 = ~n924 & n930 ;
  assign n1571 = n921 & n943 ;
  assign n1572 = ~n1570 & n1571 ;
  assign n1573 = ~n1569 & n1572 ;
  assign n1574 = ~n937 & n943 ;
  assign n1575 = n934 & n956 ;
  assign n1576 = ~n1574 & n1575 ;
  assign n1577 = ~n1573 & n1576 ;
  assign n1578 = ~n950 & n956 ;
  assign n1579 = n947 & n969 ;
  assign n1580 = ~n1578 & n1579 ;
  assign n1581 = ~n1577 & n1580 ;
  assign n1582 = ~n963 & n969 ;
  assign n1583 = n960 & n982 ;
  assign n1584 = ~n1582 & n1583 ;
  assign n1585 = ~n1581 & n1584 ;
  assign n1586 = ~n976 & n982 ;
  assign n1587 = n626 & n973 ;
  assign n1588 = ~n1586 & n1587 ;
  assign n1589 = ~n1585 & n1588 ;
  assign n1590 = n626 & ~n986 ;
  assign n1591 = ~\req[1]  & ~\req[2]  ;
  assign n1592 = ~n627 & n1591 ;
  assign n1593 = n1480 & n1592 ;
  assign n1594 = ~n1590 & n1593 ;
  assign n1595 = ~n1589 & n1594 ;
  assign n1596 = ~n1481 & ~n1595 ;
  assign n1597 = \req[5]  & ~n275 ;
  assign n1598 = ~n272 & n1597 ;
  assign n1599 = ~\priority[7]  & ~n267 ;
  assign n1600 = n1009 & ~n1599 ;
  assign n1601 = n1002 & n1023 ;
  assign n1602 = ~n1600 & n1601 ;
  assign n1603 = ~n1017 & n1023 ;
  assign n1604 = n1014 & n1036 ;
  assign n1605 = ~n1603 & n1604 ;
  assign n1606 = ~n1602 & n1605 ;
  assign n1607 = ~n1030 & n1036 ;
  assign n1608 = n1027 & n1049 ;
  assign n1609 = ~n1607 & n1608 ;
  assign n1610 = ~n1606 & n1609 ;
  assign n1611 = ~n1043 & n1049 ;
  assign n1612 = n1040 & n1062 ;
  assign n1613 = ~n1611 & n1612 ;
  assign n1614 = ~n1610 & n1613 ;
  assign n1615 = ~n1056 & n1062 ;
  assign n1616 = n1053 & n1075 ;
  assign n1617 = ~n1615 & n1616 ;
  assign n1618 = ~n1614 & n1617 ;
  assign n1619 = ~n1069 & n1075 ;
  assign n1620 = n1066 & n1088 ;
  assign n1621 = ~n1619 & n1620 ;
  assign n1622 = ~n1618 & n1621 ;
  assign n1623 = ~n1082 & n1088 ;
  assign n1624 = n1079 & n1101 ;
  assign n1625 = ~n1623 & n1624 ;
  assign n1626 = ~n1622 & n1625 ;
  assign n1627 = ~n1095 & n1101 ;
  assign n1628 = n1092 & n1114 ;
  assign n1629 = ~n1627 & n1628 ;
  assign n1630 = ~n1626 & n1629 ;
  assign n1631 = ~n1108 & n1114 ;
  assign n1632 = n1105 & n1127 ;
  assign n1633 = ~n1631 & n1632 ;
  assign n1634 = ~n1630 & n1633 ;
  assign n1635 = ~n1121 & n1127 ;
  assign n1636 = n1118 & n1140 ;
  assign n1637 = ~n1635 & n1636 ;
  assign n1638 = ~n1634 & n1637 ;
  assign n1639 = ~n1134 & n1140 ;
  assign n1640 = n1131 & n1153 ;
  assign n1641 = ~n1639 & n1640 ;
  assign n1642 = ~n1638 & n1641 ;
  assign n1643 = ~n1147 & n1153 ;
  assign n1644 = n1144 & n1166 ;
  assign n1645 = ~n1643 & n1644 ;
  assign n1646 = ~n1642 & n1645 ;
  assign n1647 = ~n1160 & n1166 ;
  assign n1648 = n1157 & n1179 ;
  assign n1649 = ~n1647 & n1648 ;
  assign n1650 = ~n1646 & n1649 ;
  assign n1651 = ~n1173 & n1179 ;
  assign n1652 = n1170 & n1192 ;
  assign n1653 = ~n1651 & n1652 ;
  assign n1654 = ~n1650 & n1653 ;
  assign n1655 = ~n1186 & n1192 ;
  assign n1656 = n1183 & n1205 ;
  assign n1657 = ~n1655 & n1656 ;
  assign n1658 = ~n1654 & n1657 ;
  assign n1659 = ~n1199 & n1205 ;
  assign n1660 = n1196 & n1218 ;
  assign n1661 = ~n1659 & n1660 ;
  assign n1662 = ~n1658 & n1661 ;
  assign n1663 = ~n1212 & n1218 ;
  assign n1664 = n1209 & n1231 ;
  assign n1665 = ~n1663 & n1664 ;
  assign n1666 = ~n1662 & n1665 ;
  assign n1667 = ~n1225 & n1231 ;
  assign n1668 = n1222 & n1244 ;
  assign n1669 = ~n1667 & n1668 ;
  assign n1670 = ~n1666 & n1669 ;
  assign n1671 = ~n1238 & n1244 ;
  assign n1672 = n1235 & n1257 ;
  assign n1673 = ~n1671 & n1672 ;
  assign n1674 = ~n1670 & n1673 ;
  assign n1675 = ~n1251 & n1257 ;
  assign n1676 = n1248 & n1270 ;
  assign n1677 = ~n1675 & n1676 ;
  assign n1678 = ~n1674 & n1677 ;
  assign n1679 = ~n1264 & n1270 ;
  assign n1680 = n1261 & n1283 ;
  assign n1681 = ~n1679 & n1680 ;
  assign n1682 = ~n1678 & n1681 ;
  assign n1683 = ~n1277 & n1283 ;
  assign n1684 = n1274 & n1296 ;
  assign n1685 = ~n1683 & n1684 ;
  assign n1686 = ~n1682 & n1685 ;
  assign n1687 = ~n1290 & n1296 ;
  assign n1688 = n1287 & n1309 ;
  assign n1689 = ~n1687 & n1688 ;
  assign n1690 = ~n1686 & n1689 ;
  assign n1691 = ~n1303 & n1309 ;
  assign n1692 = n1300 & n1322 ;
  assign n1693 = ~n1691 & n1692 ;
  assign n1694 = ~n1690 & n1693 ;
  assign n1695 = ~n1316 & n1322 ;
  assign n1696 = n1313 & n1335 ;
  assign n1697 = ~n1695 & n1696 ;
  assign n1698 = ~n1694 & n1697 ;
  assign n1699 = ~n1329 & n1335 ;
  assign n1700 = n1326 & n1348 ;
  assign n1701 = ~n1699 & n1700 ;
  assign n1702 = ~n1698 & n1701 ;
  assign n1703 = ~n1342 & n1348 ;
  assign n1704 = n993 & n1339 ;
  assign n1705 = ~n1703 & n1704 ;
  assign n1706 = ~n1702 & n1705 ;
  assign n1707 = n993 & ~n1352 ;
  assign n1708 = n265 & ~n994 ;
  assign n1709 = n1597 & n1708 ;
  assign n1710 = ~n1707 & n1709 ;
  assign n1711 = ~n1706 & n1710 ;
  assign n1712 = ~n1598 & ~n1711 ;
  assign n1713 = \req[6]  & ~n642 ;
  assign n1714 = ~n639 & n1713 ;
  assign n1715 = ~\priority[8]  & ~n634 ;
  assign n1716 = n283 & ~n1715 ;
  assign n1717 = n290 & n297 ;
  assign n1718 = ~n1716 & n1717 ;
  assign n1719 = ~n281 & n297 ;
  assign n1720 = n303 & n310 ;
  assign n1721 = ~n1719 & n1720 ;
  assign n1722 = ~n1718 & n1721 ;
  assign n1723 = ~n294 & n310 ;
  assign n1724 = n316 & n323 ;
  assign n1725 = ~n1723 & n1724 ;
  assign n1726 = ~n1722 & n1725 ;
  assign n1727 = ~n307 & n323 ;
  assign n1728 = n329 & n336 ;
  assign n1729 = ~n1727 & n1728 ;
  assign n1730 = ~n1726 & n1729 ;
  assign n1731 = ~n320 & n336 ;
  assign n1732 = n342 & n349 ;
  assign n1733 = ~n1731 & n1732 ;
  assign n1734 = ~n1730 & n1733 ;
  assign n1735 = ~n333 & n349 ;
  assign n1736 = n355 & n362 ;
  assign n1737 = ~n1735 & n1736 ;
  assign n1738 = ~n1734 & n1737 ;
  assign n1739 = ~n346 & n362 ;
  assign n1740 = n368 & n375 ;
  assign n1741 = ~n1739 & n1740 ;
  assign n1742 = ~n1738 & n1741 ;
  assign n1743 = ~n359 & n375 ;
  assign n1744 = n381 & n388 ;
  assign n1745 = ~n1743 & n1744 ;
  assign n1746 = ~n1742 & n1745 ;
  assign n1747 = ~n372 & n388 ;
  assign n1748 = n394 & n401 ;
  assign n1749 = ~n1747 & n1748 ;
  assign n1750 = ~n1746 & n1749 ;
  assign n1751 = ~n385 & n401 ;
  assign n1752 = n407 & n414 ;
  assign n1753 = ~n1751 & n1752 ;
  assign n1754 = ~n1750 & n1753 ;
  assign n1755 = ~n398 & n414 ;
  assign n1756 = n420 & n427 ;
  assign n1757 = ~n1755 & n1756 ;
  assign n1758 = ~n1754 & n1757 ;
  assign n1759 = ~n411 & n427 ;
  assign n1760 = n433 & n440 ;
  assign n1761 = ~n1759 & n1760 ;
  assign n1762 = ~n1758 & n1761 ;
  assign n1763 = ~n424 & n440 ;
  assign n1764 = n446 & n453 ;
  assign n1765 = ~n1763 & n1764 ;
  assign n1766 = ~n1762 & n1765 ;
  assign n1767 = ~n437 & n453 ;
  assign n1768 = n459 & n466 ;
  assign n1769 = ~n1767 & n1768 ;
  assign n1770 = ~n1766 & n1769 ;
  assign n1771 = ~n450 & n466 ;
  assign n1772 = n472 & n479 ;
  assign n1773 = ~n1771 & n1772 ;
  assign n1774 = ~n1770 & n1773 ;
  assign n1775 = ~n463 & n479 ;
  assign n1776 = n485 & n492 ;
  assign n1777 = ~n1775 & n1776 ;
  assign n1778 = ~n1774 & n1777 ;
  assign n1779 = ~n476 & n492 ;
  assign n1780 = n498 & n505 ;
  assign n1781 = ~n1779 & n1780 ;
  assign n1782 = ~n1778 & n1781 ;
  assign n1783 = ~n489 & n505 ;
  assign n1784 = n511 & n518 ;
  assign n1785 = ~n1783 & n1784 ;
  assign n1786 = ~n1782 & n1785 ;
  assign n1787 = ~n502 & n518 ;
  assign n1788 = n524 & n531 ;
  assign n1789 = ~n1787 & n1788 ;
  assign n1790 = ~n1786 & n1789 ;
  assign n1791 = ~n515 & n531 ;
  assign n1792 = n537 & n544 ;
  assign n1793 = ~n1791 & n1792 ;
  assign n1794 = ~n1790 & n1793 ;
  assign n1795 = ~n528 & n544 ;
  assign n1796 = n550 & n557 ;
  assign n1797 = ~n1795 & n1796 ;
  assign n1798 = ~n1794 & n1797 ;
  assign n1799 = ~n541 & n557 ;
  assign n1800 = n563 & n570 ;
  assign n1801 = ~n1799 & n1800 ;
  assign n1802 = ~n1798 & n1801 ;
  assign n1803 = ~n554 & n570 ;
  assign n1804 = n576 & n583 ;
  assign n1805 = ~n1803 & n1804 ;
  assign n1806 = ~n1802 & n1805 ;
  assign n1807 = ~n567 & n583 ;
  assign n1808 = n589 & n596 ;
  assign n1809 = ~n1807 & n1808 ;
  assign n1810 = ~n1806 & n1809 ;
  assign n1811 = ~n580 & n596 ;
  assign n1812 = n602 & n609 ;
  assign n1813 = ~n1811 & n1812 ;
  assign n1814 = ~n1810 & n1813 ;
  assign n1815 = ~n593 & n609 ;
  assign n1816 = n615 & n619 ;
  assign n1817 = ~n1815 & n1816 ;
  assign n1818 = ~n1814 & n1817 ;
  assign n1819 = ~n606 & n619 ;
  assign n1820 = n259 & n1358 ;
  assign n1821 = ~n1819 & n1820 ;
  assign n1822 = ~n1818 & n1821 ;
  assign n1823 = n1358 & ~n1472 ;
  assign n1824 = n632 & ~n1359 ;
  assign n1825 = n1713 & n1824 ;
  assign n1826 = ~n1823 & n1825 ;
  assign n1827 = ~n1822 & n1826 ;
  assign n1828 = ~n1714 & ~n1827 ;
  assign n1829 = \req[7]  & ~n1008 ;
  assign n1830 = ~n1005 & n1829 ;
  assign n1831 = ~\priority[9]  & ~n1000 ;
  assign n1832 = n650 & ~n1831 ;
  assign n1833 = n657 & n664 ;
  assign n1834 = ~n1832 & n1833 ;
  assign n1835 = ~n648 & n664 ;
  assign n1836 = n670 & n677 ;
  assign n1837 = ~n1835 & n1836 ;
  assign n1838 = ~n1834 & n1837 ;
  assign n1839 = ~n661 & n677 ;
  assign n1840 = n683 & n690 ;
  assign n1841 = ~n1839 & n1840 ;
  assign n1842 = ~n1838 & n1841 ;
  assign n1843 = ~n674 & n690 ;
  assign n1844 = n696 & n703 ;
  assign n1845 = ~n1843 & n1844 ;
  assign n1846 = ~n1842 & n1845 ;
  assign n1847 = ~n687 & n703 ;
  assign n1848 = n709 & n716 ;
  assign n1849 = ~n1847 & n1848 ;
  assign n1850 = ~n1846 & n1849 ;
  assign n1851 = ~n700 & n716 ;
  assign n1852 = n722 & n729 ;
  assign n1853 = ~n1851 & n1852 ;
  assign n1854 = ~n1850 & n1853 ;
  assign n1855 = ~n713 & n729 ;
  assign n1856 = n735 & n742 ;
  assign n1857 = ~n1855 & n1856 ;
  assign n1858 = ~n1854 & n1857 ;
  assign n1859 = ~n726 & n742 ;
  assign n1860 = n748 & n755 ;
  assign n1861 = ~n1859 & n1860 ;
  assign n1862 = ~n1858 & n1861 ;
  assign n1863 = ~n739 & n755 ;
  assign n1864 = n761 & n768 ;
  assign n1865 = ~n1863 & n1864 ;
  assign n1866 = ~n1862 & n1865 ;
  assign n1867 = ~n752 & n768 ;
  assign n1868 = n774 & n781 ;
  assign n1869 = ~n1867 & n1868 ;
  assign n1870 = ~n1866 & n1869 ;
  assign n1871 = ~n765 & n781 ;
  assign n1872 = n787 & n794 ;
  assign n1873 = ~n1871 & n1872 ;
  assign n1874 = ~n1870 & n1873 ;
  assign n1875 = ~n778 & n794 ;
  assign n1876 = n800 & n807 ;
  assign n1877 = ~n1875 & n1876 ;
  assign n1878 = ~n1874 & n1877 ;
  assign n1879 = ~n791 & n807 ;
  assign n1880 = n813 & n820 ;
  assign n1881 = ~n1879 & n1880 ;
  assign n1882 = ~n1878 & n1881 ;
  assign n1883 = ~n804 & n820 ;
  assign n1884 = n826 & n833 ;
  assign n1885 = ~n1883 & n1884 ;
  assign n1886 = ~n1882 & n1885 ;
  assign n1887 = ~n817 & n833 ;
  assign n1888 = n839 & n846 ;
  assign n1889 = ~n1887 & n1888 ;
  assign n1890 = ~n1886 & n1889 ;
  assign n1891 = ~n830 & n846 ;
  assign n1892 = n852 & n859 ;
  assign n1893 = ~n1891 & n1892 ;
  assign n1894 = ~n1890 & n1893 ;
  assign n1895 = ~n843 & n859 ;
  assign n1896 = n865 & n872 ;
  assign n1897 = ~n1895 & n1896 ;
  assign n1898 = ~n1894 & n1897 ;
  assign n1899 = ~n856 & n872 ;
  assign n1900 = n878 & n885 ;
  assign n1901 = ~n1899 & n1900 ;
  assign n1902 = ~n1898 & n1901 ;
  assign n1903 = ~n869 & n885 ;
  assign n1904 = n891 & n898 ;
  assign n1905 = ~n1903 & n1904 ;
  assign n1906 = ~n1902 & n1905 ;
  assign n1907 = ~n882 & n898 ;
  assign n1908 = n904 & n911 ;
  assign n1909 = ~n1907 & n1908 ;
  assign n1910 = ~n1906 & n1909 ;
  assign n1911 = ~n895 & n911 ;
  assign n1912 = n917 & n924 ;
  assign n1913 = ~n1911 & n1912 ;
  assign n1914 = ~n1910 & n1913 ;
  assign n1915 = ~n908 & n924 ;
  assign n1916 = n930 & n937 ;
  assign n1917 = ~n1915 & n1916 ;
  assign n1918 = ~n1914 & n1917 ;
  assign n1919 = ~n921 & n937 ;
  assign n1920 = n943 & n950 ;
  assign n1921 = ~n1919 & n1920 ;
  assign n1922 = ~n1918 & n1921 ;
  assign n1923 = ~n934 & n950 ;
  assign n1924 = n956 & n963 ;
  assign n1925 = ~n1923 & n1924 ;
  assign n1926 = ~n1922 & n1925 ;
  assign n1927 = ~n947 & n963 ;
  assign n1928 = n969 & n976 ;
  assign n1929 = ~n1927 & n1928 ;
  assign n1930 = ~n1926 & n1929 ;
  assign n1931 = ~n960 & n976 ;
  assign n1932 = n982 & n986 ;
  assign n1933 = ~n1931 & n1932 ;
  assign n1934 = ~n1930 & n1933 ;
  assign n1935 = ~n973 & n986 ;
  assign n1936 = n626 & n1478 ;
  assign n1937 = ~n1935 & n1936 ;
  assign n1938 = ~n1934 & n1937 ;
  assign n1939 = n1478 & ~n1592 ;
  assign n1940 = n998 & ~n1479 ;
  assign n1941 = n1829 & n1940 ;
  assign n1942 = ~n1939 & n1941 ;
  assign n1943 = ~n1938 & n1942 ;
  assign n1944 = ~n1830 & ~n1943 ;
  assign n1945 = \req[8]  & ~n282 ;
  assign n1946 = ~n269 & n1945 ;
  assign n1947 = ~\priority[10]  & ~n288 ;
  assign n1948 = n1016 & ~n1947 ;
  assign n1949 = n1023 & n1030 ;
  assign n1950 = ~n1948 & n1949 ;
  assign n1951 = ~n1014 & n1030 ;
  assign n1952 = n1036 & n1043 ;
  assign n1953 = ~n1951 & n1952 ;
  assign n1954 = ~n1950 & n1953 ;
  assign n1955 = ~n1027 & n1043 ;
  assign n1956 = n1049 & n1056 ;
  assign n1957 = ~n1955 & n1956 ;
  assign n1958 = ~n1954 & n1957 ;
  assign n1959 = ~n1040 & n1056 ;
  assign n1960 = n1062 & n1069 ;
  assign n1961 = ~n1959 & n1960 ;
  assign n1962 = ~n1958 & n1961 ;
  assign n1963 = ~n1053 & n1069 ;
  assign n1964 = n1075 & n1082 ;
  assign n1965 = ~n1963 & n1964 ;
  assign n1966 = ~n1962 & n1965 ;
  assign n1967 = ~n1066 & n1082 ;
  assign n1968 = n1088 & n1095 ;
  assign n1969 = ~n1967 & n1968 ;
  assign n1970 = ~n1966 & n1969 ;
  assign n1971 = ~n1079 & n1095 ;
  assign n1972 = n1101 & n1108 ;
  assign n1973 = ~n1971 & n1972 ;
  assign n1974 = ~n1970 & n1973 ;
  assign n1975 = ~n1092 & n1108 ;
  assign n1976 = n1114 & n1121 ;
  assign n1977 = ~n1975 & n1976 ;
  assign n1978 = ~n1974 & n1977 ;
  assign n1979 = ~n1105 & n1121 ;
  assign n1980 = n1127 & n1134 ;
  assign n1981 = ~n1979 & n1980 ;
  assign n1982 = ~n1978 & n1981 ;
  assign n1983 = ~n1118 & n1134 ;
  assign n1984 = n1140 & n1147 ;
  assign n1985 = ~n1983 & n1984 ;
  assign n1986 = ~n1982 & n1985 ;
  assign n1987 = ~n1131 & n1147 ;
  assign n1988 = n1153 & n1160 ;
  assign n1989 = ~n1987 & n1988 ;
  assign n1990 = ~n1986 & n1989 ;
  assign n1991 = ~n1144 & n1160 ;
  assign n1992 = n1166 & n1173 ;
  assign n1993 = ~n1991 & n1992 ;
  assign n1994 = ~n1990 & n1993 ;
  assign n1995 = ~n1157 & n1173 ;
  assign n1996 = n1179 & n1186 ;
  assign n1997 = ~n1995 & n1996 ;
  assign n1998 = ~n1994 & n1997 ;
  assign n1999 = ~n1170 & n1186 ;
  assign n2000 = n1192 & n1199 ;
  assign n2001 = ~n1999 & n2000 ;
  assign n2002 = ~n1998 & n2001 ;
  assign n2003 = ~n1183 & n1199 ;
  assign n2004 = n1205 & n1212 ;
  assign n2005 = ~n2003 & n2004 ;
  assign n2006 = ~n2002 & n2005 ;
  assign n2007 = ~n1196 & n1212 ;
  assign n2008 = n1218 & n1225 ;
  assign n2009 = ~n2007 & n2008 ;
  assign n2010 = ~n2006 & n2009 ;
  assign n2011 = ~n1209 & n1225 ;
  assign n2012 = n1231 & n1238 ;
  assign n2013 = ~n2011 & n2012 ;
  assign n2014 = ~n2010 & n2013 ;
  assign n2015 = ~n1222 & n1238 ;
  assign n2016 = n1244 & n1251 ;
  assign n2017 = ~n2015 & n2016 ;
  assign n2018 = ~n2014 & n2017 ;
  assign n2019 = ~n1235 & n1251 ;
  assign n2020 = n1257 & n1264 ;
  assign n2021 = ~n2019 & n2020 ;
  assign n2022 = ~n2018 & n2021 ;
  assign n2023 = ~n1248 & n1264 ;
  assign n2024 = n1270 & n1277 ;
  assign n2025 = ~n2023 & n2024 ;
  assign n2026 = ~n2022 & n2025 ;
  assign n2027 = ~n1261 & n1277 ;
  assign n2028 = n1283 & n1290 ;
  assign n2029 = ~n2027 & n2028 ;
  assign n2030 = ~n2026 & n2029 ;
  assign n2031 = ~n1274 & n1290 ;
  assign n2032 = n1296 & n1303 ;
  assign n2033 = ~n2031 & n2032 ;
  assign n2034 = ~n2030 & n2033 ;
  assign n2035 = ~n1287 & n1303 ;
  assign n2036 = n1309 & n1316 ;
  assign n2037 = ~n2035 & n2036 ;
  assign n2038 = ~n2034 & n2037 ;
  assign n2039 = ~n1300 & n1316 ;
  assign n2040 = n1322 & n1329 ;
  assign n2041 = ~n2039 & n2040 ;
  assign n2042 = ~n2038 & n2041 ;
  assign n2043 = ~n1313 & n1329 ;
  assign n2044 = n1335 & n1342 ;
  assign n2045 = ~n2043 & n2044 ;
  assign n2046 = ~n2042 & n2045 ;
  assign n2047 = ~n1326 & n1342 ;
  assign n2048 = n1348 & n1352 ;
  assign n2049 = ~n2047 & n2048 ;
  assign n2050 = ~n2046 & n2049 ;
  assign n2051 = ~n1339 & n1352 ;
  assign n2052 = n272 & n993 ;
  assign n2053 = ~n2051 & n2052 ;
  assign n2054 = ~n2050 & n2053 ;
  assign n2055 = n272 & ~n1708 ;
  assign n2056 = n277 & n1945 ;
  assign n2057 = ~n2055 & n2056 ;
  assign n2058 = ~n2054 & n2057 ;
  assign n2059 = ~n1946 & ~n2058 ;
  assign n2060 = \req[9]  & ~n649 ;
  assign n2061 = ~n636 & n2060 ;
  assign n2062 = ~\priority[11]  & ~n655 ;
  assign n2063 = n280 & ~n2062 ;
  assign n2064 = n298 & ~n2063 ;
  assign n2065 = n312 & ~n2064 ;
  assign n2066 = n325 & ~n2065 ;
  assign n2067 = n338 & ~n2066 ;
  assign n2068 = n351 & ~n2067 ;
  assign n2069 = n364 & ~n2068 ;
  assign n2070 = n377 & ~n2069 ;
  assign n2071 = n390 & ~n2070 ;
  assign n2072 = n403 & ~n2071 ;
  assign n2073 = n416 & ~n2072 ;
  assign n2074 = n429 & ~n2073 ;
  assign n2075 = n442 & ~n2074 ;
  assign n2076 = n455 & ~n2075 ;
  assign n2077 = n468 & ~n2076 ;
  assign n2078 = n481 & ~n2077 ;
  assign n2079 = n494 & ~n2078 ;
  assign n2080 = n507 & ~n2079 ;
  assign n2081 = n520 & ~n2080 ;
  assign n2082 = n533 & ~n2081 ;
  assign n2083 = n546 & ~n2082 ;
  assign n2084 = n559 & ~n2083 ;
  assign n2085 = n572 & ~n2084 ;
  assign n2086 = n585 & ~n2085 ;
  assign n2087 = n598 & ~n2086 ;
  assign n2088 = n611 & ~n2087 ;
  assign n2089 = n619 & n1472 ;
  assign n2090 = ~n616 & n2089 ;
  assign n2091 = ~n2088 & n2090 ;
  assign n2092 = ~n259 & n1472 ;
  assign n2093 = n639 & n1358 ;
  assign n2094 = ~n2092 & n2093 ;
  assign n2095 = ~n2091 & n2094 ;
  assign n2096 = n639 & ~n1824 ;
  assign n2097 = n644 & n2060 ;
  assign n2098 = ~n2096 & n2097 ;
  assign n2099 = ~n2095 & n2098 ;
  assign n2100 = ~n2061 & ~n2099 ;
  assign n2101 = \req[10]  & ~n1015 ;
  assign n2102 = ~n1002 & n2101 ;
  assign n2103 = ~\priority[12]  & ~n1021 ;
  assign n2104 = n647 & ~n2103 ;
  assign n2105 = n665 & ~n2104 ;
  assign n2106 = n679 & ~n2105 ;
  assign n2107 = n692 & ~n2106 ;
  assign n2108 = n705 & ~n2107 ;
  assign n2109 = n718 & ~n2108 ;
  assign n2110 = n731 & ~n2109 ;
  assign n2111 = n744 & ~n2110 ;
  assign n2112 = n757 & ~n2111 ;
  assign n2113 = n770 & ~n2112 ;
  assign n2114 = n783 & ~n2113 ;
  assign n2115 = n796 & ~n2114 ;
  assign n2116 = n809 & ~n2115 ;
  assign n2117 = ~n814 & n821 ;
  assign n2118 = ~n2116 & n2117 ;
  assign n2119 = n835 & ~n2118 ;
  assign n2120 = n848 & ~n2119 ;
  assign n2121 = n861 & ~n2120 ;
  assign n2122 = n874 & ~n2121 ;
  assign n2123 = n887 & ~n2122 ;
  assign n2124 = n900 & ~n2123 ;
  assign n2125 = n913 & ~n2124 ;
  assign n2126 = n926 & ~n2125 ;
  assign n2127 = n939 & ~n2126 ;
  assign n2128 = n952 & ~n2127 ;
  assign n2129 = n965 & ~n2128 ;
  assign n2130 = n978 & ~n2129 ;
  assign n2131 = n986 & n1592 ;
  assign n2132 = ~n983 & n2131 ;
  assign n2133 = ~n2130 & n2132 ;
  assign n2134 = ~n626 & n1592 ;
  assign n2135 = n1005 & n1478 ;
  assign n2136 = ~n2134 & n2135 ;
  assign n2137 = ~n2133 & n2136 ;
  assign n2138 = n1005 & ~n1940 ;
  assign n2139 = n1010 & n2101 ;
  assign n2140 = ~n2138 & n2139 ;
  assign n2141 = ~n2137 & n2140 ;
  assign n2142 = ~n2102 & ~n2141 ;
  assign n2143 = \req[11]  & ~n279 ;
  assign n2144 = ~n290 & n2143 ;
  assign n2145 = ~\priority[13]  & ~n295 ;
  assign n2146 = n1013 & ~n2145 ;
  assign n2147 = n1031 & ~n2146 ;
  assign n2148 = n1045 & ~n2147 ;
  assign n2149 = n1058 & ~n2148 ;
  assign n2150 = n1071 & ~n2149 ;
  assign n2151 = n1084 & ~n2150 ;
  assign n2152 = n1097 & ~n2151 ;
  assign n2153 = n1110 & ~n2152 ;
  assign n2154 = n1123 & ~n2153 ;
  assign n2155 = n1136 & ~n2154 ;
  assign n2156 = n1149 & ~n2155 ;
  assign n2157 = n1162 & ~n2156 ;
  assign n2158 = n1175 & ~n2157 ;
  assign n2159 = n1188 & ~n2158 ;
  assign n2160 = n1201 & ~n2159 ;
  assign n2161 = n1214 & ~n2160 ;
  assign n2162 = n1227 & ~n2161 ;
  assign n2163 = n1240 & ~n2162 ;
  assign n2164 = n1253 & ~n2163 ;
  assign n2165 = n1266 & ~n2164 ;
  assign n2166 = n1279 & ~n2165 ;
  assign n2167 = n1292 & ~n2166 ;
  assign n2168 = n1305 & ~n2167 ;
  assign n2169 = n1318 & ~n2168 ;
  assign n2170 = n1331 & ~n2169 ;
  assign n2171 = n1344 & ~n2170 ;
  assign n2172 = n1352 & n1708 ;
  assign n2173 = ~n1349 & n2172 ;
  assign n2174 = ~n2171 & n2173 ;
  assign n2175 = ~n993 & n1708 ;
  assign n2176 = n273 & ~n2175 ;
  assign n2177 = ~n2174 & n2176 ;
  assign n2178 = n284 & n2143 ;
  assign n2179 = ~n278 & n2178 ;
  assign n2180 = ~n2177 & n2179 ;
  assign n2181 = ~n2144 & ~n2180 ;
  assign n2182 = \req[12]  & ~n646 ;
  assign n2183 = ~n657 & n2182 ;
  assign n2184 = ~\priority[14]  & ~n662 ;
  assign n2185 = n302 & ~n2184 ;
  assign n2186 = n1371 & ~n2185 ;
  assign n2187 = n1376 & ~n2186 ;
  assign n2188 = n1380 & ~n2187 ;
  assign n2189 = n1384 & ~n2188 ;
  assign n2190 = n1388 & ~n2189 ;
  assign n2191 = n1392 & ~n2190 ;
  assign n2192 = n1396 & ~n2191 ;
  assign n2193 = n1400 & ~n2192 ;
  assign n2194 = n1404 & ~n2193 ;
  assign n2195 = n1408 & ~n2194 ;
  assign n2196 = n1412 & ~n2195 ;
  assign n2197 = n1416 & ~n2196 ;
  assign n2198 = n1420 & ~n2197 ;
  assign n2199 = n1424 & ~n2198 ;
  assign n2200 = n1428 & ~n2199 ;
  assign n2201 = n1432 & ~n2200 ;
  assign n2202 = n1436 & ~n2201 ;
  assign n2203 = n1440 & ~n2202 ;
  assign n2204 = n1444 & ~n2203 ;
  assign n2205 = n1448 & ~n2204 ;
  assign n2206 = n1452 & ~n2205 ;
  assign n2207 = n1456 & ~n2206 ;
  assign n2208 = n1460 & ~n2207 ;
  assign n2209 = n1464 & ~n2208 ;
  assign n2210 = n1468 & ~n2209 ;
  assign n2211 = n1472 & n1824 ;
  assign n2212 = ~n1470 & n2211 ;
  assign n2213 = ~n2210 & n2212 ;
  assign n2214 = ~n1358 & n1824 ;
  assign n2215 = n640 & ~n2214 ;
  assign n2216 = ~n2213 & n2215 ;
  assign n2217 = n651 & n2182 ;
  assign n2218 = ~n645 & n2217 ;
  assign n2219 = ~n2216 & n2218 ;
  assign n2220 = ~n2183 & ~n2219 ;
  assign n2221 = \req[13]  & ~n1012 ;
  assign n2222 = ~n1023 & n2221 ;
  assign n2223 = ~\priority[15]  & ~n1028 ;
  assign n2224 = n669 & ~n2223 ;
  assign n2225 = n1491 & ~n2224 ;
  assign n2226 = n1496 & ~n2225 ;
  assign n2227 = n1500 & ~n2226 ;
  assign n2228 = n1504 & ~n2227 ;
  assign n2229 = ~n1506 & n1507 ;
  assign n2230 = ~n2228 & n2229 ;
  assign n2231 = n1512 & ~n2230 ;
  assign n2232 = n1516 & ~n2231 ;
  assign n2233 = n1520 & ~n2232 ;
  assign n2234 = n1524 & ~n2233 ;
  assign n2235 = n1528 & ~n2234 ;
  assign n2236 = n1532 & ~n2235 ;
  assign n2237 = n1536 & ~n2236 ;
  assign n2238 = n1540 & ~n2237 ;
  assign n2239 = n1544 & ~n2238 ;
  assign n2240 = n1548 & ~n2239 ;
  assign n2241 = n1552 & ~n2240 ;
  assign n2242 = n1556 & ~n2241 ;
  assign n2243 = n1560 & ~n2242 ;
  assign n2244 = n1564 & ~n2243 ;
  assign n2245 = n1568 & ~n2244 ;
  assign n2246 = n1572 & ~n2245 ;
  assign n2247 = n1576 & ~n2246 ;
  assign n2248 = n1580 & ~n2247 ;
  assign n2249 = n1584 & ~n2248 ;
  assign n2250 = n1588 & ~n2249 ;
  assign n2251 = n1592 & n1940 ;
  assign n2252 = ~n1590 & n2251 ;
  assign n2253 = ~n2250 & n2252 ;
  assign n2254 = ~n1478 & n1940 ;
  assign n2255 = n1006 & ~n2254 ;
  assign n2256 = ~n2253 & n2255 ;
  assign n2257 = n1017 & n2221 ;
  assign n2258 = ~n1011 & n2257 ;
  assign n2259 = ~n2256 & n2258 ;
  assign n2260 = ~n2222 & ~n2259 ;
  assign n2261 = \req[14]  & ~n301 ;
  assign n2262 = ~n297 & n2261 ;
  assign n2263 = ~\priority[16]  & ~n292 ;
  assign n2264 = n1035 & ~n2263 ;
  assign n2265 = n1608 & ~n2264 ;
  assign n2266 = n1613 & ~n2265 ;
  assign n2267 = n1617 & ~n2266 ;
  assign n2268 = n1621 & ~n2267 ;
  assign n2269 = n1625 & ~n2268 ;
  assign n2270 = n1629 & ~n2269 ;
  assign n2271 = n1633 & ~n2270 ;
  assign n2272 = n1637 & ~n2271 ;
  assign n2273 = n1641 & ~n2272 ;
  assign n2274 = n1645 & ~n2273 ;
  assign n2275 = n1649 & ~n2274 ;
  assign n2276 = n1653 & ~n2275 ;
  assign n2277 = n1657 & ~n2276 ;
  assign n2278 = n1661 & ~n2277 ;
  assign n2279 = n1665 & ~n2278 ;
  assign n2280 = n1669 & ~n2279 ;
  assign n2281 = n1673 & ~n2280 ;
  assign n2282 = n1677 & ~n2281 ;
  assign n2283 = n1681 & ~n2282 ;
  assign n2284 = n1685 & ~n2283 ;
  assign n2285 = n1689 & ~n2284 ;
  assign n2286 = n1693 & ~n2285 ;
  assign n2287 = n1697 & ~n2286 ;
  assign n2288 = n1701 & ~n2287 ;
  assign n2289 = n1705 & ~n2288 ;
  assign n2290 = n277 & n1708 ;
  assign n2291 = ~n1707 & n2290 ;
  assign n2292 = ~n2289 & n2291 ;
  assign n2293 = ~n272 & n277 ;
  assign n2294 = n1364 & ~n2293 ;
  assign n2295 = ~n2292 & n2294 ;
  assign n2296 = n281 & n2261 ;
  assign n2297 = ~n1366 & n2296 ;
  assign n2298 = ~n2295 & n2297 ;
  assign n2299 = ~n2262 & ~n2298 ;
  assign n2300 = \req[15]  & ~n668 ;
  assign n2301 = ~n664 & n2300 ;
  assign n2302 = ~\priority[17]  & ~n659 ;
  assign n2303 = n309 & ~n2302 ;
  assign n2304 = n1724 & ~n2303 ;
  assign n2305 = n1729 & ~n2304 ;
  assign n2306 = n1733 & ~n2305 ;
  assign n2307 = n1737 & ~n2306 ;
  assign n2308 = n1741 & ~n2307 ;
  assign n2309 = n1745 & ~n2308 ;
  assign n2310 = n1749 & ~n2309 ;
  assign n2311 = n1753 & ~n2310 ;
  assign n2312 = n1757 & ~n2311 ;
  assign n2313 = n1761 & ~n2312 ;
  assign n2314 = n1765 & ~n2313 ;
  assign n2315 = n1769 & ~n2314 ;
  assign n2316 = n1773 & ~n2315 ;
  assign n2317 = n1777 & ~n2316 ;
  assign n2318 = n1781 & ~n2317 ;
  assign n2319 = n1785 & ~n2318 ;
  assign n2320 = n1789 & ~n2319 ;
  assign n2321 = n1793 & ~n2320 ;
  assign n2322 = n1797 & ~n2321 ;
  assign n2323 = n1801 & ~n2322 ;
  assign n2324 = n1805 & ~n2323 ;
  assign n2325 = n1809 & ~n2324 ;
  assign n2326 = n1813 & ~n2325 ;
  assign n2327 = n1817 & ~n2326 ;
  assign n2328 = n1821 & ~n2327 ;
  assign n2329 = n644 & n1824 ;
  assign n2330 = ~n1823 & n2329 ;
  assign n2331 = ~n2328 & n2330 ;
  assign n2332 = ~n639 & n644 ;
  assign n2333 = n1484 & ~n2332 ;
  assign n2334 = ~n2331 & n2333 ;
  assign n2335 = n648 & n2300 ;
  assign n2336 = ~n1486 & n2335 ;
  assign n2337 = ~n2334 & n2336 ;
  assign n2338 = ~n2301 & ~n2337 ;
  assign n2339 = \req[16]  & ~n1034 ;
  assign n2340 = ~n1030 & n2339 ;
  assign n2341 = ~\priority[18]  & ~n1025 ;
  assign n2342 = n676 & ~n2341 ;
  assign n2343 = n1840 & ~n2342 ;
  assign n2344 = n1845 & ~n2343 ;
  assign n2345 = n1849 & ~n2344 ;
  assign n2346 = n1853 & ~n2345 ;
  assign n2347 = n1857 & ~n2346 ;
  assign n2348 = n1861 & ~n2347 ;
  assign n2349 = n1865 & ~n2348 ;
  assign n2350 = n1869 & ~n2349 ;
  assign n2351 = n1873 & ~n2350 ;
  assign n2352 = n1877 & ~n2351 ;
  assign n2353 = n1881 & ~n2352 ;
  assign n2354 = n1885 & ~n2353 ;
  assign n2355 = n1889 & ~n2354 ;
  assign n2356 = n1893 & ~n2355 ;
  assign n2357 = n1897 & ~n2356 ;
  assign n2358 = n1901 & ~n2357 ;
  assign n2359 = n1905 & ~n2358 ;
  assign n2360 = n1909 & ~n2359 ;
  assign n2361 = n1913 & ~n2360 ;
  assign n2362 = n1917 & ~n2361 ;
  assign n2363 = n1921 & ~n2362 ;
  assign n2364 = n1925 & ~n2363 ;
  assign n2365 = n1929 & ~n2364 ;
  assign n2366 = n1933 & ~n2365 ;
  assign n2367 = n1937 & ~n2366 ;
  assign n2368 = n1010 & n1940 ;
  assign n2369 = ~n1939 & n2368 ;
  assign n2370 = ~n2367 & n2369 ;
  assign n2371 = ~n1005 & n1010 ;
  assign n2372 = n1601 & ~n2371 ;
  assign n2373 = ~n2370 & n2372 ;
  assign n2374 = n1014 & n2339 ;
  assign n2375 = ~n1603 & n2374 ;
  assign n2376 = ~n2373 & n2375 ;
  assign n2377 = ~n2340 & ~n2376 ;
  assign n2378 = \req[17]  & ~n308 ;
  assign n2379 = ~n294 & n2378 ;
  assign n2380 = ~\priority[19]  & ~n314 ;
  assign n2381 = n1042 & ~n2380 ;
  assign n2382 = n1956 & ~n2381 ;
  assign n2383 = n1961 & ~n2382 ;
  assign n2384 = n1965 & ~n2383 ;
  assign n2385 = n1969 & ~n2384 ;
  assign n2386 = n1973 & ~n2385 ;
  assign n2387 = n1977 & ~n2386 ;
  assign n2388 = n1981 & ~n2387 ;
  assign n2389 = n1985 & ~n2388 ;
  assign n2390 = n1989 & ~n2389 ;
  assign n2391 = n1993 & ~n2390 ;
  assign n2392 = n1997 & ~n2391 ;
  assign n2393 = n2001 & ~n2392 ;
  assign n2394 = n2005 & ~n2393 ;
  assign n2395 = n2009 & ~n2394 ;
  assign n2396 = n2013 & ~n2395 ;
  assign n2397 = n2017 & ~n2396 ;
  assign n2398 = n2021 & ~n2397 ;
  assign n2399 = n2025 & ~n2398 ;
  assign n2400 = n2029 & ~n2399 ;
  assign n2401 = n2033 & ~n2400 ;
  assign n2402 = n2037 & ~n2401 ;
  assign n2403 = n2041 & ~n2402 ;
  assign n2404 = n2045 & ~n2403 ;
  assign n2405 = n2049 & ~n2404 ;
  assign n2406 = n2053 & ~n2405 ;
  assign n2407 = n277 & n284 ;
  assign n2408 = ~n2055 & n2407 ;
  assign n2409 = ~n2406 & n2408 ;
  assign n2410 = ~n269 & n284 ;
  assign n2411 = n1717 & ~n2410 ;
  assign n2412 = ~n2409 & n2411 ;
  assign n2413 = n303 & n2378 ;
  assign n2414 = ~n1719 & n2413 ;
  assign n2415 = ~n2412 & n2414 ;
  assign n2416 = ~n2379 & ~n2415 ;
  assign n2417 = \req[18]  & ~n675 ;
  assign n2418 = ~n661 & n2417 ;
  assign n2419 = ~\priority[20]  & ~n681 ;
  assign n2420 = n306 & ~n2419 ;
  assign n2421 = n324 & ~n2420 ;
  assign n2422 = n338 & ~n2421 ;
  assign n2423 = n351 & ~n2422 ;
  assign n2424 = n364 & ~n2423 ;
  assign n2425 = n377 & ~n2424 ;
  assign n2426 = n390 & ~n2425 ;
  assign n2427 = n403 & ~n2426 ;
  assign n2428 = n416 & ~n2427 ;
  assign n2429 = n429 & ~n2428 ;
  assign n2430 = n442 & ~n2429 ;
  assign n2431 = n455 & ~n2430 ;
  assign n2432 = n468 & ~n2431 ;
  assign n2433 = n481 & ~n2432 ;
  assign n2434 = n494 & ~n2433 ;
  assign n2435 = n507 & ~n2434 ;
  assign n2436 = n520 & ~n2435 ;
  assign n2437 = n533 & ~n2436 ;
  assign n2438 = n546 & ~n2437 ;
  assign n2439 = n559 & ~n2438 ;
  assign n2440 = n572 & ~n2439 ;
  assign n2441 = n585 & ~n2440 ;
  assign n2442 = n598 & ~n2441 ;
  assign n2443 = n611 & ~n2442 ;
  assign n2444 = n2090 & ~n2443 ;
  assign n2445 = n2094 & ~n2444 ;
  assign n2446 = n644 & n651 ;
  assign n2447 = ~n2096 & n2446 ;
  assign n2448 = ~n2445 & n2447 ;
  assign n2449 = ~n636 & n651 ;
  assign n2450 = n1833 & ~n2449 ;
  assign n2451 = ~n2448 & n2450 ;
  assign n2452 = n670 & n2417 ;
  assign n2453 = ~n1835 & n2452 ;
  assign n2454 = ~n2451 & n2453 ;
  assign n2455 = ~n2418 & ~n2454 ;
  assign n2456 = \req[19]  & ~n1041 ;
  assign n2457 = ~n1027 & n2456 ;
  assign n2458 = ~\priority[21]  & ~n1047 ;
  assign n2459 = n673 & ~n2458 ;
  assign n2460 = n691 & ~n2459 ;
  assign n2461 = n705 & ~n2460 ;
  assign n2462 = n718 & ~n2461 ;
  assign n2463 = n731 & ~n2462 ;
  assign n2464 = n744 & ~n2463 ;
  assign n2465 = ~n749 & n756 ;
  assign n2466 = ~n2464 & n2465 ;
  assign n2467 = n770 & ~n2466 ;
  assign n2468 = n783 & ~n2467 ;
  assign n2469 = n796 & ~n2468 ;
  assign n2470 = n809 & ~n2469 ;
  assign n2471 = n2117 & ~n2470 ;
  assign n2472 = n835 & ~n2471 ;
  assign n2473 = n848 & ~n2472 ;
  assign n2474 = n861 & ~n2473 ;
  assign n2475 = n874 & ~n2474 ;
  assign n2476 = n887 & ~n2475 ;
  assign n2477 = n900 & ~n2476 ;
  assign n2478 = n913 & ~n2477 ;
  assign n2479 = n926 & ~n2478 ;
  assign n2480 = n939 & ~n2479 ;
  assign n2481 = n952 & ~n2480 ;
  assign n2482 = n965 & ~n2481 ;
  assign n2483 = n978 & ~n2482 ;
  assign n2484 = n2132 & ~n2483 ;
  assign n2485 = n2136 & ~n2484 ;
  assign n2486 = n1010 & n1017 ;
  assign n2487 = ~n2138 & n2486 ;
  assign n2488 = ~n2485 & n2487 ;
  assign n2489 = ~n1002 & n1017 ;
  assign n2490 = n1949 & ~n2489 ;
  assign n2491 = ~n2488 & n2490 ;
  assign n2492 = n1036 & n2456 ;
  assign n2493 = ~n1951 & n2492 ;
  assign n2494 = ~n2491 & n2493 ;
  assign n2495 = ~n2457 & ~n2494 ;
  assign n2496 = \req[20]  & ~n305 ;
  assign n2497 = ~n316 & n2496 ;
  assign n2498 = ~\priority[22]  & ~n321 ;
  assign n2499 = n1039 & ~n2498 ;
  assign n2500 = n1057 & ~n2499 ;
  assign n2501 = n1071 & ~n2500 ;
  assign n2502 = n1084 & ~n2501 ;
  assign n2503 = n1097 & ~n2502 ;
  assign n2504 = n1110 & ~n2503 ;
  assign n2505 = n1123 & ~n2504 ;
  assign n2506 = n1136 & ~n2505 ;
  assign n2507 = n1149 & ~n2506 ;
  assign n2508 = n1162 & ~n2507 ;
  assign n2509 = n1175 & ~n2508 ;
  assign n2510 = n1188 & ~n2509 ;
  assign n2511 = n1201 & ~n2510 ;
  assign n2512 = n1214 & ~n2511 ;
  assign n2513 = n1227 & ~n2512 ;
  assign n2514 = n1240 & ~n2513 ;
  assign n2515 = n1253 & ~n2514 ;
  assign n2516 = n1266 & ~n2515 ;
  assign n2517 = n1279 & ~n2516 ;
  assign n2518 = n1292 & ~n2517 ;
  assign n2519 = n1305 & ~n2518 ;
  assign n2520 = n1318 & ~n2519 ;
  assign n2521 = n1331 & ~n2520 ;
  assign n2522 = n1344 & ~n2521 ;
  assign n2523 = n2173 & ~n2522 ;
  assign n2524 = n2176 & ~n2523 ;
  assign n2525 = n286 & ~n2524 ;
  assign n2526 = n299 & ~n2525 ;
  assign n2527 = n310 & n2496 ;
  assign n2528 = ~n304 & n2527 ;
  assign n2529 = ~n2526 & n2528 ;
  assign n2530 = ~n2497 & ~n2529 ;
  assign n2531 = \req[21]  & ~n672 ;
  assign n2532 = ~n683 & n2531 ;
  assign n2533 = ~\priority[23]  & ~n688 ;
  assign n2534 = n328 & ~n2533 ;
  assign n2535 = n1379 & ~n2534 ;
  assign n2536 = n1384 & ~n2535 ;
  assign n2537 = n1388 & ~n2536 ;
  assign n2538 = n1392 & ~n2537 ;
  assign n2539 = n1396 & ~n2538 ;
  assign n2540 = n1400 & ~n2539 ;
  assign n2541 = n1404 & ~n2540 ;
  assign n2542 = n1408 & ~n2541 ;
  assign n2543 = n1412 & ~n2542 ;
  assign n2544 = n1416 & ~n2543 ;
  assign n2545 = n1420 & ~n2544 ;
  assign n2546 = n1424 & ~n2545 ;
  assign n2547 = n1428 & ~n2546 ;
  assign n2548 = n1432 & ~n2547 ;
  assign n2549 = n1436 & ~n2548 ;
  assign n2550 = n1440 & ~n2549 ;
  assign n2551 = n1444 & ~n2550 ;
  assign n2552 = n1448 & ~n2551 ;
  assign n2553 = n1452 & ~n2552 ;
  assign n2554 = n1456 & ~n2553 ;
  assign n2555 = n1460 & ~n2554 ;
  assign n2556 = n1464 & ~n2555 ;
  assign n2557 = n1468 & ~n2556 ;
  assign n2558 = n2212 & ~n2557 ;
  assign n2559 = n2215 & ~n2558 ;
  assign n2560 = n653 & ~n2559 ;
  assign n2561 = n666 & ~n2560 ;
  assign n2562 = n677 & n2531 ;
  assign n2563 = ~n671 & n2562 ;
  assign n2564 = ~n2561 & n2563 ;
  assign n2565 = ~n2532 & ~n2564 ;
  assign n2566 = \req[22]  & ~n1038 ;
  assign n2567 = ~n1049 & n2566 ;
  assign n2568 = ~\priority[24]  & ~n1054 ;
  assign n2569 = n695 & ~n2568 ;
  assign n2570 = n1499 & ~n2569 ;
  assign n2571 = n1504 & ~n2570 ;
  assign n2572 = n2229 & ~n2571 ;
  assign n2573 = n1512 & ~n2572 ;
  assign n2574 = n1516 & ~n2573 ;
  assign n2575 = n1520 & ~n2574 ;
  assign n2576 = n1524 & ~n2575 ;
  assign n2577 = n1528 & ~n2576 ;
  assign n2578 = n1532 & ~n2577 ;
  assign n2579 = n1536 & ~n2578 ;
  assign n2580 = n1540 & ~n2579 ;
  assign n2581 = n1544 & ~n2580 ;
  assign n2582 = n1548 & ~n2581 ;
  assign n2583 = n1552 & ~n2582 ;
  assign n2584 = n1556 & ~n2583 ;
  assign n2585 = n1560 & ~n2584 ;
  assign n2586 = n1564 & ~n2585 ;
  assign n2587 = n1568 & ~n2586 ;
  assign n2588 = n1572 & ~n2587 ;
  assign n2589 = n1576 & ~n2588 ;
  assign n2590 = n1580 & ~n2589 ;
  assign n2591 = n1584 & ~n2590 ;
  assign n2592 = n1588 & ~n2591 ;
  assign n2593 = n2252 & ~n2592 ;
  assign n2594 = n2255 & ~n2593 ;
  assign n2595 = n1019 & ~n2594 ;
  assign n2596 = n1032 & ~n2595 ;
  assign n2597 = n1043 & n2566 ;
  assign n2598 = ~n1037 & n2597 ;
  assign n2599 = ~n2596 & n2598 ;
  assign n2600 = ~n2567 & ~n2599 ;
  assign n2601 = \req[23]  & ~n327 ;
  assign n2602 = ~n323 & n2601 ;
  assign n2603 = ~\priority[25]  & ~n318 ;
  assign n2604 = n1061 & ~n2603 ;
  assign n2605 = n1616 & ~n2604 ;
  assign n2606 = n1621 & ~n2605 ;
  assign n2607 = n1625 & ~n2606 ;
  assign n2608 = n1629 & ~n2607 ;
  assign n2609 = n1633 & ~n2608 ;
  assign n2610 = n1637 & ~n2609 ;
  assign n2611 = n1641 & ~n2610 ;
  assign n2612 = n1645 & ~n2611 ;
  assign n2613 = n1649 & ~n2612 ;
  assign n2614 = n1653 & ~n2613 ;
  assign n2615 = n1657 & ~n2614 ;
  assign n2616 = n1661 & ~n2615 ;
  assign n2617 = n1665 & ~n2616 ;
  assign n2618 = n1669 & ~n2617 ;
  assign n2619 = n1673 & ~n2618 ;
  assign n2620 = n1677 & ~n2619 ;
  assign n2621 = n1681 & ~n2620 ;
  assign n2622 = n1685 & ~n2621 ;
  assign n2623 = n1689 & ~n2622 ;
  assign n2624 = n1693 & ~n2623 ;
  assign n2625 = n1697 & ~n2624 ;
  assign n2626 = n1701 & ~n2625 ;
  assign n2627 = n1705 & ~n2626 ;
  assign n2628 = n2291 & ~n2627 ;
  assign n2629 = n2294 & ~n2628 ;
  assign n2630 = n1368 & ~n2629 ;
  assign n2631 = n1372 & ~n2630 ;
  assign n2632 = n307 & n2601 ;
  assign n2633 = ~n1374 & n2632 ;
  assign n2634 = ~n2631 & n2633 ;
  assign n2635 = ~n2602 & ~n2634 ;
  assign n2636 = \req[24]  & ~n694 ;
  assign n2637 = ~n690 & n2636 ;
  assign n2638 = ~\priority[26]  & ~n685 ;
  assign n2639 = n335 & ~n2638 ;
  assign n2640 = n1732 & ~n2639 ;
  assign n2641 = n1737 & ~n2640 ;
  assign n2642 = n1741 & ~n2641 ;
  assign n2643 = n1745 & ~n2642 ;
  assign n2644 = n1749 & ~n2643 ;
  assign n2645 = n1753 & ~n2644 ;
  assign n2646 = n1757 & ~n2645 ;
  assign n2647 = n1761 & ~n2646 ;
  assign n2648 = n1765 & ~n2647 ;
  assign n2649 = n1769 & ~n2648 ;
  assign n2650 = n1773 & ~n2649 ;
  assign n2651 = n1777 & ~n2650 ;
  assign n2652 = n1781 & ~n2651 ;
  assign n2653 = n1785 & ~n2652 ;
  assign n2654 = n1789 & ~n2653 ;
  assign n2655 = n1793 & ~n2654 ;
  assign n2656 = n1797 & ~n2655 ;
  assign n2657 = n1801 & ~n2656 ;
  assign n2658 = n1805 & ~n2657 ;
  assign n2659 = n1809 & ~n2658 ;
  assign n2660 = n1813 & ~n2659 ;
  assign n2661 = n1817 & ~n2660 ;
  assign n2662 = n1821 & ~n2661 ;
  assign n2663 = n2330 & ~n2662 ;
  assign n2664 = n2333 & ~n2663 ;
  assign n2665 = n1488 & ~n2664 ;
  assign n2666 = n1492 & ~n2665 ;
  assign n2667 = n674 & n2636 ;
  assign n2668 = ~n1494 & n2667 ;
  assign n2669 = ~n2666 & n2668 ;
  assign n2670 = ~n2637 & ~n2669 ;
  assign n2671 = \req[25]  & ~n1060 ;
  assign n2672 = ~n1056 & n2671 ;
  assign n2673 = ~\priority[27]  & ~n1051 ;
  assign n2674 = n702 & ~n2673 ;
  assign n2675 = n1848 & ~n2674 ;
  assign n2676 = n1853 & ~n2675 ;
  assign n2677 = n1857 & ~n2676 ;
  assign n2678 = n1861 & ~n2677 ;
  assign n2679 = n1865 & ~n2678 ;
  assign n2680 = n1869 & ~n2679 ;
  assign n2681 = n1873 & ~n2680 ;
  assign n2682 = n1877 & ~n2681 ;
  assign n2683 = n1881 & ~n2682 ;
  assign n2684 = n1885 & ~n2683 ;
  assign n2685 = n1889 & ~n2684 ;
  assign n2686 = n1893 & ~n2685 ;
  assign n2687 = n1897 & ~n2686 ;
  assign n2688 = n1901 & ~n2687 ;
  assign n2689 = n1905 & ~n2688 ;
  assign n2690 = n1909 & ~n2689 ;
  assign n2691 = n1913 & ~n2690 ;
  assign n2692 = n1917 & ~n2691 ;
  assign n2693 = n1921 & ~n2692 ;
  assign n2694 = n1925 & ~n2693 ;
  assign n2695 = n1929 & ~n2694 ;
  assign n2696 = n1933 & ~n2695 ;
  assign n2697 = n1937 & ~n2696 ;
  assign n2698 = n2369 & ~n2697 ;
  assign n2699 = n2372 & ~n2698 ;
  assign n2700 = n1605 & ~n2699 ;
  assign n2701 = n1609 & ~n2700 ;
  assign n2702 = n1040 & n2671 ;
  assign n2703 = ~n1611 & n2702 ;
  assign n2704 = ~n2701 & n2703 ;
  assign n2705 = ~n2672 & ~n2704 ;
  assign n2706 = \req[26]  & ~n334 ;
  assign n2707 = ~n320 & n2706 ;
  assign n2708 = ~\priority[28]  & ~n340 ;
  assign n2709 = n1068 & ~n2708 ;
  assign n2710 = n1964 & ~n2709 ;
  assign n2711 = n1969 & ~n2710 ;
  assign n2712 = n1973 & ~n2711 ;
  assign n2713 = ~n1975 & n1976 ;
  assign n2714 = ~n2712 & n2713 ;
  assign n2715 = n1981 & ~n2714 ;
  assign n2716 = n1985 & ~n2715 ;
  assign n2717 = n1989 & ~n2716 ;
  assign n2718 = n1993 & ~n2717 ;
  assign n2719 = n1997 & ~n2718 ;
  assign n2720 = n2001 & ~n2719 ;
  assign n2721 = n2005 & ~n2720 ;
  assign n2722 = n2009 & ~n2721 ;
  assign n2723 = n2013 & ~n2722 ;
  assign n2724 = n2017 & ~n2723 ;
  assign n2725 = n2021 & ~n2724 ;
  assign n2726 = n2025 & ~n2725 ;
  assign n2727 = n2029 & ~n2726 ;
  assign n2728 = n2033 & ~n2727 ;
  assign n2729 = n2037 & ~n2728 ;
  assign n2730 = n2041 & ~n2729 ;
  assign n2731 = n2045 & ~n2730 ;
  assign n2732 = n2049 & ~n2731 ;
  assign n2733 = n2053 & ~n2732 ;
  assign n2734 = n2408 & ~n2733 ;
  assign n2735 = n2411 & ~n2734 ;
  assign n2736 = n1721 & ~n2735 ;
  assign n2737 = n1725 & ~n2736 ;
  assign n2738 = n329 & n2706 ;
  assign n2739 = ~n1727 & n2738 ;
  assign n2740 = ~n2737 & n2739 ;
  assign n2741 = ~n2707 & ~n2740 ;
  assign n2742 = \req[27]  & ~n701 ;
  assign n2743 = ~n687 & n2742 ;
  assign n2744 = ~\priority[29]  & ~n707 ;
  assign n2745 = n332 & ~n2744 ;
  assign n2746 = n350 & ~n2745 ;
  assign n2747 = n364 & ~n2746 ;
  assign n2748 = n377 & ~n2747 ;
  assign n2749 = n390 & ~n2748 ;
  assign n2750 = n403 & ~n2749 ;
  assign n2751 = n416 & ~n2750 ;
  assign n2752 = n429 & ~n2751 ;
  assign n2753 = n442 & ~n2752 ;
  assign n2754 = n455 & ~n2753 ;
  assign n2755 = n468 & ~n2754 ;
  assign n2756 = n481 & ~n2755 ;
  assign n2757 = n494 & ~n2756 ;
  assign n2758 = n507 & ~n2757 ;
  assign n2759 = n520 & ~n2758 ;
  assign n2760 = n533 & ~n2759 ;
  assign n2761 = n546 & ~n2760 ;
  assign n2762 = n559 & ~n2761 ;
  assign n2763 = n572 & ~n2762 ;
  assign n2764 = n585 & ~n2763 ;
  assign n2765 = n598 & ~n2764 ;
  assign n2766 = n611 & ~n2765 ;
  assign n2767 = n2090 & ~n2766 ;
  assign n2768 = n2094 & ~n2767 ;
  assign n2769 = n2447 & ~n2768 ;
  assign n2770 = n2450 & ~n2769 ;
  assign n2771 = n1837 & ~n2770 ;
  assign n2772 = n1841 & ~n2771 ;
  assign n2773 = n696 & n2742 ;
  assign n2774 = ~n1843 & n2773 ;
  assign n2775 = ~n2772 & n2774 ;
  assign n2776 = ~n2743 & ~n2775 ;
  assign n2777 = \req[28]  & ~n1067 ;
  assign n2778 = ~n1053 & n2777 ;
  assign n2779 = ~\priority[30]  & ~n1073 ;
  assign n2780 = n699 & ~n2779 ;
  assign n2781 = n717 & ~n2780 ;
  assign n2782 = n731 & ~n2781 ;
  assign n2783 = n744 & ~n2782 ;
  assign n2784 = n2465 & ~n2783 ;
  assign n2785 = n770 & ~n2784 ;
  assign n2786 = n783 & ~n2785 ;
  assign n2787 = n796 & ~n2786 ;
  assign n2788 = n809 & ~n2787 ;
  assign n2789 = n2117 & ~n2788 ;
  assign n2790 = n835 & ~n2789 ;
  assign n2791 = n848 & ~n2790 ;
  assign n2792 = n861 & ~n2791 ;
  assign n2793 = n874 & ~n2792 ;
  assign n2794 = n887 & ~n2793 ;
  assign n2795 = n900 & ~n2794 ;
  assign n2796 = n913 & ~n2795 ;
  assign n2797 = n926 & ~n2796 ;
  assign n2798 = n939 & ~n2797 ;
  assign n2799 = n952 & ~n2798 ;
  assign n2800 = n965 & ~n2799 ;
  assign n2801 = n978 & ~n2800 ;
  assign n2802 = n2132 & ~n2801 ;
  assign n2803 = n2136 & ~n2802 ;
  assign n2804 = n2487 & ~n2803 ;
  assign n2805 = n2490 & ~n2804 ;
  assign n2806 = n1953 & ~n2805 ;
  assign n2807 = n1957 & ~n2806 ;
  assign n2808 = n1062 & n2777 ;
  assign n2809 = ~n1959 & n2808 ;
  assign n2810 = ~n2807 & n2809 ;
  assign n2811 = ~n2778 & ~n2810 ;
  assign n2812 = \req[29]  & ~n331 ;
  assign n2813 = ~n342 & n2812 ;
  assign n2814 = ~\priority[31]  & ~n347 ;
  assign n2815 = n1065 & ~n2814 ;
  assign n2816 = n1083 & ~n2815 ;
  assign n2817 = n1097 & ~n2816 ;
  assign n2818 = n1110 & ~n2817 ;
  assign n2819 = n1123 & ~n2818 ;
  assign n2820 = n1136 & ~n2819 ;
  assign n2821 = n1149 & ~n2820 ;
  assign n2822 = n1162 & ~n2821 ;
  assign n2823 = n1175 & ~n2822 ;
  assign n2824 = n1188 & ~n2823 ;
  assign n2825 = n1201 & ~n2824 ;
  assign n2826 = n1214 & ~n2825 ;
  assign n2827 = n1227 & ~n2826 ;
  assign n2828 = n1240 & ~n2827 ;
  assign n2829 = n1253 & ~n2828 ;
  assign n2830 = n1266 & ~n2829 ;
  assign n2831 = n1279 & ~n2830 ;
  assign n2832 = n1292 & ~n2831 ;
  assign n2833 = n1305 & ~n2832 ;
  assign n2834 = n1318 & ~n2833 ;
  assign n2835 = n1331 & ~n2834 ;
  assign n2836 = n1344 & ~n2835 ;
  assign n2837 = n2173 & ~n2836 ;
  assign n2838 = n2176 & ~n2837 ;
  assign n2839 = n286 & ~n2838 ;
  assign n2840 = n299 & ~n2839 ;
  assign n2841 = n312 & ~n2840 ;
  assign n2842 = n325 & ~n2841 ;
  assign n2843 = n336 & n2812 ;
  assign n2844 = ~n330 & n2843 ;
  assign n2845 = ~n2842 & n2844 ;
  assign n2846 = ~n2813 & ~n2845 ;
  assign n2847 = \req[30]  & ~n698 ;
  assign n2848 = ~n709 & n2847 ;
  assign n2849 = ~\priority[32]  & ~n714 ;
  assign n2850 = n354 & ~n2849 ;
  assign n2851 = n1387 & ~n2850 ;
  assign n2852 = n1392 & ~n2851 ;
  assign n2853 = n1396 & ~n2852 ;
  assign n2854 = n1400 & ~n2853 ;
  assign n2855 = n1404 & ~n2854 ;
  assign n2856 = n1408 & ~n2855 ;
  assign n2857 = n1412 & ~n2856 ;
  assign n2858 = n1416 & ~n2857 ;
  assign n2859 = n1420 & ~n2858 ;
  assign n2860 = n1424 & ~n2859 ;
  assign n2861 = n1428 & ~n2860 ;
  assign n2862 = n1432 & ~n2861 ;
  assign n2863 = n1436 & ~n2862 ;
  assign n2864 = n1440 & ~n2863 ;
  assign n2865 = n1444 & ~n2864 ;
  assign n2866 = n1448 & ~n2865 ;
  assign n2867 = n1452 & ~n2866 ;
  assign n2868 = n1456 & ~n2867 ;
  assign n2869 = n1460 & ~n2868 ;
  assign n2870 = n1464 & ~n2869 ;
  assign n2871 = n1468 & ~n2870 ;
  assign n2872 = n2212 & ~n2871 ;
  assign n2873 = n2215 & ~n2872 ;
  assign n2874 = n653 & ~n2873 ;
  assign n2875 = n666 & ~n2874 ;
  assign n2876 = n679 & ~n2875 ;
  assign n2877 = n692 & ~n2876 ;
  assign n2878 = n703 & n2847 ;
  assign n2879 = ~n697 & n2878 ;
  assign n2880 = ~n2877 & n2879 ;
  assign n2881 = ~n2848 & ~n2880 ;
  assign n2882 = \req[31]  & ~n1064 ;
  assign n2883 = ~n1075 & n2882 ;
  assign n2884 = ~\priority[33]  & ~n1080 ;
  assign n2885 = n721 & ~n2884 ;
  assign n2886 = n1507 & ~n2885 ;
  assign n2887 = n1512 & ~n2886 ;
  assign n2888 = n1516 & ~n2887 ;
  assign n2889 = n1520 & ~n2888 ;
  assign n2890 = n1524 & ~n2889 ;
  assign n2891 = n1528 & ~n2890 ;
  assign n2892 = n1532 & ~n2891 ;
  assign n2893 = n1536 & ~n2892 ;
  assign n2894 = n1540 & ~n2893 ;
  assign n2895 = n1544 & ~n2894 ;
  assign n2896 = n1548 & ~n2895 ;
  assign n2897 = n1552 & ~n2896 ;
  assign n2898 = n1556 & ~n2897 ;
  assign n2899 = n1560 & ~n2898 ;
  assign n2900 = n1564 & ~n2899 ;
  assign n2901 = n1568 & ~n2900 ;
  assign n2902 = n1572 & ~n2901 ;
  assign n2903 = n1576 & ~n2902 ;
  assign n2904 = n1580 & ~n2903 ;
  assign n2905 = n1584 & ~n2904 ;
  assign n2906 = n1588 & ~n2905 ;
  assign n2907 = n2252 & ~n2906 ;
  assign n2908 = n2255 & ~n2907 ;
  assign n2909 = n1019 & ~n2908 ;
  assign n2910 = n1032 & ~n2909 ;
  assign n2911 = n1045 & ~n2910 ;
  assign n2912 = n1058 & ~n2911 ;
  assign n2913 = n1069 & n2882 ;
  assign n2914 = ~n1063 & n2913 ;
  assign n2915 = ~n2912 & n2914 ;
  assign n2916 = ~n2883 & ~n2915 ;
  assign n2917 = \req[32]  & ~n353 ;
  assign n2918 = ~n349 & n2917 ;
  assign n2919 = ~\priority[34]  & ~n344 ;
  assign n2920 = n1087 & ~n2919 ;
  assign n2921 = n1624 & ~n2920 ;
  assign n2922 = n1629 & ~n2921 ;
  assign n2923 = n1633 & ~n2922 ;
  assign n2924 = n1637 & ~n2923 ;
  assign n2925 = n1641 & ~n2924 ;
  assign n2926 = n1645 & ~n2925 ;
  assign n2927 = n1649 & ~n2926 ;
  assign n2928 = n1653 & ~n2927 ;
  assign n2929 = n1657 & ~n2928 ;
  assign n2930 = n1661 & ~n2929 ;
  assign n2931 = n1665 & ~n2930 ;
  assign n2932 = n1669 & ~n2931 ;
  assign n2933 = n1673 & ~n2932 ;
  assign n2934 = n1677 & ~n2933 ;
  assign n2935 = n1681 & ~n2934 ;
  assign n2936 = n1685 & ~n2935 ;
  assign n2937 = n1689 & ~n2936 ;
  assign n2938 = n1693 & ~n2937 ;
  assign n2939 = n1697 & ~n2938 ;
  assign n2940 = n1701 & ~n2939 ;
  assign n2941 = n1705 & ~n2940 ;
  assign n2942 = n2291 & ~n2941 ;
  assign n2943 = n2294 & ~n2942 ;
  assign n2944 = n1368 & ~n2943 ;
  assign n2945 = n1372 & ~n2944 ;
  assign n2946 = n1376 & ~n2945 ;
  assign n2947 = n1380 & ~n2946 ;
  assign n2948 = n333 & n2917 ;
  assign n2949 = ~n1382 & n2948 ;
  assign n2950 = ~n2947 & n2949 ;
  assign n2951 = ~n2918 & ~n2950 ;
  assign n2952 = \req[33]  & ~n720 ;
  assign n2953 = ~n716 & n2952 ;
  assign n2954 = ~\priority[35]  & ~n711 ;
  assign n2955 = n361 & ~n2954 ;
  assign n2956 = n1740 & ~n2955 ;
  assign n2957 = n1745 & ~n2956 ;
  assign n2958 = n1749 & ~n2957 ;
  assign n2959 = n1753 & ~n2958 ;
  assign n2960 = n1757 & ~n2959 ;
  assign n2961 = n1761 & ~n2960 ;
  assign n2962 = n1765 & ~n2961 ;
  assign n2963 = n1769 & ~n2962 ;
  assign n2964 = n1773 & ~n2963 ;
  assign n2965 = n1777 & ~n2964 ;
  assign n2966 = n1781 & ~n2965 ;
  assign n2967 = n1785 & ~n2966 ;
  assign n2968 = n1789 & ~n2967 ;
  assign n2969 = n1793 & ~n2968 ;
  assign n2970 = n1797 & ~n2969 ;
  assign n2971 = n1801 & ~n2970 ;
  assign n2972 = n1805 & ~n2971 ;
  assign n2973 = n1809 & ~n2972 ;
  assign n2974 = n1813 & ~n2973 ;
  assign n2975 = n1817 & ~n2974 ;
  assign n2976 = n1821 & ~n2975 ;
  assign n2977 = n2330 & ~n2976 ;
  assign n2978 = n2333 & ~n2977 ;
  assign n2979 = n1488 & ~n2978 ;
  assign n2980 = n1492 & ~n2979 ;
  assign n2981 = n1496 & ~n2980 ;
  assign n2982 = n1500 & ~n2981 ;
  assign n2983 = n700 & n2952 ;
  assign n2984 = ~n1502 & n2983 ;
  assign n2985 = ~n2982 & n2984 ;
  assign n2986 = ~n2953 & ~n2985 ;
  assign n2987 = \req[34]  & ~n1086 ;
  assign n2988 = ~n1082 & n2987 ;
  assign n2989 = ~\priority[36]  & ~n1077 ;
  assign n2990 = n728 & ~n2989 ;
  assign n2991 = n1856 & ~n2990 ;
  assign n2992 = n1861 & ~n2991 ;
  assign n2993 = n1865 & ~n2992 ;
  assign n2994 = n1869 & ~n2993 ;
  assign n2995 = n1873 & ~n2994 ;
  assign n2996 = n1877 & ~n2995 ;
  assign n2997 = n1881 & ~n2996 ;
  assign n2998 = n1885 & ~n2997 ;
  assign n2999 = n1889 & ~n2998 ;
  assign n3000 = n1893 & ~n2999 ;
  assign n3001 = n1897 & ~n3000 ;
  assign n3002 = n1901 & ~n3001 ;
  assign n3003 = n1905 & ~n3002 ;
  assign n3004 = n1909 & ~n3003 ;
  assign n3005 = n1913 & ~n3004 ;
  assign n3006 = n1917 & ~n3005 ;
  assign n3007 = n1921 & ~n3006 ;
  assign n3008 = n1925 & ~n3007 ;
  assign n3009 = n1929 & ~n3008 ;
  assign n3010 = n1933 & ~n3009 ;
  assign n3011 = n1937 & ~n3010 ;
  assign n3012 = n2369 & ~n3011 ;
  assign n3013 = n2372 & ~n3012 ;
  assign n3014 = n1605 & ~n3013 ;
  assign n3015 = n1609 & ~n3014 ;
  assign n3016 = n1613 & ~n3015 ;
  assign n3017 = n1617 & ~n3016 ;
  assign n3018 = n1066 & n2987 ;
  assign n3019 = ~n1619 & n3018 ;
  assign n3020 = ~n3017 & n3019 ;
  assign n3021 = ~n2988 & ~n3020 ;
  assign n3022 = \req[35]  & ~n360 ;
  assign n3023 = ~n346 & n3022 ;
  assign n3024 = ~\priority[37]  & ~n366 ;
  assign n3025 = n1094 & ~n3024 ;
  assign n3026 = n1972 & ~n3025 ;
  assign n3027 = n2713 & ~n3026 ;
  assign n3028 = n1981 & ~n3027 ;
  assign n3029 = n1985 & ~n3028 ;
  assign n3030 = n1989 & ~n3029 ;
  assign n3031 = n1993 & ~n3030 ;
  assign n3032 = n1997 & ~n3031 ;
  assign n3033 = n2001 & ~n3032 ;
  assign n3034 = n2005 & ~n3033 ;
  assign n3035 = n2009 & ~n3034 ;
  assign n3036 = n2013 & ~n3035 ;
  assign n3037 = n2017 & ~n3036 ;
  assign n3038 = n2021 & ~n3037 ;
  assign n3039 = n2025 & ~n3038 ;
  assign n3040 = n2029 & ~n3039 ;
  assign n3041 = n2033 & ~n3040 ;
  assign n3042 = n2037 & ~n3041 ;
  assign n3043 = n2041 & ~n3042 ;
  assign n3044 = n2045 & ~n3043 ;
  assign n3045 = n2049 & ~n3044 ;
  assign n3046 = n2053 & ~n3045 ;
  assign n3047 = n2408 & ~n3046 ;
  assign n3048 = n2411 & ~n3047 ;
  assign n3049 = n1721 & ~n3048 ;
  assign n3050 = n1725 & ~n3049 ;
  assign n3051 = n1729 & ~n3050 ;
  assign n3052 = n1733 & ~n3051 ;
  assign n3053 = n355 & n3022 ;
  assign n3054 = ~n1735 & n3053 ;
  assign n3055 = ~n3052 & n3054 ;
  assign n3056 = ~n3023 & ~n3055 ;
  assign n3057 = \req[36]  & ~n727 ;
  assign n3058 = ~n713 & n3057 ;
  assign n3059 = ~\priority[38]  & ~n733 ;
  assign n3060 = n358 & ~n3059 ;
  assign n3061 = n376 & ~n3060 ;
  assign n3062 = n390 & ~n3061 ;
  assign n3063 = n403 & ~n3062 ;
  assign n3064 = n416 & ~n3063 ;
  assign n3065 = n429 & ~n3064 ;
  assign n3066 = n442 & ~n3065 ;
  assign n3067 = n455 & ~n3066 ;
  assign n3068 = n468 & ~n3067 ;
  assign n3069 = n481 & ~n3068 ;
  assign n3070 = n494 & ~n3069 ;
  assign n3071 = n507 & ~n3070 ;
  assign n3072 = n520 & ~n3071 ;
  assign n3073 = n533 & ~n3072 ;
  assign n3074 = n546 & ~n3073 ;
  assign n3075 = n559 & ~n3074 ;
  assign n3076 = n572 & ~n3075 ;
  assign n3077 = n585 & ~n3076 ;
  assign n3078 = n598 & ~n3077 ;
  assign n3079 = n611 & ~n3078 ;
  assign n3080 = n2090 & ~n3079 ;
  assign n3081 = n2094 & ~n3080 ;
  assign n3082 = n2447 & ~n3081 ;
  assign n3083 = n2450 & ~n3082 ;
  assign n3084 = n1837 & ~n3083 ;
  assign n3085 = n1841 & ~n3084 ;
  assign n3086 = n1845 & ~n3085 ;
  assign n3087 = n1849 & ~n3086 ;
  assign n3088 = n722 & n3057 ;
  assign n3089 = ~n1851 & n3088 ;
  assign n3090 = ~n3087 & n3089 ;
  assign n3091 = ~n3058 & ~n3090 ;
  assign n3092 = \req[37]  & ~n1093 ;
  assign n3093 = ~n1079 & n3092 ;
  assign n3094 = ~\priority[39]  & ~n1099 ;
  assign n3095 = n725 & ~n3094 ;
  assign n3096 = n743 & ~n3095 ;
  assign n3097 = n2465 & ~n3096 ;
  assign n3098 = n770 & ~n3097 ;
  assign n3099 = ~n775 & n782 ;
  assign n3100 = ~n3098 & n3099 ;
  assign n3101 = n796 & ~n3100 ;
  assign n3102 = n809 & ~n3101 ;
  assign n3103 = n2117 & ~n3102 ;
  assign n3104 = n835 & ~n3103 ;
  assign n3105 = n848 & ~n3104 ;
  assign n3106 = n861 & ~n3105 ;
  assign n3107 = n874 & ~n3106 ;
  assign n3108 = n887 & ~n3107 ;
  assign n3109 = n900 & ~n3108 ;
  assign n3110 = n913 & ~n3109 ;
  assign n3111 = n926 & ~n3110 ;
  assign n3112 = n939 & ~n3111 ;
  assign n3113 = n952 & ~n3112 ;
  assign n3114 = n965 & ~n3113 ;
  assign n3115 = n978 & ~n3114 ;
  assign n3116 = n2132 & ~n3115 ;
  assign n3117 = n2136 & ~n3116 ;
  assign n3118 = n2487 & ~n3117 ;
  assign n3119 = n2490 & ~n3118 ;
  assign n3120 = n1953 & ~n3119 ;
  assign n3121 = n1957 & ~n3120 ;
  assign n3122 = n1961 & ~n3121 ;
  assign n3123 = n1965 & ~n3122 ;
  assign n3124 = n1088 & n3092 ;
  assign n3125 = ~n1967 & n3124 ;
  assign n3126 = ~n3123 & n3125 ;
  assign n3127 = ~n3093 & ~n3126 ;
  assign n3128 = \req[38]  & ~n357 ;
  assign n3129 = ~n368 & n3128 ;
  assign n3130 = ~\priority[40]  & ~n373 ;
  assign n3131 = n1091 & ~n3130 ;
  assign n3132 = n1109 & ~n3131 ;
  assign n3133 = n1123 & ~n3132 ;
  assign n3134 = n1136 & ~n3133 ;
  assign n3135 = n1149 & ~n3134 ;
  assign n3136 = n1162 & ~n3135 ;
  assign n3137 = n1175 & ~n3136 ;
  assign n3138 = n1188 & ~n3137 ;
  assign n3139 = n1201 & ~n3138 ;
  assign n3140 = n1214 & ~n3139 ;
  assign n3141 = n1227 & ~n3140 ;
  assign n3142 = n1240 & ~n3141 ;
  assign n3143 = n1253 & ~n3142 ;
  assign n3144 = n1266 & ~n3143 ;
  assign n3145 = n1279 & ~n3144 ;
  assign n3146 = n1292 & ~n3145 ;
  assign n3147 = n1305 & ~n3146 ;
  assign n3148 = ~n1310 & n1317 ;
  assign n3149 = ~n3147 & n3148 ;
  assign n3150 = n1331 & ~n3149 ;
  assign n3151 = n1344 & ~n3150 ;
  assign n3152 = n2173 & ~n3151 ;
  assign n3153 = n2176 & ~n3152 ;
  assign n3154 = n286 & ~n3153 ;
  assign n3155 = n299 & ~n3154 ;
  assign n3156 = n312 & ~n3155 ;
  assign n3157 = n325 & ~n3156 ;
  assign n3158 = n338 & ~n3157 ;
  assign n3159 = n351 & ~n3158 ;
  assign n3160 = n362 & n3128 ;
  assign n3161 = ~n356 & n3160 ;
  assign n3162 = ~n3159 & n3161 ;
  assign n3163 = ~n3129 & ~n3162 ;
  assign n3164 = \req[39]  & ~n724 ;
  assign n3165 = ~n735 & n3164 ;
  assign n3166 = ~\priority[41]  & ~n740 ;
  assign n3167 = n380 & ~n3166 ;
  assign n3168 = n1395 & ~n3167 ;
  assign n3169 = n1400 & ~n3168 ;
  assign n3170 = n1404 & ~n3169 ;
  assign n3171 = n1408 & ~n3170 ;
  assign n3172 = n1412 & ~n3171 ;
  assign n3173 = n1416 & ~n3172 ;
  assign n3174 = n1420 & ~n3173 ;
  assign n3175 = n1424 & ~n3174 ;
  assign n3176 = n1428 & ~n3175 ;
  assign n3177 = n1432 & ~n3176 ;
  assign n3178 = n1436 & ~n3177 ;
  assign n3179 = n1440 & ~n3178 ;
  assign n3180 = n1444 & ~n3179 ;
  assign n3181 = n1448 & ~n3180 ;
  assign n3182 = n1452 & ~n3181 ;
  assign n3183 = n1456 & ~n3182 ;
  assign n3184 = n1460 & ~n3183 ;
  assign n3185 = n1464 & ~n3184 ;
  assign n3186 = n1468 & ~n3185 ;
  assign n3187 = n2212 & ~n3186 ;
  assign n3188 = n2215 & ~n3187 ;
  assign n3189 = n653 & ~n3188 ;
  assign n3190 = n666 & ~n3189 ;
  assign n3191 = n679 & ~n3190 ;
  assign n3192 = n692 & ~n3191 ;
  assign n3193 = n705 & ~n3192 ;
  assign n3194 = n718 & ~n3193 ;
  assign n3195 = n729 & n3164 ;
  assign n3196 = ~n723 & n3195 ;
  assign n3197 = ~n3194 & n3196 ;
  assign n3198 = ~n3165 & ~n3197 ;
  assign n3199 = \req[40]  & ~n1090 ;
  assign n3200 = ~n1101 & n3199 ;
  assign n3201 = ~\priority[42]  & ~n1106 ;
  assign n3202 = n747 & ~n3201 ;
  assign n3203 = n1515 & ~n3202 ;
  assign n3204 = n1520 & ~n3203 ;
  assign n3205 = n1524 & ~n3204 ;
  assign n3206 = n1528 & ~n3205 ;
  assign n3207 = n1532 & ~n3206 ;
  assign n3208 = n1536 & ~n3207 ;
  assign n3209 = n1540 & ~n3208 ;
  assign n3210 = n1544 & ~n3209 ;
  assign n3211 = n1548 & ~n3210 ;
  assign n3212 = n1552 & ~n3211 ;
  assign n3213 = n1556 & ~n3212 ;
  assign n3214 = n1560 & ~n3213 ;
  assign n3215 = n1564 & ~n3214 ;
  assign n3216 = n1568 & ~n3215 ;
  assign n3217 = n1572 & ~n3216 ;
  assign n3218 = n1576 & ~n3217 ;
  assign n3219 = n1580 & ~n3218 ;
  assign n3220 = n1584 & ~n3219 ;
  assign n3221 = n1588 & ~n3220 ;
  assign n3222 = n2252 & ~n3221 ;
  assign n3223 = n2255 & ~n3222 ;
  assign n3224 = n1019 & ~n3223 ;
  assign n3225 = n1032 & ~n3224 ;
  assign n3226 = n1045 & ~n3225 ;
  assign n3227 = n1058 & ~n3226 ;
  assign n3228 = n1071 & ~n3227 ;
  assign n3229 = n1084 & ~n3228 ;
  assign n3230 = n1095 & n3199 ;
  assign n3231 = ~n1089 & n3230 ;
  assign n3232 = ~n3229 & n3231 ;
  assign n3233 = ~n3200 & ~n3232 ;
  assign n3234 = \req[41]  & ~n379 ;
  assign n3235 = ~n375 & n3234 ;
  assign n3236 = ~\priority[43]  & ~n370 ;
  assign n3237 = n1113 & ~n3236 ;
  assign n3238 = n1632 & ~n3237 ;
  assign n3239 = n1637 & ~n3238 ;
  assign n3240 = n1641 & ~n3239 ;
  assign n3241 = n1645 & ~n3240 ;
  assign n3242 = n1649 & ~n3241 ;
  assign n3243 = n1653 & ~n3242 ;
  assign n3244 = n1657 & ~n3243 ;
  assign n3245 = n1661 & ~n3244 ;
  assign n3246 = n1665 & ~n3245 ;
  assign n3247 = n1669 & ~n3246 ;
  assign n3248 = n1673 & ~n3247 ;
  assign n3249 = n1677 & ~n3248 ;
  assign n3250 = n1681 & ~n3249 ;
  assign n3251 = n1685 & ~n3250 ;
  assign n3252 = n1689 & ~n3251 ;
  assign n3253 = n1693 & ~n3252 ;
  assign n3254 = n1697 & ~n3253 ;
  assign n3255 = n1701 & ~n3254 ;
  assign n3256 = n1705 & ~n3255 ;
  assign n3257 = n2291 & ~n3256 ;
  assign n3258 = n2294 & ~n3257 ;
  assign n3259 = n1368 & ~n3258 ;
  assign n3260 = n1372 & ~n3259 ;
  assign n3261 = n1376 & ~n3260 ;
  assign n3262 = n1380 & ~n3261 ;
  assign n3263 = n1384 & ~n3262 ;
  assign n3264 = n1388 & ~n3263 ;
  assign n3265 = n359 & n3234 ;
  assign n3266 = ~n1390 & n3265 ;
  assign n3267 = ~n3264 & n3266 ;
  assign n3268 = ~n3235 & ~n3267 ;
  assign n3269 = \req[42]  & ~n746 ;
  assign n3270 = ~n742 & n3269 ;
  assign n3271 = ~\priority[44]  & ~n737 ;
  assign n3272 = n387 & ~n3271 ;
  assign n3273 = n1748 & ~n3272 ;
  assign n3274 = n1753 & ~n3273 ;
  assign n3275 = n1757 & ~n3274 ;
  assign n3276 = n1761 & ~n3275 ;
  assign n3277 = n1765 & ~n3276 ;
  assign n3278 = n1769 & ~n3277 ;
  assign n3279 = n1773 & ~n3278 ;
  assign n3280 = n1777 & ~n3279 ;
  assign n3281 = n1781 & ~n3280 ;
  assign n3282 = n1785 & ~n3281 ;
  assign n3283 = n1789 & ~n3282 ;
  assign n3284 = n1793 & ~n3283 ;
  assign n3285 = n1797 & ~n3284 ;
  assign n3286 = n1801 & ~n3285 ;
  assign n3287 = n1805 & ~n3286 ;
  assign n3288 = n1809 & ~n3287 ;
  assign n3289 = n1813 & ~n3288 ;
  assign n3290 = n1817 & ~n3289 ;
  assign n3291 = n1821 & ~n3290 ;
  assign n3292 = n2330 & ~n3291 ;
  assign n3293 = n2333 & ~n3292 ;
  assign n3294 = n1488 & ~n3293 ;
  assign n3295 = n1492 & ~n3294 ;
  assign n3296 = n1496 & ~n3295 ;
  assign n3297 = n1500 & ~n3296 ;
  assign n3298 = n1504 & ~n3297 ;
  assign n3299 = n2229 & ~n3298 ;
  assign n3300 = n726 & n3269 ;
  assign n3301 = ~n1510 & n3300 ;
  assign n3302 = ~n3299 & n3301 ;
  assign n3303 = ~n3270 & ~n3302 ;
  assign n3304 = \req[43]  & ~n1112 ;
  assign n3305 = ~n1108 & n3304 ;
  assign n3306 = ~\priority[45]  & ~n1103 ;
  assign n3307 = n754 & ~n3306 ;
  assign n3308 = n1864 & ~n3307 ;
  assign n3309 = n1869 & ~n3308 ;
  assign n3310 = n1873 & ~n3309 ;
  assign n3311 = n1877 & ~n3310 ;
  assign n3312 = n1881 & ~n3311 ;
  assign n3313 = n1885 & ~n3312 ;
  assign n3314 = n1889 & ~n3313 ;
  assign n3315 = n1893 & ~n3314 ;
  assign n3316 = n1897 & ~n3315 ;
  assign n3317 = n1901 & ~n3316 ;
  assign n3318 = n1905 & ~n3317 ;
  assign n3319 = n1909 & ~n3318 ;
  assign n3320 = n1913 & ~n3319 ;
  assign n3321 = n1917 & ~n3320 ;
  assign n3322 = n1921 & ~n3321 ;
  assign n3323 = n1925 & ~n3322 ;
  assign n3324 = n1929 & ~n3323 ;
  assign n3325 = n1933 & ~n3324 ;
  assign n3326 = n1937 & ~n3325 ;
  assign n3327 = n2369 & ~n3326 ;
  assign n3328 = n2372 & ~n3327 ;
  assign n3329 = n1605 & ~n3328 ;
  assign n3330 = n1609 & ~n3329 ;
  assign n3331 = n1613 & ~n3330 ;
  assign n3332 = n1617 & ~n3331 ;
  assign n3333 = n1621 & ~n3332 ;
  assign n3334 = n1625 & ~n3333 ;
  assign n3335 = n1092 & n3304 ;
  assign n3336 = ~n1627 & n3335 ;
  assign n3337 = ~n3334 & n3336 ;
  assign n3338 = ~n3305 & ~n3337 ;
  assign n3339 = \req[44]  & ~n386 ;
  assign n3340 = ~n372 & n3339 ;
  assign n3341 = ~\priority[46]  & ~n392 ;
  assign n3342 = n1120 & ~n3341 ;
  assign n3343 = n1980 & ~n3342 ;
  assign n3344 = n1985 & ~n3343 ;
  assign n3345 = n1989 & ~n3344 ;
  assign n3346 = n1993 & ~n3345 ;
  assign n3347 = n1997 & ~n3346 ;
  assign n3348 = n2001 & ~n3347 ;
  assign n3349 = n2005 & ~n3348 ;
  assign n3350 = n2009 & ~n3349 ;
  assign n3351 = n2013 & ~n3350 ;
  assign n3352 = n2017 & ~n3351 ;
  assign n3353 = n2021 & ~n3352 ;
  assign n3354 = n2025 & ~n3353 ;
  assign n3355 = n2029 & ~n3354 ;
  assign n3356 = n2033 & ~n3355 ;
  assign n3357 = n2037 & ~n3356 ;
  assign n3358 = n2041 & ~n3357 ;
  assign n3359 = n2045 & ~n3358 ;
  assign n3360 = n2049 & ~n3359 ;
  assign n3361 = n2053 & ~n3360 ;
  assign n3362 = n2408 & ~n3361 ;
  assign n3363 = n2411 & ~n3362 ;
  assign n3364 = n1721 & ~n3363 ;
  assign n3365 = n1725 & ~n3364 ;
  assign n3366 = n1729 & ~n3365 ;
  assign n3367 = n1733 & ~n3366 ;
  assign n3368 = n1737 & ~n3367 ;
  assign n3369 = n1741 & ~n3368 ;
  assign n3370 = n381 & n3339 ;
  assign n3371 = ~n1743 & n3370 ;
  assign n3372 = ~n3369 & n3371 ;
  assign n3373 = ~n3340 & ~n3372 ;
  assign n3374 = \req[45]  & ~n753 ;
  assign n3375 = ~n739 & n3374 ;
  assign n3376 = ~\priority[47]  & ~n759 ;
  assign n3377 = n384 & ~n3376 ;
  assign n3378 = n402 & ~n3377 ;
  assign n3379 = n416 & ~n3378 ;
  assign n3380 = n429 & ~n3379 ;
  assign n3381 = n442 & ~n3380 ;
  assign n3382 = n455 & ~n3381 ;
  assign n3383 = n468 & ~n3382 ;
  assign n3384 = n481 & ~n3383 ;
  assign n3385 = n494 & ~n3384 ;
  assign n3386 = n507 & ~n3385 ;
  assign n3387 = n520 & ~n3386 ;
  assign n3388 = n533 & ~n3387 ;
  assign n3389 = n546 & ~n3388 ;
  assign n3390 = n559 & ~n3389 ;
  assign n3391 = n572 & ~n3390 ;
  assign n3392 = n585 & ~n3391 ;
  assign n3393 = n598 & ~n3392 ;
  assign n3394 = n611 & ~n3393 ;
  assign n3395 = n2090 & ~n3394 ;
  assign n3396 = n2094 & ~n3395 ;
  assign n3397 = n2447 & ~n3396 ;
  assign n3398 = n2450 & ~n3397 ;
  assign n3399 = n1837 & ~n3398 ;
  assign n3400 = n1841 & ~n3399 ;
  assign n3401 = n1845 & ~n3400 ;
  assign n3402 = n1849 & ~n3401 ;
  assign n3403 = n1853 & ~n3402 ;
  assign n3404 = n1857 & ~n3403 ;
  assign n3405 = n748 & n3374 ;
  assign n3406 = ~n1859 & n3405 ;
  assign n3407 = ~n3404 & n3406 ;
  assign n3408 = ~n3375 & ~n3407 ;
  assign n3409 = \req[46]  & ~n1119 ;
  assign n3410 = ~n1105 & n3409 ;
  assign n3411 = ~\priority[48]  & ~n1125 ;
  assign n3412 = n751 & ~n3411 ;
  assign n3413 = n769 & ~n3412 ;
  assign n3414 = n3099 & ~n3413 ;
  assign n3415 = n796 & ~n3414 ;
  assign n3416 = n809 & ~n3415 ;
  assign n3417 = n2117 & ~n3416 ;
  assign n3418 = n835 & ~n3417 ;
  assign n3419 = n848 & ~n3418 ;
  assign n3420 = n861 & ~n3419 ;
  assign n3421 = n874 & ~n3420 ;
  assign n3422 = n887 & ~n3421 ;
  assign n3423 = n900 & ~n3422 ;
  assign n3424 = n913 & ~n3423 ;
  assign n3425 = n926 & ~n3424 ;
  assign n3426 = n939 & ~n3425 ;
  assign n3427 = n952 & ~n3426 ;
  assign n3428 = n965 & ~n3427 ;
  assign n3429 = n978 & ~n3428 ;
  assign n3430 = n2132 & ~n3429 ;
  assign n3431 = n2136 & ~n3430 ;
  assign n3432 = n2487 & ~n3431 ;
  assign n3433 = n2490 & ~n3432 ;
  assign n3434 = n1953 & ~n3433 ;
  assign n3435 = n1957 & ~n3434 ;
  assign n3436 = n1961 & ~n3435 ;
  assign n3437 = n1965 & ~n3436 ;
  assign n3438 = n1969 & ~n3437 ;
  assign n3439 = n1973 & ~n3438 ;
  assign n3440 = n1114 & n3409 ;
  assign n3441 = ~n1975 & n3440 ;
  assign n3442 = ~n3439 & n3441 ;
  assign n3443 = ~n3410 & ~n3442 ;
  assign n3444 = \req[47]  & ~n383 ;
  assign n3445 = ~n394 & n3444 ;
  assign n3446 = ~\priority[49]  & ~n399 ;
  assign n3447 = n1117 & ~n3446 ;
  assign n3448 = n1135 & ~n3447 ;
  assign n3449 = n1149 & ~n3448 ;
  assign n3450 = n1162 & ~n3449 ;
  assign n3451 = n1175 & ~n3450 ;
  assign n3452 = n1188 & ~n3451 ;
  assign n3453 = n1201 & ~n3452 ;
  assign n3454 = n1214 & ~n3453 ;
  assign n3455 = n1227 & ~n3454 ;
  assign n3456 = n1240 & ~n3455 ;
  assign n3457 = n1253 & ~n3456 ;
  assign n3458 = n1266 & ~n3457 ;
  assign n3459 = n1279 & ~n3458 ;
  assign n3460 = n1292 & ~n3459 ;
  assign n3461 = n1305 & ~n3460 ;
  assign n3462 = n3148 & ~n3461 ;
  assign n3463 = n1331 & ~n3462 ;
  assign n3464 = n1344 & ~n3463 ;
  assign n3465 = n2173 & ~n3464 ;
  assign n3466 = n2176 & ~n3465 ;
  assign n3467 = n286 & ~n3466 ;
  assign n3468 = n299 & ~n3467 ;
  assign n3469 = n312 & ~n3468 ;
  assign n3470 = n325 & ~n3469 ;
  assign n3471 = n338 & ~n3470 ;
  assign n3472 = n351 & ~n3471 ;
  assign n3473 = n364 & ~n3472 ;
  assign n3474 = n377 & ~n3473 ;
  assign n3475 = n388 & n3444 ;
  assign n3476 = ~n382 & n3475 ;
  assign n3477 = ~n3474 & n3476 ;
  assign n3478 = ~n3445 & ~n3477 ;
  assign n3479 = \req[48]  & ~n750 ;
  assign n3480 = ~n761 & n3479 ;
  assign n3481 = ~\priority[50]  & ~n766 ;
  assign n3482 = n406 & ~n3481 ;
  assign n3483 = n1403 & ~n3482 ;
  assign n3484 = n1408 & ~n3483 ;
  assign n3485 = n1412 & ~n3484 ;
  assign n3486 = n1416 & ~n3485 ;
  assign n3487 = n1420 & ~n3486 ;
  assign n3488 = n1424 & ~n3487 ;
  assign n3489 = n1428 & ~n3488 ;
  assign n3490 = n1432 & ~n3489 ;
  assign n3491 = n1436 & ~n3490 ;
  assign n3492 = n1440 & ~n3491 ;
  assign n3493 = n1444 & ~n3492 ;
  assign n3494 = n1448 & ~n3493 ;
  assign n3495 = n1452 & ~n3494 ;
  assign n3496 = n1456 & ~n3495 ;
  assign n3497 = n1460 & ~n3496 ;
  assign n3498 = n1464 & ~n3497 ;
  assign n3499 = n1468 & ~n3498 ;
  assign n3500 = n2212 & ~n3499 ;
  assign n3501 = n2215 & ~n3500 ;
  assign n3502 = n653 & ~n3501 ;
  assign n3503 = n666 & ~n3502 ;
  assign n3504 = n679 & ~n3503 ;
  assign n3505 = n692 & ~n3504 ;
  assign n3506 = n705 & ~n3505 ;
  assign n3507 = n718 & ~n3506 ;
  assign n3508 = n731 & ~n3507 ;
  assign n3509 = n744 & ~n3508 ;
  assign n3510 = n755 & n3479 ;
  assign n3511 = ~n749 & n3510 ;
  assign n3512 = ~n3509 & n3511 ;
  assign n3513 = ~n3480 & ~n3512 ;
  assign n3514 = \req[49]  & ~n1116 ;
  assign n3515 = ~n1127 & n3514 ;
  assign n3516 = ~\priority[51]  & ~n1132 ;
  assign n3517 = n773 & ~n3516 ;
  assign n3518 = n1523 & ~n3517 ;
  assign n3519 = n1528 & ~n3518 ;
  assign n3520 = n1532 & ~n3519 ;
  assign n3521 = n1536 & ~n3520 ;
  assign n3522 = n1540 & ~n3521 ;
  assign n3523 = n1544 & ~n3522 ;
  assign n3524 = n1548 & ~n3523 ;
  assign n3525 = n1552 & ~n3524 ;
  assign n3526 = n1556 & ~n3525 ;
  assign n3527 = n1560 & ~n3526 ;
  assign n3528 = n1564 & ~n3527 ;
  assign n3529 = n1568 & ~n3528 ;
  assign n3530 = n1572 & ~n3529 ;
  assign n3531 = n1576 & ~n3530 ;
  assign n3532 = n1580 & ~n3531 ;
  assign n3533 = n1584 & ~n3532 ;
  assign n3534 = n1588 & ~n3533 ;
  assign n3535 = n2252 & ~n3534 ;
  assign n3536 = n2255 & ~n3535 ;
  assign n3537 = n1019 & ~n3536 ;
  assign n3538 = n1032 & ~n3537 ;
  assign n3539 = n1045 & ~n3538 ;
  assign n3540 = n1058 & ~n3539 ;
  assign n3541 = n1071 & ~n3540 ;
  assign n3542 = n1084 & ~n3541 ;
  assign n3543 = n1097 & ~n3542 ;
  assign n3544 = n1110 & ~n3543 ;
  assign n3545 = n1121 & n3514 ;
  assign n3546 = ~n1115 & n3545 ;
  assign n3547 = ~n3544 & n3546 ;
  assign n3548 = ~n3515 & ~n3547 ;
  assign n3549 = \req[50]  & ~n405 ;
  assign n3550 = ~n401 & n3549 ;
  assign n3551 = ~\priority[52]  & ~n396 ;
  assign n3552 = n1139 & ~n3551 ;
  assign n3553 = n1640 & ~n3552 ;
  assign n3554 = n1645 & ~n3553 ;
  assign n3555 = n1649 & ~n3554 ;
  assign n3556 = n1653 & ~n3555 ;
  assign n3557 = n1657 & ~n3556 ;
  assign n3558 = n1661 & ~n3557 ;
  assign n3559 = n1665 & ~n3558 ;
  assign n3560 = n1669 & ~n3559 ;
  assign n3561 = n1673 & ~n3560 ;
  assign n3562 = n1677 & ~n3561 ;
  assign n3563 = n1681 & ~n3562 ;
  assign n3564 = n1685 & ~n3563 ;
  assign n3565 = n1689 & ~n3564 ;
  assign n3566 = n1693 & ~n3565 ;
  assign n3567 = n1697 & ~n3566 ;
  assign n3568 = n1701 & ~n3567 ;
  assign n3569 = ~n1342 & n1348 ;
  assign n3570 = n1704 & ~n3569 ;
  assign n3571 = ~n3568 & n3570 ;
  assign n3572 = n2291 & ~n3571 ;
  assign n3573 = n2294 & ~n3572 ;
  assign n3574 = n1368 & ~n3573 ;
  assign n3575 = n1372 & ~n3574 ;
  assign n3576 = n1376 & ~n3575 ;
  assign n3577 = n1380 & ~n3576 ;
  assign n3578 = n1384 & ~n3577 ;
  assign n3579 = n1388 & ~n3578 ;
  assign n3580 = n1392 & ~n3579 ;
  assign n3581 = n1396 & ~n3580 ;
  assign n3582 = n385 & n3549 ;
  assign n3583 = ~n1398 & n3582 ;
  assign n3584 = ~n3581 & n3583 ;
  assign n3585 = ~n3550 & ~n3584 ;
  assign n3586 = \req[51]  & ~n772 ;
  assign n3587 = ~n768 & n3586 ;
  assign n3588 = ~\priority[53]  & ~n763 ;
  assign n3589 = n413 & ~n3588 ;
  assign n3590 = n1756 & ~n3589 ;
  assign n3591 = n1761 & ~n3590 ;
  assign n3592 = n1765 & ~n3591 ;
  assign n3593 = n1769 & ~n3592 ;
  assign n3594 = n1773 & ~n3593 ;
  assign n3595 = n1777 & ~n3594 ;
  assign n3596 = n1781 & ~n3595 ;
  assign n3597 = n1785 & ~n3596 ;
  assign n3598 = n1789 & ~n3597 ;
  assign n3599 = n1793 & ~n3598 ;
  assign n3600 = n1797 & ~n3599 ;
  assign n3601 = n1801 & ~n3600 ;
  assign n3602 = n1805 & ~n3601 ;
  assign n3603 = n1809 & ~n3602 ;
  assign n3604 = n1813 & ~n3603 ;
  assign n3605 = n1817 & ~n3604 ;
  assign n3606 = n1821 & ~n3605 ;
  assign n3607 = n2330 & ~n3606 ;
  assign n3608 = n2333 & ~n3607 ;
  assign n3609 = n1488 & ~n3608 ;
  assign n3610 = n1492 & ~n3609 ;
  assign n3611 = n1496 & ~n3610 ;
  assign n3612 = n1500 & ~n3611 ;
  assign n3613 = n1504 & ~n3612 ;
  assign n3614 = n2229 & ~n3613 ;
  assign n3615 = n1512 & ~n3614 ;
  assign n3616 = n1516 & ~n3615 ;
  assign n3617 = n752 & n3586 ;
  assign n3618 = ~n1518 & n3617 ;
  assign n3619 = ~n3616 & n3618 ;
  assign n3620 = ~n3587 & ~n3619 ;
  assign n3621 = \req[52]  & ~n1138 ;
  assign n3622 = ~n1134 & n3621 ;
  assign n3623 = ~\priority[54]  & ~n1129 ;
  assign n3624 = n780 & ~n3623 ;
  assign n3625 = n1872 & ~n3624 ;
  assign n3626 = n1877 & ~n3625 ;
  assign n3627 = ~n1879 & n1880 ;
  assign n3628 = ~n3626 & n3627 ;
  assign n3629 = n1885 & ~n3628 ;
  assign n3630 = n1889 & ~n3629 ;
  assign n3631 = n1893 & ~n3630 ;
  assign n3632 = n1897 & ~n3631 ;
  assign n3633 = n1901 & ~n3632 ;
  assign n3634 = n1905 & ~n3633 ;
  assign n3635 = n1909 & ~n3634 ;
  assign n3636 = n1913 & ~n3635 ;
  assign n3637 = n1917 & ~n3636 ;
  assign n3638 = n1921 & ~n3637 ;
  assign n3639 = n1925 & ~n3638 ;
  assign n3640 = n1929 & ~n3639 ;
  assign n3641 = n1933 & ~n3640 ;
  assign n3642 = n1937 & ~n3641 ;
  assign n3643 = n2369 & ~n3642 ;
  assign n3644 = n2372 & ~n3643 ;
  assign n3645 = n1605 & ~n3644 ;
  assign n3646 = n1609 & ~n3645 ;
  assign n3647 = n1613 & ~n3646 ;
  assign n3648 = n1617 & ~n3647 ;
  assign n3649 = n1621 & ~n3648 ;
  assign n3650 = n1625 & ~n3649 ;
  assign n3651 = n1629 & ~n3650 ;
  assign n3652 = n1633 & ~n3651 ;
  assign n3653 = n1118 & n3621 ;
  assign n3654 = ~n1635 & n3653 ;
  assign n3655 = ~n3652 & n3654 ;
  assign n3656 = ~n3622 & ~n3655 ;
  assign n3657 = \req[53]  & ~n412 ;
  assign n3658 = ~n398 & n3657 ;
  assign n3659 = ~\priority[55]  & ~n418 ;
  assign n3660 = n1146 & ~n3659 ;
  assign n3661 = n1988 & ~n3660 ;
  assign n3662 = n1993 & ~n3661 ;
  assign n3663 = n1997 & ~n3662 ;
  assign n3664 = n2001 & ~n3663 ;
  assign n3665 = n2005 & ~n3664 ;
  assign n3666 = n2009 & ~n3665 ;
  assign n3667 = n2013 & ~n3666 ;
  assign n3668 = n2017 & ~n3667 ;
  assign n3669 = n2021 & ~n3668 ;
  assign n3670 = n2025 & ~n3669 ;
  assign n3671 = ~n2027 & n2028 ;
  assign n3672 = ~n3670 & n3671 ;
  assign n3673 = n2033 & ~n3672 ;
  assign n3674 = n2037 & ~n3673 ;
  assign n3675 = n2041 & ~n3674 ;
  assign n3676 = n2045 & ~n3675 ;
  assign n3677 = n2049 & ~n3676 ;
  assign n3678 = n2053 & ~n3677 ;
  assign n3679 = n2408 & ~n3678 ;
  assign n3680 = n2411 & ~n3679 ;
  assign n3681 = n1721 & ~n3680 ;
  assign n3682 = n1725 & ~n3681 ;
  assign n3683 = n1729 & ~n3682 ;
  assign n3684 = n1733 & ~n3683 ;
  assign n3685 = n1737 & ~n3684 ;
  assign n3686 = n1741 & ~n3685 ;
  assign n3687 = n1745 & ~n3686 ;
  assign n3688 = n1749 & ~n3687 ;
  assign n3689 = n407 & n3657 ;
  assign n3690 = ~n1751 & n3689 ;
  assign n3691 = ~n3688 & n3690 ;
  assign n3692 = ~n3658 & ~n3691 ;
  assign n3693 = \req[54]  & ~n779 ;
  assign n3694 = ~n765 & n3693 ;
  assign n3695 = ~\priority[56]  & ~n785 ;
  assign n3696 = n410 & ~n3695 ;
  assign n3697 = n428 & ~n3696 ;
  assign n3698 = n442 & ~n3697 ;
  assign n3699 = n455 & ~n3698 ;
  assign n3700 = n468 & ~n3699 ;
  assign n3701 = n481 & ~n3700 ;
  assign n3702 = n494 & ~n3701 ;
  assign n3703 = n507 & ~n3702 ;
  assign n3704 = n520 & ~n3703 ;
  assign n3705 = n533 & ~n3704 ;
  assign n3706 = n546 & ~n3705 ;
  assign n3707 = n559 & ~n3706 ;
  assign n3708 = n572 & ~n3707 ;
  assign n3709 = n585 & ~n3708 ;
  assign n3710 = n598 & ~n3709 ;
  assign n3711 = n611 & ~n3710 ;
  assign n3712 = n2090 & ~n3711 ;
  assign n3713 = n2094 & ~n3712 ;
  assign n3714 = n2447 & ~n3713 ;
  assign n3715 = n2450 & ~n3714 ;
  assign n3716 = n1837 & ~n3715 ;
  assign n3717 = n1841 & ~n3716 ;
  assign n3718 = n1845 & ~n3717 ;
  assign n3719 = n1849 & ~n3718 ;
  assign n3720 = ~n1851 & n1852 ;
  assign n3721 = ~n3719 & n3720 ;
  assign n3722 = n1857 & ~n3721 ;
  assign n3723 = n1861 & ~n3722 ;
  assign n3724 = n1865 & ~n3723 ;
  assign n3725 = n774 & n3693 ;
  assign n3726 = ~n1867 & n3725 ;
  assign n3727 = ~n3724 & n3726 ;
  assign n3728 = ~n3694 & ~n3727 ;
  assign n3729 = \req[55]  & ~n1145 ;
  assign n3730 = ~n1131 & n3729 ;
  assign n3731 = ~\priority[57]  & ~n1151 ;
  assign n3732 = n777 & ~n3731 ;
  assign n3733 = n795 & ~n3732 ;
  assign n3734 = n809 & ~n3733 ;
  assign n3735 = n2117 & ~n3734 ;
  assign n3736 = n835 & ~n3735 ;
  assign n3737 = n848 & ~n3736 ;
  assign n3738 = n861 & ~n3737 ;
  assign n3739 = n874 & ~n3738 ;
  assign n3740 = n887 & ~n3739 ;
  assign n3741 = n900 & ~n3740 ;
  assign n3742 = n913 & ~n3741 ;
  assign n3743 = n926 & ~n3742 ;
  assign n3744 = n939 & ~n3743 ;
  assign n3745 = n952 & ~n3744 ;
  assign n3746 = n965 & ~n3745 ;
  assign n3747 = n978 & ~n3746 ;
  assign n3748 = n2132 & ~n3747 ;
  assign n3749 = n2136 & ~n3748 ;
  assign n3750 = n2487 & ~n3749 ;
  assign n3751 = n2490 & ~n3750 ;
  assign n3752 = n1953 & ~n3751 ;
  assign n3753 = n1957 & ~n3752 ;
  assign n3754 = n1961 & ~n3753 ;
  assign n3755 = n1965 & ~n3754 ;
  assign n3756 = n1969 & ~n3755 ;
  assign n3757 = n1973 & ~n3756 ;
  assign n3758 = n2713 & ~n3757 ;
  assign n3759 = n1981 & ~n3758 ;
  assign n3760 = n1140 & n3729 ;
  assign n3761 = ~n1983 & n3760 ;
  assign n3762 = ~n3759 & n3761 ;
  assign n3763 = ~n3730 & ~n3762 ;
  assign n3764 = \req[56]  & ~n409 ;
  assign n3765 = ~n420 & n3764 ;
  assign n3766 = ~\priority[58]  & ~n425 ;
  assign n3767 = n1143 & ~n3766 ;
  assign n3768 = n1161 & ~n3767 ;
  assign n3769 = n1175 & ~n3768 ;
  assign n3770 = n1188 & ~n3769 ;
  assign n3771 = n1201 & ~n3770 ;
  assign n3772 = n1214 & ~n3771 ;
  assign n3773 = n1227 & ~n3772 ;
  assign n3774 = n1240 & ~n3773 ;
  assign n3775 = n1253 & ~n3774 ;
  assign n3776 = n1266 & ~n3775 ;
  assign n3777 = n1279 & ~n3776 ;
  assign n3778 = n1292 & ~n3777 ;
  assign n3779 = n1305 & ~n3778 ;
  assign n3780 = n3148 & ~n3779 ;
  assign n3781 = n1331 & ~n3780 ;
  assign n3782 = n1344 & ~n3781 ;
  assign n3783 = n2173 & ~n3782 ;
  assign n3784 = n2176 & ~n3783 ;
  assign n3785 = n286 & ~n3784 ;
  assign n3786 = n299 & ~n3785 ;
  assign n3787 = n312 & ~n3786 ;
  assign n3788 = n325 & ~n3787 ;
  assign n3789 = n338 & ~n3788 ;
  assign n3790 = n351 & ~n3789 ;
  assign n3791 = n364 & ~n3790 ;
  assign n3792 = n377 & ~n3791 ;
  assign n3793 = n390 & ~n3792 ;
  assign n3794 = n403 & ~n3793 ;
  assign n3795 = n414 & n3764 ;
  assign n3796 = ~n408 & n3795 ;
  assign n3797 = ~n3794 & n3796 ;
  assign n3798 = ~n3765 & ~n3797 ;
  assign n3799 = \req[57]  & ~n776 ;
  assign n3800 = ~n787 & n3799 ;
  assign n3801 = ~\priority[59]  & ~n792 ;
  assign n3802 = n432 & ~n3801 ;
  assign n3803 = n1411 & ~n3802 ;
  assign n3804 = n1416 & ~n3803 ;
  assign n3805 = n1420 & ~n3804 ;
  assign n3806 = n1424 & ~n3805 ;
  assign n3807 = n1428 & ~n3806 ;
  assign n3808 = n1432 & ~n3807 ;
  assign n3809 = n1436 & ~n3808 ;
  assign n3810 = n1440 & ~n3809 ;
  assign n3811 = ~n1442 & n1443 ;
  assign n3812 = ~n3810 & n3811 ;
  assign n3813 = n1448 & ~n3812 ;
  assign n3814 = n1452 & ~n3813 ;
  assign n3815 = n1456 & ~n3814 ;
  assign n3816 = n580 & n602 ;
  assign n3817 = ~n1458 & n3816 ;
  assign n3818 = ~n3815 & n3817 ;
  assign n3819 = n1464 & ~n3818 ;
  assign n3820 = n1468 & ~n3819 ;
  assign n3821 = n2212 & ~n3820 ;
  assign n3822 = n2215 & ~n3821 ;
  assign n3823 = n653 & ~n3822 ;
  assign n3824 = n666 & ~n3823 ;
  assign n3825 = n679 & ~n3824 ;
  assign n3826 = ~n684 & n691 ;
  assign n3827 = ~n3825 & n3826 ;
  assign n3828 = n705 & ~n3827 ;
  assign n3829 = n718 & ~n3828 ;
  assign n3830 = n731 & ~n3829 ;
  assign n3831 = n744 & ~n3830 ;
  assign n3832 = n2465 & ~n3831 ;
  assign n3833 = n770 & ~n3832 ;
  assign n3834 = n781 & n3799 ;
  assign n3835 = ~n775 & n3834 ;
  assign n3836 = ~n3833 & n3835 ;
  assign n3837 = ~n3800 & ~n3836 ;
  assign n3838 = \req[58]  & ~n1142 ;
  assign n3839 = ~n1153 & n3838 ;
  assign n3840 = ~\priority[60]  & ~n1158 ;
  assign n3841 = n799 & ~n3840 ;
  assign n3842 = n1531 & ~n3841 ;
  assign n3843 = n1536 & ~n3842 ;
  assign n3844 = n1540 & ~n3843 ;
  assign n3845 = n1544 & ~n3844 ;
  assign n3846 = n1548 & ~n3845 ;
  assign n3847 = n1552 & ~n3846 ;
  assign n3848 = n1556 & ~n3847 ;
  assign n3849 = n1560 & ~n3848 ;
  assign n3850 = n1564 & ~n3849 ;
  assign n3851 = n1568 & ~n3850 ;
  assign n3852 = n1572 & ~n3851 ;
  assign n3853 = n1576 & ~n3852 ;
  assign n3854 = n1580 & ~n3853 ;
  assign n3855 = n1584 & ~n3854 ;
  assign n3856 = n1588 & ~n3855 ;
  assign n3857 = n2252 & ~n3856 ;
  assign n3858 = n2255 & ~n3857 ;
  assign n3859 = n1019 & ~n3858 ;
  assign n3860 = n1032 & ~n3859 ;
  assign n3861 = ~n1037 & n1044 ;
  assign n3862 = ~n3860 & n3861 ;
  assign n3863 = n1058 & ~n3862 ;
  assign n3864 = n1071 & ~n3863 ;
  assign n3865 = n1084 & ~n3864 ;
  assign n3866 = n1097 & ~n3865 ;
  assign n3867 = n1110 & ~n3866 ;
  assign n3868 = n1123 & ~n3867 ;
  assign n3869 = n1136 & ~n3868 ;
  assign n3870 = n1147 & n3838 ;
  assign n3871 = ~n1141 & n3870 ;
  assign n3872 = ~n3869 & n3871 ;
  assign n3873 = ~n3839 & ~n3872 ;
  assign n3874 = \req[59]  & ~n431 ;
  assign n3875 = ~n427 & n3874 ;
  assign n3876 = ~\priority[61]  & ~n422 ;
  assign n3877 = n1165 & ~n3876 ;
  assign n3878 = n1648 & ~n3877 ;
  assign n3879 = n1653 & ~n3878 ;
  assign n3880 = n1657 & ~n3879 ;
  assign n3881 = n1661 & ~n3880 ;
  assign n3882 = n1665 & ~n3881 ;
  assign n3883 = n1669 & ~n3882 ;
  assign n3884 = n1673 & ~n3883 ;
  assign n3885 = n1677 & ~n3884 ;
  assign n3886 = n1681 & ~n3885 ;
  assign n3887 = n1685 & ~n3886 ;
  assign n3888 = n1689 & ~n3887 ;
  assign n3889 = n1693 & ~n3888 ;
  assign n3890 = n1697 & ~n3889 ;
  assign n3891 = n1701 & ~n3890 ;
  assign n3892 = n3570 & ~n3891 ;
  assign n3893 = n2291 & ~n3892 ;
  assign n3894 = n2294 & ~n3893 ;
  assign n3895 = n1368 & ~n3894 ;
  assign n3896 = n1372 & ~n3895 ;
  assign n3897 = n1376 & ~n3896 ;
  assign n3898 = n1380 & ~n3897 ;
  assign n3899 = n1384 & ~n3898 ;
  assign n3900 = n1388 & ~n3899 ;
  assign n3901 = n1392 & ~n3900 ;
  assign n3902 = n1396 & ~n3901 ;
  assign n3903 = n1400 & ~n3902 ;
  assign n3904 = n1404 & ~n3903 ;
  assign n3905 = n411 & n3874 ;
  assign n3906 = ~n1406 & n3905 ;
  assign n3907 = ~n3904 & n3906 ;
  assign n3908 = ~n3875 & ~n3907 ;
  assign n3909 = \req[60]  & ~n798 ;
  assign n3910 = ~n794 & n3909 ;
  assign n3911 = ~\priority[62]  & ~n789 ;
  assign n3912 = n439 & ~n3911 ;
  assign n3913 = n1764 & ~n3912 ;
  assign n3914 = n1769 & ~n3913 ;
  assign n3915 = n1773 & ~n3914 ;
  assign n3916 = n1777 & ~n3915 ;
  assign n3917 = n1781 & ~n3916 ;
  assign n3918 = n1785 & ~n3917 ;
  assign n3919 = n1789 & ~n3918 ;
  assign n3920 = ~n1791 & n1792 ;
  assign n3921 = ~n3919 & n3920 ;
  assign n3922 = n1797 & ~n3921 ;
  assign n3923 = n1801 & ~n3922 ;
  assign n3924 = n1805 & ~n3923 ;
  assign n3925 = n1809 & ~n3924 ;
  assign n3926 = n1813 & ~n3925 ;
  assign n3927 = n1817 & ~n3926 ;
  assign n3928 = n1821 & ~n3927 ;
  assign n3929 = n2330 & ~n3928 ;
  assign n3930 = n2333 & ~n3929 ;
  assign n3931 = n1488 & ~n3930 ;
  assign n3932 = n1492 & ~n3931 ;
  assign n3933 = n1496 & ~n3932 ;
  assign n3934 = n1500 & ~n3933 ;
  assign n3935 = n1504 & ~n3934 ;
  assign n3936 = n2229 & ~n3935 ;
  assign n3937 = n1512 & ~n3936 ;
  assign n3938 = n1516 & ~n3937 ;
  assign n3939 = n1520 & ~n3938 ;
  assign n3940 = n1524 & ~n3939 ;
  assign n3941 = n778 & n3909 ;
  assign n3942 = ~n1526 & n3941 ;
  assign n3943 = ~n3940 & n3942 ;
  assign n3944 = ~n3910 & ~n3943 ;
  assign n3945 = \req[61]  & ~n1164 ;
  assign n3946 = ~n1160 & n3945 ;
  assign n3947 = ~\priority[63]  & ~n1155 ;
  assign n3948 = n806 & ~n3947 ;
  assign n3949 = n1880 & ~n3948 ;
  assign n3950 = n1885 & ~n3949 ;
  assign n3951 = n1889 & ~n3950 ;
  assign n3952 = n1893 & ~n3951 ;
  assign n3953 = n1897 & ~n3952 ;
  assign n3954 = n1901 & ~n3953 ;
  assign n3955 = n1905 & ~n3954 ;
  assign n3956 = n1909 & ~n3955 ;
  assign n3957 = n1913 & ~n3956 ;
  assign n3958 = n1917 & ~n3957 ;
  assign n3959 = n1921 & ~n3958 ;
  assign n3960 = n1925 & ~n3959 ;
  assign n3961 = n1929 & ~n3960 ;
  assign n3962 = n1933 & ~n3961 ;
  assign n3963 = n1937 & ~n3962 ;
  assign n3964 = n2369 & ~n3963 ;
  assign n3965 = n2372 & ~n3964 ;
  assign n3966 = n1605 & ~n3965 ;
  assign n3967 = n1609 & ~n3966 ;
  assign n3968 = n1613 & ~n3967 ;
  assign n3969 = n1617 & ~n3968 ;
  assign n3970 = n1621 & ~n3969 ;
  assign n3971 = n1625 & ~n3970 ;
  assign n3972 = n1629 & ~n3971 ;
  assign n3973 = n1633 & ~n3972 ;
  assign n3974 = n1637 & ~n3973 ;
  assign n3975 = n1641 & ~n3974 ;
  assign n3976 = n1144 & n3945 ;
  assign n3977 = ~n1643 & n3976 ;
  assign n3978 = ~n3975 & n3977 ;
  assign n3979 = ~n3946 & ~n3978 ;
  assign n3980 = \req[62]  & ~n438 ;
  assign n3981 = ~n424 & n3980 ;
  assign n3982 = ~\priority[64]  & ~n444 ;
  assign n3983 = n1172 & ~n3982 ;
  assign n3984 = n1996 & ~n3983 ;
  assign n3985 = n2001 & ~n3984 ;
  assign n3986 = n2005 & ~n3985 ;
  assign n3987 = n2009 & ~n3986 ;
  assign n3988 = n2013 & ~n3987 ;
  assign n3989 = n2017 & ~n3988 ;
  assign n3990 = n2021 & ~n3989 ;
  assign n3991 = n2025 & ~n3990 ;
  assign n3992 = n3671 & ~n3991 ;
  assign n3993 = n2033 & ~n3992 ;
  assign n3994 = n2037 & ~n3993 ;
  assign n3995 = n2041 & ~n3994 ;
  assign n3996 = n2045 & ~n3995 ;
  assign n3997 = n2049 & ~n3996 ;
  assign n3998 = n2053 & ~n3997 ;
  assign n3999 = n2408 & ~n3998 ;
  assign n4000 = n2411 & ~n3999 ;
  assign n4001 = n1721 & ~n4000 ;
  assign n4002 = n1725 & ~n4001 ;
  assign n4003 = n1729 & ~n4002 ;
  assign n4004 = n1733 & ~n4003 ;
  assign n4005 = n1737 & ~n4004 ;
  assign n4006 = n1741 & ~n4005 ;
  assign n4007 = n1745 & ~n4006 ;
  assign n4008 = n1749 & ~n4007 ;
  assign n4009 = n1753 & ~n4008 ;
  assign n4010 = n1757 & ~n4009 ;
  assign n4011 = n433 & n3980 ;
  assign n4012 = ~n1759 & n4011 ;
  assign n4013 = ~n4010 & n4012 ;
  assign n4014 = ~n3981 & ~n4013 ;
  assign n4015 = \req[63]  & ~n805 ;
  assign n4016 = ~n791 & n4015 ;
  assign n4017 = ~\priority[65]  & ~n811 ;
  assign n4018 = n436 & ~n4017 ;
  assign n4019 = n454 & ~n4018 ;
  assign n4020 = n468 & ~n4019 ;
  assign n4021 = n481 & ~n4020 ;
  assign n4022 = n494 & ~n4021 ;
  assign n4023 = n507 & ~n4022 ;
  assign n4024 = n520 & ~n4023 ;
  assign n4025 = n533 & ~n4024 ;
  assign n4026 = n546 & ~n4025 ;
  assign n4027 = n559 & ~n4026 ;
  assign n4028 = n572 & ~n4027 ;
  assign n4029 = n585 & ~n4028 ;
  assign n4030 = n598 & ~n4029 ;
  assign n4031 = n611 & ~n4030 ;
  assign n4032 = n2090 & ~n4031 ;
  assign n4033 = n2094 & ~n4032 ;
  assign n4034 = n2447 & ~n4033 ;
  assign n4035 = n2450 & ~n4034 ;
  assign n4036 = n1837 & ~n4035 ;
  assign n4037 = n1841 & ~n4036 ;
  assign n4038 = n1845 & ~n4037 ;
  assign n4039 = n1849 & ~n4038 ;
  assign n4040 = n3720 & ~n4039 ;
  assign n4041 = n1857 & ~n4040 ;
  assign n4042 = n1861 & ~n4041 ;
  assign n4043 = n1865 & ~n4042 ;
  assign n4044 = n1869 & ~n4043 ;
  assign n4045 = n1873 & ~n4044 ;
  assign n4046 = n800 & n4015 ;
  assign n4047 = ~n1875 & n4046 ;
  assign n4048 = ~n4045 & n4047 ;
  assign n4049 = ~n4016 & ~n4048 ;
  assign n4050 = \req[64]  & ~n1171 ;
  assign n4051 = ~n1157 & n4050 ;
  assign n4052 = ~\priority[66]  & ~n1177 ;
  assign n4053 = n803 & ~n4052 ;
  assign n4054 = n821 & ~n4053 ;
  assign n4055 = n835 & ~n4054 ;
  assign n4056 = n848 & ~n4055 ;
  assign n4057 = n861 & ~n4056 ;
  assign n4058 = n874 & ~n4057 ;
  assign n4059 = n887 & ~n4058 ;
  assign n4060 = n900 & ~n4059 ;
  assign n4061 = n913 & ~n4060 ;
  assign n4062 = n926 & ~n4061 ;
  assign n4063 = n939 & ~n4062 ;
  assign n4064 = n952 & ~n4063 ;
  assign n4065 = n965 & ~n4064 ;
  assign n4066 = n978 & ~n4065 ;
  assign n4067 = n2132 & ~n4066 ;
  assign n4068 = n2136 & ~n4067 ;
  assign n4069 = n2487 & ~n4068 ;
  assign n4070 = n2490 & ~n4069 ;
  assign n4071 = n1953 & ~n4070 ;
  assign n4072 = n1957 & ~n4071 ;
  assign n4073 = n1961 & ~n4072 ;
  assign n4074 = n1965 & ~n4073 ;
  assign n4075 = n1969 & ~n4074 ;
  assign n4076 = n1973 & ~n4075 ;
  assign n4077 = n2713 & ~n4076 ;
  assign n4078 = n1981 & ~n4077 ;
  assign n4079 = n1985 & ~n4078 ;
  assign n4080 = n1989 & ~n4079 ;
  assign n4081 = n1166 & n4050 ;
  assign n4082 = ~n1991 & n4081 ;
  assign n4083 = ~n4080 & n4082 ;
  assign n4084 = ~n4051 & ~n4083 ;
  assign n4085 = \req[65]  & ~n435 ;
  assign n4086 = ~n446 & n4085 ;
  assign n4087 = ~\priority[67]  & ~n451 ;
  assign n4088 = n1169 & ~n4087 ;
  assign n4089 = n1187 & ~n4088 ;
  assign n4090 = n1201 & ~n4089 ;
  assign n4091 = n1214 & ~n4090 ;
  assign n4092 = n1227 & ~n4091 ;
  assign n4093 = n1240 & ~n4092 ;
  assign n4094 = n1253 & ~n4093 ;
  assign n4095 = n1266 & ~n4094 ;
  assign n4096 = n1279 & ~n4095 ;
  assign n4097 = n1292 & ~n4096 ;
  assign n4098 = n1305 & ~n4097 ;
  assign n4099 = n3148 & ~n4098 ;
  assign n4100 = n1331 & ~n4099 ;
  assign n4101 = n1344 & ~n4100 ;
  assign n4102 = n2173 & ~n4101 ;
  assign n4103 = n2176 & ~n4102 ;
  assign n4104 = n286 & ~n4103 ;
  assign n4105 = n299 & ~n4104 ;
  assign n4106 = n312 & ~n4105 ;
  assign n4107 = n325 & ~n4106 ;
  assign n4108 = n338 & ~n4107 ;
  assign n4109 = n351 & ~n4108 ;
  assign n4110 = n364 & ~n4109 ;
  assign n4111 = n377 & ~n4110 ;
  assign n4112 = n390 & ~n4111 ;
  assign n4113 = n403 & ~n4112 ;
  assign n4114 = n416 & ~n4113 ;
  assign n4115 = ~n421 & n428 ;
  assign n4116 = ~n4114 & n4115 ;
  assign n4117 = n440 & n4085 ;
  assign n4118 = ~n434 & n4117 ;
  assign n4119 = ~n4116 & n4118 ;
  assign n4120 = ~n4086 & ~n4119 ;
  assign n4121 = \req[66]  & ~n802 ;
  assign n4122 = ~n813 & n4121 ;
  assign n4123 = ~\priority[68]  & ~n818 ;
  assign n4124 = n458 & ~n4123 ;
  assign n4125 = n1419 & ~n4124 ;
  assign n4126 = n1424 & ~n4125 ;
  assign n4127 = n1428 & ~n4126 ;
  assign n4128 = n1432 & ~n4127 ;
  assign n4129 = n1436 & ~n4128 ;
  assign n4130 = n1440 & ~n4129 ;
  assign n4131 = n3811 & ~n4130 ;
  assign n4132 = n1448 & ~n4131 ;
  assign n4133 = n1452 & ~n4132 ;
  assign n4134 = n1456 & ~n4133 ;
  assign n4135 = n3817 & ~n4134 ;
  assign n4136 = n1464 & ~n4135 ;
  assign n4137 = n1468 & ~n4136 ;
  assign n4138 = n2212 & ~n4137 ;
  assign n4139 = n2215 & ~n4138 ;
  assign n4140 = n653 & ~n4139 ;
  assign n4141 = n666 & ~n4140 ;
  assign n4142 = n679 & ~n4141 ;
  assign n4143 = n3826 & ~n4142 ;
  assign n4144 = n705 & ~n4143 ;
  assign n4145 = n718 & ~n4144 ;
  assign n4146 = n731 & ~n4145 ;
  assign n4147 = n744 & ~n4146 ;
  assign n4148 = n2465 & ~n4147 ;
  assign n4149 = n770 & ~n4148 ;
  assign n4150 = n3099 & ~n4149 ;
  assign n4151 = n796 & ~n4150 ;
  assign n4152 = n807 & n4121 ;
  assign n4153 = ~n801 & n4152 ;
  assign n4154 = ~n4151 & n4153 ;
  assign n4155 = ~n4122 & ~n4154 ;
  assign n4156 = \req[67]  & ~n1168 ;
  assign n4157 = ~n1179 & n4156 ;
  assign n4158 = ~\priority[69]  & ~n1184 ;
  assign n4159 = n825 & ~n4158 ;
  assign n4160 = n1539 & ~n4159 ;
  assign n4161 = n1544 & ~n4160 ;
  assign n4162 = n1548 & ~n4161 ;
  assign n4163 = n1552 & ~n4162 ;
  assign n4164 = n1556 & ~n4163 ;
  assign n4165 = n1560 & ~n4164 ;
  assign n4166 = n1564 & ~n4165 ;
  assign n4167 = n1568 & ~n4166 ;
  assign n4168 = n1572 & ~n4167 ;
  assign n4169 = n1576 & ~n4168 ;
  assign n4170 = n1580 & ~n4169 ;
  assign n4171 = n1584 & ~n4170 ;
  assign n4172 = n1588 & ~n4171 ;
  assign n4173 = n2252 & ~n4172 ;
  assign n4174 = n2255 & ~n4173 ;
  assign n4175 = n1019 & ~n4174 ;
  assign n4176 = n1032 & ~n4175 ;
  assign n4177 = n3861 & ~n4176 ;
  assign n4178 = n1058 & ~n4177 ;
  assign n4179 = n1071 & ~n4178 ;
  assign n4180 = n1084 & ~n4179 ;
  assign n4181 = n1097 & ~n4180 ;
  assign n4182 = n1110 & ~n4181 ;
  assign n4183 = n1123 & ~n4182 ;
  assign n4184 = n1136 & ~n4183 ;
  assign n4185 = n1149 & ~n4184 ;
  assign n4186 = n1162 & ~n4185 ;
  assign n4187 = n1173 & n4156 ;
  assign n4188 = ~n1167 & n4187 ;
  assign n4189 = ~n4186 & n4188 ;
  assign n4190 = ~n4157 & ~n4189 ;
  assign n4191 = \req[68]  & ~n457 ;
  assign n4192 = ~n453 & n4191 ;
  assign n4193 = ~\priority[70]  & ~n448 ;
  assign n4194 = n1191 & ~n4193 ;
  assign n4195 = n1656 & ~n4194 ;
  assign n4196 = n1661 & ~n4195 ;
  assign n4197 = n1665 & ~n4196 ;
  assign n4198 = n1669 & ~n4197 ;
  assign n4199 = n1673 & ~n4198 ;
  assign n4200 = n1677 & ~n4199 ;
  assign n4201 = n1681 & ~n4200 ;
  assign n4202 = n1685 & ~n4201 ;
  assign n4203 = n1689 & ~n4202 ;
  assign n4204 = n1693 & ~n4203 ;
  assign n4205 = n1697 & ~n4204 ;
  assign n4206 = n1701 & ~n4205 ;
  assign n4207 = n3570 & ~n4206 ;
  assign n4208 = n2291 & ~n4207 ;
  assign n4209 = n2294 & ~n4208 ;
  assign n4210 = n1368 & ~n4209 ;
  assign n4211 = n1372 & ~n4210 ;
  assign n4212 = n1376 & ~n4211 ;
  assign n4213 = n1380 & ~n4212 ;
  assign n4214 = n1384 & ~n4213 ;
  assign n4215 = n1388 & ~n4214 ;
  assign n4216 = n1392 & ~n4215 ;
  assign n4217 = n1396 & ~n4216 ;
  assign n4218 = n1400 & ~n4217 ;
  assign n4219 = n1404 & ~n4218 ;
  assign n4220 = n1408 & ~n4219 ;
  assign n4221 = n1412 & ~n4220 ;
  assign n4222 = n437 & n4191 ;
  assign n4223 = ~n1414 & n4222 ;
  assign n4224 = ~n4221 & n4223 ;
  assign n4225 = ~n4192 & ~n4224 ;
  assign n4226 = \req[69]  & ~n824 ;
  assign n4227 = ~n820 & n4226 ;
  assign n4228 = ~\priority[71]  & ~n815 ;
  assign n4229 = n465 & ~n4228 ;
  assign n4230 = n1772 & ~n4229 ;
  assign n4231 = n1777 & ~n4230 ;
  assign n4232 = n1781 & ~n4231 ;
  assign n4233 = n1785 & ~n4232 ;
  assign n4234 = n1789 & ~n4233 ;
  assign n4235 = n3920 & ~n4234 ;
  assign n4236 = n1797 & ~n4235 ;
  assign n4237 = n1801 & ~n4236 ;
  assign n4238 = n1805 & ~n4237 ;
  assign n4239 = n1809 & ~n4238 ;
  assign n4240 = n1813 & ~n4239 ;
  assign n4241 = n1817 & ~n4240 ;
  assign n4242 = n1821 & ~n4241 ;
  assign n4243 = n2330 & ~n4242 ;
  assign n4244 = n2333 & ~n4243 ;
  assign n4245 = n1488 & ~n4244 ;
  assign n4246 = n1492 & ~n4245 ;
  assign n4247 = n1496 & ~n4246 ;
  assign n4248 = n1500 & ~n4247 ;
  assign n4249 = n1504 & ~n4248 ;
  assign n4250 = n2229 & ~n4249 ;
  assign n4251 = n1512 & ~n4250 ;
  assign n4252 = n1516 & ~n4251 ;
  assign n4253 = n1520 & ~n4252 ;
  assign n4254 = n1524 & ~n4253 ;
  assign n4255 = n1528 & ~n4254 ;
  assign n4256 = n1532 & ~n4255 ;
  assign n4257 = n804 & n4226 ;
  assign n4258 = ~n1534 & n4257 ;
  assign n4259 = ~n4256 & n4258 ;
  assign n4260 = ~n4227 & ~n4259 ;
  assign n4261 = \req[70]  & ~n1190 ;
  assign n4262 = ~n1186 & n4261 ;
  assign n4263 = ~\priority[72]  & ~n1181 ;
  assign n4264 = n832 & ~n4263 ;
  assign n4265 = n1888 & ~n4264 ;
  assign n4266 = n1893 & ~n4265 ;
  assign n4267 = n1897 & ~n4266 ;
  assign n4268 = n1901 & ~n4267 ;
  assign n4269 = n1905 & ~n4268 ;
  assign n4270 = n1909 & ~n4269 ;
  assign n4271 = n1913 & ~n4270 ;
  assign n4272 = n1917 & ~n4271 ;
  assign n4273 = n1921 & ~n4272 ;
  assign n4274 = n1925 & ~n4273 ;
  assign n4275 = n1929 & ~n4274 ;
  assign n4276 = n1933 & ~n4275 ;
  assign n4277 = n1937 & ~n4276 ;
  assign n4278 = n2369 & ~n4277 ;
  assign n4279 = n2372 & ~n4278 ;
  assign n4280 = n1605 & ~n4279 ;
  assign n4281 = n1609 & ~n4280 ;
  assign n4282 = n1613 & ~n4281 ;
  assign n4283 = n1617 & ~n4282 ;
  assign n4284 = n1621 & ~n4283 ;
  assign n4285 = n1625 & ~n4284 ;
  assign n4286 = n1629 & ~n4285 ;
  assign n4287 = n1633 & ~n4286 ;
  assign n4288 = n1637 & ~n4287 ;
  assign n4289 = n1641 & ~n4288 ;
  assign n4290 = n1645 & ~n4289 ;
  assign n4291 = n1649 & ~n4290 ;
  assign n4292 = n1170 & n4261 ;
  assign n4293 = ~n1651 & n4292 ;
  assign n4294 = ~n4291 & n4293 ;
  assign n4295 = ~n4262 & ~n4294 ;
  assign n4296 = \req[71]  & ~n464 ;
  assign n4297 = ~n450 & n4296 ;
  assign n4298 = ~\priority[73]  & ~n470 ;
  assign n4299 = n1198 & ~n4298 ;
  assign n4300 = n2004 & ~n4299 ;
  assign n4301 = n2009 & ~n4300 ;
  assign n4302 = n2013 & ~n4301 ;
  assign n4303 = n2017 & ~n4302 ;
  assign n4304 = n2021 & ~n4303 ;
  assign n4305 = n2025 & ~n4304 ;
  assign n4306 = n3671 & ~n4305 ;
  assign n4307 = n2033 & ~n4306 ;
  assign n4308 = n2037 & ~n4307 ;
  assign n4309 = n2041 & ~n4308 ;
  assign n4310 = n2045 & ~n4309 ;
  assign n4311 = n2049 & ~n4310 ;
  assign n4312 = n2053 & ~n4311 ;
  assign n4313 = n2408 & ~n4312 ;
  assign n4314 = n2411 & ~n4313 ;
  assign n4315 = n1721 & ~n4314 ;
  assign n4316 = n1725 & ~n4315 ;
  assign n4317 = n1729 & ~n4316 ;
  assign n4318 = n1733 & ~n4317 ;
  assign n4319 = n1737 & ~n4318 ;
  assign n4320 = n1741 & ~n4319 ;
  assign n4321 = n1745 & ~n4320 ;
  assign n4322 = n1749 & ~n4321 ;
  assign n4323 = n1753 & ~n4322 ;
  assign n4324 = n1757 & ~n4323 ;
  assign n4325 = n1761 & ~n4324 ;
  assign n4326 = n1765 & ~n4325 ;
  assign n4327 = n459 & n4296 ;
  assign n4328 = ~n1767 & n4327 ;
  assign n4329 = ~n4326 & n4328 ;
  assign n4330 = ~n4297 & ~n4329 ;
  assign n4331 = \req[72]  & ~n831 ;
  assign n4332 = ~n817 & n4331 ;
  assign n4333 = ~\priority[74]  & ~n837 ;
  assign n4334 = n462 & ~n4333 ;
  assign n4335 = n480 & ~n4334 ;
  assign n4336 = n494 & ~n4335 ;
  assign n4337 = n507 & ~n4336 ;
  assign n4338 = n520 & ~n4337 ;
  assign n4339 = n533 & ~n4338 ;
  assign n4340 = n546 & ~n4339 ;
  assign n4341 = n559 & ~n4340 ;
  assign n4342 = n572 & ~n4341 ;
  assign n4343 = n585 & ~n4342 ;
  assign n4344 = n598 & ~n4343 ;
  assign n4345 = n611 & ~n4344 ;
  assign n4346 = n2090 & ~n4345 ;
  assign n4347 = n2094 & ~n4346 ;
  assign n4348 = n2447 & ~n4347 ;
  assign n4349 = n2450 & ~n4348 ;
  assign n4350 = n1837 & ~n4349 ;
  assign n4351 = n1841 & ~n4350 ;
  assign n4352 = n1845 & ~n4351 ;
  assign n4353 = n1849 & ~n4352 ;
  assign n4354 = n3720 & ~n4353 ;
  assign n4355 = n1857 & ~n4354 ;
  assign n4356 = n1861 & ~n4355 ;
  assign n4357 = n1865 & ~n4356 ;
  assign n4358 = n1869 & ~n4357 ;
  assign n4359 = n1873 & ~n4358 ;
  assign n4360 = n1877 & ~n4359 ;
  assign n4361 = n3627 & ~n4360 ;
  assign n4362 = n826 & n4331 ;
  assign n4363 = ~n1883 & n4362 ;
  assign n4364 = ~n4361 & n4363 ;
  assign n4365 = ~n4332 & ~n4364 ;
  assign n4366 = \req[73]  & ~n1197 ;
  assign n4367 = ~n1183 & n4366 ;
  assign n4368 = ~\priority[75]  & ~n1203 ;
  assign n4369 = n829 & ~n4368 ;
  assign n4370 = n847 & ~n4369 ;
  assign n4371 = n861 & ~n4370 ;
  assign n4372 = n874 & ~n4371 ;
  assign n4373 = n887 & ~n4372 ;
  assign n4374 = n900 & ~n4373 ;
  assign n4375 = n913 & ~n4374 ;
  assign n4376 = n926 & ~n4375 ;
  assign n4377 = n939 & ~n4376 ;
  assign n4378 = n952 & ~n4377 ;
  assign n4379 = n965 & ~n4378 ;
  assign n4380 = n978 & ~n4379 ;
  assign n4381 = n2132 & ~n4380 ;
  assign n4382 = n2136 & ~n4381 ;
  assign n4383 = n2487 & ~n4382 ;
  assign n4384 = n2490 & ~n4383 ;
  assign n4385 = n1953 & ~n4384 ;
  assign n4386 = n1957 & ~n4385 ;
  assign n4387 = n1961 & ~n4386 ;
  assign n4388 = n1965 & ~n4387 ;
  assign n4389 = n1969 & ~n4388 ;
  assign n4390 = n1973 & ~n4389 ;
  assign n4391 = n2713 & ~n4390 ;
  assign n4392 = n1981 & ~n4391 ;
  assign n4393 = n1985 & ~n4392 ;
  assign n4394 = n1989 & ~n4393 ;
  assign n4395 = n1993 & ~n4394 ;
  assign n4396 = n1997 & ~n4395 ;
  assign n4397 = n1192 & n4366 ;
  assign n4398 = ~n1999 & n4397 ;
  assign n4399 = ~n4396 & n4398 ;
  assign n4400 = ~n4367 & ~n4399 ;
  assign n4401 = \req[74]  & ~n461 ;
  assign n4402 = ~n472 & n4401 ;
  assign n4403 = ~\priority[76]  & ~n477 ;
  assign n4404 = n1195 & ~n4403 ;
  assign n4405 = n1213 & ~n4404 ;
  assign n4406 = n1227 & ~n4405 ;
  assign n4407 = n1240 & ~n4406 ;
  assign n4408 = n1253 & ~n4407 ;
  assign n4409 = ~n1258 & n1265 ;
  assign n4410 = ~n4408 & n4409 ;
  assign n4411 = n1279 & ~n4410 ;
  assign n4412 = n1292 & ~n4411 ;
  assign n4413 = n1305 & ~n4412 ;
  assign n4414 = n3148 & ~n4413 ;
  assign n4415 = n1331 & ~n4414 ;
  assign n4416 = n1344 & ~n4415 ;
  assign n4417 = n2173 & ~n4416 ;
  assign n4418 = n2176 & ~n4417 ;
  assign n4419 = n286 & ~n4418 ;
  assign n4420 = n299 & ~n4419 ;
  assign n4421 = n312 & ~n4420 ;
  assign n4422 = n325 & ~n4421 ;
  assign n4423 = n338 & ~n4422 ;
  assign n4424 = n351 & ~n4423 ;
  assign n4425 = n364 & ~n4424 ;
  assign n4426 = n377 & ~n4425 ;
  assign n4427 = n390 & ~n4426 ;
  assign n4428 = n403 & ~n4427 ;
  assign n4429 = n416 & ~n4428 ;
  assign n4430 = n4115 & ~n4429 ;
  assign n4431 = n442 & ~n4430 ;
  assign n4432 = n455 & ~n4431 ;
  assign n4433 = n466 & n4401 ;
  assign n4434 = ~n460 & n4433 ;
  assign n4435 = ~n4432 & n4434 ;
  assign n4436 = ~n4402 & ~n4435 ;
  assign n4437 = \req[75]  & ~n828 ;
  assign n4438 = ~n839 & n4437 ;
  assign n4439 = ~\priority[77]  & ~n844 ;
  assign n4440 = n484 & ~n4439 ;
  assign n4441 = n1427 & ~n4440 ;
  assign n4442 = n1432 & ~n4441 ;
  assign n4443 = n1436 & ~n4442 ;
  assign n4444 = n1440 & ~n4443 ;
  assign n4445 = n3811 & ~n4444 ;
  assign n4446 = n1448 & ~n4445 ;
  assign n4447 = n1452 & ~n4446 ;
  assign n4448 = n1456 & ~n4447 ;
  assign n4449 = n3817 & ~n4448 ;
  assign n4450 = n1464 & ~n4449 ;
  assign n4451 = n1468 & ~n4450 ;
  assign n4452 = n2212 & ~n4451 ;
  assign n4453 = n640 & ~n2214 ;
  assign n4454 = ~n4452 & n4453 ;
  assign n4455 = n653 & ~n4454 ;
  assign n4456 = n666 & ~n4455 ;
  assign n4457 = n679 & ~n4456 ;
  assign n4458 = n3826 & ~n4457 ;
  assign n4459 = ~n697 & n704 ;
  assign n4460 = ~n4458 & n4459 ;
  assign n4461 = n718 & ~n4460 ;
  assign n4462 = n731 & ~n4461 ;
  assign n4463 = n739 & n742 ;
  assign n4464 = ~n736 & n4463 ;
  assign n4465 = ~n4462 & n4464 ;
  assign n4466 = n2465 & ~n4465 ;
  assign n4467 = n770 & ~n4466 ;
  assign n4468 = n3099 & ~n4467 ;
  assign n4469 = n796 & ~n4468 ;
  assign n4470 = n809 & ~n4469 ;
  assign n4471 = n2117 & ~n4470 ;
  assign n4472 = n833 & n4437 ;
  assign n4473 = ~n827 & n4472 ;
  assign n4474 = ~n4471 & n4473 ;
  assign n4475 = ~n4438 & ~n4474 ;
  assign n4476 = \req[76]  & ~n1194 ;
  assign n4477 = ~n1205 & n4476 ;
  assign n4478 = ~\priority[78]  & ~n1210 ;
  assign n4479 = n851 & ~n4478 ;
  assign n4480 = n1547 & ~n4479 ;
  assign n4481 = n1552 & ~n4480 ;
  assign n4482 = n1556 & ~n4481 ;
  assign n4483 = n1560 & ~n4482 ;
  assign n4484 = n1564 & ~n4483 ;
  assign n4485 = n1568 & ~n4484 ;
  assign n4486 = n1572 & ~n4485 ;
  assign n4487 = n1576 & ~n4486 ;
  assign n4488 = n1580 & ~n4487 ;
  assign n4489 = n1584 & ~n4488 ;
  assign n4490 = n1588 & ~n4489 ;
  assign n4491 = n2252 & ~n4490 ;
  assign n4492 = n2255 & ~n4491 ;
  assign n4493 = n1019 & ~n4492 ;
  assign n4494 = n1032 & ~n4493 ;
  assign n4495 = n3861 & ~n4494 ;
  assign n4496 = n1058 & ~n4495 ;
  assign n4497 = n1071 & ~n4496 ;
  assign n4498 = n1084 & ~n4497 ;
  assign n4499 = n1097 & ~n4498 ;
  assign n4500 = n1110 & ~n4499 ;
  assign n4501 = n1123 & ~n4500 ;
  assign n4502 = n1136 & ~n4501 ;
  assign n4503 = n1149 & ~n4502 ;
  assign n4504 = n1162 & ~n4503 ;
  assign n4505 = n1175 & ~n4504 ;
  assign n4506 = n1188 & ~n4505 ;
  assign n4507 = n1199 & n4476 ;
  assign n4508 = ~n1193 & n4507 ;
  assign n4509 = ~n4506 & n4508 ;
  assign n4510 = ~n4477 & ~n4509 ;
  assign n4511 = \req[77]  & ~n483 ;
  assign n4512 = ~n479 & n4511 ;
  assign n4513 = ~\priority[79]  & ~n474 ;
  assign n4514 = n1217 & ~n4513 ;
  assign n4515 = n1664 & ~n4514 ;
  assign n4516 = n1669 & ~n4515 ;
  assign n4517 = n1673 & ~n4516 ;
  assign n4518 = n1677 & ~n4517 ;
  assign n4519 = n1681 & ~n4518 ;
  assign n4520 = n1685 & ~n4519 ;
  assign n4521 = n1689 & ~n4520 ;
  assign n4522 = n1693 & ~n4521 ;
  assign n4523 = n1697 & ~n4522 ;
  assign n4524 = n1701 & ~n4523 ;
  assign n4525 = n3570 & ~n4524 ;
  assign n4526 = n2291 & ~n4525 ;
  assign n4527 = n2294 & ~n4526 ;
  assign n4528 = n1368 & ~n4527 ;
  assign n4529 = n1372 & ~n4528 ;
  assign n4530 = n1376 & ~n4529 ;
  assign n4531 = n1380 & ~n4530 ;
  assign n4532 = n1384 & ~n4531 ;
  assign n4533 = n1388 & ~n4532 ;
  assign n4534 = n1392 & ~n4533 ;
  assign n4535 = n1396 & ~n4534 ;
  assign n4536 = n1400 & ~n4535 ;
  assign n4537 = n1404 & ~n4536 ;
  assign n4538 = n1408 & ~n4537 ;
  assign n4539 = n1412 & ~n4538 ;
  assign n4540 = n1416 & ~n4539 ;
  assign n4541 = n1420 & ~n4540 ;
  assign n4542 = n463 & n4511 ;
  assign n4543 = ~n1422 & n4542 ;
  assign n4544 = ~n4541 & n4543 ;
  assign n4545 = ~n4512 & ~n4544 ;
  assign n4546 = \req[78]  & ~n850 ;
  assign n4547 = ~n846 & n4546 ;
  assign n4548 = ~\priority[80]  & ~n841 ;
  assign n4549 = n491 & ~n4548 ;
  assign n4550 = n1780 & ~n4549 ;
  assign n4551 = n1785 & ~n4550 ;
  assign n4552 = n1789 & ~n4551 ;
  assign n4553 = n3920 & ~n4552 ;
  assign n4554 = n1797 & ~n4553 ;
  assign n4555 = n1801 & ~n4554 ;
  assign n4556 = n1805 & ~n4555 ;
  assign n4557 = n589 & n596 ;
  assign n4558 = ~n1807 & n4557 ;
  assign n4559 = ~n4556 & n4558 ;
  assign n4560 = n1813 & ~n4559 ;
  assign n4561 = n1817 & ~n4560 ;
  assign n4562 = n1821 & ~n4561 ;
  assign n4563 = n2330 & ~n4562 ;
  assign n4564 = n2333 & ~n4563 ;
  assign n4565 = n1488 & ~n4564 ;
  assign n4566 = n1492 & ~n4565 ;
  assign n4567 = n1496 & ~n4566 ;
  assign n4568 = n1500 & ~n4567 ;
  assign n4569 = n1504 & ~n4568 ;
  assign n4570 = n2229 & ~n4569 ;
  assign n4571 = n1512 & ~n4570 ;
  assign n4572 = n1516 & ~n4571 ;
  assign n4573 = n1520 & ~n4572 ;
  assign n4574 = n1524 & ~n4573 ;
  assign n4575 = n1528 & ~n4574 ;
  assign n4576 = n1532 & ~n4575 ;
  assign n4577 = n1536 & ~n4576 ;
  assign n4578 = n1540 & ~n4577 ;
  assign n4579 = n830 & n4546 ;
  assign n4580 = ~n1542 & n4579 ;
  assign n4581 = ~n4578 & n4580 ;
  assign n4582 = ~n4547 & ~n4581 ;
  assign n4583 = \req[79]  & ~n1216 ;
  assign n4584 = ~n1212 & n4583 ;
  assign n4585 = ~\priority[81]  & ~n1207 ;
  assign n4586 = n858 & ~n4585 ;
  assign n4587 = n1896 & ~n4586 ;
  assign n4588 = n1901 & ~n4587 ;
  assign n4589 = n1905 & ~n4588 ;
  assign n4590 = n1909 & ~n4589 ;
  assign n4591 = ~n895 & n911 ;
  assign n4592 = n1912 & ~n4591 ;
  assign n4593 = ~n4590 & n4592 ;
  assign n4594 = n1917 & ~n4593 ;
  assign n4595 = n1921 & ~n4594 ;
  assign n4596 = n1925 & ~n4595 ;
  assign n4597 = n1929 & ~n4596 ;
  assign n4598 = n1933 & ~n4597 ;
  assign n4599 = n1937 & ~n4598 ;
  assign n4600 = n2369 & ~n4599 ;
  assign n4601 = n2372 & ~n4600 ;
  assign n4602 = n1605 & ~n4601 ;
  assign n4603 = n1609 & ~n4602 ;
  assign n4604 = n1613 & ~n4603 ;
  assign n4605 = n1617 & ~n4604 ;
  assign n4606 = n1621 & ~n4605 ;
  assign n4607 = n1625 & ~n4606 ;
  assign n4608 = n1629 & ~n4607 ;
  assign n4609 = n1633 & ~n4608 ;
  assign n4610 = n1637 & ~n4609 ;
  assign n4611 = n1641 & ~n4610 ;
  assign n4612 = n1645 & ~n4611 ;
  assign n4613 = n1649 & ~n4612 ;
  assign n4614 = ~n1651 & n1652 ;
  assign n4615 = ~n4613 & n4614 ;
  assign n4616 = n1657 & ~n4615 ;
  assign n4617 = n1196 & n4583 ;
  assign n4618 = ~n1659 & n4617 ;
  assign n4619 = ~n4616 & n4618 ;
  assign n4620 = ~n4584 & ~n4619 ;
  assign n4621 = \req[80]  & ~n490 ;
  assign n4622 = ~n476 & n4621 ;
  assign n4623 = ~\priority[82]  & ~n496 ;
  assign n4624 = n1224 & ~n4623 ;
  assign n4625 = n2012 & ~n4624 ;
  assign n4626 = n2017 & ~n4625 ;
  assign n4627 = n2021 & ~n4626 ;
  assign n4628 = n2025 & ~n4627 ;
  assign n4629 = n3671 & ~n4628 ;
  assign n4630 = n2033 & ~n4629 ;
  assign n4631 = n2037 & ~n4630 ;
  assign n4632 = n2041 & ~n4631 ;
  assign n4633 = n2045 & ~n4632 ;
  assign n4634 = n2049 & ~n4633 ;
  assign n4635 = n2053 & ~n4634 ;
  assign n4636 = n2408 & ~n4635 ;
  assign n4637 = n2411 & ~n4636 ;
  assign n4638 = n1721 & ~n4637 ;
  assign n4639 = n1725 & ~n4638 ;
  assign n4640 = n1729 & ~n4639 ;
  assign n4641 = n1733 & ~n4640 ;
  assign n4642 = n1737 & ~n4641 ;
  assign n4643 = n1741 & ~n4642 ;
  assign n4644 = n1745 & ~n4643 ;
  assign n4645 = n1749 & ~n4644 ;
  assign n4646 = n1753 & ~n4645 ;
  assign n4647 = n1757 & ~n4646 ;
  assign n4648 = n1761 & ~n4647 ;
  assign n4649 = n1765 & ~n4648 ;
  assign n4650 = n1769 & ~n4649 ;
  assign n4651 = n1773 & ~n4650 ;
  assign n4652 = n485 & n4621 ;
  assign n4653 = ~n1775 & n4652 ;
  assign n4654 = ~n4651 & n4653 ;
  assign n4655 = ~n4622 & ~n4654 ;
  assign n4656 = \req[81]  & ~n857 ;
  assign n4657 = ~n843 & n4656 ;
  assign n4658 = ~\priority[83]  & ~n863 ;
  assign n4659 = n488 & ~n4658 ;
  assign n4660 = n506 & ~n4659 ;
  assign n4661 = n520 & ~n4660 ;
  assign n4662 = n533 & ~n4661 ;
  assign n4663 = n546 & ~n4662 ;
  assign n4664 = n559 & ~n4663 ;
  assign n4665 = n572 & ~n4664 ;
  assign n4666 = n585 & ~n4665 ;
  assign n4667 = n598 & ~n4666 ;
  assign n4668 = n611 & ~n4667 ;
  assign n4669 = n2090 & ~n4668 ;
  assign n4670 = n2094 & ~n4669 ;
  assign n4671 = n2447 & ~n4670 ;
  assign n4672 = n2450 & ~n4671 ;
  assign n4673 = n1837 & ~n4672 ;
  assign n4674 = n1841 & ~n4673 ;
  assign n4675 = n1845 & ~n4674 ;
  assign n4676 = n1849 & ~n4675 ;
  assign n4677 = n3720 & ~n4676 ;
  assign n4678 = n1857 & ~n4677 ;
  assign n4679 = n1861 & ~n4678 ;
  assign n4680 = n1865 & ~n4679 ;
  assign n4681 = n1869 & ~n4680 ;
  assign n4682 = n1873 & ~n4681 ;
  assign n4683 = n1877 & ~n4682 ;
  assign n4684 = n3627 & ~n4683 ;
  assign n4685 = n1885 & ~n4684 ;
  assign n4686 = n1889 & ~n4685 ;
  assign n4687 = n852 & n4656 ;
  assign n4688 = ~n1891 & n4687 ;
  assign n4689 = ~n4686 & n4688 ;
  assign n4690 = ~n4657 & ~n4689 ;
  assign n4691 = \req[82]  & ~n1223 ;
  assign n4692 = ~n1209 & n4691 ;
  assign n4693 = ~\priority[84]  & ~n1229 ;
  assign n4694 = n855 & ~n4693 ;
  assign n4695 = n873 & ~n4694 ;
  assign n4696 = n887 & ~n4695 ;
  assign n4697 = n900 & ~n4696 ;
  assign n4698 = n913 & ~n4697 ;
  assign n4699 = n926 & ~n4698 ;
  assign n4700 = n939 & ~n4699 ;
  assign n4701 = n952 & ~n4700 ;
  assign n4702 = n965 & ~n4701 ;
  assign n4703 = n978 & ~n4702 ;
  assign n4704 = n2132 & ~n4703 ;
  assign n4705 = n2136 & ~n4704 ;
  assign n4706 = n2487 & ~n4705 ;
  assign n4707 = n2490 & ~n4706 ;
  assign n4708 = n1953 & ~n4707 ;
  assign n4709 = n1957 & ~n4708 ;
  assign n4710 = n1961 & ~n4709 ;
  assign n4711 = n1965 & ~n4710 ;
  assign n4712 = n1969 & ~n4711 ;
  assign n4713 = n1973 & ~n4712 ;
  assign n4714 = n2713 & ~n4713 ;
  assign n4715 = n1981 & ~n4714 ;
  assign n4716 = n1985 & ~n4715 ;
  assign n4717 = n1989 & ~n4716 ;
  assign n4718 = n1993 & ~n4717 ;
  assign n4719 = n1997 & ~n4718 ;
  assign n4720 = n2001 & ~n4719 ;
  assign n4721 = n2005 & ~n4720 ;
  assign n4722 = n1218 & n4691 ;
  assign n4723 = ~n2007 & n4722 ;
  assign n4724 = ~n4721 & n4723 ;
  assign n4725 = ~n4692 & ~n4724 ;
  assign n4726 = \req[83]  & ~n487 ;
  assign n4727 = ~n498 & n4726 ;
  assign n4728 = ~\priority[85]  & ~n503 ;
  assign n4729 = n1221 & ~n4728 ;
  assign n4730 = n1239 & ~n4729 ;
  assign n4731 = n1253 & ~n4730 ;
  assign n4732 = n4409 & ~n4731 ;
  assign n4733 = n1279 & ~n4732 ;
  assign n4734 = n1292 & ~n4733 ;
  assign n4735 = n1305 & ~n4734 ;
  assign n4736 = n3148 & ~n4735 ;
  assign n4737 = n1331 & ~n4736 ;
  assign n4738 = n1344 & ~n4737 ;
  assign n4739 = n2173 & ~n4738 ;
  assign n4740 = n2176 & ~n4739 ;
  assign n4741 = n286 & ~n4740 ;
  assign n4742 = n299 & ~n4741 ;
  assign n4743 = n312 & ~n4742 ;
  assign n4744 = n325 & ~n4743 ;
  assign n4745 = n338 & ~n4744 ;
  assign n4746 = n351 & ~n4745 ;
  assign n4747 = n364 & ~n4746 ;
  assign n4748 = n377 & ~n4747 ;
  assign n4749 = n390 & ~n4748 ;
  assign n4750 = n403 & ~n4749 ;
  assign n4751 = n416 & ~n4750 ;
  assign n4752 = n4115 & ~n4751 ;
  assign n4753 = n442 & ~n4752 ;
  assign n4754 = n455 & ~n4753 ;
  assign n4755 = n468 & ~n4754 ;
  assign n4756 = n481 & ~n4755 ;
  assign n4757 = n492 & n4726 ;
  assign n4758 = ~n486 & n4757 ;
  assign n4759 = ~n4756 & n4758 ;
  assign n4760 = ~n4727 & ~n4759 ;
  assign n4761 = \req[84]  & ~n854 ;
  assign n4762 = ~n865 & n4761 ;
  assign n4763 = ~\priority[86]  & ~n870 ;
  assign n4764 = n510 & ~n4763 ;
  assign n4765 = n1435 & ~n4764 ;
  assign n4766 = n1440 & ~n4765 ;
  assign n4767 = n3811 & ~n4766 ;
  assign n4768 = n1448 & ~n4767 ;
  assign n4769 = n1452 & ~n4768 ;
  assign n4770 = n1456 & ~n4769 ;
  assign n4771 = n3817 & ~n4770 ;
  assign n4772 = n1464 & ~n4771 ;
  assign n4773 = n1468 & ~n4772 ;
  assign n4774 = n2212 & ~n4773 ;
  assign n4775 = n4453 & ~n4774 ;
  assign n4776 = n653 & ~n4775 ;
  assign n4777 = n666 & ~n4776 ;
  assign n4778 = n679 & ~n4777 ;
  assign n4779 = n3826 & ~n4778 ;
  assign n4780 = n4459 & ~n4779 ;
  assign n4781 = n718 & ~n4780 ;
  assign n4782 = n731 & ~n4781 ;
  assign n4783 = n4464 & ~n4782 ;
  assign n4784 = n2465 & ~n4783 ;
  assign n4785 = n770 & ~n4784 ;
  assign n4786 = n3099 & ~n4785 ;
  assign n4787 = n796 & ~n4786 ;
  assign n4788 = n809 & ~n4787 ;
  assign n4789 = n2117 & ~n4788 ;
  assign n4790 = n835 & ~n4789 ;
  assign n4791 = n848 & ~n4790 ;
  assign n4792 = n859 & n4761 ;
  assign n4793 = ~n853 & n4792 ;
  assign n4794 = ~n4791 & n4793 ;
  assign n4795 = ~n4762 & ~n4794 ;
  assign n4796 = \req[85]  & ~n1220 ;
  assign n4797 = ~n1231 & n4796 ;
  assign n4798 = ~\priority[87]  & ~n1236 ;
  assign n4799 = n877 & ~n4798 ;
  assign n4800 = n1555 & ~n4799 ;
  assign n4801 = n1560 & ~n4800 ;
  assign n4802 = n1564 & ~n4801 ;
  assign n4803 = n1568 & ~n4802 ;
  assign n4804 = n1572 & ~n4803 ;
  assign n4805 = n1576 & ~n4804 ;
  assign n4806 = n1580 & ~n4805 ;
  assign n4807 = n1584 & ~n4806 ;
  assign n4808 = n1588 & ~n4807 ;
  assign n4809 = n2252 & ~n4808 ;
  assign n4810 = n2255 & ~n4809 ;
  assign n4811 = n1019 & ~n4810 ;
  assign n4812 = n1032 & ~n4811 ;
  assign n4813 = n3861 & ~n4812 ;
  assign n4814 = n1058 & ~n4813 ;
  assign n4815 = n1071 & ~n4814 ;
  assign n4816 = n1084 & ~n4815 ;
  assign n4817 = n1097 & ~n4816 ;
  assign n4818 = n1110 & ~n4817 ;
  assign n4819 = n1123 & ~n4818 ;
  assign n4820 = n1136 & ~n4819 ;
  assign n4821 = n1149 & ~n4820 ;
  assign n4822 = n1162 & ~n4821 ;
  assign n4823 = n1175 & ~n4822 ;
  assign n4824 = n1188 & ~n4823 ;
  assign n4825 = n1201 & ~n4824 ;
  assign n4826 = n1214 & ~n4825 ;
  assign n4827 = n1225 & n4796 ;
  assign n4828 = ~n1219 & n4827 ;
  assign n4829 = ~n4826 & n4828 ;
  assign n4830 = ~n4797 & ~n4829 ;
  assign n4831 = \req[86]  & ~n509 ;
  assign n4832 = ~n505 & n4831 ;
  assign n4833 = ~\priority[88]  & ~n500 ;
  assign n4834 = n1243 & ~n4833 ;
  assign n4835 = n1672 & ~n4834 ;
  assign n4836 = n1677 & ~n4835 ;
  assign n4837 = n1681 & ~n4836 ;
  assign n4838 = n1685 & ~n4837 ;
  assign n4839 = n1689 & ~n4838 ;
  assign n4840 = n1693 & ~n4839 ;
  assign n4841 = n1697 & ~n4840 ;
  assign n4842 = n1701 & ~n4841 ;
  assign n4843 = n3570 & ~n4842 ;
  assign n4844 = n2291 & ~n4843 ;
  assign n4845 = n2294 & ~n4844 ;
  assign n4846 = n1368 & ~n4845 ;
  assign n4847 = n1372 & ~n4846 ;
  assign n4848 = n1376 & ~n4847 ;
  assign n4849 = n1380 & ~n4848 ;
  assign n4850 = n1384 & ~n4849 ;
  assign n4851 = n1388 & ~n4850 ;
  assign n4852 = n1392 & ~n4851 ;
  assign n4853 = n1396 & ~n4852 ;
  assign n4854 = n1400 & ~n4853 ;
  assign n4855 = n1404 & ~n4854 ;
  assign n4856 = n1408 & ~n4855 ;
  assign n4857 = n1412 & ~n4856 ;
  assign n4858 = n1416 & ~n4857 ;
  assign n4859 = n1420 & ~n4858 ;
  assign n4860 = n1424 & ~n4859 ;
  assign n4861 = n1428 & ~n4860 ;
  assign n4862 = n489 & n4831 ;
  assign n4863 = ~n1430 & n4862 ;
  assign n4864 = ~n4861 & n4863 ;
  assign n4865 = ~n4832 & ~n4864 ;
  assign n4866 = \req[87]  & ~n876 ;
  assign n4867 = ~n872 & n4866 ;
  assign n4868 = ~\priority[89]  & ~n867 ;
  assign n4869 = n517 & ~n4868 ;
  assign n4870 = n1788 & ~n4869 ;
  assign n4871 = n3920 & ~n4870 ;
  assign n4872 = n1797 & ~n4871 ;
  assign n4873 = n1801 & ~n4872 ;
  assign n4874 = n1805 & ~n4873 ;
  assign n4875 = n4558 & ~n4874 ;
  assign n4876 = n1813 & ~n4875 ;
  assign n4877 = n1817 & ~n4876 ;
  assign n4878 = n1821 & ~n4877 ;
  assign n4879 = n2330 & ~n4878 ;
  assign n4880 = n2333 & ~n4879 ;
  assign n4881 = n1488 & ~n4880 ;
  assign n4882 = n1492 & ~n4881 ;
  assign n4883 = n1496 & ~n4882 ;
  assign n4884 = n1500 & ~n4883 ;
  assign n4885 = n1504 & ~n4884 ;
  assign n4886 = n2229 & ~n4885 ;
  assign n4887 = n1512 & ~n4886 ;
  assign n4888 = n1516 & ~n4887 ;
  assign n4889 = n1520 & ~n4888 ;
  assign n4890 = n1524 & ~n4889 ;
  assign n4891 = n1528 & ~n4890 ;
  assign n4892 = n1532 & ~n4891 ;
  assign n4893 = n1536 & ~n4892 ;
  assign n4894 = n1540 & ~n4893 ;
  assign n4895 = n1544 & ~n4894 ;
  assign n4896 = n1548 & ~n4895 ;
  assign n4897 = n856 & n4866 ;
  assign n4898 = ~n1550 & n4897 ;
  assign n4899 = ~n4896 & n4898 ;
  assign n4900 = ~n4867 & ~n4899 ;
  assign n4901 = \req[88]  & ~n1242 ;
  assign n4902 = ~n1238 & n4901 ;
  assign n4903 = ~\priority[90]  & ~n1233 ;
  assign n4904 = n884 & ~n4903 ;
  assign n4905 = n1904 & ~n4904 ;
  assign n4906 = n1909 & ~n4905 ;
  assign n4907 = n4592 & ~n4906 ;
  assign n4908 = n1917 & ~n4907 ;
  assign n4909 = n1921 & ~n4908 ;
  assign n4910 = n1925 & ~n4909 ;
  assign n4911 = n1929 & ~n4910 ;
  assign n4912 = n1933 & ~n4911 ;
  assign n4913 = n1937 & ~n4912 ;
  assign n4914 = n2369 & ~n4913 ;
  assign n4915 = n2372 & ~n4914 ;
  assign n4916 = n1605 & ~n4915 ;
  assign n4917 = n1609 & ~n4916 ;
  assign n4918 = n1613 & ~n4917 ;
  assign n4919 = n1617 & ~n4918 ;
  assign n4920 = n1621 & ~n4919 ;
  assign n4921 = n1625 & ~n4920 ;
  assign n4922 = n1629 & ~n4921 ;
  assign n4923 = n1633 & ~n4922 ;
  assign n4924 = n1637 & ~n4923 ;
  assign n4925 = n1641 & ~n4924 ;
  assign n4926 = n1645 & ~n4925 ;
  assign n4927 = n1649 & ~n4926 ;
  assign n4928 = n4614 & ~n4927 ;
  assign n4929 = n1657 & ~n4928 ;
  assign n4930 = ~n1659 & n1660 ;
  assign n4931 = ~n4929 & n4930 ;
  assign n4932 = n1665 & ~n4931 ;
  assign n4933 = n1222 & n4901 ;
  assign n4934 = ~n1667 & n4933 ;
  assign n4935 = ~n4932 & n4934 ;
  assign n4936 = ~n4902 & ~n4935 ;
  assign n4937 = \req[89]  & ~n516 ;
  assign n4938 = ~n502 & n4937 ;
  assign n4939 = ~\priority[91]  & ~n522 ;
  assign n4940 = n1250 & ~n4939 ;
  assign n4941 = n2020 & ~n4940 ;
  assign n4942 = n2025 & ~n4941 ;
  assign n4943 = n3671 & ~n4942 ;
  assign n4944 = n2033 & ~n4943 ;
  assign n4945 = n2037 & ~n4944 ;
  assign n4946 = n2041 & ~n4945 ;
  assign n4947 = n2045 & ~n4946 ;
  assign n4948 = n2049 & ~n4947 ;
  assign n4949 = n2053 & ~n4948 ;
  assign n4950 = n2408 & ~n4949 ;
  assign n4951 = n2411 & ~n4950 ;
  assign n4952 = n1721 & ~n4951 ;
  assign n4953 = n1725 & ~n4952 ;
  assign n4954 = n1729 & ~n4953 ;
  assign n4955 = n1733 & ~n4954 ;
  assign n4956 = n1737 & ~n4955 ;
  assign n4957 = n1741 & ~n4956 ;
  assign n4958 = n1745 & ~n4957 ;
  assign n4959 = n1749 & ~n4958 ;
  assign n4960 = n1753 & ~n4959 ;
  assign n4961 = n1757 & ~n4960 ;
  assign n4962 = n1761 & ~n4961 ;
  assign n4963 = n1765 & ~n4962 ;
  assign n4964 = n1769 & ~n4963 ;
  assign n4965 = n1773 & ~n4964 ;
  assign n4966 = n1777 & ~n4965 ;
  assign n4967 = n1781 & ~n4966 ;
  assign n4968 = n511 & n4937 ;
  assign n4969 = ~n1783 & n4968 ;
  assign n4970 = ~n4967 & n4969 ;
  assign n4971 = ~n4938 & ~n4970 ;
  assign n4972 = \req[90]  & ~n883 ;
  assign n4973 = ~n869 & n4972 ;
  assign n4974 = ~\priority[92]  & ~n889 ;
  assign n4975 = n514 & ~n4974 ;
  assign n4976 = n532 & ~n4975 ;
  assign n4977 = n546 & ~n4976 ;
  assign n4978 = n559 & ~n4977 ;
  assign n4979 = n572 & ~n4978 ;
  assign n4980 = n585 & ~n4979 ;
  assign n4981 = n598 & ~n4980 ;
  assign n4982 = n611 & ~n4981 ;
  assign n4983 = n2090 & ~n4982 ;
  assign n4984 = n2094 & ~n4983 ;
  assign n4985 = n2447 & ~n4984 ;
  assign n4986 = n2450 & ~n4985 ;
  assign n4987 = n1837 & ~n4986 ;
  assign n4988 = n1841 & ~n4987 ;
  assign n4989 = n1845 & ~n4988 ;
  assign n4990 = n1849 & ~n4989 ;
  assign n4991 = n3720 & ~n4990 ;
  assign n4992 = n1857 & ~n4991 ;
  assign n4993 = n1861 & ~n4992 ;
  assign n4994 = n1865 & ~n4993 ;
  assign n4995 = n1869 & ~n4994 ;
  assign n4996 = n1873 & ~n4995 ;
  assign n4997 = n1877 & ~n4996 ;
  assign n4998 = n3627 & ~n4997 ;
  assign n4999 = n1885 & ~n4998 ;
  assign n5000 = n1889 & ~n4999 ;
  assign n5001 = n1893 & ~n5000 ;
  assign n5002 = n1897 & ~n5001 ;
  assign n5003 = n878 & n4972 ;
  assign n5004 = ~n1899 & n5003 ;
  assign n5005 = ~n5002 & n5004 ;
  assign n5006 = ~n4973 & ~n5005 ;
  assign n5007 = \req[91]  & ~n1249 ;
  assign n5008 = ~n1235 & n5007 ;
  assign n5009 = ~\priority[93]  & ~n1255 ;
  assign n5010 = n881 & ~n5009 ;
  assign n5011 = n899 & ~n5010 ;
  assign n5012 = n913 & ~n5011 ;
  assign n5013 = n926 & ~n5012 ;
  assign n5014 = n939 & ~n5013 ;
  assign n5015 = n952 & ~n5014 ;
  assign n5016 = n965 & ~n5015 ;
  assign n5017 = n978 & ~n5016 ;
  assign n5018 = n2132 & ~n5017 ;
  assign n5019 = n2136 & ~n5018 ;
  assign n5020 = n2487 & ~n5019 ;
  assign n5021 = n2490 & ~n5020 ;
  assign n5022 = n1953 & ~n5021 ;
  assign n5023 = n1957 & ~n5022 ;
  assign n5024 = n1961 & ~n5023 ;
  assign n5025 = n1965 & ~n5024 ;
  assign n5026 = n1969 & ~n5025 ;
  assign n5027 = n1973 & ~n5026 ;
  assign n5028 = n2713 & ~n5027 ;
  assign n5029 = n1981 & ~n5028 ;
  assign n5030 = n1985 & ~n5029 ;
  assign n5031 = n1989 & ~n5030 ;
  assign n5032 = n1993 & ~n5031 ;
  assign n5033 = n1997 & ~n5032 ;
  assign n5034 = n2001 & ~n5033 ;
  assign n5035 = n2005 & ~n5034 ;
  assign n5036 = n2009 & ~n5035 ;
  assign n5037 = n2013 & ~n5036 ;
  assign n5038 = n1244 & n5007 ;
  assign n5039 = ~n2015 & n5038 ;
  assign n5040 = ~n5037 & n5039 ;
  assign n5041 = ~n5008 & ~n5040 ;
  assign n5042 = \req[92]  & ~n513 ;
  assign n5043 = ~n524 & n5042 ;
  assign n5044 = ~\priority[94]  & ~n529 ;
  assign n5045 = n1247 & ~n5044 ;
  assign n5046 = n1265 & ~n5045 ;
  assign n5047 = n1279 & ~n5046 ;
  assign n5048 = n1292 & ~n5047 ;
  assign n5049 = n1305 & ~n5048 ;
  assign n5050 = n3148 & ~n5049 ;
  assign n5051 = n1331 & ~n5050 ;
  assign n5052 = n1344 & ~n5051 ;
  assign n5053 = n2173 & ~n5052 ;
  assign n5054 = n2176 & ~n5053 ;
  assign n5055 = n286 & ~n5054 ;
  assign n5056 = n299 & ~n5055 ;
  assign n5057 = n312 & ~n5056 ;
  assign n5058 = n325 & ~n5057 ;
  assign n5059 = n338 & ~n5058 ;
  assign n5060 = n351 & ~n5059 ;
  assign n5061 = n364 & ~n5060 ;
  assign n5062 = n377 & ~n5061 ;
  assign n5063 = n390 & ~n5062 ;
  assign n5064 = ~n395 & n402 ;
  assign n5065 = ~n5063 & n5064 ;
  assign n5066 = n416 & ~n5065 ;
  assign n5067 = n4115 & ~n5066 ;
  assign n5068 = n442 & ~n5067 ;
  assign n5069 = n455 & ~n5068 ;
  assign n5070 = n468 & ~n5069 ;
  assign n5071 = n481 & ~n5070 ;
  assign n5072 = n494 & ~n5071 ;
  assign n5073 = n507 & ~n5072 ;
  assign n5074 = n518 & n5042 ;
  assign n5075 = ~n512 & n5074 ;
  assign n5076 = ~n5073 & n5075 ;
  assign n5077 = ~n5043 & ~n5076 ;
  assign n5078 = \req[93]  & ~n880 ;
  assign n5079 = ~n891 & n5078 ;
  assign n5080 = ~\priority[95]  & ~n896 ;
  assign n5081 = n536 & ~n5080 ;
  assign n5082 = n1443 & ~n5081 ;
  assign n5083 = n1448 & ~n5082 ;
  assign n5084 = n1452 & ~n5083 ;
  assign n5085 = n1456 & ~n5084 ;
  assign n5086 = n3817 & ~n5085 ;
  assign n5087 = n1464 & ~n5086 ;
  assign n5088 = n1468 & ~n5087 ;
  assign n5089 = n2212 & ~n5088 ;
  assign n5090 = n4453 & ~n5089 ;
  assign n5091 = n653 & ~n5090 ;
  assign n5092 = n666 & ~n5091 ;
  assign n5093 = n679 & ~n5092 ;
  assign n5094 = n3826 & ~n5093 ;
  assign n5095 = n4459 & ~n5094 ;
  assign n5096 = n718 & ~n5095 ;
  assign n5097 = n731 & ~n5096 ;
  assign n5098 = n4464 & ~n5097 ;
  assign n5099 = n2465 & ~n5098 ;
  assign n5100 = n770 & ~n5099 ;
  assign n5101 = n3099 & ~n5100 ;
  assign n5102 = n796 & ~n5101 ;
  assign n5103 = n809 & ~n5102 ;
  assign n5104 = n2117 & ~n5103 ;
  assign n5105 = n835 & ~n5104 ;
  assign n5106 = n848 & ~n5105 ;
  assign n5107 = ~n853 & n860 ;
  assign n5108 = ~n5106 & n5107 ;
  assign n5109 = n874 & ~n5108 ;
  assign n5110 = n885 & n5078 ;
  assign n5111 = ~n879 & n5110 ;
  assign n5112 = ~n5109 & n5111 ;
  assign n5113 = ~n5079 & ~n5112 ;
  assign n5114 = \req[94]  & ~n1246 ;
  assign n5115 = ~n1257 & n5114 ;
  assign n5116 = ~\priority[96]  & ~n1262 ;
  assign n5117 = n903 & ~n5116 ;
  assign n5118 = n1563 & ~n5117 ;
  assign n5119 = n1568 & ~n5118 ;
  assign n5120 = n1572 & ~n5119 ;
  assign n5121 = n1576 & ~n5120 ;
  assign n5122 = n1580 & ~n5121 ;
  assign n5123 = n1584 & ~n5122 ;
  assign n5124 = n1588 & ~n5123 ;
  assign n5125 = n2252 & ~n5124 ;
  assign n5126 = n2255 & ~n5125 ;
  assign n5127 = n1019 & ~n5126 ;
  assign n5128 = n1032 & ~n5127 ;
  assign n5129 = n3861 & ~n5128 ;
  assign n5130 = n1058 & ~n5129 ;
  assign n5131 = n1071 & ~n5130 ;
  assign n5132 = n1084 & ~n5131 ;
  assign n5133 = n1097 & ~n5132 ;
  assign n5134 = n1110 & ~n5133 ;
  assign n5135 = n1123 & ~n5134 ;
  assign n5136 = n1136 & ~n5135 ;
  assign n5137 = ~n1141 & n1148 ;
  assign n5138 = ~n5136 & n5137 ;
  assign n5139 = n1162 & ~n5138 ;
  assign n5140 = n1175 & ~n5139 ;
  assign n5141 = n1188 & ~n5140 ;
  assign n5142 = n1201 & ~n5141 ;
  assign n5143 = n1214 & ~n5142 ;
  assign n5144 = n1227 & ~n5143 ;
  assign n5145 = n1240 & ~n5144 ;
  assign n5146 = n1251 & n5114 ;
  assign n5147 = ~n1245 & n5146 ;
  assign n5148 = ~n5145 & n5147 ;
  assign n5149 = ~n5115 & ~n5148 ;
  assign n5150 = \req[95]  & ~n535 ;
  assign n5151 = ~n531 & n5150 ;
  assign n5152 = ~\priority[97]  & ~n526 ;
  assign n5153 = n1269 & ~n5152 ;
  assign n5154 = n1680 & ~n5153 ;
  assign n5155 = n1685 & ~n5154 ;
  assign n5156 = n1689 & ~n5155 ;
  assign n5157 = n1693 & ~n5156 ;
  assign n5158 = n1697 & ~n5157 ;
  assign n5159 = n1701 & ~n5158 ;
  assign n5160 = n3570 & ~n5159 ;
  assign n5161 = n2291 & ~n5160 ;
  assign n5162 = n2294 & ~n5161 ;
  assign n5163 = n1368 & ~n5162 ;
  assign n5164 = n1372 & ~n5163 ;
  assign n5165 = n1376 & ~n5164 ;
  assign n5166 = n1380 & ~n5165 ;
  assign n5167 = n1384 & ~n5166 ;
  assign n5168 = n1388 & ~n5167 ;
  assign n5169 = n1392 & ~n5168 ;
  assign n5170 = n1396 & ~n5169 ;
  assign n5171 = n1400 & ~n5170 ;
  assign n5172 = n1404 & ~n5171 ;
  assign n5173 = n1408 & ~n5172 ;
  assign n5174 = n1412 & ~n5173 ;
  assign n5175 = n1416 & ~n5174 ;
  assign n5176 = n1420 & ~n5175 ;
  assign n5177 = n1424 & ~n5176 ;
  assign n5178 = n1428 & ~n5177 ;
  assign n5179 = n1432 & ~n5178 ;
  assign n5180 = n1436 & ~n5179 ;
  assign n5181 = n515 & n5150 ;
  assign n5182 = ~n1438 & n5181 ;
  assign n5183 = ~n5180 & n5182 ;
  assign n5184 = ~n5151 & ~n5183 ;
  assign n5185 = \req[96]  & ~n902 ;
  assign n5186 = ~n898 & n5185 ;
  assign n5187 = ~\priority[98]  & ~n893 ;
  assign n5188 = n543 & ~n5187 ;
  assign n5189 = n1796 & ~n5188 ;
  assign n5190 = n1801 & ~n5189 ;
  assign n5191 = n1805 & ~n5190 ;
  assign n5192 = n4558 & ~n5191 ;
  assign n5193 = n1813 & ~n5192 ;
  assign n5194 = n1817 & ~n5193 ;
  assign n5195 = n1821 & ~n5194 ;
  assign n5196 = n2330 & ~n5195 ;
  assign n5197 = n2333 & ~n5196 ;
  assign n5198 = n1488 & ~n5197 ;
  assign n5199 = n1492 & ~n5198 ;
  assign n5200 = n1496 & ~n5199 ;
  assign n5201 = n1500 & ~n5200 ;
  assign n5202 = n1504 & ~n5201 ;
  assign n5203 = n2229 & ~n5202 ;
  assign n5204 = n1512 & ~n5203 ;
  assign n5205 = n1516 & ~n5204 ;
  assign n5206 = n1520 & ~n5205 ;
  assign n5207 = n1524 & ~n5206 ;
  assign n5208 = n1528 & ~n5207 ;
  assign n5209 = n1532 & ~n5208 ;
  assign n5210 = n1536 & ~n5209 ;
  assign n5211 = n1540 & ~n5210 ;
  assign n5212 = n1544 & ~n5211 ;
  assign n5213 = n1548 & ~n5212 ;
  assign n5214 = n1552 & ~n5213 ;
  assign n5215 = n1556 & ~n5214 ;
  assign n5216 = n882 & n5185 ;
  assign n5217 = ~n1558 & n5216 ;
  assign n5218 = ~n5215 & n5217 ;
  assign n5219 = ~n5186 & ~n5218 ;
  assign n5220 = \req[97]  & ~n1268 ;
  assign n5221 = ~n1264 & n5220 ;
  assign n5222 = ~\priority[99]  & ~n1259 ;
  assign n5223 = n910 & ~n5222 ;
  assign n5224 = n1912 & ~n5223 ;
  assign n5225 = n1917 & ~n5224 ;
  assign n5226 = n1921 & ~n5225 ;
  assign n5227 = n1925 & ~n5226 ;
  assign n5228 = n1929 & ~n5227 ;
  assign n5229 = n1933 & ~n5228 ;
  assign n5230 = n1937 & ~n5229 ;
  assign n5231 = n2369 & ~n5230 ;
  assign n5232 = n2372 & ~n5231 ;
  assign n5233 = n1605 & ~n5232 ;
  assign n5234 = n1609 & ~n5233 ;
  assign n5235 = n1613 & ~n5234 ;
  assign n5236 = n1617 & ~n5235 ;
  assign n5237 = n1621 & ~n5236 ;
  assign n5238 = n1625 & ~n5237 ;
  assign n5239 = n1629 & ~n5238 ;
  assign n5240 = n1633 & ~n5239 ;
  assign n5241 = n1637 & ~n5240 ;
  assign n5242 = n1641 & ~n5241 ;
  assign n5243 = n1645 & ~n5242 ;
  assign n5244 = n1649 & ~n5243 ;
  assign n5245 = n4614 & ~n5244 ;
  assign n5246 = n1657 & ~n5245 ;
  assign n5247 = n4930 & ~n5246 ;
  assign n5248 = n1665 & ~n5247 ;
  assign n5249 = n1669 & ~n5248 ;
  assign n5250 = n1673 & ~n5249 ;
  assign n5251 = n1248 & n5220 ;
  assign n5252 = ~n1675 & n5251 ;
  assign n5253 = ~n5250 & n5252 ;
  assign n5254 = ~n5221 & ~n5253 ;
  assign n5255 = \req[98]  & ~n542 ;
  assign n5256 = ~n528 & n5255 ;
  assign n5257 = ~\priority[100]  & ~n548 ;
  assign n5258 = n1276 & ~n5257 ;
  assign n5259 = n2028 & ~n5258 ;
  assign n5260 = n2033 & ~n5259 ;
  assign n5261 = n2037 & ~n5260 ;
  assign n5262 = n2041 & ~n5261 ;
  assign n5263 = n2045 & ~n5262 ;
  assign n5264 = n2049 & ~n5263 ;
  assign n5265 = n2053 & ~n5264 ;
  assign n5266 = n2408 & ~n5265 ;
  assign n5267 = n2411 & ~n5266 ;
  assign n5268 = n1721 & ~n5267 ;
  assign n5269 = n1725 & ~n5268 ;
  assign n5270 = n1729 & ~n5269 ;
  assign n5271 = n1733 & ~n5270 ;
  assign n5272 = n1737 & ~n5271 ;
  assign n5273 = n1741 & ~n5272 ;
  assign n5274 = n1745 & ~n5273 ;
  assign n5275 = n1749 & ~n5274 ;
  assign n5276 = n1753 & ~n5275 ;
  assign n5277 = n1757 & ~n5276 ;
  assign n5278 = n1761 & ~n5277 ;
  assign n5279 = n1765 & ~n5278 ;
  assign n5280 = n1769 & ~n5279 ;
  assign n5281 = n1773 & ~n5280 ;
  assign n5282 = n1777 & ~n5281 ;
  assign n5283 = n1781 & ~n5282 ;
  assign n5284 = n1785 & ~n5283 ;
  assign n5285 = n1789 & ~n5284 ;
  assign n5286 = n537 & n5255 ;
  assign n5287 = ~n1791 & n5286 ;
  assign n5288 = ~n5285 & n5287 ;
  assign n5289 = ~n5256 & ~n5288 ;
  assign n5290 = \req[99]  & ~n909 ;
  assign n5291 = ~n895 & n5290 ;
  assign n5292 = ~\priority[101]  & ~n915 ;
  assign n5293 = n540 & ~n5292 ;
  assign n5294 = n558 & ~n5293 ;
  assign n5295 = n572 & ~n5294 ;
  assign n5296 = n585 & ~n5295 ;
  assign n5297 = n598 & ~n5296 ;
  assign n5298 = n611 & ~n5297 ;
  assign n5299 = n2090 & ~n5298 ;
  assign n5300 = n2094 & ~n5299 ;
  assign n5301 = n2447 & ~n5300 ;
  assign n5302 = n2450 & ~n5301 ;
  assign n5303 = n1837 & ~n5302 ;
  assign n5304 = n1841 & ~n5303 ;
  assign n5305 = n1845 & ~n5304 ;
  assign n5306 = n1849 & ~n5305 ;
  assign n5307 = n3720 & ~n5306 ;
  assign n5308 = n1857 & ~n5307 ;
  assign n5309 = n1861 & ~n5308 ;
  assign n5310 = n1865 & ~n5309 ;
  assign n5311 = n1869 & ~n5310 ;
  assign n5312 = n1873 & ~n5311 ;
  assign n5313 = n1877 & ~n5312 ;
  assign n5314 = n3627 & ~n5313 ;
  assign n5315 = n1885 & ~n5314 ;
  assign n5316 = n1889 & ~n5315 ;
  assign n5317 = n1893 & ~n5316 ;
  assign n5318 = n1897 & ~n5317 ;
  assign n5319 = n1901 & ~n5318 ;
  assign n5320 = n1905 & ~n5319 ;
  assign n5321 = n904 & n5290 ;
  assign n5322 = ~n1907 & n5321 ;
  assign n5323 = ~n5320 & n5322 ;
  assign n5324 = ~n5291 & ~n5323 ;
  assign n5325 = \req[100]  & ~n1275 ;
  assign n5326 = ~n1261 & n5325 ;
  assign n5327 = ~\priority[102]  & ~n1281 ;
  assign n5328 = n907 & ~n5327 ;
  assign n5329 = n925 & ~n5328 ;
  assign n5330 = n939 & ~n5329 ;
  assign n5331 = n952 & ~n5330 ;
  assign n5332 = n965 & ~n5331 ;
  assign n5333 = n978 & ~n5332 ;
  assign n5334 = n2132 & ~n5333 ;
  assign n5335 = n2136 & ~n5334 ;
  assign n5336 = n2487 & ~n5335 ;
  assign n5337 = n2490 & ~n5336 ;
  assign n5338 = n1953 & ~n5337 ;
  assign n5339 = n1957 & ~n5338 ;
  assign n5340 = n1961 & ~n5339 ;
  assign n5341 = n1965 & ~n5340 ;
  assign n5342 = n1969 & ~n5341 ;
  assign n5343 = n1973 & ~n5342 ;
  assign n5344 = n2713 & ~n5343 ;
  assign n5345 = n1981 & ~n5344 ;
  assign n5346 = n1985 & ~n5345 ;
  assign n5347 = n1989 & ~n5346 ;
  assign n5348 = n1993 & ~n5347 ;
  assign n5349 = n1997 & ~n5348 ;
  assign n5350 = n2001 & ~n5349 ;
  assign n5351 = n2005 & ~n5350 ;
  assign n5352 = n2009 & ~n5351 ;
  assign n5353 = n2013 & ~n5352 ;
  assign n5354 = n2017 & ~n5353 ;
  assign n5355 = n2021 & ~n5354 ;
  assign n5356 = n1270 & n5325 ;
  assign n5357 = ~n2023 & n5356 ;
  assign n5358 = ~n5355 & n5357 ;
  assign n5359 = ~n5326 & ~n5358 ;
  assign n5360 = \req[101]  & ~n539 ;
  assign n5361 = ~n550 & n5360 ;
  assign n5362 = ~\priority[103]  & ~n555 ;
  assign n5363 = n1273 & ~n5362 ;
  assign n5364 = n1291 & ~n5363 ;
  assign n5365 = n1305 & ~n5364 ;
  assign n5366 = n3148 & ~n5365 ;
  assign n5367 = n1331 & ~n5366 ;
  assign n5368 = n1344 & ~n5367 ;
  assign n5369 = n2173 & ~n5368 ;
  assign n5370 = n2176 & ~n5369 ;
  assign n5371 = n286 & ~n5370 ;
  assign n5372 = n294 & n297 ;
  assign n5373 = ~n291 & n5372 ;
  assign n5374 = ~n5371 & n5373 ;
  assign n5375 = n312 & ~n5374 ;
  assign n5376 = n325 & ~n5375 ;
  assign n5377 = n338 & ~n5376 ;
  assign n5378 = n346 & n349 ;
  assign n5379 = ~n343 & n5378 ;
  assign n5380 = ~n5377 & n5379 ;
  assign n5381 = n364 & ~n5380 ;
  assign n5382 = n377 & ~n5381 ;
  assign n5383 = n390 & ~n5382 ;
  assign n5384 = n5064 & ~n5383 ;
  assign n5385 = n416 & ~n5384 ;
  assign n5386 = n4115 & ~n5385 ;
  assign n5387 = n442 & ~n5386 ;
  assign n5388 = n455 & ~n5387 ;
  assign n5389 = n468 & ~n5388 ;
  assign n5390 = n481 & ~n5389 ;
  assign n5391 = n494 & ~n5390 ;
  assign n5392 = n507 & ~n5391 ;
  assign n5393 = n520 & ~n5392 ;
  assign n5394 = n533 & ~n5393 ;
  assign n5395 = n544 & n5360 ;
  assign n5396 = ~n538 & n5395 ;
  assign n5397 = ~n5394 & n5396 ;
  assign n5398 = ~n5361 & ~n5397 ;
  assign n5399 = \req[102]  & ~n906 ;
  assign n5400 = ~n917 & n5399 ;
  assign n5401 = ~\priority[104]  & ~n922 ;
  assign n5402 = n562 & ~n5401 ;
  assign n5403 = n1451 & ~n5402 ;
  assign n5404 = n1456 & ~n5403 ;
  assign n5405 = n3817 & ~n5404 ;
  assign n5406 = n1464 & ~n5405 ;
  assign n5407 = n1468 & ~n5406 ;
  assign n5408 = n2212 & ~n5407 ;
  assign n5409 = n4453 & ~n5408 ;
  assign n5410 = ~n645 & n652 ;
  assign n5411 = ~n5409 & n5410 ;
  assign n5412 = n666 & ~n5411 ;
  assign n5413 = n679 & ~n5412 ;
  assign n5414 = n3826 & ~n5413 ;
  assign n5415 = n4459 & ~n5414 ;
  assign n5416 = n718 & ~n5415 ;
  assign n5417 = n731 & ~n5416 ;
  assign n5418 = n4464 & ~n5417 ;
  assign n5419 = n2465 & ~n5418 ;
  assign n5420 = n770 & ~n5419 ;
  assign n5421 = n3099 & ~n5420 ;
  assign n5422 = n796 & ~n5421 ;
  assign n5423 = n809 & ~n5422 ;
  assign n5424 = n2117 & ~n5423 ;
  assign n5425 = n835 & ~n5424 ;
  assign n5426 = n848 & ~n5425 ;
  assign n5427 = n5107 & ~n5426 ;
  assign n5428 = n874 & ~n5427 ;
  assign n5429 = n887 & ~n5428 ;
  assign n5430 = n900 & ~n5429 ;
  assign n5431 = n911 & n5399 ;
  assign n5432 = ~n905 & n5431 ;
  assign n5433 = ~n5430 & n5432 ;
  assign n5434 = ~n5400 & ~n5433 ;
  assign n5435 = \req[103]  & ~n1272 ;
  assign n5436 = ~n1283 & n5435 ;
  assign n5437 = ~\priority[105]  & ~n1288 ;
  assign n5438 = n929 & ~n5437 ;
  assign n5439 = n1571 & ~n5438 ;
  assign n5440 = ~n937 & n943 ;
  assign n5441 = n1575 & ~n5440 ;
  assign n5442 = ~n5439 & n5441 ;
  assign n5443 = n1580 & ~n5442 ;
  assign n5444 = n1584 & ~n5443 ;
  assign n5445 = n1588 & ~n5444 ;
  assign n5446 = n2252 & ~n5445 ;
  assign n5447 = n2255 & ~n5446 ;
  assign n5448 = n1019 & ~n5447 ;
  assign n5449 = n1032 & ~n5448 ;
  assign n5450 = n3861 & ~n5449 ;
  assign n5451 = n1058 & ~n5450 ;
  assign n5452 = n1071 & ~n5451 ;
  assign n5453 = n1084 & ~n5452 ;
  assign n5454 = n1097 & ~n5453 ;
  assign n5455 = n1110 & ~n5454 ;
  assign n5456 = n1123 & ~n5455 ;
  assign n5457 = n1136 & ~n5456 ;
  assign n5458 = n5137 & ~n5457 ;
  assign n5459 = n1162 & ~n5458 ;
  assign n5460 = n1175 & ~n5459 ;
  assign n5461 = n1188 & ~n5460 ;
  assign n5462 = n1201 & ~n5461 ;
  assign n5463 = n1214 & ~n5462 ;
  assign n5464 = n1227 & ~n5463 ;
  assign n5465 = n1240 & ~n5464 ;
  assign n5466 = n1253 & ~n5465 ;
  assign n5467 = n4409 & ~n5466 ;
  assign n5468 = n1277 & n5435 ;
  assign n5469 = ~n1271 & n5468 ;
  assign n5470 = ~n5467 & n5469 ;
  assign n5471 = ~n5436 & ~n5470 ;
  assign n5472 = \req[104]  & ~n561 ;
  assign n5473 = ~n557 & n5472 ;
  assign n5474 = ~\priority[106]  & ~n552 ;
  assign n5475 = n1295 & ~n5474 ;
  assign n5476 = n1688 & ~n5475 ;
  assign n5477 = n1693 & ~n5476 ;
  assign n5478 = n1697 & ~n5477 ;
  assign n5479 = n1701 & ~n5478 ;
  assign n5480 = n3570 & ~n5479 ;
  assign n5481 = n2291 & ~n5480 ;
  assign n5482 = n2294 & ~n5481 ;
  assign n5483 = n1368 & ~n5482 ;
  assign n5484 = n1372 & ~n5483 ;
  assign n5485 = n1376 & ~n5484 ;
  assign n5486 = n1380 & ~n5485 ;
  assign n5487 = n1384 & ~n5486 ;
  assign n5488 = n1388 & ~n5487 ;
  assign n5489 = n1392 & ~n5488 ;
  assign n5490 = n1396 & ~n5489 ;
  assign n5491 = ~n1398 & n1399 ;
  assign n5492 = ~n5490 & n5491 ;
  assign n5493 = n1404 & ~n5492 ;
  assign n5494 = n1408 & ~n5493 ;
  assign n5495 = n1412 & ~n5494 ;
  assign n5496 = n1416 & ~n5495 ;
  assign n5497 = n1420 & ~n5496 ;
  assign n5498 = n1424 & ~n5497 ;
  assign n5499 = n1428 & ~n5498 ;
  assign n5500 = n1432 & ~n5499 ;
  assign n5501 = ~n1434 & n1435 ;
  assign n5502 = ~n5500 & n5501 ;
  assign n5503 = n1440 & ~n5502 ;
  assign n5504 = n3811 & ~n5503 ;
  assign n5505 = n541 & n5472 ;
  assign n5506 = ~n1446 & n5505 ;
  assign n5507 = ~n5504 & n5506 ;
  assign n5508 = ~n5473 & ~n5507 ;
  assign n5509 = \req[105]  & ~n928 ;
  assign n5510 = ~n924 & n5509 ;
  assign n5511 = ~\priority[107]  & ~n919 ;
  assign n5512 = n569 & ~n5511 ;
  assign n5513 = n1804 & ~n5512 ;
  assign n5514 = n4558 & ~n5513 ;
  assign n5515 = n1813 & ~n5514 ;
  assign n5516 = n1817 & ~n5515 ;
  assign n5517 = n1821 & ~n5516 ;
  assign n5518 = n2330 & ~n5517 ;
  assign n5519 = n2333 & ~n5518 ;
  assign n5520 = n1488 & ~n5519 ;
  assign n5521 = n1492 & ~n5520 ;
  assign n5522 = n1496 & ~n5521 ;
  assign n5523 = n1500 & ~n5522 ;
  assign n5524 = n1504 & ~n5523 ;
  assign n5525 = n2229 & ~n5524 ;
  assign n5526 = n1512 & ~n5525 ;
  assign n5527 = n1516 & ~n5526 ;
  assign n5528 = n1520 & ~n5527 ;
  assign n5529 = n1524 & ~n5528 ;
  assign n5530 = n1528 & ~n5529 ;
  assign n5531 = n1532 & ~n5530 ;
  assign n5532 = n1536 & ~n5531 ;
  assign n5533 = n1540 & ~n5532 ;
  assign n5534 = n1544 & ~n5533 ;
  assign n5535 = n1548 & ~n5534 ;
  assign n5536 = n1552 & ~n5535 ;
  assign n5537 = n1556 & ~n5536 ;
  assign n5538 = ~n1558 & n1559 ;
  assign n5539 = ~n5537 & n5538 ;
  assign n5540 = n1564 & ~n5539 ;
  assign n5541 = n908 & n5509 ;
  assign n5542 = ~n1566 & n5541 ;
  assign n5543 = ~n5540 & n5542 ;
  assign n5544 = ~n5510 & ~n5543 ;
  assign n5545 = \req[106]  & ~n1294 ;
  assign n5546 = ~n1290 & n5545 ;
  assign n5547 = ~\priority[108]  & ~n1285 ;
  assign n5548 = n936 & ~n5547 ;
  assign n5549 = n1920 & ~n5548 ;
  assign n5550 = n1925 & ~n5549 ;
  assign n5551 = n1929 & ~n5550 ;
  assign n5552 = n1933 & ~n5551 ;
  assign n5553 = n1937 & ~n5552 ;
  assign n5554 = n2369 & ~n5553 ;
  assign n5555 = n2372 & ~n5554 ;
  assign n5556 = n1605 & ~n5555 ;
  assign n5557 = n1609 & ~n5556 ;
  assign n5558 = n1613 & ~n5557 ;
  assign n5559 = n1617 & ~n5558 ;
  assign n5560 = n1621 & ~n5559 ;
  assign n5561 = n1625 & ~n5560 ;
  assign n5562 = n1629 & ~n5561 ;
  assign n5563 = n1633 & ~n5562 ;
  assign n5564 = ~n1635 & n1636 ;
  assign n5565 = ~n5563 & n5564 ;
  assign n5566 = n1641 & ~n5565 ;
  assign n5567 = n1645 & ~n5566 ;
  assign n5568 = n1649 & ~n5567 ;
  assign n5569 = n4614 & ~n5568 ;
  assign n5570 = n1657 & ~n5569 ;
  assign n5571 = n4930 & ~n5570 ;
  assign n5572 = n1665 & ~n5571 ;
  assign n5573 = n1669 & ~n5572 ;
  assign n5574 = n1673 & ~n5573 ;
  assign n5575 = n1677 & ~n5574 ;
  assign n5576 = n1681 & ~n5575 ;
  assign n5577 = n1274 & n5545 ;
  assign n5578 = ~n1683 & n5577 ;
  assign n5579 = ~n5576 & n5578 ;
  assign n5580 = ~n5546 & ~n5579 ;
  assign n5581 = \req[107]  & ~n568 ;
  assign n5582 = ~n554 & n5581 ;
  assign n5583 = ~\priority[109]  & ~n574 ;
  assign n5584 = n1302 & ~n5583 ;
  assign n5585 = n2036 & ~n5584 ;
  assign n5586 = n2041 & ~n5585 ;
  assign n5587 = n2045 & ~n5586 ;
  assign n5588 = n2049 & ~n5587 ;
  assign n5589 = n2053 & ~n5588 ;
  assign n5590 = n2408 & ~n5589 ;
  assign n5591 = n2411 & ~n5590 ;
  assign n5592 = n1721 & ~n5591 ;
  assign n5593 = n1725 & ~n5592 ;
  assign n5594 = n1729 & ~n5593 ;
  assign n5595 = n1733 & ~n5594 ;
  assign n5596 = n1737 & ~n5595 ;
  assign n5597 = n1741 & ~n5596 ;
  assign n5598 = n1745 & ~n5597 ;
  assign n5599 = n1749 & ~n5598 ;
  assign n5600 = n1753 & ~n5599 ;
  assign n5601 = n1757 & ~n5600 ;
  assign n5602 = n1761 & ~n5601 ;
  assign n5603 = n1765 & ~n5602 ;
  assign n5604 = n1769 & ~n5603 ;
  assign n5605 = n1773 & ~n5604 ;
  assign n5606 = n1777 & ~n5605 ;
  assign n5607 = n1781 & ~n5606 ;
  assign n5608 = n1785 & ~n5607 ;
  assign n5609 = n1789 & ~n5608 ;
  assign n5610 = n3920 & ~n5609 ;
  assign n5611 = n1797 & ~n5610 ;
  assign n5612 = n563 & n5581 ;
  assign n5613 = ~n1799 & n5612 ;
  assign n5614 = ~n5611 & n5613 ;
  assign n5615 = ~n5582 & ~n5614 ;
  assign n5616 = \req[108]  & ~n935 ;
  assign n5617 = ~n921 & n5616 ;
  assign n5618 = ~\priority[110]  & ~n941 ;
  assign n5619 = n566 & ~n5618 ;
  assign n5620 = n584 & ~n5619 ;
  assign n5621 = n598 & ~n5620 ;
  assign n5622 = n611 & ~n5621 ;
  assign n5623 = n2090 & ~n5622 ;
  assign n5624 = n2094 & ~n5623 ;
  assign n5625 = n2447 & ~n5624 ;
  assign n5626 = n2450 & ~n5625 ;
  assign n5627 = n1837 & ~n5626 ;
  assign n5628 = n1841 & ~n5627 ;
  assign n5629 = n1845 & ~n5628 ;
  assign n5630 = n1849 & ~n5629 ;
  assign n5631 = n3720 & ~n5630 ;
  assign n5632 = n1857 & ~n5631 ;
  assign n5633 = n1861 & ~n5632 ;
  assign n5634 = n1865 & ~n5633 ;
  assign n5635 = n1869 & ~n5634 ;
  assign n5636 = n1873 & ~n5635 ;
  assign n5637 = n1877 & ~n5636 ;
  assign n5638 = n3627 & ~n5637 ;
  assign n5639 = n1885 & ~n5638 ;
  assign n5640 = n1889 & ~n5639 ;
  assign n5641 = n1893 & ~n5640 ;
  assign n5642 = n1897 & ~n5641 ;
  assign n5643 = n1901 & ~n5642 ;
  assign n5644 = n1905 & ~n5643 ;
  assign n5645 = n1909 & ~n5644 ;
  assign n5646 = n4592 & ~n5645 ;
  assign n5647 = ~n908 & n924 ;
  assign n5648 = n930 & n5616 ;
  assign n5649 = ~n5647 & n5648 ;
  assign n5650 = ~n5646 & n5649 ;
  assign n5651 = ~n5617 & ~n5650 ;
  assign n5652 = \req[109]  & ~n1301 ;
  assign n5653 = ~n1287 & n5652 ;
  assign n5654 = ~\priority[111]  & ~n1307 ;
  assign n5655 = n933 & ~n5654 ;
  assign n5656 = n951 & ~n5655 ;
  assign n5657 = n965 & ~n5656 ;
  assign n5658 = n978 & ~n5657 ;
  assign n5659 = n2132 & ~n5658 ;
  assign n5660 = n2136 & ~n5659 ;
  assign n5661 = n2487 & ~n5660 ;
  assign n5662 = n2490 & ~n5661 ;
  assign n5663 = n1953 & ~n5662 ;
  assign n5664 = n1957 & ~n5663 ;
  assign n5665 = n1961 & ~n5664 ;
  assign n5666 = n1965 & ~n5665 ;
  assign n5667 = n1969 & ~n5666 ;
  assign n5668 = n1973 & ~n5667 ;
  assign n5669 = n2713 & ~n5668 ;
  assign n5670 = n1981 & ~n5669 ;
  assign n5671 = n1985 & ~n5670 ;
  assign n5672 = n1989 & ~n5671 ;
  assign n5673 = n1993 & ~n5672 ;
  assign n5674 = n1997 & ~n5673 ;
  assign n5675 = n2001 & ~n5674 ;
  assign n5676 = n2005 & ~n5675 ;
  assign n5677 = n2009 & ~n5676 ;
  assign n5678 = n2013 & ~n5677 ;
  assign n5679 = n2017 & ~n5678 ;
  assign n5680 = n2021 & ~n5679 ;
  assign n5681 = n2025 & ~n5680 ;
  assign n5682 = n3671 & ~n5681 ;
  assign n5683 = n1296 & n5652 ;
  assign n5684 = ~n2031 & n5683 ;
  assign n5685 = ~n5682 & n5684 ;
  assign n5686 = ~n5653 & ~n5685 ;
  assign n5687 = \req[110]  & ~n565 ;
  assign n5688 = ~n576 & n5687 ;
  assign n5689 = ~\priority[112]  & ~n581 ;
  assign n5690 = n1299 & ~n5689 ;
  assign n5691 = n1317 & ~n5690 ;
  assign n5692 = n1331 & ~n5691 ;
  assign n5693 = n1344 & ~n5692 ;
  assign n5694 = n2173 & ~n5693 ;
  assign n5695 = n2176 & ~n5694 ;
  assign n5696 = n286 & ~n5695 ;
  assign n5697 = n5373 & ~n5696 ;
  assign n5698 = n312 & ~n5697 ;
  assign n5699 = n325 & ~n5698 ;
  assign n5700 = n338 & ~n5699 ;
  assign n5701 = n5379 & ~n5700 ;
  assign n5702 = n364 & ~n5701 ;
  assign n5703 = n377 & ~n5702 ;
  assign n5704 = n390 & ~n5703 ;
  assign n5705 = n398 & n401 ;
  assign n5706 = ~n395 & n5705 ;
  assign n5707 = ~n5704 & n5706 ;
  assign n5708 = n416 & ~n5707 ;
  assign n5709 = n4115 & ~n5708 ;
  assign n5710 = n442 & ~n5709 ;
  assign n5711 = n455 & ~n5710 ;
  assign n5712 = n468 & ~n5711 ;
  assign n5713 = ~n473 & n480 ;
  assign n5714 = ~n5712 & n5713 ;
  assign n5715 = n494 & ~n5714 ;
  assign n5716 = n507 & ~n5715 ;
  assign n5717 = n520 & ~n5716 ;
  assign n5718 = n533 & ~n5717 ;
  assign n5719 = n546 & ~n5718 ;
  assign n5720 = n559 & ~n5719 ;
  assign n5721 = n570 & n5687 ;
  assign n5722 = ~n564 & n5721 ;
  assign n5723 = ~n5720 & n5722 ;
  assign n5724 = ~n5688 & ~n5723 ;
  assign n5725 = \req[111]  & ~n932 ;
  assign n5726 = ~n943 & n5725 ;
  assign n5727 = ~\priority[113]  & ~n948 ;
  assign n5728 = n588 & ~n5727 ;
  assign n5729 = n3816 & ~n5728 ;
  assign n5730 = n1464 & ~n5729 ;
  assign n5731 = n1468 & ~n5730 ;
  assign n5732 = n2212 & ~n5731 ;
  assign n5733 = n4453 & ~n5732 ;
  assign n5734 = n5410 & ~n5733 ;
  assign n5735 = n666 & ~n5734 ;
  assign n5736 = n679 & ~n5735 ;
  assign n5737 = n3826 & ~n5736 ;
  assign n5738 = n4459 & ~n5737 ;
  assign n5739 = n718 & ~n5738 ;
  assign n5740 = n731 & ~n5739 ;
  assign n5741 = n4464 & ~n5740 ;
  assign n5742 = n2465 & ~n5741 ;
  assign n5743 = n770 & ~n5742 ;
  assign n5744 = n3099 & ~n5743 ;
  assign n5745 = n796 & ~n5744 ;
  assign n5746 = n809 & ~n5745 ;
  assign n5747 = n2117 & ~n5746 ;
  assign n5748 = n835 & ~n5747 ;
  assign n5749 = n848 & ~n5748 ;
  assign n5750 = n5107 & ~n5749 ;
  assign n5751 = n874 & ~n5750 ;
  assign n5752 = n887 & ~n5751 ;
  assign n5753 = n900 & ~n5752 ;
  assign n5754 = n913 & ~n5753 ;
  assign n5755 = n926 & ~n5754 ;
  assign n5756 = n937 & n5725 ;
  assign n5757 = ~n931 & n5756 ;
  assign n5758 = ~n5755 & n5757 ;
  assign n5759 = ~n5726 & ~n5758 ;
  assign n5760 = \req[112]  & ~n1298 ;
  assign n5761 = ~n1309 & n5760 ;
  assign n5762 = ~\priority[114]  & ~n1314 ;
  assign n5763 = n955 & ~n5762 ;
  assign n5764 = n1579 & ~n5763 ;
  assign n5765 = n1584 & ~n5764 ;
  assign n5766 = n1588 & ~n5765 ;
  assign n5767 = n2252 & ~n5766 ;
  assign n5768 = n2255 & ~n5767 ;
  assign n5769 = n1019 & ~n5768 ;
  assign n5770 = n1032 & ~n5769 ;
  assign n5771 = n3861 & ~n5770 ;
  assign n5772 = n1058 & ~n5771 ;
  assign n5773 = n1071 & ~n5772 ;
  assign n5774 = n1084 & ~n5773 ;
  assign n5775 = n1097 & ~n5774 ;
  assign n5776 = n1110 & ~n5775 ;
  assign n5777 = n1123 & ~n5776 ;
  assign n5778 = n1136 & ~n5777 ;
  assign n5779 = n5137 & ~n5778 ;
  assign n5780 = n1162 & ~n5779 ;
  assign n5781 = n1175 & ~n5780 ;
  assign n5782 = n1188 & ~n5781 ;
  assign n5783 = n1201 & ~n5782 ;
  assign n5784 = n1214 & ~n5783 ;
  assign n5785 = n1227 & ~n5784 ;
  assign n5786 = n1240 & ~n5785 ;
  assign n5787 = n1253 & ~n5786 ;
  assign n5788 = n4409 & ~n5787 ;
  assign n5789 = n1279 & ~n5788 ;
  assign n5790 = n1292 & ~n5789 ;
  assign n5791 = n1303 & n5760 ;
  assign n5792 = ~n1297 & n5791 ;
  assign n5793 = ~n5790 & n5792 ;
  assign n5794 = ~n5761 & ~n5793 ;
  assign n5795 = \req[113]  & ~n587 ;
  assign n5796 = ~n583 & n5795 ;
  assign n5797 = ~\priority[115]  & ~n578 ;
  assign n5798 = n1321 & ~n5797 ;
  assign n5799 = n1696 & ~n5798 ;
  assign n5800 = n1701 & ~n5799 ;
  assign n5801 = n3570 & ~n5800 ;
  assign n5802 = n2291 & ~n5801 ;
  assign n5803 = n2294 & ~n5802 ;
  assign n5804 = n1368 & ~n5803 ;
  assign n5805 = n1372 & ~n5804 ;
  assign n5806 = n1376 & ~n5805 ;
  assign n5807 = n1380 & ~n5806 ;
  assign n5808 = n1384 & ~n5807 ;
  assign n5809 = n1388 & ~n5808 ;
  assign n5810 = n1392 & ~n5809 ;
  assign n5811 = n1396 & ~n5810 ;
  assign n5812 = n5491 & ~n5811 ;
  assign n5813 = n1404 & ~n5812 ;
  assign n5814 = n1408 & ~n5813 ;
  assign n5815 = n1412 & ~n5814 ;
  assign n5816 = n1416 & ~n5815 ;
  assign n5817 = n1420 & ~n5816 ;
  assign n5818 = n1424 & ~n5817 ;
  assign n5819 = n1428 & ~n5818 ;
  assign n5820 = n1432 & ~n5819 ;
  assign n5821 = n5501 & ~n5820 ;
  assign n5822 = n1440 & ~n5821 ;
  assign n5823 = n3811 & ~n5822 ;
  assign n5824 = n1448 & ~n5823 ;
  assign n5825 = n1452 & ~n5824 ;
  assign n5826 = n567 & n5795 ;
  assign n5827 = ~n1454 & n5826 ;
  assign n5828 = ~n5825 & n5827 ;
  assign n5829 = ~n5796 & ~n5828 ;
  assign n5830 = \req[114]  & ~n954 ;
  assign n5831 = ~n950 & n5830 ;
  assign n5832 = ~\priority[116]  & ~n945 ;
  assign n5833 = n595 & ~n5832 ;
  assign n5834 = n1812 & ~n5833 ;
  assign n5835 = n1817 & ~n5834 ;
  assign n5836 = n1821 & ~n5835 ;
  assign n5837 = n2330 & ~n5836 ;
  assign n5838 = n2333 & ~n5837 ;
  assign n5839 = n1488 & ~n5838 ;
  assign n5840 = n1492 & ~n5839 ;
  assign n5841 = n1496 & ~n5840 ;
  assign n5842 = n1500 & ~n5841 ;
  assign n5843 = n1504 & ~n5842 ;
  assign n5844 = n2229 & ~n5843 ;
  assign n5845 = n1512 & ~n5844 ;
  assign n5846 = n1516 & ~n5845 ;
  assign n5847 = n1520 & ~n5846 ;
  assign n5848 = n1524 & ~n5847 ;
  assign n5849 = n1528 & ~n5848 ;
  assign n5850 = n1532 & ~n5849 ;
  assign n5851 = n1536 & ~n5850 ;
  assign n5852 = n1540 & ~n5851 ;
  assign n5853 = n1544 & ~n5852 ;
  assign n5854 = n1548 & ~n5853 ;
  assign n5855 = n1552 & ~n5854 ;
  assign n5856 = n1556 & ~n5855 ;
  assign n5857 = n5538 & ~n5856 ;
  assign n5858 = n1564 & ~n5857 ;
  assign n5859 = n1568 & ~n5858 ;
  assign n5860 = ~n1570 & n1571 ;
  assign n5861 = ~n5859 & n5860 ;
  assign n5862 = n934 & n5830 ;
  assign n5863 = ~n5440 & n5862 ;
  assign n5864 = ~n5861 & n5863 ;
  assign n5865 = ~n5831 & ~n5864 ;
  assign n5866 = \req[115]  & ~n1320 ;
  assign n5867 = ~n1316 & n5866 ;
  assign n5868 = ~\priority[117]  & ~n1311 ;
  assign n5869 = n962 & ~n5868 ;
  assign n5870 = n1928 & ~n5869 ;
  assign n5871 = n1933 & ~n5870 ;
  assign n5872 = n1937 & ~n5871 ;
  assign n5873 = n2369 & ~n5872 ;
  assign n5874 = n2372 & ~n5873 ;
  assign n5875 = n1605 & ~n5874 ;
  assign n5876 = n1609 & ~n5875 ;
  assign n5877 = n1613 & ~n5876 ;
  assign n5878 = n1617 & ~n5877 ;
  assign n5879 = n1621 & ~n5878 ;
  assign n5880 = n1625 & ~n5879 ;
  assign n5881 = n1629 & ~n5880 ;
  assign n5882 = n1633 & ~n5881 ;
  assign n5883 = n5564 & ~n5882 ;
  assign n5884 = n1641 & ~n5883 ;
  assign n5885 = n1645 & ~n5884 ;
  assign n5886 = n1649 & ~n5885 ;
  assign n5887 = n4614 & ~n5886 ;
  assign n5888 = n1657 & ~n5887 ;
  assign n5889 = n4930 & ~n5888 ;
  assign n5890 = n1665 & ~n5889 ;
  assign n5891 = n1669 & ~n5890 ;
  assign n5892 = n1673 & ~n5891 ;
  assign n5893 = n1677 & ~n5892 ;
  assign n5894 = n1681 & ~n5893 ;
  assign n5895 = n1685 & ~n5894 ;
  assign n5896 = n1689 & ~n5895 ;
  assign n5897 = n1300 & n5866 ;
  assign n5898 = ~n1691 & n5897 ;
  assign n5899 = ~n5896 & n5898 ;
  assign n5900 = ~n5867 & ~n5899 ;
  assign n5901 = \req[116]  & ~n594 ;
  assign n5902 = ~n580 & n5901 ;
  assign n5903 = ~\priority[118]  & ~n600 ;
  assign n5904 = n1328 & ~n5903 ;
  assign n5905 = n2044 & ~n5904 ;
  assign n5906 = n2049 & ~n5905 ;
  assign n5907 = n2053 & ~n5906 ;
  assign n5908 = n2408 & ~n5907 ;
  assign n5909 = n2411 & ~n5908 ;
  assign n5910 = n1721 & ~n5909 ;
  assign n5911 = n1725 & ~n5910 ;
  assign n5912 = n1729 & ~n5911 ;
  assign n5913 = n1733 & ~n5912 ;
  assign n5914 = n1737 & ~n5913 ;
  assign n5915 = n1741 & ~n5914 ;
  assign n5916 = n1745 & ~n5915 ;
  assign n5917 = n1749 & ~n5916 ;
  assign n5918 = n1753 & ~n5917 ;
  assign n5919 = n1757 & ~n5918 ;
  assign n5920 = n433 & n440 ;
  assign n5921 = ~n1759 & n5920 ;
  assign n5922 = ~n5919 & n5921 ;
  assign n5923 = n1765 & ~n5922 ;
  assign n5924 = n1769 & ~n5923 ;
  assign n5925 = n1773 & ~n5924 ;
  assign n5926 = n1777 & ~n5925 ;
  assign n5927 = n1781 & ~n5926 ;
  assign n5928 = n1785 & ~n5927 ;
  assign n5929 = ~n1787 & n1788 ;
  assign n5930 = ~n5928 & n5929 ;
  assign n5931 = n3920 & ~n5930 ;
  assign n5932 = n1797 & ~n5931 ;
  assign n5933 = n1801 & ~n5932 ;
  assign n5934 = n1805 & ~n5933 ;
  assign n5935 = n589 & n5901 ;
  assign n5936 = ~n1807 & n5935 ;
  assign n5937 = ~n5934 & n5936 ;
  assign n5938 = ~n5902 & ~n5937 ;
  assign n5939 = \req[117]  & ~n961 ;
  assign n5940 = ~n947 & n5939 ;
  assign n5941 = ~\priority[119]  & ~n967 ;
  assign n5942 = n592 & ~n5941 ;
  assign n5943 = n610 & ~n5942 ;
  assign n5944 = n2090 & ~n5943 ;
  assign n5945 = n2094 & ~n5944 ;
  assign n5946 = n2447 & ~n5945 ;
  assign n5947 = n2450 & ~n5946 ;
  assign n5948 = n1837 & ~n5947 ;
  assign n5949 = n1841 & ~n5948 ;
  assign n5950 = n1845 & ~n5949 ;
  assign n5951 = n1849 & ~n5950 ;
  assign n5952 = n3720 & ~n5951 ;
  assign n5953 = n1857 & ~n5952 ;
  assign n5954 = n1861 & ~n5953 ;
  assign n5955 = n1865 & ~n5954 ;
  assign n5956 = n1869 & ~n5955 ;
  assign n5957 = n1873 & ~n5956 ;
  assign n5958 = n1877 & ~n5957 ;
  assign n5959 = n3627 & ~n5958 ;
  assign n5960 = n1885 & ~n5959 ;
  assign n5961 = n1889 & ~n5960 ;
  assign n5962 = n1893 & ~n5961 ;
  assign n5963 = n1897 & ~n5962 ;
  assign n5964 = n1901 & ~n5963 ;
  assign n5965 = n1905 & ~n5964 ;
  assign n5966 = n1909 & ~n5965 ;
  assign n5967 = n4592 & ~n5966 ;
  assign n5968 = n1916 & ~n5647 ;
  assign n5969 = ~n5967 & n5968 ;
  assign n5970 = n1921 & ~n5969 ;
  assign n5971 = n956 & n5939 ;
  assign n5972 = ~n1923 & n5971 ;
  assign n5973 = ~n5970 & n5972 ;
  assign n5974 = ~n5940 & ~n5973 ;
  assign n5975 = \req[118]  & ~n1327 ;
  assign n5976 = ~n1313 & n5975 ;
  assign n5977 = ~\priority[120]  & ~n1333 ;
  assign n5978 = n959 & ~n5977 ;
  assign n5979 = n977 & ~n5978 ;
  assign n5980 = n2132 & ~n5979 ;
  assign n5981 = n2136 & ~n5980 ;
  assign n5982 = n2487 & ~n5981 ;
  assign n5983 = n2490 & ~n5982 ;
  assign n5984 = n1953 & ~n5983 ;
  assign n5985 = n1957 & ~n5984 ;
  assign n5986 = n1961 & ~n5985 ;
  assign n5987 = n1965 & ~n5986 ;
  assign n5988 = n1969 & ~n5987 ;
  assign n5989 = n1973 & ~n5988 ;
  assign n5990 = n2713 & ~n5989 ;
  assign n5991 = n1981 & ~n5990 ;
  assign n5992 = n1985 & ~n5991 ;
  assign n5993 = n1989 & ~n5992 ;
  assign n5994 = n1993 & ~n5993 ;
  assign n5995 = n1997 & ~n5994 ;
  assign n5996 = n2001 & ~n5995 ;
  assign n5997 = n2005 & ~n5996 ;
  assign n5998 = n2009 & ~n5997 ;
  assign n5999 = n2013 & ~n5998 ;
  assign n6000 = n2017 & ~n5999 ;
  assign n6001 = n2021 & ~n6000 ;
  assign n6002 = n2025 & ~n6001 ;
  assign n6003 = n3671 & ~n6002 ;
  assign n6004 = n2033 & ~n6003 ;
  assign n6005 = n2037 & ~n6004 ;
  assign n6006 = n1322 & n5975 ;
  assign n6007 = ~n2039 & n6006 ;
  assign n6008 = ~n6005 & n6007 ;
  assign n6009 = ~n5976 & ~n6008 ;
  assign n6010 = \req[119]  & ~n591 ;
  assign n6011 = ~n602 & n6010 ;
  assign n6012 = ~\priority[121]  & ~n607 ;
  assign n6013 = n1325 & ~n6012 ;
  assign n6014 = n1343 & ~n6013 ;
  assign n6015 = n2173 & ~n6014 ;
  assign n6016 = n2176 & ~n6015 ;
  assign n6017 = n286 & ~n6016 ;
  assign n6018 = n5373 & ~n6017 ;
  assign n6019 = n312 & ~n6018 ;
  assign n6020 = n325 & ~n6019 ;
  assign n6021 = n338 & ~n6020 ;
  assign n6022 = n5379 & ~n6021 ;
  assign n6023 = n364 & ~n6022 ;
  assign n6024 = n377 & ~n6023 ;
  assign n6025 = n390 & ~n6024 ;
  assign n6026 = n5706 & ~n6025 ;
  assign n6027 = n416 & ~n6026 ;
  assign n6028 = n4115 & ~n6027 ;
  assign n6029 = n424 & ~n433 ;
  assign n6030 = n441 & ~n6029 ;
  assign n6031 = ~n6028 & n6030 ;
  assign n6032 = n455 & ~n6031 ;
  assign n6033 = n468 & ~n6032 ;
  assign n6034 = n5713 & ~n6033 ;
  assign n6035 = n494 & ~n6034 ;
  assign n6036 = n507 & ~n6035 ;
  assign n6037 = n520 & ~n6036 ;
  assign n6038 = n533 & ~n6037 ;
  assign n6039 = n546 & ~n6038 ;
  assign n6040 = n559 & ~n6039 ;
  assign n6041 = n572 & ~n6040 ;
  assign n6042 = n585 & ~n6041 ;
  assign n6043 = n596 & n6010 ;
  assign n6044 = ~n590 & n6043 ;
  assign n6045 = ~n6042 & n6044 ;
  assign n6046 = ~n6011 & ~n6045 ;
  assign n6047 = \req[120]  & ~n958 ;
  assign n6048 = ~n969 & n6047 ;
  assign n6049 = ~\priority[122]  & ~n974 ;
  assign n6050 = n614 & ~n6049 ;
  assign n6051 = n1467 & ~n6050 ;
  assign n6052 = n2212 & ~n6051 ;
  assign n6053 = n4453 & ~n6052 ;
  assign n6054 = n5410 & ~n6053 ;
  assign n6055 = n666 & ~n6054 ;
  assign n6056 = n679 & ~n6055 ;
  assign n6057 = n3826 & ~n6056 ;
  assign n6058 = n4459 & ~n6057 ;
  assign n6059 = n718 & ~n6058 ;
  assign n6060 = n731 & ~n6059 ;
  assign n6061 = n4464 & ~n6060 ;
  assign n6062 = n2465 & ~n6061 ;
  assign n6063 = n770 & ~n6062 ;
  assign n6064 = n3099 & ~n6063 ;
  assign n6065 = n796 & ~n6064 ;
  assign n6066 = n809 & ~n6065 ;
  assign n6067 = n2117 & ~n6066 ;
  assign n6068 = n835 & ~n6067 ;
  assign n6069 = n848 & ~n6068 ;
  assign n6070 = n5107 & ~n6069 ;
  assign n6071 = n874 & ~n6070 ;
  assign n6072 = ~n879 & n886 ;
  assign n6073 = ~n6071 & n6072 ;
  assign n6074 = n900 & ~n6073 ;
  assign n6075 = n913 & ~n6074 ;
  assign n6076 = n926 & ~n6075 ;
  assign n6077 = n939 & ~n6076 ;
  assign n6078 = n952 & ~n6077 ;
  assign n6079 = n963 & n6047 ;
  assign n6080 = ~n957 & n6079 ;
  assign n6081 = ~n6078 & n6080 ;
  assign n6082 = ~n6048 & ~n6081 ;
  assign n6083 = \req[121]  & ~n1324 ;
  assign n6084 = ~n1335 & n6083 ;
  assign n6085 = ~\priority[123]  & ~n1340 ;
  assign n6086 = n981 & ~n6085 ;
  assign n6087 = n1587 & ~n6086 ;
  assign n6088 = n2252 & ~n6087 ;
  assign n6089 = n2255 & ~n6088 ;
  assign n6090 = n1019 & ~n6089 ;
  assign n6091 = n1032 & ~n6090 ;
  assign n6092 = n3861 & ~n6091 ;
  assign n6093 = n1058 & ~n6092 ;
  assign n6094 = n1071 & ~n6093 ;
  assign n6095 = n1084 & ~n6094 ;
  assign n6096 = n1097 & ~n6095 ;
  assign n6097 = n1110 & ~n6096 ;
  assign n6098 = n1123 & ~n6097 ;
  assign n6099 = n1136 & ~n6098 ;
  assign n6100 = n5137 & ~n6099 ;
  assign n6101 = n1162 & ~n6100 ;
  assign n6102 = n1175 & ~n6101 ;
  assign n6103 = n1188 & ~n6102 ;
  assign n6104 = n1201 & ~n6103 ;
  assign n6105 = n1214 & ~n6104 ;
  assign n6106 = n1227 & ~n6105 ;
  assign n6107 = n1240 & ~n6106 ;
  assign n6108 = n1253 & ~n6107 ;
  assign n6109 = n4409 & ~n6108 ;
  assign n6110 = n1279 & ~n6109 ;
  assign n6111 = n1292 & ~n6110 ;
  assign n6112 = n1305 & ~n6111 ;
  assign n6113 = n3148 & ~n6112 ;
  assign n6114 = n1329 & n6083 ;
  assign n6115 = ~n1323 & n6114 ;
  assign n6116 = ~n6113 & n6115 ;
  assign n6117 = ~n6084 & ~n6116 ;
  assign n6118 = \req[122]  & ~n613 ;
  assign n6119 = ~n609 & n6118 ;
  assign n6120 = ~\priority[124]  & ~n604 ;
  assign n6121 = n1347 & ~n6120 ;
  assign n6122 = n1704 & ~n6121 ;
  assign n6123 = n2291 & ~n6122 ;
  assign n6124 = n2294 & ~n6123 ;
  assign n6125 = n1368 & ~n6124 ;
  assign n6126 = n1372 & ~n6125 ;
  assign n6127 = n1376 & ~n6126 ;
  assign n6128 = n1380 & ~n6127 ;
  assign n6129 = n1384 & ~n6128 ;
  assign n6130 = n1388 & ~n6129 ;
  assign n6131 = n1392 & ~n6130 ;
  assign n6132 = n1396 & ~n6131 ;
  assign n6133 = n5491 & ~n6132 ;
  assign n6134 = n1404 & ~n6133 ;
  assign n6135 = n1408 & ~n6134 ;
  assign n6136 = n1412 & ~n6135 ;
  assign n6137 = n1416 & ~n6136 ;
  assign n6138 = n1420 & ~n6137 ;
  assign n6139 = n1424 & ~n6138 ;
  assign n6140 = n1428 & ~n6139 ;
  assign n6141 = n1432 & ~n6140 ;
  assign n6142 = n5501 & ~n6141 ;
  assign n6143 = n1440 & ~n6142 ;
  assign n6144 = n3811 & ~n6143 ;
  assign n6145 = n1448 & ~n6144 ;
  assign n6146 = n1452 & ~n6145 ;
  assign n6147 = n1456 & ~n6146 ;
  assign n6148 = n3817 & ~n6147 ;
  assign n6149 = n593 & n6118 ;
  assign n6150 = ~n1462 & n6149 ;
  assign n6151 = ~n6148 & n6150 ;
  assign n6152 = ~n6119 & ~n6151 ;
  assign n6153 = \req[123]  & ~n980 ;
  assign n6154 = ~n976 & n6153 ;
  assign n6155 = ~\priority[125]  & ~n971 ;
  assign n6156 = n618 & ~n6155 ;
  assign n6157 = n1820 & ~n6156 ;
  assign n6158 = n2330 & ~n6157 ;
  assign n6159 = n2333 & ~n6158 ;
  assign n6160 = n1488 & ~n6159 ;
  assign n6161 = n1492 & ~n6160 ;
  assign n6162 = n1496 & ~n6161 ;
  assign n6163 = n1500 & ~n6162 ;
  assign n6164 = n1504 & ~n6163 ;
  assign n6165 = n2229 & ~n6164 ;
  assign n6166 = n1512 & ~n6165 ;
  assign n6167 = n1516 & ~n6166 ;
  assign n6168 = n1520 & ~n6167 ;
  assign n6169 = n1524 & ~n6168 ;
  assign n6170 = n1528 & ~n6169 ;
  assign n6171 = n1532 & ~n6170 ;
  assign n6172 = n1536 & ~n6171 ;
  assign n6173 = n1540 & ~n6172 ;
  assign n6174 = n1544 & ~n6173 ;
  assign n6175 = n1548 & ~n6174 ;
  assign n6176 = n1552 & ~n6175 ;
  assign n6177 = n1556 & ~n6176 ;
  assign n6178 = n5538 & ~n6177 ;
  assign n6179 = n1564 & ~n6178 ;
  assign n6180 = n1568 & ~n6179 ;
  assign n6181 = n5860 & ~n6180 ;
  assign n6182 = n5441 & ~n6181 ;
  assign n6183 = n1580 & ~n6182 ;
  assign n6184 = n960 & n6153 ;
  assign n6185 = ~n1582 & n6184 ;
  assign n6186 = ~n6183 & n6185 ;
  assign n6187 = ~n6154 & ~n6186 ;
  assign n6188 = \req[124]  & ~n1346 ;
  assign n6189 = ~n1342 & n6188 ;
  assign n6190 = ~\priority[126]  & ~n1337 ;
  assign n6191 = n985 & ~n6190 ;
  assign n6192 = n1936 & ~n6191 ;
  assign n6193 = n2369 & ~n6192 ;
  assign n6194 = n2372 & ~n6193 ;
  assign n6195 = n1605 & ~n6194 ;
  assign n6196 = n1609 & ~n6195 ;
  assign n6197 = n1613 & ~n6196 ;
  assign n6198 = n1617 & ~n6197 ;
  assign n6199 = ~n1619 & n1620 ;
  assign n6200 = ~n6198 & n6199 ;
  assign n6201 = n1625 & ~n6200 ;
  assign n6202 = n1629 & ~n6201 ;
  assign n6203 = n1633 & ~n6202 ;
  assign n6204 = n5564 & ~n6203 ;
  assign n6205 = n1641 & ~n6204 ;
  assign n6206 = n1645 & ~n6205 ;
  assign n6207 = n1649 & ~n6206 ;
  assign n6208 = n4614 & ~n6207 ;
  assign n6209 = n1657 & ~n6208 ;
  assign n6210 = n4930 & ~n6209 ;
  assign n6211 = n1665 & ~n6210 ;
  assign n6212 = n1669 & ~n6211 ;
  assign n6213 = n1673 & ~n6212 ;
  assign n6214 = n1677 & ~n6213 ;
  assign n6215 = n1681 & ~n6214 ;
  assign n6216 = n1685 & ~n6215 ;
  assign n6217 = n1689 & ~n6216 ;
  assign n6218 = n1693 & ~n6217 ;
  assign n6219 = n1697 & ~n6218 ;
  assign n6220 = n1326 & n6188 ;
  assign n6221 = ~n1699 & n6220 ;
  assign n6222 = ~n6219 & n6221 ;
  assign n6223 = ~n6189 & ~n6222 ;
  assign n6224 = \req[125]  & ~n617 ;
  assign n6225 = ~n606 & n6224 ;
  assign n6226 = ~\priority[127]  & ~n257 ;
  assign n6227 = n1351 & ~n6226 ;
  assign n6228 = n2052 & ~n6227 ;
  assign n6229 = n2408 & ~n6228 ;
  assign n6230 = n2411 & ~n6229 ;
  assign n6231 = n1721 & ~n6230 ;
  assign n6232 = n1725 & ~n6231 ;
  assign n6233 = n1729 & ~n6232 ;
  assign n6234 = n1733 & ~n6233 ;
  assign n6235 = n1737 & ~n6234 ;
  assign n6236 = n1741 & ~n6235 ;
  assign n6237 = n1745 & ~n6236 ;
  assign n6238 = n1749 & ~n6237 ;
  assign n6239 = n1753 & ~n6238 ;
  assign n6240 = n1757 & ~n6239 ;
  assign n6241 = n5921 & ~n6240 ;
  assign n6242 = n1765 & ~n6241 ;
  assign n6243 = n1769 & ~n6242 ;
  assign n6244 = n1773 & ~n6243 ;
  assign n6245 = n1777 & ~n6244 ;
  assign n6246 = n1781 & ~n6245 ;
  assign n6247 = n1785 & ~n6246 ;
  assign n6248 = n5929 & ~n6247 ;
  assign n6249 = n3920 & ~n6248 ;
  assign n6250 = n1797 & ~n6249 ;
  assign n6251 = n1801 & ~n6250 ;
  assign n6252 = n1805 & ~n6251 ;
  assign n6253 = n4558 & ~n6252 ;
  assign n6254 = n1813 & ~n6253 ;
  assign n6255 = n615 & n6224 ;
  assign n6256 = ~n1815 & n6255 ;
  assign n6257 = ~n6254 & n6256 ;
  assign n6258 = ~n6225 & ~n6257 ;
  assign n6259 = \req[126]  & ~n984 ;
  assign n6260 = ~n973 & n6259 ;
  assign n6261 = ~\priority[0]  & ~n624 ;
  assign n6262 = n1471 & ~n6261 ;
  assign n6263 = n2093 & ~n6262 ;
  assign n6264 = n2447 & ~n6263 ;
  assign n6265 = n2450 & ~n6264 ;
  assign n6266 = n1837 & ~n6265 ;
  assign n6267 = n1841 & ~n6266 ;
  assign n6268 = n1845 & ~n6267 ;
  assign n6269 = n1849 & ~n6268 ;
  assign n6270 = n3720 & ~n6269 ;
  assign n6271 = n1857 & ~n6270 ;
  assign n6272 = n1861 & ~n6271 ;
  assign n6273 = n1865 & ~n6272 ;
  assign n6274 = n1869 & ~n6273 ;
  assign n6275 = n1873 & ~n6274 ;
  assign n6276 = n1877 & ~n6275 ;
  assign n6277 = n3627 & ~n6276 ;
  assign n6278 = n1885 & ~n6277 ;
  assign n6279 = n1889 & ~n6278 ;
  assign n6280 = n1893 & ~n6279 ;
  assign n6281 = n1897 & ~n6280 ;
  assign n6282 = n1901 & ~n6281 ;
  assign n6283 = n1905 & ~n6282 ;
  assign n6284 = n1909 & ~n6283 ;
  assign n6285 = n4592 & ~n6284 ;
  assign n6286 = n5968 & ~n6285 ;
  assign n6287 = n1921 & ~n6286 ;
  assign n6288 = n1925 & ~n6287 ;
  assign n6289 = n1929 & ~n6288 ;
  assign n6290 = n982 & n6259 ;
  assign n6291 = ~n1931 & n6290 ;
  assign n6292 = ~n6289 & n6291 ;
  assign n6293 = ~n6260 & ~n6292 ;
  assign n6294 = \req[127]  & ~n1350 ;
  assign n6295 = ~n1339 & n6294 ;
  assign n6296 = ~\priority[1]  & ~n991 ;
  assign n6297 = n1591 & ~n6296 ;
  assign n6298 = n2135 & ~n6297 ;
  assign n6299 = n2487 & ~n6298 ;
  assign n6300 = n2490 & ~n6299 ;
  assign n6301 = n1953 & ~n6300 ;
  assign n6302 = n1957 & ~n6301 ;
  assign n6303 = n1961 & ~n6302 ;
  assign n6304 = n1965 & ~n6303 ;
  assign n6305 = n1969 & ~n6304 ;
  assign n6306 = n1973 & ~n6305 ;
  assign n6307 = n2713 & ~n6306 ;
  assign n6308 = n1981 & ~n6307 ;
  assign n6309 = n1985 & ~n6308 ;
  assign n6310 = n1989 & ~n6309 ;
  assign n6311 = n1993 & ~n6310 ;
  assign n6312 = n1997 & ~n6311 ;
  assign n6313 = n2001 & ~n6312 ;
  assign n6314 = n2005 & ~n6313 ;
  assign n6315 = n2009 & ~n6314 ;
  assign n6316 = n2013 & ~n6315 ;
  assign n6317 = n2017 & ~n6316 ;
  assign n6318 = n2021 & ~n6317 ;
  assign n6319 = n2025 & ~n6318 ;
  assign n6320 = n3671 & ~n6319 ;
  assign n6321 = n2033 & ~n6320 ;
  assign n6322 = n2037 & ~n6321 ;
  assign n6323 = n2041 & ~n6322 ;
  assign n6324 = n2045 & ~n6323 ;
  assign n6325 = n1348 & n6294 ;
  assign n6326 = ~n2047 & n6325 ;
  assign n6327 = ~n6324 & n6326 ;
  assign n6328 = ~n6295 & ~n6327 ;
  assign n6329 = n614 & n643 ;
  assign n6330 = n647 & n676 ;
  assign n6331 = n6329 & n6330 ;
  assign n6332 = n543 & n562 ;
  assign n6333 = n566 & n595 ;
  assign n6334 = n6332 & n6333 ;
  assign n6335 = n6331 & n6334 ;
  assign n6336 = n751 & n780 ;
  assign n6337 = n799 & n803 ;
  assign n6338 = n6336 & n6337 ;
  assign n6339 = n695 & n699 ;
  assign n6340 = n728 & n747 ;
  assign n6341 = n6339 & n6340 ;
  assign n6342 = n6338 & n6341 ;
  assign n6343 = n6335 & n6342 ;
  assign n6344 = n335 & n354 ;
  assign n6345 = n358 & n387 ;
  assign n6346 = n6344 & n6345 ;
  assign n6347 = n265 & n283 ;
  assign n6348 = n302 & n306 ;
  assign n6349 = n6347 & n6348 ;
  assign n6350 = n6346 & n6349 ;
  assign n6351 = n462 & n491 ;
  assign n6352 = n510 & n514 ;
  assign n6353 = n6351 & n6352 ;
  assign n6354 = n406 & n410 ;
  assign n6355 = n439 & n458 ;
  assign n6356 = n6354 & n6355 ;
  assign n6357 = n6353 & n6356 ;
  assign n6358 = n6350 & n6357 ;
  assign n6359 = n6343 & n6358 ;
  assign n6360 = n1172 & n1191 ;
  assign n6361 = n1195 & n1224 ;
  assign n6362 = n6360 & n6361 ;
  assign n6363 = n1091 & n1120 ;
  assign n6364 = n1139 & n1143 ;
  assign n6365 = n6363 & n6364 ;
  assign n6366 = n6362 & n6365 ;
  assign n6367 = n1299 & n1328 ;
  assign n6368 = n1347 & n1471 ;
  assign n6369 = n6367 & n6368 ;
  assign n6370 = n1243 & n1247 ;
  assign n6371 = n1276 & n1295 ;
  assign n6372 = n6370 & n6371 ;
  assign n6373 = n6369 & n6372 ;
  assign n6374 = n6366 & n6373 ;
  assign n6375 = n903 & n907 ;
  assign n6376 = n936 & n955 ;
  assign n6377 = n6375 & n6376 ;
  assign n6378 = n832 & n851 ;
  assign n6379 = n855 & n884 ;
  assign n6380 = n6378 & n6379 ;
  assign n6381 = n6377 & n6380 ;
  assign n6382 = n1035 & n1039 ;
  assign n6383 = n1068 & n1087 ;
  assign n6384 = n6382 & n6383 ;
  assign n6385 = n959 & n985 ;
  assign n6386 = n998 & n1016 ;
  assign n6387 = n6385 & n6386 ;
  assign n6388 = n6384 & n6387 ;
  assign n6389 = n6381 & n6388 ;
  assign n6390 = n6374 & n6389 ;
  assign n6391 = n6359 & n6390 ;
  assign \grant[0]  = ~n623 ;
  assign \grant[1]  = ~n990 ;
  assign \grant[2]  = ~n1356 ;
  assign \grant[3]  = ~n1476 ;
  assign \grant[4]  = ~n1596 ;
  assign \grant[5]  = ~n1712 ;
  assign \grant[6]  = ~n1828 ;
  assign \grant[7]  = ~n1944 ;
  assign \grant[8]  = ~n2059 ;
  assign \grant[9]  = ~n2100 ;
  assign \grant[10]  = ~n2142 ;
  assign \grant[11]  = ~n2181 ;
  assign \grant[12]  = ~n2220 ;
  assign \grant[13]  = ~n2260 ;
  assign \grant[14]  = ~n2299 ;
  assign \grant[15]  = ~n2338 ;
  assign \grant[16]  = ~n2377 ;
  assign \grant[17]  = ~n2416 ;
  assign \grant[18]  = ~n2455 ;
  assign \grant[19]  = ~n2495 ;
  assign \grant[20]  = ~n2530 ;
  assign \grant[21]  = ~n2565 ;
  assign \grant[22]  = ~n2600 ;
  assign \grant[23]  = ~n2635 ;
  assign \grant[24]  = ~n2670 ;
  assign \grant[25]  = ~n2705 ;
  assign \grant[26]  = ~n2741 ;
  assign \grant[27]  = ~n2776 ;
  assign \grant[28]  = ~n2811 ;
  assign \grant[29]  = ~n2846 ;
  assign \grant[30]  = ~n2881 ;
  assign \grant[31]  = ~n2916 ;
  assign \grant[32]  = ~n2951 ;
  assign \grant[33]  = ~n2986 ;
  assign \grant[34]  = ~n3021 ;
  assign \grant[35]  = ~n3056 ;
  assign \grant[36]  = ~n3091 ;
  assign \grant[37]  = ~n3127 ;
  assign \grant[38]  = ~n3163 ;
  assign \grant[39]  = ~n3198 ;
  assign \grant[40]  = ~n3233 ;
  assign \grant[41]  = ~n3268 ;
  assign \grant[42]  = ~n3303 ;
  assign \grant[43]  = ~n3338 ;
  assign \grant[44]  = ~n3373 ;
  assign \grant[45]  = ~n3408 ;
  assign \grant[46]  = ~n3443 ;
  assign \grant[47]  = ~n3478 ;
  assign \grant[48]  = ~n3513 ;
  assign \grant[49]  = ~n3548 ;
  assign \grant[50]  = ~n3585 ;
  assign \grant[51]  = ~n3620 ;
  assign \grant[52]  = ~n3656 ;
  assign \grant[53]  = ~n3692 ;
  assign \grant[54]  = ~n3728 ;
  assign \grant[55]  = ~n3763 ;
  assign \grant[56]  = ~n3798 ;
  assign \grant[57]  = ~n3837 ;
  assign \grant[58]  = ~n3873 ;
  assign \grant[59]  = ~n3908 ;
  assign \grant[60]  = ~n3944 ;
  assign \grant[61]  = ~n3979 ;
  assign \grant[62]  = ~n4014 ;
  assign \grant[63]  = ~n4049 ;
  assign \grant[64]  = ~n4084 ;
  assign \grant[65]  = ~n4120 ;
  assign \grant[66]  = ~n4155 ;
  assign \grant[67]  = ~n4190 ;
  assign \grant[68]  = ~n4225 ;
  assign \grant[69]  = ~n4260 ;
  assign \grant[70]  = ~n4295 ;
  assign \grant[71]  = ~n4330 ;
  assign \grant[72]  = ~n4365 ;
  assign \grant[73]  = ~n4400 ;
  assign \grant[74]  = ~n4436 ;
  assign \grant[75]  = ~n4475 ;
  assign \grant[76]  = ~n4510 ;
  assign \grant[77]  = ~n4545 ;
  assign \grant[78]  = ~n4582 ;
  assign \grant[79]  = ~n4620 ;
  assign \grant[80]  = ~n4655 ;
  assign \grant[81]  = ~n4690 ;
  assign \grant[82]  = ~n4725 ;
  assign \grant[83]  = ~n4760 ;
  assign \grant[84]  = ~n4795 ;
  assign \grant[85]  = ~n4830 ;
  assign \grant[86]  = ~n4865 ;
  assign \grant[87]  = ~n4900 ;
  assign \grant[88]  = ~n4936 ;
  assign \grant[89]  = ~n4971 ;
  assign \grant[90]  = ~n5006 ;
  assign \grant[91]  = ~n5041 ;
  assign \grant[92]  = ~n5077 ;
  assign \grant[93]  = ~n5113 ;
  assign \grant[94]  = ~n5149 ;
  assign \grant[95]  = ~n5184 ;
  assign \grant[96]  = ~n5219 ;
  assign \grant[97]  = ~n5254 ;
  assign \grant[98]  = ~n5289 ;
  assign \grant[99]  = ~n5324 ;
  assign \grant[100]  = ~n5359 ;
  assign \grant[101]  = ~n5398 ;
  assign \grant[102]  = ~n5434 ;
  assign \grant[103]  = ~n5471 ;
  assign \grant[104]  = ~n5508 ;
  assign \grant[105]  = ~n5544 ;
  assign \grant[106]  = ~n5580 ;
  assign \grant[107]  = ~n5615 ;
  assign \grant[108]  = ~n5651 ;
  assign \grant[109]  = ~n5686 ;
  assign \grant[110]  = ~n5724 ;
  assign \grant[111]  = ~n5759 ;
  assign \grant[112]  = ~n5794 ;
  assign \grant[113]  = ~n5829 ;
  assign \grant[114]  = ~n5865 ;
  assign \grant[115]  = ~n5900 ;
  assign \grant[116]  = ~n5938 ;
  assign \grant[117]  = ~n5974 ;
  assign \grant[118]  = ~n6009 ;
  assign \grant[119]  = ~n6046 ;
  assign \grant[120]  = ~n6082 ;
  assign \grant[121]  = ~n6117 ;
  assign \grant[122]  = ~n6152 ;
  assign \grant[123]  = ~n6187 ;
  assign \grant[124]  = ~n6223 ;
  assign \grant[125]  = ~n6258 ;
  assign \grant[126]  = ~n6293 ;
  assign \grant[127]  = ~n6328 ;
  assign anyGrant = ~n6391 ;
endmodule
