module top( \cont_reg[0]/NET0131  , \cont_reg[1]/NET0131  , \cont_reg[2]/NET0131  , \cont_reg[3]/NET0131  , \cont_reg[4]/NET0131  , \cont_reg[5]/NET0131  , \cont_reg[6]/NET0131  , \cont_reg[7]/NET0131  , \mar_reg[0]/NET0131  , \mar_reg[1]/NET0131  , \mar_reg[2]/NET0131  , \mar_reg[3]/NET0131  , \punti_retta[3]_pad  , \punti_retta[4]_pad  , \punti_retta[6]_pad  , \punti_retta[7]_pad  , \punti_retta_reg[0]/NET0131  , \punti_retta_reg[1]/NET0131  , \punti_retta_reg[2]/NET0131  , \punti_retta_reg[5]/NET0131  , start_pad , \stato_reg[0]/NET0131  , \stato_reg[1]/NET0131  , \stato_reg[2]/NET0131  , \t_reg[1]/NET0131  , \t_reg[2]/NET0131  , \t_reg[3]/NET0131  , \t_reg[4]/NET0131  , \t_reg[5]/NET0131  , \t_reg[6]/NET0131  , \x_reg[0]/NET0131  , \x_reg[1]/NET0131  , \x_reg[2]/NET0131  , \x_reg[3]/NET0131  , \x_reg[4]/NET0131  , \x_reg[5]/NET0131  , \x_reg[6]/NET0131  , \x_reg[7]/NET0131  , \y_reg[0]/NET0131  , \y_reg[1]/NET0131  , \y_reg[2]/NET0131  , \y_reg[3]/NET0131  , \_al_n0  , \_al_n1  , \g2119/_0_  , \g2123/_0_  , \g2129/_0_  , \g2133/_0_  , \g2136/_0_  , \g2140/_0_  , \g2141/_0_  , \g2151/_0_  , \g2152/_0_  , \g2166/_0_  , \g2167/_0_  , \g2180/_0_  , \g2181/_0_  , \g2199/_0_  , \g2225/_0_  , \g2227/_0_  , \g2242/_0_  , \g2243/_0_  , \g2272/_0_  , \g2273/_0_  , \g2274/_0_  , \g2275/_0_  , \g2284/_0_  , \g2289/_0_  , \g2303/_0_  , \g2304/_0_  , \g2308/_0_  , \g2309/_0_  , \g2310/_0_  , \g2311/_0_  , \g2312/_0_  , \g2346/_0_  , \g2973/_0_  , \g2984/_0_  , \g3052/_0_  , \g3176/_0_  , \g3277/_0_  , \g3306/_0_  , \g3366/_0_  , \g3371/_0_  , \g3398/_0_  );
  input \cont_reg[0]/NET0131  ;
  input \cont_reg[1]/NET0131  ;
  input \cont_reg[2]/NET0131  ;
  input \cont_reg[3]/NET0131  ;
  input \cont_reg[4]/NET0131  ;
  input \cont_reg[5]/NET0131  ;
  input \cont_reg[6]/NET0131  ;
  input \cont_reg[7]/NET0131  ;
  input \mar_reg[0]/NET0131  ;
  input \mar_reg[1]/NET0131  ;
  input \mar_reg[2]/NET0131  ;
  input \mar_reg[3]/NET0131  ;
  input \punti_retta[3]_pad  ;
  input \punti_retta[4]_pad  ;
  input \punti_retta[6]_pad  ;
  input \punti_retta[7]_pad  ;
  input \punti_retta_reg[0]/NET0131  ;
  input \punti_retta_reg[1]/NET0131  ;
  input \punti_retta_reg[2]/NET0131  ;
  input \punti_retta_reg[5]/NET0131  ;
  input start_pad ;
  input \stato_reg[0]/NET0131  ;
  input \stato_reg[1]/NET0131  ;
  input \stato_reg[2]/NET0131  ;
  input \t_reg[1]/NET0131  ;
  input \t_reg[2]/NET0131  ;
  input \t_reg[3]/NET0131  ;
  input \t_reg[4]/NET0131  ;
  input \t_reg[5]/NET0131  ;
  input \t_reg[6]/NET0131  ;
  input \x_reg[0]/NET0131  ;
  input \x_reg[1]/NET0131  ;
  input \x_reg[2]/NET0131  ;
  input \x_reg[3]/NET0131  ;
  input \x_reg[4]/NET0131  ;
  input \x_reg[5]/NET0131  ;
  input \x_reg[6]/NET0131  ;
  input \x_reg[7]/NET0131  ;
  input \y_reg[0]/NET0131  ;
  input \y_reg[1]/NET0131  ;
  input \y_reg[2]/NET0131  ;
  input \y_reg[3]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g2119/_0_  ;
  output \g2123/_0_  ;
  output \g2129/_0_  ;
  output \g2133/_0_  ;
  output \g2136/_0_  ;
  output \g2140/_0_  ;
  output \g2141/_0_  ;
  output \g2151/_0_  ;
  output \g2152/_0_  ;
  output \g2166/_0_  ;
  output \g2167/_0_  ;
  output \g2180/_0_  ;
  output \g2181/_0_  ;
  output \g2199/_0_  ;
  output \g2225/_0_  ;
  output \g2227/_0_  ;
  output \g2242/_0_  ;
  output \g2243/_0_  ;
  output \g2272/_0_  ;
  output \g2273/_0_  ;
  output \g2274/_0_  ;
  output \g2275/_0_  ;
  output \g2284/_0_  ;
  output \g2289/_0_  ;
  output \g2303/_0_  ;
  output \g2304/_0_  ;
  output \g2308/_0_  ;
  output \g2309/_0_  ;
  output \g2310/_0_  ;
  output \g2311/_0_  ;
  output \g2312/_0_  ;
  output \g2346/_0_  ;
  output \g2973/_0_  ;
  output \g2984/_0_  ;
  output \g3052/_0_  ;
  output \g3176/_0_  ;
  output \g3277/_0_  ;
  output \g3306/_0_  ;
  output \g3366/_0_  ;
  output \g3371/_0_  ;
  output \g3398/_0_  ;
  wire n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 ;
  assign n43 = ~\stato_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n44 = \stato_reg[2]/NET0131  & n43 ;
  assign n47 = ~\x_reg[4]/NET0131  & ~\x_reg[5]/NET0131  ;
  assign n48 = ~\x_reg[6]/NET0131  & ~\x_reg[7]/NET0131  ;
  assign n49 = n47 & n48 ;
  assign n45 = ~\x_reg[0]/NET0131  & \x_reg[1]/NET0131  ;
  assign n46 = ~\x_reg[2]/NET0131  & ~\x_reg[3]/NET0131  ;
  assign n50 = n45 & n46 ;
  assign n51 = n49 & n50 ;
  assign n52 = \cont_reg[0]/NET0131  & \cont_reg[1]/NET0131  ;
  assign n53 = \cont_reg[2]/NET0131  & \cont_reg[3]/NET0131  ;
  assign n54 = n52 & n53 ;
  assign n55 = n51 & n54 ;
  assign n56 = \cont_reg[4]/NET0131  & n55 ;
  assign n57 = \cont_reg[5]/NET0131  & n56 ;
  assign n58 = \mar_reg[0]/NET0131  & \mar_reg[1]/NET0131  ;
  assign n59 = \mar_reg[2]/NET0131  & n58 ;
  assign n60 = \mar_reg[3]/NET0131  & n59 ;
  assign n61 = n57 & ~n60 ;
  assign n62 = n44 & n61 ;
  assign n63 = ~\cont_reg[6]/NET0131  & ~n62 ;
  assign n64 = n44 & ~n61 ;
  assign n65 = ~\stato_reg[1]/NET0131  & ~\stato_reg[2]/NET0131  ;
  assign n66 = \stato_reg[0]/NET0131  & n65 ;
  assign n67 = ~start_pad & n66 ;
  assign n68 = \stato_reg[1]/NET0131  & \stato_reg[2]/NET0131  ;
  assign n69 = ~n66 & ~n68 ;
  assign n70 = ~n67 & ~n69 ;
  assign n71 = \cont_reg[6]/NET0131  & n70 ;
  assign n72 = ~n64 & n71 ;
  assign n73 = ~n63 & ~n72 ;
  assign n74 = ~\cont_reg[4]/NET0131  & ~n55 ;
  assign n75 = ~n56 & ~n74 ;
  assign n76 = ~n60 & ~n75 ;
  assign n77 = ~\cont_reg[4]/NET0131  & n60 ;
  assign n78 = n44 & ~n77 ;
  assign n79 = ~n76 & n78 ;
  assign n80 = \cont_reg[4]/NET0131  & ~n70 ;
  assign n81 = ~n79 & ~n80 ;
  assign n82 = \cont_reg[7]/NET0131  & ~n70 ;
  assign n84 = \cont_reg[5]/NET0131  & \cont_reg[6]/NET0131  ;
  assign n85 = n56 & n84 ;
  assign n86 = ~\cont_reg[7]/NET0131  & ~n85 ;
  assign n87 = \cont_reg[7]/NET0131  & n85 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = ~n60 & ~n88 ;
  assign n83 = ~\cont_reg[7]/NET0131  & n60 ;
  assign n90 = n44 & ~n83 ;
  assign n91 = ~n89 & n90 ;
  assign n92 = ~n82 & ~n91 ;
  assign n93 = start_pad & n66 ;
  assign n94 = ~n69 & ~n93 ;
  assign n95 = ~start_pad & n60 ;
  assign n96 = n44 & ~n95 ;
  assign n97 = n94 & ~n96 ;
  assign n98 = \punti_retta[6]_pad  & ~n97 ;
  assign n99 = ~\cont_reg[6]/NET0131  & ~n57 ;
  assign n100 = n44 & n95 ;
  assign n101 = ~n85 & n100 ;
  assign n102 = ~n99 & n101 ;
  assign n103 = ~n98 & ~n102 ;
  assign n104 = \cont_reg[3]/NET0131  & ~n70 ;
  assign n106 = \cont_reg[0]/NET0131  & n51 ;
  assign n107 = \cont_reg[1]/NET0131  & n106 ;
  assign n108 = \cont_reg[2]/NET0131  & n107 ;
  assign n109 = ~\cont_reg[3]/NET0131  & ~n108 ;
  assign n110 = ~n55 & ~n109 ;
  assign n111 = ~n60 & ~n110 ;
  assign n105 = ~\cont_reg[3]/NET0131  & n60 ;
  assign n112 = n44 & ~n105 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = ~n104 & ~n113 ;
  assign n115 = \punti_retta_reg[2]/NET0131  & ~n94 ;
  assign n118 = ~\cont_reg[2]/NET0131  & ~n107 ;
  assign n119 = ~n108 & ~n118 ;
  assign n120 = ~start_pad & n119 ;
  assign n117 = \punti_retta_reg[2]/NET0131  & start_pad ;
  assign n121 = n60 & ~n117 ;
  assign n122 = ~n120 & n121 ;
  assign n116 = ~\punti_retta_reg[2]/NET0131  & ~n60 ;
  assign n123 = n44 & ~n116 ;
  assign n124 = ~n122 & n123 ;
  assign n125 = ~n115 & ~n124 ;
  assign n128 = ~\cont_reg[5]/NET0131  & ~n56 ;
  assign n129 = ~n57 & ~n128 ;
  assign n130 = ~start_pad & n129 ;
  assign n127 = \punti_retta_reg[5]/NET0131  & start_pad ;
  assign n131 = n60 & ~n127 ;
  assign n132 = ~n130 & n131 ;
  assign n126 = ~\punti_retta_reg[5]/NET0131  & ~n60 ;
  assign n133 = n44 & ~n126 ;
  assign n134 = ~n132 & n133 ;
  assign n135 = \punti_retta_reg[5]/NET0131  & ~n94 ;
  assign n136 = ~n134 & ~n135 ;
  assign n137 = ~\cont_reg[0]/NET0131  & ~n51 ;
  assign n138 = ~n106 & ~n137 ;
  assign n139 = n95 & ~n138 ;
  assign n140 = n44 & ~n139 ;
  assign n141 = n94 & ~n140 ;
  assign n142 = \punti_retta_reg[0]/NET0131  & ~n141 ;
  assign n143 = n95 & n140 ;
  assign n144 = ~n142 & ~n143 ;
  assign n145 = \punti_retta_reg[1]/NET0131  & ~n97 ;
  assign n146 = ~\cont_reg[1]/NET0131  & ~n106 ;
  assign n147 = n100 & ~n107 ;
  assign n148 = ~n146 & n147 ;
  assign n149 = ~n145 & ~n148 ;
  assign n150 = ~n60 & ~n129 ;
  assign n151 = ~\cont_reg[5]/NET0131  & n60 ;
  assign n152 = n44 & ~n151 ;
  assign n153 = ~n150 & n152 ;
  assign n154 = \cont_reg[5]/NET0131  & ~n70 ;
  assign n155 = ~n153 & ~n154 ;
  assign n156 = ~n60 & ~n119 ;
  assign n157 = ~\cont_reg[2]/NET0131  & n60 ;
  assign n158 = n44 & ~n157 ;
  assign n159 = ~n156 & n158 ;
  assign n160 = \cont_reg[2]/NET0131  & ~n70 ;
  assign n161 = ~n159 & ~n160 ;
  assign n162 = ~n60 & n106 ;
  assign n163 = n44 & ~n162 ;
  assign n164 = n70 & ~n163 ;
  assign n165 = \cont_reg[1]/NET0131  & ~n164 ;
  assign n166 = ~\cont_reg[1]/NET0131  & n44 ;
  assign n167 = n162 & n166 ;
  assign n168 = ~n165 & ~n167 ;
  assign n169 = ~n60 & ~n138 ;
  assign n170 = ~\cont_reg[0]/NET0131  & n60 ;
  assign n171 = n44 & ~n170 ;
  assign n172 = ~n169 & n171 ;
  assign n173 = \cont_reg[0]/NET0131  & ~n70 ;
  assign n174 = ~n172 & ~n173 ;
  assign n175 = \stato_reg[1]/NET0131  & ~\stato_reg[2]/NET0131  ;
  assign n176 = \stato_reg[0]/NET0131  & n175 ;
  assign n177 = ~n60 & n176 ;
  assign n178 = ~n44 & ~n177 ;
  assign n179 = n59 & ~n178 ;
  assign n180 = ~\mar_reg[3]/NET0131  & ~n179 ;
  assign n181 = ~\stato_reg[1]/NET0131  & \stato_reg[2]/NET0131  ;
  assign n182 = ~\stato_reg[0]/NET0131  & ~\stato_reg[2]/NET0131  ;
  assign n183 = ~n181 & ~n182 ;
  assign n184 = ~n67 & n183 ;
  assign n185 = n178 & n184 ;
  assign n186 = ~n180 & ~n185 ;
  assign n190 = \mar_reg[0]/NET0131  & ~n184 ;
  assign n187 = ~n44 & ~n176 ;
  assign n188 = ~\mar_reg[0]/NET0131  & ~n187 ;
  assign n189 = n44 & n60 ;
  assign n191 = ~n188 & ~n189 ;
  assign n192 = ~n190 & n191 ;
  assign n193 = ~\stato_reg[0]/NET0131  & n181 ;
  assign n194 = \t_reg[1]/NET0131  & \x_reg[1]/NET0131  ;
  assign n195 = ~\t_reg[1]/NET0131  & ~\x_reg[1]/NET0131  ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = n193 & n196 ;
  assign n198 = ~\stato_reg[0]/NET0131  & n175 ;
  assign n199 = \mar_reg[1]/NET0131  & ~\mar_reg[2]/NET0131  ;
  assign n200 = \mar_reg[3]/NET0131  & n199 ;
  assign n201 = ~\mar_reg[0]/NET0131  & n200 ;
  assign n202 = \mar_reg[2]/NET0131  & \mar_reg[3]/NET0131  ;
  assign n203 = \mar_reg[1]/NET0131  & ~n202 ;
  assign n204 = \mar_reg[0]/NET0131  & ~n203 ;
  assign n205 = ~n201 & ~n204 ;
  assign n206 = n198 & ~n205 ;
  assign n218 = ~n197 & ~n206 ;
  assign n207 = ~n65 & n187 ;
  assign n208 = \x_reg[1]/NET0131  & ~n207 ;
  assign n210 = \x_reg[0]/NET0131  & \y_reg[0]/NET0131  ;
  assign n211 = \x_reg[1]/NET0131  & \y_reg[1]/NET0131  ;
  assign n212 = ~\x_reg[1]/NET0131  & ~\y_reg[1]/NET0131  ;
  assign n213 = ~n211 & ~n212 ;
  assign n215 = n210 & n213 ;
  assign n209 = \stato_reg[0]/NET0131  & n181 ;
  assign n214 = ~n210 & ~n213 ;
  assign n216 = n209 & ~n214 ;
  assign n217 = ~n215 & n216 ;
  assign n219 = ~n208 & ~n217 ;
  assign n220 = n218 & n219 ;
  assign n224 = \mar_reg[1]/NET0131  & ~n184 ;
  assign n221 = ~\mar_reg[0]/NET0131  & ~\mar_reg[1]/NET0131  ;
  assign n222 = ~n58 & ~n221 ;
  assign n223 = ~n187 & n222 ;
  assign n225 = ~n189 & ~n223 ;
  assign n226 = ~n224 & n225 ;
  assign n230 = \mar_reg[2]/NET0131  & ~n184 ;
  assign n227 = ~\mar_reg[2]/NET0131  & ~n58 ;
  assign n228 = ~n59 & ~n227 ;
  assign n229 = ~n187 & n228 ;
  assign n231 = ~n189 & ~n229 ;
  assign n232 = ~n230 & n231 ;
  assign n237 = ~n193 & n207 ;
  assign n238 = \x_reg[0]/NET0131  & ~n237 ;
  assign n233 = ~\mar_reg[1]/NET0131  & ~\mar_reg[2]/NET0131  ;
  assign n234 = ~\mar_reg[3]/NET0131  & n233 ;
  assign n235 = ~n200 & ~n234 ;
  assign n236 = n198 & ~n235 ;
  assign n239 = ~\x_reg[0]/NET0131  & ~\y_reg[0]/NET0131  ;
  assign n240 = ~n210 & ~n239 ;
  assign n241 = n209 & n240 ;
  assign n242 = ~n236 & ~n241 ;
  assign n243 = ~n238 & n242 ;
  assign n244 = n193 & ~n205 ;
  assign n245 = \stato_reg[2]/NET0131  & ~n43 ;
  assign n246 = ~n209 & n245 ;
  assign n247 = \y_reg[1]/NET0131  & ~n246 ;
  assign n248 = ~n244 & ~n247 ;
  assign n249 = ~\stato_reg[0]/NET0131  & ~n68 ;
  assign n250 = n60 & n68 ;
  assign n251 = ~n65 & ~n250 ;
  assign n252 = ~start_pad & ~n251 ;
  assign n253 = ~n249 & ~n252 ;
  assign n254 = n68 & ~n95 ;
  assign n255 = ~n198 & ~n209 ;
  assign n256 = ~n93 & n255 ;
  assign n257 = ~n254 & n256 ;
  assign n258 = \x_reg[5]/NET0131  & n176 ;
  assign n259 = \stato_reg[1]/NET0131  & ~n44 ;
  assign n260 = ~n198 & n259 ;
  assign n261 = \t_reg[6]/NET0131  & ~n260 ;
  assign n262 = ~n258 & ~n261 ;
  assign n263 = \x_reg[4]/NET0131  & n176 ;
  assign n264 = \t_reg[5]/NET0131  & ~n260 ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = \mar_reg[0]/NET0131  & n234 ;
  assign n267 = ~n200 & ~n266 ;
  assign n268 = n193 & ~n267 ;
  assign n269 = \y_reg[2]/NET0131  & ~n246 ;
  assign n270 = ~n268 & ~n269 ;
  assign n271 = ~n201 & ~n266 ;
  assign n272 = n193 & ~n271 ;
  assign n273 = \y_reg[3]/NET0131  & ~n246 ;
  assign n274 = ~n272 & ~n273 ;
  assign n275 = start_pad & n250 ;
  assign n276 = ~n176 & ~n181 ;
  assign n277 = ~n275 & n276 ;
  assign n278 = \x_reg[0]/NET0131  & n176 ;
  assign n279 = \t_reg[1]/NET0131  & ~n260 ;
  assign n280 = ~n278 & ~n279 ;
  assign n281 = \x_reg[1]/NET0131  & n176 ;
  assign n282 = \t_reg[2]/NET0131  & ~n260 ;
  assign n283 = ~n281 & ~n282 ;
  assign n284 = \x_reg[2]/NET0131  & n176 ;
  assign n285 = \t_reg[3]/NET0131  & ~n260 ;
  assign n286 = ~n284 & ~n285 ;
  assign n287 = \x_reg[3]/NET0131  & n176 ;
  assign n288 = \t_reg[4]/NET0131  & ~n260 ;
  assign n289 = ~n287 & ~n288 ;
  assign n290 = n193 & ~n235 ;
  assign n291 = \y_reg[0]/NET0131  & ~n246 ;
  assign n292 = ~n290 & ~n291 ;
  assign n293 = \punti_retta[4]_pad  & ~n94 ;
  assign n296 = ~start_pad & n75 ;
  assign n295 = \punti_retta[4]_pad  & start_pad ;
  assign n297 = n60 & ~n295 ;
  assign n298 = ~n296 & n297 ;
  assign n294 = ~\punti_retta[4]_pad  & ~n60 ;
  assign n299 = n44 & ~n294 ;
  assign n300 = ~n298 & n299 ;
  assign n301 = ~n293 & ~n300 ;
  assign n304 = ~\x_reg[4]/NET0131  & ~\y_reg[3]/NET0131  ;
  assign n305 = \x_reg[2]/NET0131  & \y_reg[2]/NET0131  ;
  assign n306 = ~\x_reg[2]/NET0131  & ~\y_reg[2]/NET0131  ;
  assign n307 = ~n210 & ~n211 ;
  assign n308 = ~n212 & ~n307 ;
  assign n309 = ~n306 & n308 ;
  assign n310 = ~n305 & ~n309 ;
  assign n311 = ~\x_reg[3]/NET0131  & ~\y_reg[3]/NET0131  ;
  assign n312 = ~n310 & ~n311 ;
  assign n313 = ~n304 & n312 ;
  assign n302 = ~\x_reg[6]/NET0131  & ~\y_reg[3]/NET0131  ;
  assign n303 = ~\x_reg[5]/NET0131  & ~\y_reg[3]/NET0131  ;
  assign n314 = ~n302 & ~n303 ;
  assign n315 = n313 & n314 ;
  assign n317 = \x_reg[4]/NET0131  & \y_reg[3]/NET0131  ;
  assign n318 = \x_reg[3]/NET0131  & \y_reg[3]/NET0131  ;
  assign n319 = ~n317 & ~n318 ;
  assign n316 = \x_reg[5]/NET0131  & \y_reg[3]/NET0131  ;
  assign n320 = \x_reg[6]/NET0131  & \y_reg[3]/NET0131  ;
  assign n321 = ~n316 & ~n320 ;
  assign n322 = n319 & n321 ;
  assign n323 = ~n315 & n322 ;
  assign n324 = n209 & ~n323 ;
  assign n327 = ~\t_reg[5]/NET0131  & ~\x_reg[5]/NET0131  ;
  assign n328 = ~\t_reg[4]/NET0131  & ~\x_reg[4]/NET0131  ;
  assign n329 = ~\t_reg[2]/NET0131  & ~\x_reg[2]/NET0131  ;
  assign n330 = n194 & ~n329 ;
  assign n331 = \t_reg[2]/NET0131  & \x_reg[2]/NET0131  ;
  assign n332 = ~n330 & ~n331 ;
  assign n333 = ~\t_reg[3]/NET0131  & ~\x_reg[3]/NET0131  ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = \t_reg[3]/NET0131  & \x_reg[3]/NET0131  ;
  assign n336 = \t_reg[4]/NET0131  & \x_reg[4]/NET0131  ;
  assign n337 = ~n335 & ~n336 ;
  assign n338 = ~n334 & n337 ;
  assign n339 = ~n328 & ~n338 ;
  assign n340 = ~n327 & n339 ;
  assign n325 = \t_reg[6]/NET0131  & \x_reg[6]/NET0131  ;
  assign n326 = \t_reg[5]/NET0131  & \x_reg[5]/NET0131  ;
  assign n341 = ~n325 & ~n326 ;
  assign n342 = ~n340 & n341 ;
  assign n343 = ~\t_reg[6]/NET0131  & ~\x_reg[6]/NET0131  ;
  assign n344 = n193 & ~n343 ;
  assign n345 = ~n342 & n344 ;
  assign n346 = \x_reg[7]/NET0131  & ~n207 ;
  assign n347 = n198 & ~n271 ;
  assign n348 = ~n346 & ~n347 ;
  assign n349 = ~n345 & n348 ;
  assign n350 = ~n324 & n349 ;
  assign n358 = ~n305 & ~n306 ;
  assign n360 = n308 & n358 ;
  assign n359 = ~n308 & ~n358 ;
  assign n361 = n209 & ~n359 ;
  assign n362 = ~n360 & n361 ;
  assign n353 = ~n329 & ~n331 ;
  assign n355 = n194 & n353 ;
  assign n354 = ~n194 & ~n353 ;
  assign n356 = n193 & ~n354 ;
  assign n357 = ~n355 & n356 ;
  assign n351 = \x_reg[2]/NET0131  & ~n207 ;
  assign n352 = n198 & ~n267 ;
  assign n363 = ~n351 & ~n352 ;
  assign n364 = ~n357 & n363 ;
  assign n365 = ~n362 & n364 ;
  assign n372 = ~n311 & ~n318 ;
  assign n374 = ~n310 & n372 ;
  assign n373 = n310 & ~n372 ;
  assign n375 = n209 & ~n373 ;
  assign n376 = ~n374 & n375 ;
  assign n367 = ~n333 & ~n335 ;
  assign n369 = ~n332 & n367 ;
  assign n368 = n332 & ~n367 ;
  assign n370 = n193 & ~n368 ;
  assign n371 = ~n369 & n370 ;
  assign n366 = \x_reg[3]/NET0131  & ~n207 ;
  assign n377 = ~n347 & ~n366 ;
  assign n378 = ~n371 & n377 ;
  assign n379 = ~n376 & n378 ;
  assign n380 = ~n303 & ~n316 ;
  assign n381 = ~n313 & n319 ;
  assign n383 = ~n380 & n381 ;
  assign n382 = n380 & ~n381 ;
  assign n384 = n209 & ~n382 ;
  assign n385 = ~n383 & n384 ;
  assign n389 = ~n326 & n340 ;
  assign n387 = ~n326 & ~n327 ;
  assign n388 = ~n339 & ~n387 ;
  assign n390 = n193 & ~n388 ;
  assign n391 = ~n389 & n390 ;
  assign n386 = \x_reg[5]/NET0131  & ~n207 ;
  assign n392 = ~n347 & ~n386 ;
  assign n393 = ~n391 & n392 ;
  assign n394 = ~n385 & n393 ;
  assign n395 = ~start_pad & n88 ;
  assign n396 = \punti_retta[7]_pad  & start_pad ;
  assign n397 = n60 & ~n396 ;
  assign n398 = ~n395 & n397 ;
  assign n399 = ~\punti_retta[7]_pad  & ~n60 ;
  assign n400 = n44 & ~n399 ;
  assign n401 = ~n398 & n400 ;
  assign n402 = \punti_retta[7]_pad  & ~n94 ;
  assign n403 = ~n401 & ~n402 ;
  assign n417 = ~n304 & ~n311 ;
  assign n418 = n309 & n417 ;
  assign n419 = n305 & ~n311 ;
  assign n420 = n319 & ~n419 ;
  assign n421 = ~n304 & ~n420 ;
  assign n422 = ~n418 & ~n421 ;
  assign n423 = ~n303 & ~n422 ;
  assign n424 = ~n316 & ~n423 ;
  assign n425 = ~n302 & ~n320 ;
  assign n427 = n424 & ~n425 ;
  assign n426 = ~n424 & n425 ;
  assign n428 = n209 & ~n426 ;
  assign n429 = ~n427 & n428 ;
  assign n405 = ~n325 & ~n343 ;
  assign n406 = ~n331 & ~n335 ;
  assign n407 = ~n330 & n406 ;
  assign n408 = ~n333 & ~n407 ;
  assign n409 = ~n336 & ~n408 ;
  assign n410 = ~n327 & ~n328 ;
  assign n411 = ~n409 & n410 ;
  assign n412 = ~n326 & ~n411 ;
  assign n414 = ~n405 & n412 ;
  assign n413 = n405 & ~n412 ;
  assign n415 = n193 & ~n413 ;
  assign n416 = ~n414 & n415 ;
  assign n404 = \x_reg[6]/NET0131  & ~n207 ;
  assign n430 = ~n347 & ~n404 ;
  assign n431 = ~n416 & n430 ;
  assign n432 = ~n429 & n431 ;
  assign n433 = \punti_retta[3]_pad  & ~n94 ;
  assign n434 = ~start_pad & n110 ;
  assign n435 = \punti_retta[3]_pad  & start_pad ;
  assign n436 = n60 & ~n435 ;
  assign n437 = ~n434 & n436 ;
  assign n438 = ~\punti_retta[3]_pad  & ~n60 ;
  assign n439 = n44 & ~n438 ;
  assign n440 = ~n437 & n439 ;
  assign n441 = ~n433 & ~n440 ;
  assign n443 = ~n304 & ~n317 ;
  assign n444 = ~n312 & ~n318 ;
  assign n446 = n443 & ~n444 ;
  assign n445 = ~n443 & n444 ;
  assign n447 = n209 & ~n445 ;
  assign n448 = ~n446 & n447 ;
  assign n449 = ~n328 & ~n336 ;
  assign n451 = ~n408 & ~n449 ;
  assign n450 = n408 & n449 ;
  assign n452 = n193 & ~n450 ;
  assign n453 = ~n451 & n452 ;
  assign n442 = \x_reg[4]/NET0131  & ~n207 ;
  assign n454 = ~n347 & ~n442 ;
  assign n455 = ~n453 & n454 ;
  assign n456 = ~n448 & n455 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g2119/_0_  = n73 ;
  assign \g2123/_0_  = ~n81 ;
  assign \g2129/_0_  = ~n92 ;
  assign \g2133/_0_  = ~n103 ;
  assign \g2136/_0_  = ~n114 ;
  assign \g2140/_0_  = ~n125 ;
  assign \g2141/_0_  = ~n136 ;
  assign \g2151/_0_  = ~n144 ;
  assign \g2152/_0_  = ~n149 ;
  assign \g2166/_0_  = ~n155 ;
  assign \g2167/_0_  = ~n161 ;
  assign \g2180/_0_  = ~n168 ;
  assign \g2181/_0_  = ~n174 ;
  assign \g2199/_0_  = n186 ;
  assign \g2225/_0_  = ~n192 ;
  assign \g2227/_0_  = ~n220 ;
  assign \g2242/_0_  = ~n226 ;
  assign \g2243/_0_  = ~n232 ;
  assign \g2272/_0_  = ~n243 ;
  assign \g2273/_0_  = ~n248 ;
  assign \g2274/_0_  = ~n253 ;
  assign \g2275/_0_  = ~n257 ;
  assign \g2284/_0_  = ~n262 ;
  assign \g2289/_0_  = ~n265 ;
  assign \g2303/_0_  = ~n270 ;
  assign \g2304/_0_  = ~n274 ;
  assign \g2308/_0_  = ~n277 ;
  assign \g2309/_0_  = ~n280 ;
  assign \g2310/_0_  = ~n283 ;
  assign \g2311/_0_  = ~n286 ;
  assign \g2312/_0_  = ~n289 ;
  assign \g2346/_0_  = ~n292 ;
  assign \g2973/_0_  = ~n301 ;
  assign \g2984/_0_  = ~n350 ;
  assign \g3052/_0_  = ~n365 ;
  assign \g3176/_0_  = ~n379 ;
  assign \g3277/_0_  = ~n394 ;
  assign \g3306/_0_  = ~n403 ;
  assign \g3366/_0_  = ~n432 ;
  assign \g3371/_0_  = ~n441 ;
  assign \g3398/_0_  = ~n456 ;
endmodule
