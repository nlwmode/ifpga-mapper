module top (\g100_reg/NET0131 , \g1037_reg/NET0131 , \g103_reg/NET0131 , \g1041_reg/NET0131 , \g1045_reg/NET0131 , \g1049_reg/NET0131 , \g104_reg/NET0131 , \g1053_reg/NET0131 , \g1057_reg/NET0131 , \g1061_reg/NET0131 , \g1065_reg/NET0131 , \g1069_reg/NET0131 , \g1073_reg/NET0131 , \g1077_reg/NET0131 , \g1080_pad , \g1087_reg/NET0131 , \g1092_reg/NET0131 , \g1097_reg/NET0131 , \g1098_reg/NET0131 , \g1102_reg/NET0131 , \g1106_reg/NET0131 , \g1110_reg/NET0131 , \g1114_reg/NET0131 , \g1118_reg/NET0131 , \g1122_reg/NET0131 , \g1126_reg/NET0131 , \g1130_reg/NET0131 , \g1134_reg/NET0131 , \g1138_reg/NET0131 , \g1142_reg/NET0131 , \g1148_reg/NET0131 , \g1149_reg/NET0131 , \g1158_reg/NET0131 , \g1166_reg/NET0131 , \g1176_reg/NET0131 , \g1179_reg/NET0131 , \g1189_reg/NET0131 , \g1207_reg/NET0131 , \g1211_reg/NET0131 , \g1214_reg/NET0131 , \g1217_reg/NET0131 , \g1220_reg/NET0131 , \g1223_reg/NET0131 , \g1224_reg/NET0131 , \g1225_reg/NET0131 , \g1226_reg/NET0131 , \g1227_reg/NET0131 , \g1228_reg/NET0131 , \g1229_reg/NET0131 , \g1230_reg/NET0131 , \g1231_reg/NET0131 , \g1247_reg/NET0131 , \g1251_reg/NET0131 , \g1252_reg/NET0131 , \g1253_reg/NET0131 , \g1257_reg/NET0131 , \g1260_reg/NET0131 , \g1263_reg/NET0131 , \g1266_reg/NET0131 , \g1268_reg/NET0131 , \g1269_reg/NET0131 , \g1272_reg/NET0131 , \g1276_reg/NET0131 , \g1280_reg/NET0131 , \g1284_reg/NET0131 , \g1288_reg/NET0131 , \g1292_reg/NET0131 , \g1296_reg/NET0131 , \g1300_reg/NET0131 , \g1304_reg/NET0131 , \g1307_reg/NET0131 , \g1313_reg/NET0131 , \g1317_reg/NET0131 , \g1318_reg/NET0131 , \g1319_reg/NET0131 , \g1320_reg/NET0131 , \g1321_reg/NET0131 , \g1322_reg/NET0131 , \g1323_reg/NET0131 , \g1324_reg/NET0131 , \g1325_reg/NET0131 , \g1326_reg/NET0131 , \g1327_reg/NET0131 , \g1328_reg/NET0131 , \g1329_reg/NET0131 , \g1330_reg/NET0131 , \g1333_reg/NET0131 , \g1336_reg/NET0131 , \g1339_reg/NET0131 , \g1342_reg/NET0131 , \g1345_reg/NET0131 , \g1348_reg/NET0131 , \g1351_reg/NET0131 , \g1354_reg/NET0131 , \g1357_reg/NET0131 , \g1360_reg/NET0131 , \g1363_reg/NET0131 , \g1364_reg/NET0131 , \g1365_reg/NET0131 , \g1366_reg/NET0131 , \g1367_reg/NET0131 , \g1368_reg/NET0131 , \g1369_reg/NET0131 , \g1370_reg/NET0131 , \g1371_reg/NET0131 , \g1372_reg/NET0131 , \g1373_reg/NET0131 , \g1374_reg/NET0131 , \g1375_reg/NET0131 , \g1405_reg/NET0131 , \g1408_reg/NET0131 , \g1412_reg/NET0131 , \g1415_reg/NET0131 , \g1416_reg/NET0131 , \g1421_reg/NET0131 , \g1428_reg/NET0131 , \g1430_reg/NET0131 , \g1432_reg/NET0131 , \g1435_reg/NET0131 , \g1439_reg/NET0131 , \g1444_reg/NET0131 , \g1450_reg/NET0131 , \g1454_reg/NET0131 , \g1462_reg/NET0131 , \g1467_reg/NET0131 , \g1472_reg/NET0131 , \g1481_reg/NET0131 , \g1486_reg/NET0131 , \g1489_reg/NET0131 , \g1494_reg/NET0131 , \g1499_reg/NET0131 , \g1504_reg/NET0131 , \g1509_reg/NET0131 , \g1514_reg/NET0131 , \g1519_reg/NET0131 , \g1944_pad , \g2662_pad , \g2888_pad , \g2_reg/NET0131 , \g4370_pad , \g4371_pad , \g4372_pad , \g4373_pad , \g43_pad , \g652_reg/NET0131 , \g7423_pad , \g7424_pad , \g7425_pad , \g7504_pad , \g7505_pad , \g7507_pad , \g7508_pad , \g785_pad , \g866_reg/NET0131 , \g871_reg/NET0131 , \g889_reg/NET0131 , \g929_reg/NET0131 , \g933_reg/NET0131 , \g936_reg/NET0131 , \g940_reg/NET0131 , \g942_reg/NET0131 , \g943_reg/NET0131 , \g944_reg/NET0131 , \g950_reg/NET0131 , \g951_reg/NET0131 , \g952_reg/NET0131 , \g953_reg/NET0131 , \g954_reg/NET0131 , \g962_pad , \g1006_pad , \g1158_reg/P0001 , \g1252_reg/P0001 , \g1260_reg/P0001 , \g1416_reg/NET0131_syn_2 , \g17/_0_ , \g19189/_0_ , \g19252/_0_ , \g19253/_0_ , \g19273/_3_ , \g19284/_0_ , \g19285/_0_ , \g19295/_3_ , \g19302/_0_ , \g19303/_0_ , \g19304/_0_ , \g19308/_0_ , \g19309/_0_ , \g19310/_0_ , \g19321/_0_ , \g19326/_3_ , \g19331/_0_ , \g19341/_0_ , \g19366/_0_ , \g19372/_3_ , \g19385/_0_ , \g19386/_0_ , \g19387/_0_ , \g19388/_0_ , \g19389/_0_ , \g19390/_0_ , \g19392/_0_ , \g19393/_0_ , \g19394/_0_ , \g19398/_0_ , \g19399/_0_ , \g19400/_0_ , \g19401/_0_ , \g19403/_0_ , \g19405/_0_ , \g19406/_0_ , \g19437/_0_ , \g19438/_0_ , \g19445/_0_ , \g19446/_0_ , \g19450/_3_ , \g19472/_0_ , \g19473/_0_ , \g19474/_0_ , \g19476/_0_ , \g19484/_0_ , \g19485/_0_ , \g19492/_0_ , \g19493/_0_ , \g19499/_0_ , \g19500/_0_ , \g19501/_0_ , \g19502/_0_ , \g19503/_0_ , \g19504/_0_ , \g19507/_3_ , \g19508/_3_ , \g19512/_3_ , \g19513/_3_ , \g19514/_3_ , \g19528/_0_ , \g19529/_0_ , \g19534/_0_ , \g19535/_0_ , \g19536/_0_ , \g19538/_0_ , \g19542/_0_ , \g19560/_0_ , \g19563/_0_ , \g19565/_0_ , \g19567/_0_ , \g19569/_1_ , \g19572/_0_ , \g19574/_3_ , \g19614/_0_ , \g19615/_0_ , \g19620/_0_ , \g19626/_0_ , \g19629/_0_ , \g19631/_0_ , \g19666/_0_ , \g19667/_0_ , \g19669/_0_ , \g19677/_0_ , \g19690/_3_ , \g19721/_0_ , \g19723/_0_ , \g19723/_1_ , \g19725/_2_ , \g19751/_0_ , \g19752/_0_ , \g19753/_0_ , \g19755/_0_ , \g19815/_0_ , \g19821/_0_ , \g19822/_0_ , \g19833/_0_ , \g19877/_0_ , \g19898/_0_ , \g19899/_0_ , \g19900/_0_ , \g19901/_0_ , \g19908/_0_ , \g19927/_0_ , \g19928/_0_ , \g19930/_0_ , \g19931/_0_ , \g19932/_0_ , \g19934/_0_ , \g19992/_0_ , \g19993/_0_ , \g20002/_0_ , \g20008/_0_ , \g20010/_0_ , \g20016/_0_ , \g20110/_0_ , \g20117/_0_ , \g20118/_0_ , \g20131/_0_ , \g20246/_0_ , \g20704/_0_ , \g20722/_0_ , \g20731/_0_ , \g20732/_2_ , \g20870/_0_ , \g20883/_0_ , \g20931/_0_ , \g20951/_0_ , \g20969/_0_ , \g20989/_0_ , \g21/_2_ , \g21070/_0_ , \g21108/_0_ , \g21122/_0_ , \g21152/_0_ , \g21191/_0_ , \g21279/_0_ , \g21316/_0_ , \g21323/_0_ , \g21349/_3_ , \g21352/_3_ , \g21464/_0_ , \g21472/_0_ , \g21484/_0_ , \g21510/_0_ , \g21517/_0_ , \g21608/_0_ , \g21625/_0_ , \g21644/_1_ , \g4655_pad , \g6850_pad , \g6895_pad , \g7048_pad , \g7103_pad , \g7731_pad , \g7732_pad , \g8219_pad , \g8663_pad );
	input \g100_reg/NET0131  ;
	input \g1037_reg/NET0131  ;
	input \g103_reg/NET0131  ;
	input \g1041_reg/NET0131  ;
	input \g1045_reg/NET0131  ;
	input \g1049_reg/NET0131  ;
	input \g104_reg/NET0131  ;
	input \g1053_reg/NET0131  ;
	input \g1057_reg/NET0131  ;
	input \g1061_reg/NET0131  ;
	input \g1065_reg/NET0131  ;
	input \g1069_reg/NET0131  ;
	input \g1073_reg/NET0131  ;
	input \g1077_reg/NET0131  ;
	input \g1080_pad  ;
	input \g1087_reg/NET0131  ;
	input \g1092_reg/NET0131  ;
	input \g1097_reg/NET0131  ;
	input \g1098_reg/NET0131  ;
	input \g1102_reg/NET0131  ;
	input \g1106_reg/NET0131  ;
	input \g1110_reg/NET0131  ;
	input \g1114_reg/NET0131  ;
	input \g1118_reg/NET0131  ;
	input \g1122_reg/NET0131  ;
	input \g1126_reg/NET0131  ;
	input \g1130_reg/NET0131  ;
	input \g1134_reg/NET0131  ;
	input \g1138_reg/NET0131  ;
	input \g1142_reg/NET0131  ;
	input \g1148_reg/NET0131  ;
	input \g1149_reg/NET0131  ;
	input \g1158_reg/NET0131  ;
	input \g1166_reg/NET0131  ;
	input \g1176_reg/NET0131  ;
	input \g1179_reg/NET0131  ;
	input \g1189_reg/NET0131  ;
	input \g1207_reg/NET0131  ;
	input \g1211_reg/NET0131  ;
	input \g1214_reg/NET0131  ;
	input \g1217_reg/NET0131  ;
	input \g1220_reg/NET0131  ;
	input \g1223_reg/NET0131  ;
	input \g1224_reg/NET0131  ;
	input \g1225_reg/NET0131  ;
	input \g1226_reg/NET0131  ;
	input \g1227_reg/NET0131  ;
	input \g1228_reg/NET0131  ;
	input \g1229_reg/NET0131  ;
	input \g1230_reg/NET0131  ;
	input \g1231_reg/NET0131  ;
	input \g1247_reg/NET0131  ;
	input \g1251_reg/NET0131  ;
	input \g1252_reg/NET0131  ;
	input \g1253_reg/NET0131  ;
	input \g1257_reg/NET0131  ;
	input \g1260_reg/NET0131  ;
	input \g1263_reg/NET0131  ;
	input \g1266_reg/NET0131  ;
	input \g1268_reg/NET0131  ;
	input \g1269_reg/NET0131  ;
	input \g1272_reg/NET0131  ;
	input \g1276_reg/NET0131  ;
	input \g1280_reg/NET0131  ;
	input \g1284_reg/NET0131  ;
	input \g1288_reg/NET0131  ;
	input \g1292_reg/NET0131  ;
	input \g1296_reg/NET0131  ;
	input \g1300_reg/NET0131  ;
	input \g1304_reg/NET0131  ;
	input \g1307_reg/NET0131  ;
	input \g1313_reg/NET0131  ;
	input \g1317_reg/NET0131  ;
	input \g1318_reg/NET0131  ;
	input \g1319_reg/NET0131  ;
	input \g1320_reg/NET0131  ;
	input \g1321_reg/NET0131  ;
	input \g1322_reg/NET0131  ;
	input \g1323_reg/NET0131  ;
	input \g1324_reg/NET0131  ;
	input \g1325_reg/NET0131  ;
	input \g1326_reg/NET0131  ;
	input \g1327_reg/NET0131  ;
	input \g1328_reg/NET0131  ;
	input \g1329_reg/NET0131  ;
	input \g1330_reg/NET0131  ;
	input \g1333_reg/NET0131  ;
	input \g1336_reg/NET0131  ;
	input \g1339_reg/NET0131  ;
	input \g1342_reg/NET0131  ;
	input \g1345_reg/NET0131  ;
	input \g1348_reg/NET0131  ;
	input \g1351_reg/NET0131  ;
	input \g1354_reg/NET0131  ;
	input \g1357_reg/NET0131  ;
	input \g1360_reg/NET0131  ;
	input \g1363_reg/NET0131  ;
	input \g1364_reg/NET0131  ;
	input \g1365_reg/NET0131  ;
	input \g1366_reg/NET0131  ;
	input \g1367_reg/NET0131  ;
	input \g1368_reg/NET0131  ;
	input \g1369_reg/NET0131  ;
	input \g1370_reg/NET0131  ;
	input \g1371_reg/NET0131  ;
	input \g1372_reg/NET0131  ;
	input \g1373_reg/NET0131  ;
	input \g1374_reg/NET0131  ;
	input \g1375_reg/NET0131  ;
	input \g1405_reg/NET0131  ;
	input \g1408_reg/NET0131  ;
	input \g1412_reg/NET0131  ;
	input \g1415_reg/NET0131  ;
	input \g1416_reg/NET0131  ;
	input \g1421_reg/NET0131  ;
	input \g1428_reg/NET0131  ;
	input \g1430_reg/NET0131  ;
	input \g1432_reg/NET0131  ;
	input \g1435_reg/NET0131  ;
	input \g1439_reg/NET0131  ;
	input \g1444_reg/NET0131  ;
	input \g1450_reg/NET0131  ;
	input \g1454_reg/NET0131  ;
	input \g1462_reg/NET0131  ;
	input \g1467_reg/NET0131  ;
	input \g1472_reg/NET0131  ;
	input \g1481_reg/NET0131  ;
	input \g1486_reg/NET0131  ;
	input \g1489_reg/NET0131  ;
	input \g1494_reg/NET0131  ;
	input \g1499_reg/NET0131  ;
	input \g1504_reg/NET0131  ;
	input \g1509_reg/NET0131  ;
	input \g1514_reg/NET0131  ;
	input \g1519_reg/NET0131  ;
	input \g1944_pad  ;
	input \g2662_pad  ;
	input \g2888_pad  ;
	input \g2_reg/NET0131  ;
	input \g4370_pad  ;
	input \g4371_pad  ;
	input \g4372_pad  ;
	input \g4373_pad  ;
	input \g43_pad  ;
	input \g652_reg/NET0131  ;
	input \g7423_pad  ;
	input \g7424_pad  ;
	input \g7425_pad  ;
	input \g7504_pad  ;
	input \g7505_pad  ;
	input \g7507_pad  ;
	input \g7508_pad  ;
	input \g785_pad  ;
	input \g866_reg/NET0131  ;
	input \g871_reg/NET0131  ;
	input \g889_reg/NET0131  ;
	input \g929_reg/NET0131  ;
	input \g933_reg/NET0131  ;
	input \g936_reg/NET0131  ;
	input \g940_reg/NET0131  ;
	input \g942_reg/NET0131  ;
	input \g943_reg/NET0131  ;
	input \g944_reg/NET0131  ;
	input \g950_reg/NET0131  ;
	input \g951_reg/NET0131  ;
	input \g952_reg/NET0131  ;
	input \g953_reg/NET0131  ;
	input \g954_reg/NET0131  ;
	input \g962_pad  ;
	output \g1006_pad  ;
	output \g1158_reg/P0001  ;
	output \g1252_reg/P0001  ;
	output \g1260_reg/P0001  ;
	output \g1416_reg/NET0131_syn_2  ;
	output \g17/_0_  ;
	output \g19189/_0_  ;
	output \g19252/_0_  ;
	output \g19253/_0_  ;
	output \g19273/_3_  ;
	output \g19284/_0_  ;
	output \g19285/_0_  ;
	output \g19295/_3_  ;
	output \g19302/_0_  ;
	output \g19303/_0_  ;
	output \g19304/_0_  ;
	output \g19308/_0_  ;
	output \g19309/_0_  ;
	output \g19310/_0_  ;
	output \g19321/_0_  ;
	output \g19326/_3_  ;
	output \g19331/_0_  ;
	output \g19341/_0_  ;
	output \g19366/_0_  ;
	output \g19372/_3_  ;
	output \g19385/_0_  ;
	output \g19386/_0_  ;
	output \g19387/_0_  ;
	output \g19388/_0_  ;
	output \g19389/_0_  ;
	output \g19390/_0_  ;
	output \g19392/_0_  ;
	output \g19393/_0_  ;
	output \g19394/_0_  ;
	output \g19398/_0_  ;
	output \g19399/_0_  ;
	output \g19400/_0_  ;
	output \g19401/_0_  ;
	output \g19403/_0_  ;
	output \g19405/_0_  ;
	output \g19406/_0_  ;
	output \g19437/_0_  ;
	output \g19438/_0_  ;
	output \g19445/_0_  ;
	output \g19446/_0_  ;
	output \g19450/_3_  ;
	output \g19472/_0_  ;
	output \g19473/_0_  ;
	output \g19474/_0_  ;
	output \g19476/_0_  ;
	output \g19484/_0_  ;
	output \g19485/_0_  ;
	output \g19492/_0_  ;
	output \g19493/_0_  ;
	output \g19499/_0_  ;
	output \g19500/_0_  ;
	output \g19501/_0_  ;
	output \g19502/_0_  ;
	output \g19503/_0_  ;
	output \g19504/_0_  ;
	output \g19507/_3_  ;
	output \g19508/_3_  ;
	output \g19512/_3_  ;
	output \g19513/_3_  ;
	output \g19514/_3_  ;
	output \g19528/_0_  ;
	output \g19529/_0_  ;
	output \g19534/_0_  ;
	output \g19535/_0_  ;
	output \g19536/_0_  ;
	output \g19538/_0_  ;
	output \g19542/_0_  ;
	output \g19560/_0_  ;
	output \g19563/_0_  ;
	output \g19565/_0_  ;
	output \g19567/_0_  ;
	output \g19569/_1_  ;
	output \g19572/_0_  ;
	output \g19574/_3_  ;
	output \g19614/_0_  ;
	output \g19615/_0_  ;
	output \g19620/_0_  ;
	output \g19626/_0_  ;
	output \g19629/_0_  ;
	output \g19631/_0_  ;
	output \g19666/_0_  ;
	output \g19667/_0_  ;
	output \g19669/_0_  ;
	output \g19677/_0_  ;
	output \g19690/_3_  ;
	output \g19721/_0_  ;
	output \g19723/_0_  ;
	output \g19723/_1_  ;
	output \g19725/_2_  ;
	output \g19751/_0_  ;
	output \g19752/_0_  ;
	output \g19753/_0_  ;
	output \g19755/_0_  ;
	output \g19815/_0_  ;
	output \g19821/_0_  ;
	output \g19822/_0_  ;
	output \g19833/_0_  ;
	output \g19877/_0_  ;
	output \g19898/_0_  ;
	output \g19899/_0_  ;
	output \g19900/_0_  ;
	output \g19901/_0_  ;
	output \g19908/_0_  ;
	output \g19927/_0_  ;
	output \g19928/_0_  ;
	output \g19930/_0_  ;
	output \g19931/_0_  ;
	output \g19932/_0_  ;
	output \g19934/_0_  ;
	output \g19992/_0_  ;
	output \g19993/_0_  ;
	output \g20002/_0_  ;
	output \g20008/_0_  ;
	output \g20010/_0_  ;
	output \g20016/_0_  ;
	output \g20110/_0_  ;
	output \g20117/_0_  ;
	output \g20118/_0_  ;
	output \g20131/_0_  ;
	output \g20246/_0_  ;
	output \g20704/_0_  ;
	output \g20722/_0_  ;
	output \g20731/_0_  ;
	output \g20732/_2_  ;
	output \g20870/_0_  ;
	output \g20883/_0_  ;
	output \g20931/_0_  ;
	output \g20951/_0_  ;
	output \g20969/_0_  ;
	output \g20989/_0_  ;
	output \g21/_2_  ;
	output \g21070/_0_  ;
	output \g21108/_0_  ;
	output \g21122/_0_  ;
	output \g21152/_0_  ;
	output \g21191/_0_  ;
	output \g21279/_0_  ;
	output \g21316/_0_  ;
	output \g21323/_0_  ;
	output \g21349/_3_  ;
	output \g21352/_3_  ;
	output \g21464/_0_  ;
	output \g21472/_0_  ;
	output \g21484/_0_  ;
	output \g21510/_0_  ;
	output \g21517/_0_  ;
	output \g21608/_0_  ;
	output \g21625/_0_  ;
	output \g21644/_1_  ;
	output \g4655_pad  ;
	output \g6850_pad  ;
	output \g6895_pad  ;
	output \g7048_pad  ;
	output \g7103_pad  ;
	output \g7731_pad  ;
	output \g7732_pad  ;
	output \g8219_pad  ;
	output \g8663_pad  ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w292_ ;
	wire _w35_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w194_ ;
	wire _w262_ ;
	wire _w135_ ;
	wire _w392_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w193_ ;
	wire _w188_ ;
	wire _w61_ ;
	wire _w318_ ;
	wire _w246_ ;
	wire _w119_ ;
	wire _w376_ ;
	wire _w195_ ;
	wire _w293_ ;
	wire _w166_ ;
	wire _w423_ ;
	wire _w225_ ;
	wire _w184_ ;
	wire _w57_ ;
	wire _w314_ ;
	wire _w173_ ;
	wire _w289_ ;
	wire _w212_ ;
	wire _w180_ ;
	wire _w279_ ;
	wire _w152_ ;
	wire _w409_ ;
	wire _w211_ ;
	wire _w181_ ;
	wire _w251_ ;
	wire _w124_ ;
	wire _w381_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\g1158_reg/NET0131 ,
		_w35_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\g1252_reg/NET0131 ,
		_w57_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\g1260_reg/NET0131 ,
		_w61_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\g1416_reg/NET0131 ,
		_w119_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\g1432_reg/NET0131 ,
		_w124_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\g1486_reg/NET0131 ,
		_w135_
	);
	LUT1 #(
		.INIT('h1)
	) name6 (
		\g43_pad ,
		_w152_
	);
	LUT1 #(
		.INIT('h1)
	) name7 (
		\g929_reg/NET0131 ,
		_w166_
	);
	LUT1 #(
		.INIT('h1)
	) name8 (
		\g944_reg/NET0131 ,
		_w173_
	);
	LUT3 #(
		.INIT('h80)
	) name9 (
		\g1330_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1336_reg/NET0131 ,
		_w180_
	);
	LUT4 #(
		.INIT('h8000)
	) name10 (
		\g1330_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1336_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w181_
	);
	LUT3 #(
		.INIT('h80)
	) name11 (
		\g1342_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w181_,
		_w182_
	);
	LUT4 #(
		.INIT('h8000)
	) name12 (
		\g1342_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g1348_reg/NET0131 ,
		_w181_,
		_w183_
	);
	LUT3 #(
		.INIT('h28)
	) name13 (
		\g1247_reg/NET0131 ,
		\g1348_reg/NET0131 ,
		_w182_,
		_w184_
	);
	LUT2 #(
		.INIT('h2)
	) name14 (
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		_w185_
	);
	LUT3 #(
		.INIT('h04)
	) name15 (
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\g1092_reg/NET0131 ,
		\g1130_reg/NET0131 ,
		_w187_
	);
	LUT3 #(
		.INIT('h80)
	) name17 (
		\g1092_reg/NET0131 ,
		\g1130_reg/NET0131 ,
		\g1134_reg/NET0131 ,
		_w188_
	);
	LUT4 #(
		.INIT('h8000)
	) name18 (
		\g1092_reg/NET0131 ,
		\g1130_reg/NET0131 ,
		\g1134_reg/NET0131 ,
		\g1138_reg/NET0131 ,
		_w189_
	);
	LUT3 #(
		.INIT('h80)
	) name19 (
		\g1037_reg/NET0131 ,
		\g1041_reg/NET0131 ,
		\g1045_reg/NET0131 ,
		_w190_
	);
	LUT3 #(
		.INIT('h80)
	) name20 (
		\g1149_reg/NET0131 ,
		_w189_,
		_w190_,
		_w191_
	);
	LUT4 #(
		.INIT('h8000)
	) name21 (
		\g1049_reg/NET0131 ,
		\g1053_reg/NET0131 ,
		\g1057_reg/NET0131 ,
		\g1061_reg/NET0131 ,
		_w192_
	);
	LUT4 #(
		.INIT('h8000)
	) name22 (
		\g1149_reg/NET0131 ,
		_w189_,
		_w190_,
		_w192_,
		_w193_
	);
	LUT4 #(
		.INIT('h8000)
	) name23 (
		\g1065_reg/NET0131 ,
		\g1069_reg/NET0131 ,
		_w186_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('he)
	) name24 (
		_w185_,
		_w194_,
		_w195_
	);
	LUT3 #(
		.INIT('h26)
	) name25 (
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		\g943_reg/NET0131 ,
		_w196_
	);
	LUT3 #(
		.INIT('h73)
	) name26 (
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w197_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name27 (
		\g1049_reg/NET0131 ,
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w198_
	);
	LUT4 #(
		.INIT('h8000)
	) name28 (
		\g1049_reg/NET0131 ,
		\g1149_reg/NET0131 ,
		_w189_,
		_w190_,
		_w199_
	);
	LUT4 #(
		.INIT('hff48)
	) name29 (
		\g1049_reg/NET0131 ,
		_w186_,
		_w191_,
		_w198_,
		_w200_
	);
	LUT4 #(
		.INIT('hfb08)
	) name30 (
		\g2_reg/NET0131 ,
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		\g954_reg/NET0131 ,
		_w201_
	);
	LUT4 #(
		.INIT('h4000)
	) name31 (
		\g1251_reg/NET0131 ,
		\g1481_reg/NET0131 ,
		\g1489_reg/NET0131 ,
		\g1494_reg/NET0131 ,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\g1499_reg/NET0131 ,
		\g1504_reg/NET0131 ,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w202_,
		_w203_,
		_w204_
	);
	LUT3 #(
		.INIT('h80)
	) name34 (
		\g1509_reg/NET0131 ,
		_w202_,
		_w203_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\g1514_reg/NET0131 ,
		\g1519_reg/NET0131 ,
		_w206_
	);
	LUT4 #(
		.INIT('h8000)
	) name36 (
		\g1462_reg/NET0131 ,
		\g1467_reg/NET0131 ,
		\g1472_reg/NET0131 ,
		\g1499_reg/NET0131 ,
		_w207_
	);
	LUT3 #(
		.INIT('h80)
	) name37 (
		_w202_,
		_w206_,
		_w207_,
		_w208_
	);
	LUT3 #(
		.INIT('h12)
	) name38 (
		\g1514_reg/NET0131 ,
		_w208_,
		_w205_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\g1087_reg/NET0131 ,
		\g1098_reg/NET0131 ,
		_w210_
	);
	LUT3 #(
		.INIT('h80)
	) name40 (
		\g1087_reg/NET0131 ,
		\g1098_reg/NET0131 ,
		\g1102_reg/NET0131 ,
		_w211_
	);
	LUT4 #(
		.INIT('h8000)
	) name41 (
		\g1087_reg/NET0131 ,
		\g1098_reg/NET0131 ,
		\g1102_reg/NET0131 ,
		\g1106_reg/NET0131 ,
		_w212_
	);
	LUT3 #(
		.INIT('h80)
	) name42 (
		\g1110_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w212_,
		_w213_
	);
	LUT4 #(
		.INIT('h8000)
	) name43 (
		\g1110_reg/NET0131 ,
		\g1114_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w212_,
		_w214_
	);
	LUT3 #(
		.INIT('hbe)
	) name44 (
		\g1097_reg/NET0131 ,
		\g1118_reg/NET0131 ,
		_w214_,
		_w215_
	);
	LUT4 #(
		.INIT('hfb08)
	) name45 (
		\g2_reg/NET0131 ,
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		\g953_reg/NET0131 ,
		_w216_
	);
	LUT4 #(
		.INIT('hbeee)
	) name46 (
		\g1097_reg/NET0131 ,
		\g1106_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w211_,
		_w217_
	);
	LUT4 #(
		.INIT('hbeee)
	) name47 (
		\g1097_reg/NET0131 ,
		\g1110_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w212_,
		_w218_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name48 (
		\g1110_reg/NET0131 ,
		\g1114_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w212_,
		_w219_
	);
	LUT2 #(
		.INIT('he)
	) name49 (
		\g1097_reg/NET0131 ,
		_w219_,
		_w220_
	);
	LUT3 #(
		.INIT('h12)
	) name50 (
		\g1509_reg/NET0131 ,
		_w208_,
		_w204_,
		_w221_
	);
	LUT4 #(
		.INIT('h1230)
	) name51 (
		\g1087_reg/NET0131 ,
		\g1097_reg/NET0131 ,
		\g1098_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w222_
	);
	LUT4 #(
		.INIT('h1444)
	) name52 (
		\g1097_reg/NET0131 ,
		\g1102_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w210_,
		_w223_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name53 (
		\g1037_reg/NET0131 ,
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w224_
	);
	LUT3 #(
		.INIT('h80)
	) name54 (
		\g1037_reg/NET0131 ,
		\g1149_reg/NET0131 ,
		_w189_,
		_w225_
	);
	LUT4 #(
		.INIT('h60a0)
	) name55 (
		\g1037_reg/NET0131 ,
		\g1149_reg/NET0131 ,
		_w186_,
		_w189_,
		_w226_
	);
	LUT2 #(
		.INIT('he)
	) name56 (
		_w224_,
		_w226_,
		_w227_
	);
	LUT4 #(
		.INIT('hfb08)
	) name57 (
		\g2_reg/NET0131 ,
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		\g952_reg/NET0131 ,
		_w228_
	);
	LUT3 #(
		.INIT('h12)
	) name58 (
		\g1087_reg/NET0131 ,
		\g1097_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w229_
	);
	LUT3 #(
		.INIT('h13)
	) name59 (
		\g1499_reg/NET0131 ,
		\g1504_reg/NET0131 ,
		_w202_,
		_w230_
	);
	LUT4 #(
		.INIT('h557f)
	) name60 (
		_w202_,
		_w206_,
		_w207_,
		_w203_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w230_,
		_w231_,
		_w232_
	);
	LUT4 #(
		.INIT('h4c0c)
	) name62 (
		\g1073_reg/NET0131 ,
		\g1149_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w233_
	);
	LUT4 #(
		.INIT('hff48)
	) name63 (
		\g1149_reg/NET0131 ,
		_w186_,
		_w189_,
		_w233_,
		_w234_
	);
	LUT4 #(
		.INIT('hfb08)
	) name64 (
		\g2_reg/NET0131 ,
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		\g951_reg/NET0131 ,
		_w235_
	);
	LUT4 #(
		.INIT('h4c1c)
	) name65 (
		\g1073_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\g100_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w237_
	);
	LUT4 #(
		.INIT('h0078)
	) name67 (
		\g1313_reg/NET0131 ,
		\g1317_reg/NET0131 ,
		\g1318_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w238_
	);
	LUT2 #(
		.INIT('he)
	) name68 (
		_w237_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h9)
	) name69 (
		\g1251_reg/NET0131 ,
		\g1481_reg/NET0131 ,
		_w240_
	);
	LUT3 #(
		.INIT('hb4)
	) name70 (
		\g1251_reg/NET0131 ,
		\g1481_reg/NET0131 ,
		\g1489_reg/NET0131 ,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\g103_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w242_
	);
	LUT4 #(
		.INIT('h8000)
	) name72 (
		\g1313_reg/NET0131 ,
		\g1317_reg/NET0131 ,
		\g1318_reg/NET0131 ,
		\g1319_reg/NET0131 ,
		_w243_
	);
	LUT3 #(
		.INIT('h80)
	) name73 (
		\g1320_reg/NET0131 ,
		\g1321_reg/NET0131 ,
		\g1322_reg/NET0131 ,
		_w244_
	);
	LUT3 #(
		.INIT('h80)
	) name74 (
		\g1323_reg/NET0131 ,
		_w243_,
		_w244_,
		_w245_
	);
	LUT4 #(
		.INIT('h8000)
	) name75 (
		\g1323_reg/NET0131 ,
		\g1324_reg/NET0131 ,
		_w243_,
		_w244_,
		_w246_
	);
	LUT4 #(
		.INIT('ha3ac)
	) name76 (
		\g103_reg/NET0131 ,
		\g1324_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w245_,
		_w247_
	);
	LUT4 #(
		.INIT('h8000)
	) name77 (
		\g1342_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g1348_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		_w248_
	);
	LUT4 #(
		.INIT('h2888)
	) name78 (
		\g1247_reg/NET0131 ,
		\g1354_reg/NET0131 ,
		_w181_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\g1363_reg/NET0131 ,
		\g1364_reg/NET0131 ,
		_w250_
	);
	LUT4 #(
		.INIT('h0001)
	) name80 (
		\g1365_reg/NET0131 ,
		\g1366_reg/NET0131 ,
		\g1367_reg/NET0131 ,
		\g1368_reg/NET0131 ,
		_w251_
	);
	LUT3 #(
		.INIT('h01)
	) name81 (
		\g1373_reg/NET0131 ,
		\g1374_reg/NET0131 ,
		\g1375_reg/NET0131 ,
		_w252_
	);
	LUT4 #(
		.INIT('h0001)
	) name82 (
		\g1369_reg/NET0131 ,
		\g1370_reg/NET0131 ,
		\g1371_reg/NET0131 ,
		\g1372_reg/NET0131 ,
		_w253_
	);
	LUT4 #(
		.INIT('h8000)
	) name83 (
		_w250_,
		_w252_,
		_w253_,
		_w251_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\g1325_reg/NET0131 ,
		\g1326_reg/NET0131 ,
		_w255_
	);
	LUT3 #(
		.INIT('h80)
	) name85 (
		\g1325_reg/NET0131 ,
		\g1326_reg/NET0131 ,
		\g1327_reg/NET0131 ,
		_w256_
	);
	LUT4 #(
		.INIT('h1333)
	) name86 (
		\g1328_reg/NET0131 ,
		\g7504_pad ,
		_w246_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\g1329_reg/NET0131 ,
		_w257_,
		_w258_
	);
	LUT3 #(
		.INIT('h80)
	) name88 (
		\g871_reg/NET0131 ,
		\g929_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w259_
	);
	LUT4 #(
		.INIT('h2000)
	) name89 (
		\g871_reg/NET0131 ,
		\g889_reg/NET0131 ,
		\g929_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		\g785_pad ,
		_w260_,
		_w261_
	);
	LUT4 #(
		.INIT('h040c)
	) name91 (
		\g1325_reg/NET0131 ,
		\g1326_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w246_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\g1326_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w263_
	);
	LUT4 #(
		.INIT('h1333)
	) name93 (
		\g1325_reg/NET0131 ,
		_w242_,
		_w246_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('hb)
	) name94 (
		_w262_,
		_w264_,
		_w265_
	);
	LUT4 #(
		.INIT('h4c0c)
	) name95 (
		\g1073_reg/NET0131 ,
		\g1134_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w266_
	);
	LUT4 #(
		.INIT('hff48)
	) name96 (
		\g1134_reg/NET0131 ,
		_w186_,
		_w187_,
		_w266_,
		_w267_
	);
	LUT4 #(
		.INIT('h060c)
	) name97 (
		\g1320_reg/NET0131 ,
		\g1321_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w243_,
		_w268_
	);
	LUT2 #(
		.INIT('he)
	) name98 (
		_w237_,
		_w268_,
		_w269_
	);
	LUT4 #(
		.INIT('h4c0c)
	) name99 (
		\g1073_reg/NET0131 ,
		\g1138_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w270_
	);
	LUT4 #(
		.INIT('hff48)
	) name100 (
		\g1138_reg/NET0131 ,
		_w186_,
		_w188_,
		_w270_,
		_w271_
	);
	LUT4 #(
		.INIT('h4c0c)
	) name101 (
		\g1073_reg/NET0131 ,
		\g1130_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w272_
	);
	LUT2 #(
		.INIT('h6)
	) name102 (
		\g1092_reg/NET0131 ,
		\g1130_reg/NET0131 ,
		_w273_
	);
	LUT3 #(
		.INIT('hec)
	) name103 (
		_w186_,
		_w272_,
		_w273_,
		_w274_
	);
	LUT4 #(
		.INIT('h0015)
	) name104 (
		\g1231_reg/NET0131 ,
		\g1405_reg/NET0131 ,
		\g1408_reg/NET0131 ,
		\g1428_reg/NET0131 ,
		_w275_
	);
	LUT4 #(
		.INIT('h0015)
	) name105 (
		\g1231_reg/NET0131 ,
		\g1412_reg/NET0131 ,
		\g1415_reg/NET0131 ,
		\g1430_reg/NET0131 ,
		_w276_
	);
	LUT3 #(
		.INIT('h80)
	) name106 (
		\g1272_reg/NET0131 ,
		\g1276_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w277_
	);
	LUT4 #(
		.INIT('h8000)
	) name107 (
		\g1272_reg/NET0131 ,
		\g1276_reg/NET0131 ,
		\g1280_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w278_
	);
	LUT3 #(
		.INIT('h12)
	) name108 (
		\g1280_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		_w277_,
		_w279_
	);
	LUT4 #(
		.INIT('h8000)
	) name109 (
		\g1272_reg/NET0131 ,
		\g1276_reg/NET0131 ,
		\g1280_reg/NET0131 ,
		\g1284_reg/NET0131 ,
		_w280_
	);
	LUT3 #(
		.INIT('h80)
	) name110 (
		\g1288_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w280_,
		_w281_
	);
	LUT4 #(
		.INIT('h8000)
	) name111 (
		\g1288_reg/NET0131 ,
		\g1292_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w280_,
		_w282_
	);
	LUT3 #(
		.INIT('h12)
	) name112 (
		\g1292_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		_w281_,
		_w283_
	);
	LUT4 #(
		.INIT('h060a)
	) name113 (
		\g1296_reg/NET0131 ,
		\g1300_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		_w282_,
		_w284_
	);
	LUT3 #(
		.INIT('h12)
	) name114 (
		\g1300_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		_w282_,
		_w285_
	);
	LUT4 #(
		.INIT('h060c)
	) name115 (
		\g1272_reg/NET0131 ,
		\g1276_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w286_
	);
	LUT4 #(
		.INIT('hefaf)
	) name116 (
		\g1430_reg/NET0131 ,
		\g1432_reg/NET0131 ,
		\g1435_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		_w287_
	);
	LUT4 #(
		.INIT('h0150)
	) name117 (
		\g1430_reg/NET0131 ,
		\g1432_reg/NET0131 ,
		\g1435_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		_w288_
	);
	LUT3 #(
		.INIT('h08)
	) name118 (
		\g1432_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		\g7507_pad ,
		_w289_
	);
	LUT4 #(
		.INIT('hbfea)
	) name119 (
		\g1430_reg/NET0131 ,
		\g1432_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		\g7507_pad ,
		_w290_
	);
	LUT4 #(
		.INIT('h1044)
	) name120 (
		\g1430_reg/NET0131 ,
		\g1432_reg/NET0131 ,
		\g1435_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\g1284_reg/NET0131 ,
		_w278_,
		_w292_
	);
	LUT3 #(
		.INIT('h15)
	) name122 (
		\g1304_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w280_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		_w292_,
		_w293_,
		_w294_
	);
	LUT3 #(
		.INIT('h6a)
	) name124 (
		\g1288_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w280_,
		_w295_
	);
	LUT4 #(
		.INIT('h8000)
	) name125 (
		\g1288_reg/NET0131 ,
		\g1292_reg/NET0131 ,
		\g1296_reg/NET0131 ,
		\g1300_reg/NET0131 ,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		\g1304_reg/NET0131 ,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('hb)
	) name127 (
		_w295_,
		_w297_,
		_w298_
	);
	LUT3 #(
		.INIT('h80)
	) name128 (
		\g1207_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w299_
	);
	LUT4 #(
		.INIT('h8000)
	) name129 (
		\g1207_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		\g1217_reg/NET0131 ,
		_w300_
	);
	LUT4 #(
		.INIT('hf6fc)
	) name130 (
		\g1220_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		\g1231_reg/NET0131 ,
		_w300_,
		_w301_
	);
	LUT3 #(
		.INIT('h12)
	) name131 (
		\g1272_reg/NET0131 ,
		\g1304_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w302_
	);
	LUT3 #(
		.INIT('ha3)
	) name132 (
		\g100_reg/NET0131 ,
		\g1313_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w303_
	);
	LUT4 #(
		.INIT('h070f)
	) name133 (
		\g1320_reg/NET0131 ,
		\g1321_reg/NET0131 ,
		\g1322_reg/NET0131 ,
		_w243_,
		_w304_
	);
	LUT3 #(
		.INIT('h15)
	) name134 (
		\g1329_reg/NET0131 ,
		_w243_,
		_w244_,
		_w305_
	);
	LUT3 #(
		.INIT('hba)
	) name135 (
		_w237_,
		_w304_,
		_w305_,
		_w306_
	);
	LUT4 #(
		.INIT('h1222)
	) name136 (
		\g1323_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w243_,
		_w244_,
		_w307_
	);
	LUT2 #(
		.INIT('he)
	) name137 (
		_w237_,
		_w307_,
		_w308_
	);
	LUT4 #(
		.INIT('ha3ac)
	) name138 (
		\g103_reg/NET0131 ,
		\g1325_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w246_,
		_w309_
	);
	LUT4 #(
		.INIT('h007f)
	) name139 (
		\g1313_reg/NET0131 ,
		\g1317_reg/NET0131 ,
		\g1318_reg/NET0131 ,
		\g1319_reg/NET0131 ,
		_w310_
	);
	LUT4 #(
		.INIT('h888b)
	) name140 (
		\g100_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w243_,
		_w310_,
		_w311_
	);
	LUT4 #(
		.INIT('h1222)
	) name141 (
		\g1327_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w246_,
		_w255_,
		_w312_
	);
	LUT2 #(
		.INIT('he)
	) name142 (
		_w242_,
		_w312_,
		_w313_
	);
	LUT4 #(
		.INIT('hbf40)
	) name143 (
		\g1251_reg/NET0131 ,
		\g1481_reg/NET0131 ,
		\g1489_reg/NET0131 ,
		\g1494_reg/NET0131 ,
		_w314_
	);
	LUT2 #(
		.INIT('h6)
	) name144 (
		\g1499_reg/NET0131 ,
		_w202_,
		_w315_
	);
	LUT4 #(
		.INIT('haa3c)
	) name145 (
		\g100_reg/NET0131 ,
		\g1313_reg/NET0131 ,
		\g1317_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w316_
	);
	LUT4 #(
		.INIT('hfb08)
	) name146 (
		\g2_reg/NET0131 ,
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		\g950_reg/NET0131 ,
		_w317_
	);
	LUT4 #(
		.INIT('ha3ac)
	) name147 (
		\g100_reg/NET0131 ,
		\g1320_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w243_,
		_w318_
	);
	LUT4 #(
		.INIT('hfbbb)
	) name148 (
		\g1307_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		\g1450_reg/NET0131 ,
		\g1454_reg/NET0131 ,
		_w319_
	);
	LUT3 #(
		.INIT('h04)
	) name149 (
		\g1444_reg/NET0131 ,
		\g1450_reg/NET0131 ,
		\g1454_reg/NET0131 ,
		_w320_
	);
	LUT4 #(
		.INIT('h0414)
	) name150 (
		\g1307_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		\g1450_reg/NET0131 ,
		\g1454_reg/NET0131 ,
		_w321_
	);
	LUT3 #(
		.INIT('hfe)
	) name151 (
		\g1231_reg/NET0131 ,
		\g1405_reg/NET0131 ,
		\g1428_reg/NET0131 ,
		_w322_
	);
	LUT3 #(
		.INIT('hfe)
	) name152 (
		\g1231_reg/NET0131 ,
		\g1412_reg/NET0131 ,
		\g1430_reg/NET0131 ,
		_w323_
	);
	LUT3 #(
		.INIT('h04)
	) name153 (
		\g1307_reg/NET0131 ,
		\g1416_reg/NET0131 ,
		\g1421_reg/NET0131 ,
		_w324_
	);
	LUT4 #(
		.INIT('h0540)
	) name154 (
		\g1307_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		\g1450_reg/NET0131 ,
		\g1454_reg/NET0131 ,
		_w325_
	);
	LUT3 #(
		.INIT('hbe)
	) name155 (
		\g1430_reg/NET0131 ,
		\g7508_pad ,
		_w289_,
		_w326_
	);
	LUT3 #(
		.INIT('h01)
	) name156 (
		\g1354_reg/NET0131 ,
		\g1357_reg/NET0131 ,
		\g1360_reg/NET0131 ,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		\g104_reg/NET0131 ,
		\g1336_reg/NET0131 ,
		_w328_
	);
	LUT4 #(
		.INIT('h0001)
	) name158 (
		\g1342_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g1348_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		_w329_
	);
	LUT3 #(
		.INIT('h80)
	) name159 (
		_w328_,
		_w327_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\g1354_reg/NET0131 ,
		\g1357_reg/NET0131 ,
		_w331_
	);
	LUT3 #(
		.INIT('h80)
	) name161 (
		\g104_reg/NET0131 ,
		\g1336_reg/NET0131 ,
		\g1360_reg/NET0131 ,
		_w332_
	);
	LUT3 #(
		.INIT('h80)
	) name162 (
		_w248_,
		_w331_,
		_w332_,
		_w333_
	);
	LUT4 #(
		.INIT('h8001)
	) name163 (
		\g104_reg/NET0131 ,
		\g1330_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w334_
	);
	LUT3 #(
		.INIT('h1f)
	) name164 (
		_w330_,
		_w333_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\g1077_reg/NET0131 ,
		\g2888_pad ,
		_w336_
	);
	LUT3 #(
		.INIT('h80)
	) name166 (
		\g1158_reg/NET0131 ,
		\g1176_reg/NET0131 ,
		\g652_reg/NET0131 ,
		_w337_
	);
	LUT2 #(
		.INIT('he)
	) name167 (
		_w336_,
		_w337_,
		_w338_
	);
	LUT3 #(
		.INIT('h28)
	) name168 (
		\g1247_reg/NET0131 ,
		\g1330_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		_w339_
	);
	LUT3 #(
		.INIT('h2a)
	) name169 (
		\g1247_reg/NET0131 ,
		_w181_,
		_w248_,
		_w340_
	);
	LUT3 #(
		.INIT('he0)
	) name170 (
		\g1351_reg/NET0131 ,
		_w183_,
		_w340_,
		_w341_
	);
	LUT3 #(
		.INIT('h40)
	) name171 (
		\g785_pad ,
		\g866_reg/NET0131 ,
		\g889_reg/NET0131 ,
		_w342_
	);
	LUT4 #(
		.INIT('h870f)
	) name172 (
		\g1158_reg/NET0131 ,
		\g1179_reg/NET0131 ,
		\g2888_pad ,
		\g652_reg/NET0131 ,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w336_,
		_w343_,
		_w344_
	);
	LUT3 #(
		.INIT('h3a)
	) name174 (
		\g1080_pad ,
		\g1176_reg/NET0131 ,
		\g1944_pad ,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		\g1223_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		_w346_
	);
	LUT3 #(
		.INIT('h80)
	) name176 (
		\g1220_reg/NET0131 ,
		_w300_,
		_w346_,
		_w347_
	);
	LUT4 #(
		.INIT('h78f0)
	) name177 (
		\g1220_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		_w300_,
		_w348_
	);
	LUT2 #(
		.INIT('he)
	) name178 (
		\g1231_reg/NET0131 ,
		_w348_,
		_w349_
	);
	LUT4 #(
		.INIT('h0201)
	) name179 (
		\g104_reg/NET0131 ,
		\g1330_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w350_
	);
	LUT3 #(
		.INIT('h1f)
	) name180 (
		_w330_,
		_w333_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		\g1257_reg/NET0131 ,
		\g1263_reg/NET0131 ,
		_w352_
	);
	LUT3 #(
		.INIT('h80)
	) name182 (
		\g1223_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		\g1225_reg/NET0131 ,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		\g1227_reg/NET0131 ,
		\g1228_reg/NET0131 ,
		_w354_
	);
	LUT3 #(
		.INIT('h20)
	) name184 (
		\g1226_reg/NET0131 ,
		\g1229_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		_w355_
	);
	LUT4 #(
		.INIT('h4000)
	) name185 (
		_w352_,
		_w353_,
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		\g1247_reg/NET0131 ,
		_w356_,
		_w357_
	);
	LUT3 #(
		.INIT('h3b)
	) name187 (
		\g1247_reg/NET0131 ,
		\g1253_reg/NET0131 ,
		_w356_,
		_w358_
	);
	LUT3 #(
		.INIT('h28)
	) name188 (
		\g1247_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w180_,
		_w359_
	);
	LUT3 #(
		.INIT('hde)
	) name189 (
		\g1220_reg/NET0131 ,
		\g1231_reg/NET0131 ,
		_w300_,
		_w360_
	);
	LUT3 #(
		.INIT('hab)
	) name190 (
		\g1307_reg/NET0131 ,
		\g1416_reg/NET0131 ,
		\g1421_reg/NET0131 ,
		_w361_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		\g1247_reg/NET0131 ,
		\g1330_reg/NET0131 ,
		_w362_
	);
	LUT4 #(
		.INIT('h2a80)
	) name192 (
		\g1247_reg/NET0131 ,
		\g1330_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1336_reg/NET0131 ,
		_w363_
	);
	LUT3 #(
		.INIT('h28)
	) name193 (
		\g1247_reg/NET0131 ,
		\g1342_reg/NET0131 ,
		_w181_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w280_,
		_w296_,
		_w365_
	);
	LUT3 #(
		.INIT('h80)
	) name195 (
		\g104_reg/NET0131 ,
		_w280_,
		_w296_,
		_w366_
	);
	LUT3 #(
		.INIT('h01)
	) name196 (
		\g1292_reg/NET0131 ,
		\g1296_reg/NET0131 ,
		\g1300_reg/NET0131 ,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		\g104_reg/NET0131 ,
		\g1272_reg/NET0131 ,
		_w368_
	);
	LUT4 #(
		.INIT('h0001)
	) name198 (
		\g1276_reg/NET0131 ,
		\g1280_reg/NET0131 ,
		\g1284_reg/NET0131 ,
		\g1288_reg/NET0131 ,
		_w369_
	);
	LUT3 #(
		.INIT('h80)
	) name199 (
		_w368_,
		_w367_,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w366_,
		_w370_,
		_w371_
	);
	LUT4 #(
		.INIT('haaca)
	) name201 (
		\g104_reg/NET0131 ,
		\g2_reg/NET0131 ,
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\g1268_reg/NET0131 ,
		\g1269_reg/NET0131 ,
		_w373_
	);
	LUT2 #(
		.INIT('h9)
	) name203 (
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		_w374_
	);
	LUT2 #(
		.INIT('h6)
	) name204 (
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w259_,
		_w374_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		\g1073_reg/NET0131 ,
		\g1179_reg/NET0131 ,
		_w377_
	);
	LUT4 #(
		.INIT('h0001)
	) name207 (
		\g4370_pad ,
		\g4371_pad ,
		\g4372_pad ,
		\g4373_pad ,
		_w378_
	);
	LUT2 #(
		.INIT('h7)
	) name208 (
		_w377_,
		_w378_,
		_w379_
	);
	LUT4 #(
		.INIT('h7fff)
	) name209 (
		\g1263_reg/NET0131 ,
		_w353_,
		_w354_,
		_w355_,
		_w380_
	);
	LUT4 #(
		.INIT('h7fff)
	) name210 (
		\g1257_reg/NET0131 ,
		_w353_,
		_w354_,
		_w355_,
		_w381_
	);
	LUT4 #(
		.INIT('h7fff)
	) name211 (
		\g1266_reg/NET0131 ,
		_w353_,
		_w354_,
		_w355_,
		_w382_
	);
	LUT4 #(
		.INIT('h7f80)
	) name212 (
		\g1207_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		\g1217_reg/NET0131 ,
		_w383_
	);
	LUT2 #(
		.INIT('he)
	) name213 (
		\g1231_reg/NET0131 ,
		_w383_,
		_w384_
	);
	LUT4 #(
		.INIT('h0001)
	) name214 (
		\g1227_reg/NET0131 ,
		\g1228_reg/NET0131 ,
		\g1229_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		_w385_
	);
	LUT4 #(
		.INIT('h0001)
	) name215 (
		\g1223_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		\g1225_reg/NET0131 ,
		\g1226_reg/NET0131 ,
		_w386_
	);
	LUT2 #(
		.INIT('h7)
	) name216 (
		_w385_,
		_w386_,
		_w387_
	);
	LUT3 #(
		.INIT('hf6)
	) name217 (
		\g1207_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1231_reg/NET0131 ,
		_w388_
	);
	LUT3 #(
		.INIT('h07)
	) name218 (
		\g1207_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w389_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		\g1231_reg/NET0131 ,
		\g2662_pad ,
		_w390_
	);
	LUT3 #(
		.INIT('h04)
	) name220 (
		_w299_,
		_w390_,
		_w389_,
		_w391_
	);
	LUT3 #(
		.INIT('h6a)
	) name221 (
		\g871_reg/NET0131 ,
		\g929_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w392_
	);
	LUT2 #(
		.INIT('hd)
	) name222 (
		\g1207_reg/NET0131 ,
		\g1231_reg/NET0131 ,
		_w393_
	);
	LUT2 #(
		.INIT('h6)
	) name223 (
		\g104_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		_w394_
	);
	LUT2 #(
		.INIT('h6)
	) name224 (
		\g104_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w395_
	);
	LUT2 #(
		.INIT('h6)
	) name225 (
		\g104_reg/NET0131 ,
		\g1220_reg/NET0131 ,
		_w396_
	);
	LUT2 #(
		.INIT('h6)
	) name226 (
		\g104_reg/NET0131 ,
		\g1207_reg/NET0131 ,
		_w397_
	);
	LUT2 #(
		.INIT('h6)
	) name227 (
		\g104_reg/NET0131 ,
		\g1225_reg/NET0131 ,
		_w398_
	);
	LUT2 #(
		.INIT('h6)
	) name228 (
		\g104_reg/NET0131 ,
		\g1227_reg/NET0131 ,
		_w399_
	);
	LUT2 #(
		.INIT('h6)
	) name229 (
		\g104_reg/NET0131 ,
		\g1228_reg/NET0131 ,
		_w400_
	);
	LUT2 #(
		.INIT('h6)
	) name230 (
		\g104_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		_w401_
	);
	LUT2 #(
		.INIT('h6)
	) name231 (
		\g104_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		_w402_
	);
	LUT2 #(
		.INIT('h6)
	) name232 (
		\g104_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		_w403_
	);
	LUT2 #(
		.INIT('h6)
	) name233 (
		\g104_reg/NET0131 ,
		\g1226_reg/NET0131 ,
		_w404_
	);
	LUT3 #(
		.INIT('h40)
	) name234 (
		\g1211_reg/NET0131 ,
		\g1217_reg/NET0131 ,
		\g1220_reg/NET0131 ,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\g1207_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w405_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		\g1207_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		_w405_,
		_w408_,
		_w409_
	);
	LUT3 #(
		.INIT('h80)
	) name239 (
		\g1211_reg/NET0131 ,
		\g1217_reg/NET0131 ,
		\g1220_reg/NET0131 ,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w408_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h6)
	) name241 (
		\g104_reg/NET0131 ,
		\g1217_reg/NET0131 ,
		_w412_
	);
	LUT2 #(
		.INIT('h6)
	) name242 (
		\g104_reg/NET0131 ,
		\g1229_reg/NET0131 ,
		_w413_
	);
	LUT2 #(
		.INIT('h6)
	) name243 (
		\g929_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w414_
	);
	LUT4 #(
		.INIT('hfff7)
	) name244 (
		\g1211_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		\g1217_reg/NET0131 ,
		\g1220_reg/NET0131 ,
		_w415_
	);
	LUT3 #(
		.INIT('h20)
	) name245 (
		\g1444_reg/NET0131 ,
		\g1450_reg/NET0131 ,
		\g1454_reg/NET0131 ,
		_w416_
	);
	LUT3 #(
		.INIT('hb0)
	) name246 (
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		\g942_reg/NET0131 ,
		_w417_
	);
	LUT3 #(
		.INIT('h80)
	) name247 (
		\g1114_reg/NET0131 ,
		\g1118_reg/NET0131 ,
		\g1122_reg/NET0131 ,
		_w418_
	);
	LUT4 #(
		.INIT('h8000)
	) name248 (
		\g1110_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w212_,
		_w418_,
		_w419_
	);
	LUT4 #(
		.INIT('h78f0)
	) name249 (
		\g1114_reg/NET0131 ,
		\g1118_reg/NET0131 ,
		\g1122_reg/NET0131 ,
		_w213_,
		_w420_
	);
	LUT2 #(
		.INIT('he)
	) name250 (
		\g1097_reg/NET0131 ,
		_w420_,
		_w421_
	);
	LUT3 #(
		.INIT('hbe)
	) name251 (
		\g1097_reg/NET0131 ,
		\g1126_reg/NET0131 ,
		_w419_,
		_w422_
	);
	LUT3 #(
		.INIT('h80)
	) name252 (
		\g1110_reg/NET0131 ,
		\g1126_reg/NET0131 ,
		\g1142_reg/NET0131 ,
		_w423_
	);
	LUT3 #(
		.INIT('h80)
	) name253 (
		_w212_,
		_w418_,
		_w423_,
		_w424_
	);
	LUT4 #(
		.INIT('h0001)
	) name254 (
		\g1166_reg/NET0131 ,
		\g7423_pad ,
		\g7424_pad ,
		\g7425_pad ,
		_w425_
	);
	LUT4 #(
		.INIT('h80ff)
	) name255 (
		_w212_,
		_w418_,
		_w423_,
		_w425_,
		_w426_
	);
	LUT4 #(
		.INIT('h8000)
	) name256 (
		\g1226_reg/NET0131 ,
		_w353_,
		_w406_,
		_w410_,
		_w427_
	);
	LUT4 #(
		.INIT('hf6fc)
	) name257 (
		\g1227_reg/NET0131 ,
		\g1228_reg/NET0131 ,
		\g1231_reg/NET0131 ,
		_w427_,
		_w428_
	);
	LUT3 #(
		.INIT('h80)
	) name258 (
		\g1227_reg/NET0131 ,
		\g1228_reg/NET0131 ,
		\g1229_reg/NET0131 ,
		_w429_
	);
	LUT4 #(
		.INIT('h60a0)
	) name259 (
		\g1229_reg/NET0131 ,
		_w354_,
		_w390_,
		_w427_,
		_w430_
	);
	LUT4 #(
		.INIT('h8000)
	) name260 (
		\g1509_reg/NET0131 ,
		_w202_,
		_w206_,
		_w203_,
		_w431_
	);
	LUT3 #(
		.INIT('h80)
	) name261 (
		\g1462_reg/NET0131 ,
		\g1467_reg/NET0131 ,
		_w431_,
		_w432_
	);
	LUT4 #(
		.INIT('h060c)
	) name262 (
		\g1462_reg/NET0131 ,
		\g1467_reg/NET0131 ,
		_w208_,
		_w431_,
		_w433_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name263 (
		\g1486_reg/NET0131 ,
		_w202_,
		_w206_,
		_w207_,
		_w434_
	);
	LUT3 #(
		.INIT('hde)
	) name264 (
		\g1227_reg/NET0131 ,
		\g1231_reg/NET0131 ,
		_w427_,
		_w435_
	);
	LUT4 #(
		.INIT('h060c)
	) name265 (
		\g1514_reg/NET0131 ,
		\g1519_reg/NET0131 ,
		_w208_,
		_w205_,
		_w436_
	);
	LUT3 #(
		.INIT('h12)
	) name266 (
		\g1462_reg/NET0131 ,
		_w208_,
		_w431_,
		_w437_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name267 (
		\g1226_reg/NET0131 ,
		_w353_,
		_w406_,
		_w410_,
		_w438_
	);
	LUT2 #(
		.INIT('he)
	) name268 (
		\g1231_reg/NET0131 ,
		_w438_,
		_w439_
	);
	LUT3 #(
		.INIT('hde)
	) name269 (
		\g1225_reg/NET0131 ,
		\g1231_reg/NET0131 ,
		_w347_,
		_w440_
	);
	LUT4 #(
		.INIT('h4888)
	) name270 (
		\g1230_reg/NET0131 ,
		\g2662_pad ,
		_w427_,
		_w429_,
		_w441_
	);
	LUT2 #(
		.INIT('he)
	) name271 (
		\g1231_reg/NET0131 ,
		_w441_,
		_w442_
	);
	LUT4 #(
		.INIT('h1333)
	) name272 (
		\g1354_reg/NET0131 ,
		\g1357_reg/NET0131 ,
		_w181_,
		_w248_,
		_w443_
	);
	LUT3 #(
		.INIT('h80)
	) name273 (
		_w181_,
		_w248_,
		_w331_,
		_w444_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name274 (
		\g1247_reg/NET0131 ,
		_w181_,
		_w248_,
		_w331_,
		_w445_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		_w443_,
		_w445_,
		_w446_
	);
	LUT4 #(
		.INIT('h8000)
	) name276 (
		\g1037_reg/NET0131 ,
		\g1041_reg/NET0131 ,
		\g1149_reg/NET0131 ,
		_w189_,
		_w447_
	);
	LUT4 #(
		.INIT('he4a8)
	) name277 (
		\g1045_reg/NET0131 ,
		_w186_,
		_w197_,
		_w447_,
		_w448_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name278 (
		\g1065_reg/NET0131 ,
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w449_
	);
	LUT4 #(
		.INIT('hff48)
	) name279 (
		\g1065_reg/NET0131 ,
		_w186_,
		_w193_,
		_w449_,
		_w450_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name280 (
		\g1053_reg/NET0131 ,
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w451_
	);
	LUT4 #(
		.INIT('hff48)
	) name281 (
		\g1053_reg/NET0131 ,
		_w186_,
		_w199_,
		_w451_,
		_w452_
	);
	LUT4 #(
		.INIT('h28a0)
	) name282 (
		\g1247_reg/NET0131 ,
		\g1342_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w181_,
		_w453_
	);
	LUT4 #(
		.INIT('h1450)
	) name283 (
		\g1097_reg/NET0131 ,
		\g1126_reg/NET0131 ,
		\g1142_reg/NET0131 ,
		_w419_,
		_w454_
	);
	LUT4 #(
		.INIT('h1333)
	) name284 (
		\g1065_reg/NET0131 ,
		\g1069_reg/NET0131 ,
		_w186_,
		_w193_,
		_w455_
	);
	LUT4 #(
		.INIT('h80a0)
	) name285 (
		\g1069_reg/NET0131 ,
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w456_
	);
	LUT4 #(
		.INIT('hb300)
	) name286 (
		\g1065_reg/NET0131 ,
		_w186_,
		_w193_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w455_,
		_w457_,
		_w458_
	);
	LUT4 #(
		.INIT('h0020)
	) name288 (
		\g1061_reg/NET0131 ,
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w459_
	);
	LUT4 #(
		.INIT('h7f00)
	) name289 (
		\g1053_reg/NET0131 ,
		\g1057_reg/NET0131 ,
		_w199_,
		_w459_,
		_w460_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name290 (
		\g1061_reg/NET0131 ,
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w461_
	);
	LUT2 #(
		.INIT('h2)
	) name291 (
		\g1057_reg/NET0131 ,
		\g1061_reg/NET0131 ,
		_w462_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w186_,
		_w462_,
		_w463_
	);
	LUT4 #(
		.INIT('h070f)
	) name293 (
		\g1053_reg/NET0131 ,
		_w199_,
		_w461_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('hb)
	) name294 (
		_w460_,
		_w464_,
		_w465_
	);
	LUT3 #(
		.INIT('h28)
	) name295 (
		\g1247_reg/NET0131 ,
		\g1360_reg/NET0131 ,
		_w444_,
		_w466_
	);
	LUT4 #(
		.INIT('h1333)
	) name296 (
		\g1053_reg/NET0131 ,
		\g1057_reg/NET0131 ,
		_w186_,
		_w199_,
		_w467_
	);
	LUT4 #(
		.INIT('h80a0)
	) name297 (
		\g1057_reg/NET0131 ,
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w468_
	);
	LUT4 #(
		.INIT('hb300)
	) name298 (
		\g1053_reg/NET0131 ,
		_w186_,
		_w199_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w467_,
		_w469_,
		_w470_
	);
	LUT4 #(
		.INIT('h1222)
	) name300 (
		\g1328_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w246_,
		_w256_,
		_w471_
	);
	LUT2 #(
		.INIT('he)
	) name301 (
		_w242_,
		_w471_,
		_w472_
	);
	LUT4 #(
		.INIT('he4a8)
	) name302 (
		\g1041_reg/NET0131 ,
		_w186_,
		_w197_,
		_w225_,
		_w473_
	);
	LUT3 #(
		.INIT('h12)
	) name303 (
		\g1472_reg/NET0131 ,
		_w208_,
		_w432_,
		_w474_
	);
	LUT2 #(
		.INIT('he)
	) name304 (
		\g2_reg/NET0131 ,
		\g962_pad ,
		_w475_
	);
	LUT2 #(
		.INIT('he)
	) name305 (
		\g1189_reg/NET0131 ,
		\g7505_pad ,
		_w476_
	);
	LUT2 #(
		.INIT('h7)
	) name306 (
		\g1405_reg/NET0131 ,
		\g1412_reg/NET0131 ,
		_w477_
	);
	assign \g1006_pad  = 1'b0;
	assign \g1158_reg/P0001  = _w35_ ;
	assign \g1252_reg/P0001  = _w57_ ;
	assign \g1260_reg/P0001  = _w61_ ;
	assign \g1416_reg/NET0131_syn_2  = _w119_ ;
	assign \g17/_0_  = _w184_ ;
	assign \g19189/_0_  = _w195_ ;
	assign \g19252/_0_  = _w196_ ;
	assign \g19253/_0_  = _w200_ ;
	assign \g19273/_3_  = _w201_ ;
	assign \g19284/_0_  = _w209_ ;
	assign \g19285/_0_  = _w215_ ;
	assign \g19295/_3_  = _w216_ ;
	assign \g19302/_0_  = _w217_ ;
	assign \g19303/_0_  = _w218_ ;
	assign \g19304/_0_  = _w220_ ;
	assign \g19308/_0_  = _w221_ ;
	assign \g19309/_0_  = _w222_ ;
	assign \g19310/_0_  = _w223_ ;
	assign \g19321/_0_  = _w227_ ;
	assign \g19326/_3_  = _w228_ ;
	assign \g19331/_0_  = _w229_ ;
	assign \g19341/_0_  = _w232_ ;
	assign \g19366/_0_  = _w234_ ;
	assign \g19372/_3_  = _w235_ ;
	assign \g19385/_0_  = _w236_ ;
	assign \g19386/_0_  = _w239_ ;
	assign \g19387/_0_  = _w240_ ;
	assign \g19388/_0_  = _w241_ ;
	assign \g19389/_0_  = _w247_ ;
	assign \g19390/_0_  = _w249_ ;
	assign \g19392/_0_  = _w254_ ;
	assign \g19393/_0_  = _w258_ ;
	assign \g19394/_0_  = _w261_ ;
	assign \g19398/_0_  = _w265_ ;
	assign \g19399/_0_  = _w267_ ;
	assign \g19400/_0_  = _w269_ ;
	assign \g19401/_0_  = _w271_ ;
	assign \g19403/_0_  = _w274_ ;
	assign \g19405/_0_  = _w275_ ;
	assign \g19406/_0_  = _w276_ ;
	assign \g19437/_0_  = _w279_ ;
	assign \g19438/_0_  = _w283_ ;
	assign \g19445/_0_  = _w284_ ;
	assign \g19446/_0_  = _w285_ ;
	assign \g19450/_3_  = _w286_ ;
	assign \g19472/_0_  = _w287_ ;
	assign \g19473/_0_  = _w288_ ;
	assign \g19474/_0_  = _w290_ ;
	assign \g19476/_0_  = _w291_ ;
	assign \g19484/_0_  = _w294_ ;
	assign \g19485/_0_  = _w298_ ;
	assign \g19492/_0_  = _w301_ ;
	assign \g19493/_0_  = _w302_ ;
	assign \g19499/_0_  = _w303_ ;
	assign \g19500/_0_  = _w306_ ;
	assign \g19501/_0_  = _w308_ ;
	assign \g19502/_0_  = _w309_ ;
	assign \g19503/_0_  = _w311_ ;
	assign \g19504/_0_  = _w313_ ;
	assign \g19507/_3_  = _w314_ ;
	assign \g19508/_3_  = _w315_ ;
	assign \g19512/_3_  = _w316_ ;
	assign \g19513/_3_  = _w317_ ;
	assign \g19514/_3_  = _w318_ ;
	assign \g19528/_0_  = _w319_ ;
	assign \g19529/_0_  = _w321_ ;
	assign \g19534/_0_  = _w322_ ;
	assign \g19535/_0_  = _w323_ ;
	assign \g19536/_0_  = _w324_ ;
	assign \g19538/_0_  = _w325_ ;
	assign \g19542/_0_  = _w326_ ;
	assign \g19560/_0_  = _w335_ ;
	assign \g19563/_0_  = _w338_ ;
	assign \g19565/_0_  = _w339_ ;
	assign \g19567/_0_  = _w341_ ;
	assign \g19569/_1_  = _w342_ ;
	assign \g19572/_0_  = _w344_ ;
	assign \g19574/_3_  = _w345_ ;
	assign \g19614/_0_  = _w349_ ;
	assign \g19615/_0_  = _w351_ ;
	assign \g19620/_0_  = _w358_ ;
	assign \g19626/_0_  = _w359_ ;
	assign \g19629/_0_  = _w360_ ;
	assign \g19631/_0_  = _w361_ ;
	assign \g19666/_0_  = _w362_ ;
	assign \g19667/_0_  = _w363_ ;
	assign \g19669/_0_  = _w364_ ;
	assign \g19677/_0_  = _w371_ ;
	assign \g19690/_3_  = _w372_ ;
	assign \g19721/_0_  = _w373_ ;
	assign \g19723/_0_  = _w376_ ;
	assign \g19723/_1_  = _w259_ ;
	assign \g19725/_2_  = _w379_ ;
	assign \g19751/_0_  = _w380_ ;
	assign \g19752/_0_  = _w381_ ;
	assign \g19753/_0_  = _w382_ ;
	assign \g19755/_0_  = _w384_ ;
	assign \g19815/_0_  = _w387_ ;
	assign \g19821/_0_  = _w388_ ;
	assign \g19822/_0_  = _w391_ ;
	assign \g19833/_0_  = _w392_ ;
	assign \g19877/_0_  = _w393_ ;
	assign \g19898/_0_  = _w394_ ;
	assign \g19899/_0_  = _w395_ ;
	assign \g19900/_0_  = _w396_ ;
	assign \g19901/_0_  = _w397_ ;
	assign \g19908/_0_  = _w398_ ;
	assign \g19927/_0_  = _w399_ ;
	assign \g19928/_0_  = _w400_ ;
	assign \g19930/_0_  = _w401_ ;
	assign \g19931/_0_  = _w402_ ;
	assign \g19932/_0_  = _w403_ ;
	assign \g19934/_0_  = _w404_ ;
	assign \g19992/_0_  = _w407_ ;
	assign \g19993/_0_  = _w409_ ;
	assign \g20002/_0_  = _w411_ ;
	assign \g20008/_0_  = _w412_ ;
	assign \g20010/_0_  = _w413_ ;
	assign \g20016/_0_  = _w414_ ;
	assign \g20110/_0_  = _w415_ ;
	assign \g20117/_0_  = _w320_ ;
	assign \g20118/_0_  = _w416_ ;
	assign \g20131/_0_  = _w417_ ;
	assign \g20246/_0_  = _w166_ ;
	assign \g20704/_0_  = _w421_ ;
	assign \g20722/_0_  = _w422_ ;
	assign \g20731/_0_  = _w426_ ;
	assign \g20732/_2_  = _w424_ ;
	assign \g20870/_0_  = _w428_ ;
	assign \g20883/_0_  = _w430_ ;
	assign \g20931/_0_  = _w433_ ;
	assign \g20951/_0_  = _w434_ ;
	assign \g20969/_0_  = _w435_ ;
	assign \g20989/_0_  = _w357_ ;
	assign \g21/_2_  = _w436_ ;
	assign \g21070/_0_  = _w437_ ;
	assign \g21108/_0_  = _w439_ ;
	assign \g21122/_0_  = _w440_ ;
	assign \g21152/_0_  = _w442_ ;
	assign \g21191/_0_  = _w446_ ;
	assign \g21279/_0_  = _w448_ ;
	assign \g21316/_0_  = _w450_ ;
	assign \g21323/_0_  = _w452_ ;
	assign \g21349/_3_  = _w365_ ;
	assign \g21352/_3_  = _w453_ ;
	assign \g21464/_0_  = _w454_ ;
	assign \g21472/_0_  = _w458_ ;
	assign \g21484/_0_  = _w465_ ;
	assign \g21510/_0_  = _w466_ ;
	assign \g21517/_0_  = _w470_ ;
	assign \g21608/_0_  = _w472_ ;
	assign \g21625/_0_  = _w473_ ;
	assign \g21644/_1_  = _w474_ ;
	assign \g4655_pad  = _w375_ ;
	assign \g6850_pad  = _w152_ ;
	assign \g6895_pad  = 1'b1;
	assign \g7048_pad  = _w173_ ;
	assign \g7103_pad  = _w475_ ;
	assign \g7731_pad  = _w476_ ;
	assign \g7732_pad  = _w135_ ;
	assign \g8219_pad  = _w124_ ;
	assign \g8663_pad  = _w477_ ;
endmodule;