module top( \a0_pad  , \a1_pad  , \a2_pad  , \a3_pad  , \a4_pad  , a_pad , \b0_pad  , \b1_pad  , \b2_pad  , \b3_pad  , \b4_pad  , b_pad , \c0_pad  , \c1_pad  , \c2_pad  , \c3_pad  , \c4_pad  , c_pad , \d0_pad  , \d1_pad  , \d2_pad  , \d3_pad  , \d4_pad  , d_pad , \e0_pad  , \e1_pad  , \e2_pad  , \e3_pad  , \e4_pad  , e_pad , \f0_pad  , \f1_pad  , \f2_pad  , \f3_pad  , \f4_pad  , f_pad , \g0_pad  , \g1_pad  , \g2_pad  , \g3_pad  , \g4_pad  , g_pad , \h0_pad  , \h1_pad  , \h2_pad  , \h3_pad  , \h4_pad  , h_pad , \i0_pad  , \i1_pad  , \i2_pad  , \i3_pad  , \i4_pad  , i_pad , \j0_pad  , \j1_pad  , \j2_pad  , \j3_pad  , \j4_pad  , j_pad , \k0_pad  , \k1_pad  , \k2_pad  , \k3_pad  , k_pad , \l0_pad  , \l1_pad  , \l2_pad  , \l3_pad  , \l4_pad  , l_pad , \m0_pad  , \m1_pad  , \m2_pad  , \m3_pad  , \m6_pad  , m_pad , \n0_pad  , \n1_pad  , \n2_pad  , \n3_pad  , \n4_pad  , n_pad , \o0_pad  , \o1_pad  , \o2_pad  , \o3_pad  , o_pad , \p0_pad  , \p1_pad  , \p2_pad  , \p3_pad  , p_pad , \q0_pad  , \q1_pad  , \q2_pad  , \q3_pad  , q_pad , \r1_pad  , \r2_pad  , \r3_pad  , r_pad , \s0_pad  , \s1_pad  , \s2_pad  , \s3_pad  , s_pad , \t0_pad  , \t1_pad  , \t2_pad  , \t3_pad  , \t4_pad  , t_pad , \u0_pad  , \u1_pad  , \u2_pad  , \u4_pad  , u_pad , \v0_pad  , \v1_pad  , \v2_pad  , v_pad , \w0_pad  , \w1_pad  , \w2_pad  , \w3_pad  , w_pad , \x0_pad  , \x1_pad  , \x2_pad  , \x3_pad  , x_pad , \y0_pad  , \y1_pad  , \y2_pad  , \y3_pad  , y_pad , \z0_pad  , \z1_pad  , \z2_pad  , \z3_pad  , z_pad , \a5_pad  , \a6_pad  , \a7_pad  , \a8_pad  , \a9_pad  , \b5_pad  , \b6_pad  , \b7_pad  , \b8_pad  , \b9_pad  , \c5_pad  , \c6_pad  , \c7_pad  , \c8_pad  , \c9_pad  , \d5_pad  , \d6_pad  , \d7_pad  , \d8_pad  , \d9_pad  , \e5_pad  , \e6_pad  , \e7_pad  , \e8_pad  , \e9_pad  , \f5_pad  , \f6_pad  , \f7_pad  , \f8_pad  , \f9_pad  , \g5_pad  , \g6_pad  , \g7_pad  , \g8_pad  , \g9_pad  , \h5_pad  , \h6_pad  , \h7_pad  , \h8_pad  , \h9_pad  , \i5_pad  , \i6_pad  , \i7_pad  , \i8_pad  , \i9_pad  , \j5_pad  , \j6_pad  , \j7_pad  , \j8_pad  , \j9_pad  , \k5_pad  , \k6_pad  , \k7_pad  , \k8_pad  , \k9_pad  , \l5_pad  , \l6_pad  , \l7_pad  , \l8_pad  , \l9_pad  , \m7_pad  , \m8_pad  , \m9_pad  , \n5_pad  , \n6_pad  , \n7_pad  , \n8_pad  , \n9_pad  , \o4_pad  , \o5_pad  , \o6_pad  , \o7_pad  , \o8_pad  , \o9_pad  , \p4_pad  , \p5_pad  , \p6_pad  , \p7_pad  , \p8_pad  , \p9_pad  , \q4_pad  , \q5_pad  , \q6_pad  , \q7_pad  , \q8_pad  , \q9_pad  , \r4_pad  , \r5_pad  , \r6_pad  , \r7_pad  , \r8_pad  , \r9_pad  , \s4_pad  , \s6_pad  , \s7_pad  , \s8_pad  , \s9_pad  , \t6_pad  , \t7_pad  , \t8_pad  , \t9_pad  , \u6_pad  , \u7_pad  , \u8_pad  , \u9_pad  , \v4_pad  , \v6_pad  , \v7_pad  , \v8_pad  , \v9_pad  , \w4_pad  , \w5_pad  , \w6_pad  , \w7_pad  , \w8_pad  , \w9_pad  , \x4_pad  , \x5_pad  , \x6_pad  , \x7_pad  , \x8_pad  , \y4_pad  , \y5_pad  , \y6_pad  , \y7_pad  , \y8_pad  , \z4_pad  , \z5_pad  , \z6_pad  , \z7_pad  , \z8_pad  );
  input \a0_pad  ;
  input \a1_pad  ;
  input \a2_pad  ;
  input \a3_pad  ;
  input \a4_pad  ;
  input a_pad ;
  input \b0_pad  ;
  input \b1_pad  ;
  input \b2_pad  ;
  input \b3_pad  ;
  input \b4_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input \c1_pad  ;
  input \c2_pad  ;
  input \c3_pad  ;
  input \c4_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input \d1_pad  ;
  input \d2_pad  ;
  input \d3_pad  ;
  input \d4_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input \e1_pad  ;
  input \e2_pad  ;
  input \e3_pad  ;
  input \e4_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input \f1_pad  ;
  input \f2_pad  ;
  input \f3_pad  ;
  input \f4_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input \g1_pad  ;
  input \g2_pad  ;
  input \g3_pad  ;
  input \g4_pad  ;
  input g_pad ;
  input \h0_pad  ;
  input \h1_pad  ;
  input \h2_pad  ;
  input \h3_pad  ;
  input \h4_pad  ;
  input h_pad ;
  input \i0_pad  ;
  input \i1_pad  ;
  input \i2_pad  ;
  input \i3_pad  ;
  input \i4_pad  ;
  input i_pad ;
  input \j0_pad  ;
  input \j1_pad  ;
  input \j2_pad  ;
  input \j3_pad  ;
  input \j4_pad  ;
  input j_pad ;
  input \k0_pad  ;
  input \k1_pad  ;
  input \k2_pad  ;
  input \k3_pad  ;
  input k_pad ;
  input \l0_pad  ;
  input \l1_pad  ;
  input \l2_pad  ;
  input \l3_pad  ;
  input \l4_pad  ;
  input l_pad ;
  input \m0_pad  ;
  input \m1_pad  ;
  input \m2_pad  ;
  input \m3_pad  ;
  input \m6_pad  ;
  input m_pad ;
  input \n0_pad  ;
  input \n1_pad  ;
  input \n2_pad  ;
  input \n3_pad  ;
  input \n4_pad  ;
  input n_pad ;
  input \o0_pad  ;
  input \o1_pad  ;
  input \o2_pad  ;
  input \o3_pad  ;
  input o_pad ;
  input \p0_pad  ;
  input \p1_pad  ;
  input \p2_pad  ;
  input \p3_pad  ;
  input p_pad ;
  input \q0_pad  ;
  input \q1_pad  ;
  input \q2_pad  ;
  input \q3_pad  ;
  input q_pad ;
  input \r1_pad  ;
  input \r2_pad  ;
  input \r3_pad  ;
  input r_pad ;
  input \s0_pad  ;
  input \s1_pad  ;
  input \s2_pad  ;
  input \s3_pad  ;
  input s_pad ;
  input \t0_pad  ;
  input \t1_pad  ;
  input \t2_pad  ;
  input \t3_pad  ;
  input \t4_pad  ;
  input t_pad ;
  input \u0_pad  ;
  input \u1_pad  ;
  input \u2_pad  ;
  input \u4_pad  ;
  input u_pad ;
  input \v0_pad  ;
  input \v1_pad  ;
  input \v2_pad  ;
  input v_pad ;
  input \w0_pad  ;
  input \w1_pad  ;
  input \w2_pad  ;
  input \w3_pad  ;
  input w_pad ;
  input \x0_pad  ;
  input \x1_pad  ;
  input \x2_pad  ;
  input \x3_pad  ;
  input x_pad ;
  input \y0_pad  ;
  input \y1_pad  ;
  input \y2_pad  ;
  input \y3_pad  ;
  input y_pad ;
  input \z0_pad  ;
  input \z1_pad  ;
  input \z2_pad  ;
  input \z3_pad  ;
  input z_pad ;
  output \a5_pad  ;
  output \a6_pad  ;
  output \a7_pad  ;
  output \a8_pad  ;
  output \a9_pad  ;
  output \b5_pad  ;
  output \b6_pad  ;
  output \b7_pad  ;
  output \b8_pad  ;
  output \b9_pad  ;
  output \c5_pad  ;
  output \c6_pad  ;
  output \c7_pad  ;
  output \c8_pad  ;
  output \c9_pad  ;
  output \d5_pad  ;
  output \d6_pad  ;
  output \d7_pad  ;
  output \d8_pad  ;
  output \d9_pad  ;
  output \e5_pad  ;
  output \e6_pad  ;
  output \e7_pad  ;
  output \e8_pad  ;
  output \e9_pad  ;
  output \f5_pad  ;
  output \f6_pad  ;
  output \f7_pad  ;
  output \f8_pad  ;
  output \f9_pad  ;
  output \g5_pad  ;
  output \g6_pad  ;
  output \g7_pad  ;
  output \g8_pad  ;
  output \g9_pad  ;
  output \h5_pad  ;
  output \h6_pad  ;
  output \h7_pad  ;
  output \h8_pad  ;
  output \h9_pad  ;
  output \i5_pad  ;
  output \i6_pad  ;
  output \i7_pad  ;
  output \i8_pad  ;
  output \i9_pad  ;
  output \j5_pad  ;
  output \j6_pad  ;
  output \j7_pad  ;
  output \j8_pad  ;
  output \j9_pad  ;
  output \k5_pad  ;
  output \k6_pad  ;
  output \k7_pad  ;
  output \k8_pad  ;
  output \k9_pad  ;
  output \l5_pad  ;
  output \l6_pad  ;
  output \l7_pad  ;
  output \l8_pad  ;
  output \l9_pad  ;
  output \m7_pad  ;
  output \m8_pad  ;
  output \m9_pad  ;
  output \n5_pad  ;
  output \n6_pad  ;
  output \n7_pad  ;
  output \n8_pad  ;
  output \n9_pad  ;
  output \o4_pad  ;
  output \o5_pad  ;
  output \o6_pad  ;
  output \o7_pad  ;
  output \o8_pad  ;
  output \o9_pad  ;
  output \p4_pad  ;
  output \p5_pad  ;
  output \p6_pad  ;
  output \p7_pad  ;
  output \p8_pad  ;
  output \p9_pad  ;
  output \q4_pad  ;
  output \q5_pad  ;
  output \q6_pad  ;
  output \q7_pad  ;
  output \q8_pad  ;
  output \q9_pad  ;
  output \r4_pad  ;
  output \r5_pad  ;
  output \r6_pad  ;
  output \r7_pad  ;
  output \r8_pad  ;
  output \r9_pad  ;
  output \s4_pad  ;
  output \s6_pad  ;
  output \s7_pad  ;
  output \s8_pad  ;
  output \s9_pad  ;
  output \t6_pad  ;
  output \t7_pad  ;
  output \t8_pad  ;
  output \t9_pad  ;
  output \u6_pad  ;
  output \u7_pad  ;
  output \u8_pad  ;
  output \u9_pad  ;
  output \v4_pad  ;
  output \v6_pad  ;
  output \v7_pad  ;
  output \v8_pad  ;
  output \v9_pad  ;
  output \w4_pad  ;
  output \w5_pad  ;
  output \w6_pad  ;
  output \w7_pad  ;
  output \w8_pad  ;
  output \w9_pad  ;
  output \x4_pad  ;
  output \x5_pad  ;
  output \x6_pad  ;
  output \x7_pad  ;
  output \x8_pad  ;
  output \y4_pad  ;
  output \y5_pad  ;
  output \y6_pad  ;
  output \y7_pad  ;
  output \y8_pad  ;
  output \z4_pad  ;
  output \z5_pad  ;
  output \z6_pad  ;
  output \z7_pad  ;
  output \z8_pad  ;
  wire n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 ;
  assign n143 = \k0_pad  & ~\l0_pad  ;
  assign n144 = ~\k0_pad  & \l0_pad  ;
  assign n145 = ~n143 & ~n144 ;
  assign n147 = ~\j3_pad  & n145 ;
  assign n146 = ~\r3_pad  & ~n145 ;
  assign n148 = \m0_pad  & ~n146 ;
  assign n149 = ~n147 & n148 ;
  assign n150 = \m1_pad  & ~\m6_pad  ;
  assign n151 = \k1_pad  & n150 ;
  assign n152 = \o0_pad  & ~\q0_pad  ;
  assign n153 = ~\k1_pad  & ~\l1_pad  ;
  assign n154 = ~\j1_pad  & n153 ;
  assign n155 = ~\h1_pad  & ~\i1_pad  ;
  assign n156 = n154 & n155 ;
  assign n157 = ~\n0_pad  & n156 ;
  assign n158 = \f0_pad  & n157 ;
  assign n159 = \y3_pad  & \z3_pad  ;
  assign n160 = ~\a4_pad  & ~\b4_pad  ;
  assign n161 = ~\c4_pad  & n160 ;
  assign n162 = n159 & n161 ;
  assign n163 = ~\x3_pad  & n162 ;
  assign n164 = \l4_pad  & ~n163 ;
  assign n166 = ~\s1_pad  & n164 ;
  assign n165 = ~\r1_pad  & ~n164 ;
  assign n167 = ~n157 & ~n165 ;
  assign n168 = ~n166 & n167 ;
  assign n169 = ~n158 & ~n168 ;
  assign n170 = n152 & ~n169 ;
  assign n171 = ~\m0_pad  & n157 ;
  assign n172 = ~h_pad & ~n143 ;
  assign n173 = ~p_pad & n143 ;
  assign n174 = ~n172 & ~n173 ;
  assign n175 = n171 & n174 ;
  assign n177 = ~\s2_pad  & n164 ;
  assign n176 = ~\r2_pad  & ~n164 ;
  assign n178 = ~n171 & ~n176 ;
  assign n179 = ~n177 & n178 ;
  assign n180 = ~n175 & ~n179 ;
  assign n181 = n152 & ~n180 ;
  assign n187 = \e4_pad  & \f4_pad  ;
  assign n188 = ~\g4_pad  & n187 ;
  assign n189 = ~\h4_pad  & n188 ;
  assign n190 = \h1_pad  & ~\x0_pad  ;
  assign n191 = \j1_pad  & ~\z0_pad  ;
  assign n195 = ~n190 & ~n191 ;
  assign n194 = ~\a1_pad  & \k1_pad  ;
  assign n192 = ~\b1_pad  & \l1_pad  ;
  assign n193 = \i1_pad  & ~\y0_pad  ;
  assign n196 = ~n192 & ~n193 ;
  assign n197 = ~n194 & n196 ;
  assign n198 = n195 & n197 ;
  assign n199 = ~n189 & ~n198 ;
  assign n200 = \m6_pad  & n199 ;
  assign n182 = \k1_pad  & \l1_pad  ;
  assign n183 = \j1_pad  & ~n153 ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = n155 & n184 ;
  assign n186 = ~n154 & ~n185 ;
  assign n201 = \h1_pad  & \i1_pad  ;
  assign n202 = ~n156 & ~n201 ;
  assign n203 = ~n186 & n202 ;
  assign n204 = n200 & n203 ;
  assign n206 = ~\s3_pad  & n204 ;
  assign n205 = ~\r3_pad  & ~n204 ;
  assign n207 = n152 & ~n205 ;
  assign n208 = ~n206 & n207 ;
  assign n210 = ~\k3_pad  & n145 ;
  assign n209 = ~\s3_pad  & ~n145 ;
  assign n211 = \m0_pad  & ~n209 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = \l1_pad  & n150 ;
  assign n214 = \e0_pad  & n157 ;
  assign n216 = ~\t1_pad  & n164 ;
  assign n215 = ~\s1_pad  & ~n164 ;
  assign n217 = ~n157 & ~n215 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = ~n214 & ~n218 ;
  assign n220 = n152 & ~n219 ;
  assign n221 = n145 & n171 ;
  assign n223 = ~\s2_pad  & ~n164 ;
  assign n224 = ~\t2_pad  & n164 ;
  assign n225 = ~n223 & ~n224 ;
  assign n226 = ~n221 & ~n225 ;
  assign n222 = ~i_pad & n221 ;
  assign n227 = n152 & ~n222 ;
  assign n228 = ~n226 & n227 ;
  assign n230 = ~\t3_pad  & n204 ;
  assign n229 = ~\s3_pad  & ~n204 ;
  assign n231 = n152 & ~n229 ;
  assign n232 = ~n230 & n231 ;
  assign n234 = ~\l3_pad  & n145 ;
  assign n233 = ~\t3_pad  & ~n145 ;
  assign n235 = \m0_pad  & ~n233 ;
  assign n236 = ~n234 & n235 ;
  assign n237 = \h1_pad  & \l4_pad  ;
  assign n238 = \d0_pad  & n157 ;
  assign n240 = ~\u1_pad  & n164 ;
  assign n239 = ~\t1_pad  & ~n164 ;
  assign n241 = ~n157 & ~n239 ;
  assign n242 = ~n240 & n241 ;
  assign n243 = ~n238 & ~n242 ;
  assign n244 = n152 & ~n243 ;
  assign n246 = ~\t2_pad  & ~n164 ;
  assign n247 = ~\u2_pad  & n164 ;
  assign n248 = ~n246 & ~n247 ;
  assign n249 = ~n221 & ~n248 ;
  assign n245 = ~j_pad & n221 ;
  assign n250 = n152 & ~n245 ;
  assign n251 = ~n249 & n250 ;
  assign n253 = ~\t4_pad  & n204 ;
  assign n252 = ~\t3_pad  & ~n204 ;
  assign n254 = n152 & ~n252 ;
  assign n255 = ~n253 & n254 ;
  assign n256 = \m0_pad  & \m3_pad  ;
  assign n257 = \i1_pad  & \l4_pad  ;
  assign n258 = n152 & ~n171 ;
  assign n260 = \v1_pad  & n164 ;
  assign n259 = \u1_pad  & ~n164 ;
  assign n261 = ~n157 & ~n259 ;
  assign n262 = ~n260 & n261 ;
  assign n263 = n258 & ~n262 ;
  assign n265 = ~\u2_pad  & ~n164 ;
  assign n266 = ~\v2_pad  & n164 ;
  assign n267 = ~n265 & ~n266 ;
  assign n268 = ~n221 & ~n267 ;
  assign n264 = ~k_pad & n221 ;
  assign n269 = n152 & ~n264 ;
  assign n270 = ~n268 & n269 ;
  assign n272 = ~\u4_pad  & n204 ;
  assign n271 = ~\t4_pad  & ~n204 ;
  assign n273 = n152 & ~n271 ;
  assign n274 = ~n272 & n273 ;
  assign n275 = \m0_pad  & \n3_pad  ;
  assign n276 = \j1_pad  & \l4_pad  ;
  assign n278 = ~\v1_pad  & ~n164 ;
  assign n279 = ~\w1_pad  & n164 ;
  assign n280 = ~n278 & ~n279 ;
  assign n281 = ~n157 & ~n280 ;
  assign n277 = ~\k0_pad  & n157 ;
  assign n282 = n152 & ~n277 ;
  assign n283 = ~n281 & n282 ;
  assign n285 = ~\v2_pad  & ~n164 ;
  assign n286 = ~\w2_pad  & n164 ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = ~n221 & ~n287 ;
  assign n284 = ~l_pad & n221 ;
  assign n289 = n152 & ~n284 ;
  assign n290 = ~n288 & n289 ;
  assign n292 = ~\w3_pad  & n204 ;
  assign n291 = ~\u4_pad  & ~n204 ;
  assign n293 = n152 & ~n291 ;
  assign n294 = ~n292 & n293 ;
  assign n295 = \m0_pad  & \o3_pad  ;
  assign n296 = \k1_pad  & \l4_pad  ;
  assign n298 = ~\w1_pad  & ~n164 ;
  assign n299 = ~\x1_pad  & n164 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = ~n157 & ~n300 ;
  assign n297 = ~\l0_pad  & n157 ;
  assign n302 = n152 & ~n297 ;
  assign n303 = ~n301 & n302 ;
  assign n305 = ~\w2_pad  & ~n164 ;
  assign n306 = ~\x2_pad  & n164 ;
  assign n307 = ~n305 & ~n306 ;
  assign n308 = ~n221 & ~n307 ;
  assign n304 = ~m_pad & n221 ;
  assign n309 = n152 & ~n304 ;
  assign n310 = ~n308 & n309 ;
  assign n311 = \w3_pad  & ~n204 ;
  assign n312 = \h1_pad  & ~\i1_pad  ;
  assign n313 = \s0_pad  & n312 ;
  assign n314 = n154 & n313 ;
  assign n325 = \t0_pad  & n154 ;
  assign n326 = \i1_pad  & ~n325 ;
  assign n318 = ~\l1_pad  & \u0_pad  ;
  assign n319 = ~\j1_pad  & \w0_pad  ;
  assign n320 = ~n318 & ~n319 ;
  assign n315 = ~\j1_pad  & ~\l1_pad  ;
  assign n321 = ~\k1_pad  & ~n315 ;
  assign n322 = ~n320 & n321 ;
  assign n316 = \k1_pad  & \v0_pad  ;
  assign n317 = n315 & n316 ;
  assign n323 = ~\i1_pad  & ~n317 ;
  assign n324 = ~n322 & n323 ;
  assign n327 = ~\h1_pad  & ~n324 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = ~n314 & ~n328 ;
  assign n330 = n200 & ~n329 ;
  assign n331 = ~n311 & ~n330 ;
  assign n332 = n152 & ~n331 ;
  assign n333 = \m0_pad  & \p3_pad  ;
  assign n334 = \l1_pad  & \l4_pad  ;
  assign n335 = q_pad & n157 ;
  assign n337 = ~\y1_pad  & n164 ;
  assign n336 = ~\x1_pad  & ~n164 ;
  assign n338 = ~n157 & ~n336 ;
  assign n339 = ~n337 & n338 ;
  assign n340 = ~n335 & ~n339 ;
  assign n341 = n152 & ~n340 ;
  assign n343 = ~\x2_pad  & ~n164 ;
  assign n344 = ~\y2_pad  & n164 ;
  assign n345 = ~n343 & ~n344 ;
  assign n346 = ~n221 & ~n345 ;
  assign n342 = ~n_pad & n221 ;
  assign n347 = n152 & ~n342 ;
  assign n348 = ~n346 & n347 ;
  assign n349 = n152 & ~n157 ;
  assign n350 = ~\l4_pad  & \x3_pad  ;
  assign n351 = \l4_pad  & ~\x3_pad  ;
  assign n352 = ~n162 & n351 ;
  assign n353 = ~n350 & ~n352 ;
  assign n354 = n349 & ~n353 ;
  assign n355 = \m0_pad  & \q3_pad  ;
  assign n356 = r_pad & n157 ;
  assign n358 = ~\z1_pad  & n164 ;
  assign n357 = ~\y1_pad  & ~n164 ;
  assign n359 = ~n157 & ~n357 ;
  assign n360 = ~n358 & n359 ;
  assign n361 = ~n356 & ~n360 ;
  assign n362 = n152 & ~n361 ;
  assign n364 = ~\y2_pad  & ~n164 ;
  assign n365 = ~\z2_pad  & n164 ;
  assign n366 = ~n364 & ~n365 ;
  assign n367 = ~n221 & ~n366 ;
  assign n363 = ~o_pad & n221 ;
  assign n368 = n152 & ~n363 ;
  assign n369 = ~n367 & n368 ;
  assign n370 = \y3_pad  & n352 ;
  assign n371 = ~\y3_pad  & ~n351 ;
  assign n372 = ~n370 & ~n371 ;
  assign n373 = n349 & ~n372 ;
  assign n374 = \m0_pad  & \r3_pad  ;
  assign n375 = s_pad & n157 ;
  assign n377 = ~\a2_pad  & n164 ;
  assign n376 = ~\z1_pad  & ~n164 ;
  assign n378 = ~n157 & ~n376 ;
  assign n379 = ~n377 & n378 ;
  assign n380 = ~n375 & ~n379 ;
  assign n381 = n152 & ~n380 ;
  assign n382 = p_pad & n221 ;
  assign n383 = \z2_pad  & ~n164 ;
  assign n384 = ~n221 & n383 ;
  assign n385 = ~n382 & ~n384 ;
  assign n386 = n152 & ~n385 ;
  assign n387 = ~\z3_pad  & ~n370 ;
  assign n388 = n159 & n351 ;
  assign n389 = ~n161 & n388 ;
  assign n390 = ~n387 & ~n389 ;
  assign n391 = n349 & ~n390 ;
  assign n392 = \m0_pad  & \s3_pad  ;
  assign n393 = t_pad & n157 ;
  assign n395 = ~\b2_pad  & n164 ;
  assign n394 = ~\a2_pad  & ~n164 ;
  assign n396 = ~n157 & ~n394 ;
  assign n397 = ~n395 & n396 ;
  assign n398 = ~n393 & ~n397 ;
  assign n399 = n152 & ~n398 ;
  assign n401 = ~\b3_pad  & n204 ;
  assign n400 = ~\a3_pad  & ~n204 ;
  assign n402 = n152 & ~n400 ;
  assign n403 = ~n401 & n402 ;
  assign n408 = ~n145 & n171 ;
  assign n404 = ~\a4_pad  & n389 ;
  assign n405 = \a4_pad  & ~n388 ;
  assign n406 = ~n157 & ~n405 ;
  assign n407 = ~n404 & n406 ;
  assign n409 = n152 & ~n407 ;
  assign n410 = ~n408 & n409 ;
  assign n411 = \m0_pad  & \t3_pad  ;
  assign n412 = u_pad & n157 ;
  assign n414 = ~\c2_pad  & n164 ;
  assign n413 = ~\b2_pad  & ~n164 ;
  assign n415 = ~n157 & ~n413 ;
  assign n416 = ~n414 & n415 ;
  assign n417 = ~n412 & ~n416 ;
  assign n418 = n152 & ~n417 ;
  assign n420 = ~\c3_pad  & n204 ;
  assign n419 = ~\b3_pad  & ~n204 ;
  assign n421 = n152 & ~n419 ;
  assign n422 = ~n420 & n421 ;
  assign n423 = \b4_pad  & ~n404 ;
  assign n424 = n160 & n389 ;
  assign n425 = ~n157 & ~n424 ;
  assign n426 = ~n423 & n425 ;
  assign n427 = n258 & ~n426 ;
  assign n428 = \g1_pad  & ~\j4_pad  ;
  assign n429 = v_pad & n157 ;
  assign n431 = ~\d2_pad  & n164 ;
  assign n430 = ~\c2_pad  & ~n164 ;
  assign n432 = ~n157 & ~n430 ;
  assign n433 = ~n431 & n432 ;
  assign n434 = ~n429 & ~n433 ;
  assign n435 = n152 & ~n434 ;
  assign n437 = ~\d3_pad  & n204 ;
  assign n436 = ~\c3_pad  & ~n204 ;
  assign n438 = n152 & ~n436 ;
  assign n439 = ~n437 & n438 ;
  assign n440 = \c4_pad  & n425 ;
  assign n441 = ~n171 & ~n440 ;
  assign n442 = n152 & ~n441 ;
  assign n443 = w_pad & n157 ;
  assign n445 = ~\e2_pad  & n164 ;
  assign n444 = ~\d2_pad  & ~n164 ;
  assign n446 = ~n157 & ~n444 ;
  assign n447 = ~n445 & n446 ;
  assign n448 = ~n443 & ~n447 ;
  assign n449 = n152 & ~n448 ;
  assign n451 = ~\e3_pad  & n204 ;
  assign n450 = ~\d3_pad  & ~n204 ;
  assign n452 = n152 & ~n450 ;
  assign n453 = ~n451 & n452 ;
  assign n454 = ~\q0_pad  & n157 ;
  assign n455 = ~\g1_pad  & ~\q0_pad  ;
  assign n456 = \d4_pad  & ~n200 ;
  assign n457 = ~\d4_pad  & n200 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = n455 & ~n458 ;
  assign n460 = ~n454 & ~n459 ;
  assign n461 = \o0_pad  & ~n460 ;
  assign n462 = \h1_pad  & ~\m6_pad  ;
  assign n463 = ~\n0_pad  & n462 ;
  assign n464 = ~\f1_pad  & ~\i4_pad  ;
  assign n465 = \f1_pad  & \i4_pad  ;
  assign n466 = ~n464 & ~n465 ;
  assign n467 = x_pad & n157 ;
  assign n469 = ~\f2_pad  & n164 ;
  assign n468 = ~\e2_pad  & ~n164 ;
  assign n470 = ~n157 & ~n468 ;
  assign n471 = ~n469 & n470 ;
  assign n472 = ~n467 & ~n471 ;
  assign n473 = n152 & ~n472 ;
  assign n475 = ~\f3_pad  & n204 ;
  assign n474 = ~\e3_pad  & ~n204 ;
  assign n476 = n152 & ~n474 ;
  assign n477 = ~n475 & n476 ;
  assign n478 = \e4_pad  & n457 ;
  assign n479 = ~\d4_pad  & ~n157 ;
  assign n480 = n200 & n479 ;
  assign n481 = ~\e4_pad  & ~n480 ;
  assign n482 = ~n478 & ~n481 ;
  assign n483 = \o0_pad  & n455 ;
  assign n484 = ~n157 & n483 ;
  assign n485 = ~n482 & n484 ;
  assign n486 = \i1_pad  & ~\m6_pad  ;
  assign n487 = ~\n0_pad  & n486 ;
  assign n488 = \x3_pad  & n162 ;
  assign n489 = y_pad & n157 ;
  assign n491 = ~\g2_pad  & n164 ;
  assign n490 = ~\f2_pad  & ~n164 ;
  assign n492 = ~n157 & ~n490 ;
  assign n493 = ~n491 & n492 ;
  assign n494 = ~n489 & ~n493 ;
  assign n495 = n152 & ~n494 ;
  assign n497 = ~\g3_pad  & n204 ;
  assign n496 = ~\f3_pad  & ~n204 ;
  assign n498 = n152 & ~n496 ;
  assign n499 = ~n497 & n498 ;
  assign n502 = \f4_pad  & ~n478 ;
  assign n500 = \e4_pad  & ~\f4_pad  ;
  assign n501 = n480 & n500 ;
  assign n503 = n484 & ~n501 ;
  assign n504 = ~n502 & n503 ;
  assign n505 = ~\l3_pad  & ~n145 ;
  assign n506 = ~\d3_pad  & n145 ;
  assign n507 = ~n505 & ~n506 ;
  assign n508 = \m0_pad  & ~n507 ;
  assign n509 = ~\m0_pad  & ~\t3_pad  ;
  assign n510 = ~n508 & ~n509 ;
  assign n511 = \j1_pad  & ~\m6_pad  ;
  assign n512 = ~\n0_pad  & n511 ;
  assign n513 = \n4_pad  & ~n189 ;
  assign n514 = n198 & n513 ;
  assign n515 = \d4_pad  & ~\g1_pad  ;
  assign n516 = n189 & n515 ;
  assign n517 = ~n514 & ~n516 ;
  assign n518 = n152 & ~n517 ;
  assign n519 = z_pad & n157 ;
  assign n521 = ~\h2_pad  & n164 ;
  assign n520 = ~\g2_pad  & ~n164 ;
  assign n522 = ~n157 & ~n520 ;
  assign n523 = ~n521 & n522 ;
  assign n524 = ~n519 & ~n523 ;
  assign n525 = n152 & ~n524 ;
  assign n527 = ~\h3_pad  & n204 ;
  assign n526 = ~\g3_pad  & ~n204 ;
  assign n528 = n152 & ~n526 ;
  assign n529 = ~n527 & n528 ;
  assign n538 = n187 & n480 ;
  assign n539 = \g4_pad  & n484 ;
  assign n540 = ~n538 & n539 ;
  assign n530 = \m0_pad  & ~n145 ;
  assign n531 = n152 & n157 ;
  assign n532 = ~n530 & n531 ;
  assign n533 = ~\g1_pad  & \m6_pad  ;
  assign n534 = ~\d4_pad  & n533 ;
  assign n535 = n188 & n534 ;
  assign n536 = n199 & n535 ;
  assign n537 = n349 & n536 ;
  assign n541 = ~n532 & ~n537 ;
  assign n542 = ~n540 & n541 ;
  assign n543 = ~\k3_pad  & ~n145 ;
  assign n544 = ~\c3_pad  & n145 ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = \m0_pad  & ~n545 ;
  assign n547 = ~\m0_pad  & ~\s3_pad  ;
  assign n548 = ~n546 & ~n547 ;
  assign n549 = \k1_pad  & ~\m6_pad  ;
  assign n550 = ~\n0_pad  & n549 ;
  assign n551 = \h1_pad  & n483 ;
  assign n552 = ~\e1_pad  & n157 ;
  assign n553 = ~\c1_pad  & ~\d1_pad  ;
  assign n554 = n152 & n553 ;
  assign n555 = n552 & n554 ;
  assign n556 = ~n551 & ~n555 ;
  assign n557 = \a0_pad  & n157 ;
  assign n559 = ~\i2_pad  & n164 ;
  assign n558 = ~\h2_pad  & ~n164 ;
  assign n560 = ~n157 & ~n558 ;
  assign n561 = ~n559 & n560 ;
  assign n562 = ~n557 & ~n561 ;
  assign n563 = n152 & ~n562 ;
  assign n565 = ~\i3_pad  & n204 ;
  assign n564 = ~\h3_pad  & ~n204 ;
  assign n566 = n152 & ~n564 ;
  assign n567 = ~n565 & n566 ;
  assign n568 = \m0_pad  & n531 ;
  assign n569 = ~\g4_pad  & n538 ;
  assign n570 = \h4_pad  & n484 ;
  assign n571 = ~n569 & n570 ;
  assign n572 = ~n568 & ~n571 ;
  assign n573 = ~\j3_pad  & ~n145 ;
  assign n574 = ~\b3_pad  & n145 ;
  assign n575 = ~n573 & ~n574 ;
  assign n576 = \m0_pad  & ~n575 ;
  assign n577 = ~\m0_pad  & ~\r3_pad  ;
  assign n578 = ~n576 & ~n577 ;
  assign n579 = \l1_pad  & ~\m6_pad  ;
  assign n580 = ~\n0_pad  & n579 ;
  assign n581 = \e1_pad  & ~n553 ;
  assign n582 = n157 & ~n581 ;
  assign n583 = ~\g1_pad  & ~n582 ;
  assign n584 = \i1_pad  & n583 ;
  assign n585 = \c1_pad  & ~\d1_pad  ;
  assign n586 = n552 & n585 ;
  assign n587 = ~n584 & ~n586 ;
  assign n588 = n152 & ~n587 ;
  assign n589 = \b0_pad  & n157 ;
  assign n591 = ~\j2_pad  & n164 ;
  assign n590 = ~\i2_pad  & ~n164 ;
  assign n592 = ~n157 & ~n590 ;
  assign n593 = ~n591 & n592 ;
  assign n594 = ~n589 & ~n593 ;
  assign n595 = n152 & ~n594 ;
  assign n597 = ~\j3_pad  & n204 ;
  assign n596 = ~\i3_pad  & ~n204 ;
  assign n598 = n152 & ~n596 ;
  assign n599 = ~n597 & n598 ;
  assign n600 = \i4_pad  & ~\n1_pad  ;
  assign n601 = ~\i4_pad  & \n1_pad  ;
  assign n602 = ~n600 & ~n601 ;
  assign n603 = n152 & ~n602 ;
  assign n604 = n164 & n603 ;
  assign n605 = ~\i3_pad  & ~n145 ;
  assign n606 = ~\a3_pad  & n145 ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = \m0_pad  & ~n607 ;
  assign n609 = ~\m0_pad  & ~\q3_pad  ;
  assign n610 = ~n608 & ~n609 ;
  assign n611 = \j1_pad  & n583 ;
  assign n612 = ~\c1_pad  & \d1_pad  ;
  assign n613 = n552 & n612 ;
  assign n614 = ~n611 & ~n613 ;
  assign n615 = n152 & ~n614 ;
  assign n616 = \c0_pad  & n157 ;
  assign n618 = ~\k2_pad  & n164 ;
  assign n617 = ~\j2_pad  & ~n164 ;
  assign n619 = ~n157 & ~n617 ;
  assign n620 = ~n618 & n619 ;
  assign n621 = ~n616 & ~n620 ;
  assign n622 = n152 & ~n621 ;
  assign n624 = ~\k3_pad  & n204 ;
  assign n623 = ~\j3_pad  & ~n204 ;
  assign n625 = n152 & ~n623 ;
  assign n626 = ~n624 & n625 ;
  assign n634 = ~\u0_pad  & n153 ;
  assign n635 = n155 & n634 ;
  assign n636 = \m6_pad  & \n4_pad  ;
  assign n637 = n184 & n636 ;
  assign n638 = ~n635 & n637 ;
  assign n639 = ~n326 & n638 ;
  assign n627 = ~\k1_pad  & ~\w0_pad  ;
  assign n628 = \l1_pad  & ~n627 ;
  assign n629 = ~\i1_pad  & ~\j1_pad  ;
  assign n630 = ~n316 & n629 ;
  assign n631 = ~n628 & n630 ;
  assign n632 = ~\h1_pad  & ~n631 ;
  assign n633 = ~n314 & ~n632 ;
  assign n640 = n199 & ~n633 ;
  assign n641 = n639 & n640 ;
  assign n642 = \j4_pad  & n483 ;
  assign n643 = ~n641 & n642 ;
  assign n644 = ~\j4_pad  & \n4_pad  ;
  assign n645 = n152 & n644 ;
  assign n646 = n533 & n645 ;
  assign n647 = n199 & n646 ;
  assign n648 = ~n329 & n647 ;
  assign n649 = ~n643 & ~n648 ;
  assign n650 = ~\k1_pad  & ~n552 ;
  assign n651 = n583 & ~n650 ;
  assign n652 = \c1_pad  & \d1_pad  ;
  assign n653 = n552 & n652 ;
  assign n654 = ~n651 & ~n653 ;
  assign n655 = n152 & ~n654 ;
  assign n656 = ~a_pad & ~n143 ;
  assign n657 = ~i_pad & n143 ;
  assign n658 = ~n656 & ~n657 ;
  assign n659 = n171 & n658 ;
  assign n661 = ~\l2_pad  & n164 ;
  assign n660 = ~\k2_pad  & ~n164 ;
  assign n662 = ~n171 & ~n660 ;
  assign n663 = ~n661 & n662 ;
  assign n664 = ~n659 & ~n663 ;
  assign n665 = n152 & ~n664 ;
  assign n667 = ~\l3_pad  & n204 ;
  assign n666 = ~\k3_pad  & ~n204 ;
  assign n668 = n152 & ~n666 ;
  assign n669 = ~n667 & n668 ;
  assign n670 = \m1_pad  & n152 ;
  assign n671 = n162 & n670 ;
  assign n672 = n157 & n553 ;
  assign n673 = ~\g1_pad  & \l1_pad  ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = n152 & ~n552 ;
  assign n676 = ~n674 & n675 ;
  assign n677 = ~b_pad & ~n143 ;
  assign n678 = ~j_pad & n143 ;
  assign n679 = ~n677 & ~n678 ;
  assign n680 = n171 & n679 ;
  assign n682 = ~\m2_pad  & n164 ;
  assign n681 = ~\l2_pad  & ~n164 ;
  assign n683 = ~n171 & ~n681 ;
  assign n684 = ~n682 & n683 ;
  assign n685 = ~n680 & ~n684 ;
  assign n686 = n152 & ~n685 ;
  assign n688 = ~\m3_pad  & n204 ;
  assign n687 = ~\l3_pad  & ~n204 ;
  assign n689 = n152 & ~n687 ;
  assign n690 = ~n688 & n689 ;
  assign n691 = ~n163 & n670 ;
  assign n693 = ~\e3_pad  & n145 ;
  assign n692 = ~\m3_pad  & ~n145 ;
  assign n694 = \m0_pad  & ~n692 ;
  assign n695 = ~n693 & n694 ;
  assign n698 = \m1_pad  & ~n517 ;
  assign n696 = ~\n0_pad  & \p0_pad  ;
  assign n697 = ~\m1_pad  & ~n696 ;
  assign n699 = n152 & ~n697 ;
  assign n700 = ~n698 & n699 ;
  assign n701 = ~c_pad & ~n143 ;
  assign n702 = ~k_pad & n143 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = n171 & n703 ;
  assign n706 = ~\n2_pad  & n164 ;
  assign n705 = ~\m2_pad  & ~n164 ;
  assign n707 = ~n171 & ~n705 ;
  assign n708 = ~n706 & n707 ;
  assign n709 = ~n704 & ~n708 ;
  assign n710 = n152 & ~n709 ;
  assign n712 = ~\n3_pad  & n204 ;
  assign n711 = ~\m3_pad  & ~n204 ;
  assign n713 = n152 & ~n711 ;
  assign n714 = ~n712 & n713 ;
  assign n715 = n198 & ~n513 ;
  assign n716 = n518 & ~n715 ;
  assign n718 = ~\f3_pad  & n145 ;
  assign n717 = ~\n3_pad  & ~n145 ;
  assign n719 = \m0_pad  & ~n717 ;
  assign n720 = ~n718 & n719 ;
  assign n721 = n162 & ~n466 ;
  assign n722 = \n1_pad  & ~n162 ;
  assign n723 = ~n721 & ~n722 ;
  assign n724 = \j0_pad  & n157 ;
  assign n726 = ~\o1_pad  & n164 ;
  assign n725 = ~\n1_pad  & ~n164 ;
  assign n727 = ~n157 & ~n725 ;
  assign n728 = ~n726 & n727 ;
  assign n729 = ~n724 & ~n728 ;
  assign n730 = n152 & ~n729 ;
  assign n731 = ~d_pad & ~n143 ;
  assign n732 = ~l_pad & n143 ;
  assign n733 = ~n731 & ~n732 ;
  assign n734 = n171 & n733 ;
  assign n736 = ~\o2_pad  & n164 ;
  assign n735 = ~\n2_pad  & ~n164 ;
  assign n737 = ~n171 & ~n735 ;
  assign n738 = ~n736 & n737 ;
  assign n739 = ~n734 & ~n738 ;
  assign n740 = n152 & ~n739 ;
  assign n742 = ~\o3_pad  & n204 ;
  assign n741 = ~\n3_pad  & ~n204 ;
  assign n743 = n152 & ~n741 ;
  assign n744 = ~n742 & n743 ;
  assign n745 = \m6_pad  & n152 ;
  assign n746 = ~n198 & n745 ;
  assign n748 = ~\g3_pad  & n145 ;
  assign n747 = ~\o3_pad  & ~n145 ;
  assign n749 = \m0_pad  & ~n747 ;
  assign n750 = ~n748 & n749 ;
  assign n751 = \h1_pad  & n150 ;
  assign n752 = \i0_pad  & n157 ;
  assign n754 = ~\p1_pad  & n164 ;
  assign n753 = ~\o1_pad  & ~n164 ;
  assign n755 = ~n157 & ~n753 ;
  assign n756 = ~n754 & n755 ;
  assign n757 = ~n752 & ~n756 ;
  assign n758 = n152 & ~n757 ;
  assign n759 = ~e_pad & ~n143 ;
  assign n760 = ~m_pad & n143 ;
  assign n761 = ~n759 & ~n760 ;
  assign n762 = n171 & n761 ;
  assign n764 = ~\p2_pad  & n164 ;
  assign n763 = ~\o2_pad  & ~n164 ;
  assign n765 = ~n171 & ~n763 ;
  assign n766 = ~n764 & n765 ;
  assign n767 = ~n762 & ~n766 ;
  assign n768 = n152 & ~n767 ;
  assign n770 = ~\p3_pad  & n204 ;
  assign n769 = ~\o3_pad  & ~n204 ;
  assign n771 = n152 & ~n769 ;
  assign n772 = ~n770 & n771 ;
  assign n774 = ~\h3_pad  & n145 ;
  assign n773 = ~\p3_pad  & ~n145 ;
  assign n775 = \m0_pad  & ~n773 ;
  assign n776 = ~n774 & n775 ;
  assign n777 = \i1_pad  & n150 ;
  assign n778 = \h0_pad  & n157 ;
  assign n780 = ~\q1_pad  & n164 ;
  assign n779 = ~\p1_pad  & ~n164 ;
  assign n781 = ~n157 & ~n779 ;
  assign n782 = ~n780 & n781 ;
  assign n783 = ~n778 & ~n782 ;
  assign n784 = n152 & ~n783 ;
  assign n785 = ~f_pad & ~n143 ;
  assign n786 = ~n_pad & n143 ;
  assign n787 = ~n785 & ~n786 ;
  assign n788 = n171 & n787 ;
  assign n790 = ~\q2_pad  & n164 ;
  assign n789 = ~\p2_pad  & ~n164 ;
  assign n791 = ~n171 & ~n789 ;
  assign n792 = ~n790 & n791 ;
  assign n793 = ~n788 & ~n792 ;
  assign n794 = n152 & ~n793 ;
  assign n796 = ~\q3_pad  & n204 ;
  assign n795 = ~\p3_pad  & ~n204 ;
  assign n797 = n152 & ~n795 ;
  assign n798 = ~n796 & n797 ;
  assign n800 = ~\i3_pad  & n145 ;
  assign n799 = ~\q3_pad  & ~n145 ;
  assign n801 = \m0_pad  & ~n799 ;
  assign n802 = ~n800 & n801 ;
  assign n803 = \j1_pad  & n150 ;
  assign n804 = \g0_pad  & n157 ;
  assign n806 = ~\r1_pad  & n164 ;
  assign n805 = ~\q1_pad  & ~n164 ;
  assign n807 = ~n157 & ~n805 ;
  assign n808 = ~n806 & n807 ;
  assign n809 = ~n804 & ~n808 ;
  assign n810 = n152 & ~n809 ;
  assign n811 = ~g_pad & ~n143 ;
  assign n812 = ~o_pad & n143 ;
  assign n813 = ~n811 & ~n812 ;
  assign n814 = n171 & n813 ;
  assign n816 = ~\r2_pad  & n164 ;
  assign n815 = ~\q2_pad  & ~n164 ;
  assign n817 = ~n171 & ~n815 ;
  assign n818 = ~n816 & n817 ;
  assign n819 = ~n814 & ~n818 ;
  assign n820 = n152 & ~n819 ;
  assign n822 = ~\r3_pad  & n204 ;
  assign n821 = ~\q3_pad  & ~n204 ;
  assign n823 = n152 & ~n821 ;
  assign n824 = ~n822 & n823 ;
  assign \a5_pad  = n149 ;
  assign \a6_pad  = ~n151 ;
  assign \a7_pad  = n170 ;
  assign \a8_pad  = n181 ;
  assign \a9_pad  = n208 ;
  assign \b5_pad  = n212 ;
  assign \b6_pad  = ~n213 ;
  assign \b7_pad  = n220 ;
  assign \b8_pad  = n228 ;
  assign \b9_pad  = n232 ;
  assign \c5_pad  = n236 ;
  assign \c6_pad  = ~n237 ;
  assign \c7_pad  = n244 ;
  assign \c8_pad  = n251 ;
  assign \c9_pad  = n255 ;
  assign \d5_pad  = n256 ;
  assign \d6_pad  = ~n257 ;
  assign \d7_pad  = n263 ;
  assign \d8_pad  = n270 ;
  assign \d9_pad  = n274 ;
  assign \e5_pad  = n275 ;
  assign \e6_pad  = ~n276 ;
  assign \e7_pad  = n283 ;
  assign \e8_pad  = n290 ;
  assign \e9_pad  = n294 ;
  assign \f5_pad  = n295 ;
  assign \f6_pad  = ~n296 ;
  assign \f7_pad  = n303 ;
  assign \f8_pad  = n310 ;
  assign \f9_pad  = n332 ;
  assign \g5_pad  = n333 ;
  assign \g6_pad  = ~n334 ;
  assign \g7_pad  = n341 ;
  assign \g8_pad  = n348 ;
  assign \g9_pad  = n354 ;
  assign \h5_pad  = n355 ;
  assign \h6_pad  = ~\h1_pad  ;
  assign \h7_pad  = n362 ;
  assign \h8_pad  = n369 ;
  assign \h9_pad  = ~n373 ;
  assign \i5_pad  = n374 ;
  assign \i6_pad  = ~\i1_pad  ;
  assign \i7_pad  = n381 ;
  assign \i8_pad  = n386 ;
  assign \i9_pad  = ~n391 ;
  assign \j5_pad  = n392 ;
  assign \j6_pad  = ~\j1_pad  ;
  assign \j7_pad  = n399 ;
  assign \j8_pad  = n403 ;
  assign \j9_pad  = n410 ;
  assign \k5_pad  = n411 ;
  assign \k6_pad  = ~\k1_pad  ;
  assign \k7_pad  = n418 ;
  assign \k8_pad  = n422 ;
  assign \k9_pad  = n427 ;
  assign \l5_pad  = n428 ;
  assign \l6_pad  = ~\l1_pad  ;
  assign \l7_pad  = n435 ;
  assign \l8_pad  = n439 ;
  assign \l9_pad  = n442 ;
  assign \m7_pad  = n449 ;
  assign \m8_pad  = n453 ;
  assign \m9_pad  = n461 ;
  assign \n5_pad  = ~n463 ;
  assign \n6_pad  = ~n466 ;
  assign \n7_pad  = n473 ;
  assign \n8_pad  = n477 ;
  assign \n9_pad  = ~n485 ;
  assign \o4_pad  = ~\g1_pad  ;
  assign \o5_pad  = ~n487 ;
  assign \o6_pad  = n488 ;
  assign \o7_pad  = n495 ;
  assign \o8_pad  = n499 ;
  assign \o9_pad  = ~n504 ;
  assign \p4_pad  = n510 ;
  assign \p5_pad  = ~n512 ;
  assign \p6_pad  = n518 ;
  assign \p7_pad  = n525 ;
  assign \p8_pad  = n529 ;
  assign \p9_pad  = ~n542 ;
  assign \q4_pad  = n548 ;
  assign \q5_pad  = ~n550 ;
  assign \q6_pad  = ~n556 ;
  assign \q7_pad  = n563 ;
  assign \q8_pad  = n567 ;
  assign \q9_pad  = ~n572 ;
  assign \r4_pad  = n578 ;
  assign \r5_pad  = ~n580 ;
  assign \r6_pad  = n588 ;
  assign \r7_pad  = n595 ;
  assign \r8_pad  = n599 ;
  assign \r9_pad  = n604 ;
  assign \s4_pad  = n610 ;
  assign \s6_pad  = n615 ;
  assign \s7_pad  = n622 ;
  assign \s8_pad  = n626 ;
  assign \s9_pad  = ~n649 ;
  assign \t6_pad  = n655 ;
  assign \t7_pad  = n665 ;
  assign \t8_pad  = n669 ;
  assign \t9_pad  = n671 ;
  assign \u6_pad  = n676 ;
  assign \u7_pad  = n686 ;
  assign \u8_pad  = n690 ;
  assign \u9_pad  = n691 ;
  assign \v4_pad  = n695 ;
  assign \v6_pad  = n700 ;
  assign \v7_pad  = n710 ;
  assign \v8_pad  = n714 ;
  assign \v9_pad  = n716 ;
  assign \w4_pad  = n720 ;
  assign \w5_pad  = ~n723 ;
  assign \w6_pad  = n730 ;
  assign \w7_pad  = n740 ;
  assign \w8_pad  = n744 ;
  assign \w9_pad  = n746 ;
  assign \x4_pad  = n750 ;
  assign \x5_pad  = ~n751 ;
  assign \x6_pad  = n758 ;
  assign \x7_pad  = n768 ;
  assign \x8_pad  = n772 ;
  assign \y4_pad  = n776 ;
  assign \y5_pad  = ~n777 ;
  assign \y6_pad  = n784 ;
  assign \y7_pad  = n794 ;
  assign \y8_pad  = n798 ;
  assign \z4_pad  = n802 ;
  assign \z5_pad  = ~n803 ;
  assign \z6_pad  = n810 ;
  assign \z7_pad  = n820 ;
  assign \z8_pad  = n824 ;
endmodule
