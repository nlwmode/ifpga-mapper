module top (\101GAT(25)_pad , \106GAT(26)_pad , \111GAT(27)_pad , \116GAT(28)_pad , \121GAT(29)_pad , \126GAT(30)_pad , \130GAT(31)_pad , \135GAT(32)_pad , \138GAT(33)_pad , \13GAT(2)_pad , \143GAT(34)_pad , \146GAT(35)_pad , \149GAT(36)_pad , \152GAT(37)_pad , \153GAT(38)_pad , \156GAT(39)_pad , \159GAT(40)_pad , \165GAT(41)_pad , \171GAT(42)_pad , \177GAT(43)_pad , \17GAT(3)_pad , \183GAT(44)_pad , \189GAT(45)_pad , \195GAT(46)_pad , \1GAT(0)_pad , \201GAT(47)_pad , \207GAT(48)_pad , \210GAT(49)_pad , \219GAT(50)_pad , \228GAT(51)_pad , \237GAT(52)_pad , \246GAT(53)_pad , \255GAT(54)_pad , \259GAT(55)_pad , \260GAT(56)_pad , \261GAT(57)_pad , \267GAT(58)_pad , \268GAT(59)_pad , \26GAT(4)_pad , \29GAT(5)_pad , \36GAT(6)_pad , \42GAT(7)_pad , \51GAT(8)_pad , \55GAT(9)_pad , \59GAT(10)_pad , \68GAT(11)_pad , \72GAT(12)_pad , \73GAT(13)_pad , \74GAT(14)_pad , \75GAT(15)_pad , \80GAT(16)_pad , \85GAT(17)_pad , \86GAT(18)_pad , \87GAT(19)_pad , \88GAT(20)_pad , \89GAT(21)_pad , \8GAT(1)_pad , \90GAT(22)_pad , \91GAT(23)_pad , \96GAT(24)_pad , \273GAT(103) , \388GAT(133)_pad , \389GAT(132)_pad , \391GAT(124)_pad , \393GAT(165) , \418GAT(168)_pad , \419GAT(164)_pad , \420GAT(158)_pad , \421GAT(162)_pad , \422GAT(161)_pad , \423GAT(155)_pad , \446GAT(183)_pad , \448GAT(179)_pad , \449GAT(176)_pad , \450GAT(173)_pad , \767GAT(349)_pad , \768GAT(334)_pad , \811GAT(378) , \837GAT(396) , \838GAT(395) , \839GAT(394) , \854GAT(419) , \866GAT(426)_pad , \867GAT(432) , \868GAT(431) , \869GAT(430) );
	input \101GAT(25)_pad  ;
	input \106GAT(26)_pad  ;
	input \111GAT(27)_pad  ;
	input \116GAT(28)_pad  ;
	input \121GAT(29)_pad  ;
	input \126GAT(30)_pad  ;
	input \130GAT(31)_pad  ;
	input \135GAT(32)_pad  ;
	input \138GAT(33)_pad  ;
	input \13GAT(2)_pad  ;
	input \143GAT(34)_pad  ;
	input \146GAT(35)_pad  ;
	input \149GAT(36)_pad  ;
	input \152GAT(37)_pad  ;
	input \153GAT(38)_pad  ;
	input \156GAT(39)_pad  ;
	input \159GAT(40)_pad  ;
	input \165GAT(41)_pad  ;
	input \171GAT(42)_pad  ;
	input \177GAT(43)_pad  ;
	input \17GAT(3)_pad  ;
	input \183GAT(44)_pad  ;
	input \189GAT(45)_pad  ;
	input \195GAT(46)_pad  ;
	input \1GAT(0)_pad  ;
	input \201GAT(47)_pad  ;
	input \207GAT(48)_pad  ;
	input \210GAT(49)_pad  ;
	input \219GAT(50)_pad  ;
	input \228GAT(51)_pad  ;
	input \237GAT(52)_pad  ;
	input \246GAT(53)_pad  ;
	input \255GAT(54)_pad  ;
	input \259GAT(55)_pad  ;
	input \260GAT(56)_pad  ;
	input \261GAT(57)_pad  ;
	input \267GAT(58)_pad  ;
	input \268GAT(59)_pad  ;
	input \26GAT(4)_pad  ;
	input \29GAT(5)_pad  ;
	input \36GAT(6)_pad  ;
	input \42GAT(7)_pad  ;
	input \51GAT(8)_pad  ;
	input \55GAT(9)_pad  ;
	input \59GAT(10)_pad  ;
	input \68GAT(11)_pad  ;
	input \72GAT(12)_pad  ;
	input \73GAT(13)_pad  ;
	input \74GAT(14)_pad  ;
	input \75GAT(15)_pad  ;
	input \80GAT(16)_pad  ;
	input \85GAT(17)_pad  ;
	input \86GAT(18)_pad  ;
	input \87GAT(19)_pad  ;
	input \88GAT(20)_pad  ;
	input \89GAT(21)_pad  ;
	input \8GAT(1)_pad  ;
	input \90GAT(22)_pad  ;
	input \91GAT(23)_pad  ;
	input \96GAT(24)_pad  ;
	output \273GAT(103)  ;
	output \388GAT(133)_pad  ;
	output \389GAT(132)_pad  ;
	output \391GAT(124)_pad  ;
	output \393GAT(165)  ;
	output \418GAT(168)_pad  ;
	output \419GAT(164)_pad  ;
	output \420GAT(158)_pad  ;
	output \421GAT(162)_pad  ;
	output \422GAT(161)_pad  ;
	output \423GAT(155)_pad  ;
	output \446GAT(183)_pad  ;
	output \448GAT(179)_pad  ;
	output \449GAT(176)_pad  ;
	output \450GAT(173)_pad  ;
	output \767GAT(349)_pad  ;
	output \768GAT(334)_pad  ;
	output \811GAT(378)  ;
	output \837GAT(396)  ;
	output \838GAT(395)  ;
	output \839GAT(394)  ;
	output \854GAT(419)  ;
	output \866GAT(426)_pad  ;
	output \867GAT(432)  ;
	output \868GAT(431)  ;
	output \869GAT(430)  ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	LUT3 #(
		.INIT('h80)
	) name0 (
		\29GAT(5)_pad ,
		\36GAT(6)_pad ,
		\42GAT(7)_pad ,
		_w62_
	);
	LUT3 #(
		.INIT('h80)
	) name1 (
		\29GAT(5)_pad ,
		\42GAT(7)_pad ,
		\75GAT(15)_pad ,
		_w63_
	);
	LUT3 #(
		.INIT('h80)
	) name2 (
		\29GAT(5)_pad ,
		\36GAT(6)_pad ,
		\80GAT(16)_pad ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\85GAT(17)_pad ,
		\86GAT(18)_pad ,
		_w65_
	);
	LUT3 #(
		.INIT('h80)
	) name4 (
		\1GAT(0)_pad ,
		\26GAT(4)_pad ,
		\51GAT(8)_pad ,
		_w66_
	);
	LUT4 #(
		.INIT('h8000)
	) name5 (
		\13GAT(2)_pad ,
		\17GAT(3)_pad ,
		\1GAT(0)_pad ,
		\8GAT(1)_pad ,
		_w67_
	);
	LUT4 #(
		.INIT('h8000)
	) name6 (
		\13GAT(2)_pad ,
		\17GAT(3)_pad ,
		\1GAT(0)_pad ,
		\26GAT(4)_pad ,
		_w68_
	);
	LUT2 #(
		.INIT('hb)
	) name7 (
		_w62_,
		_w68_,
		_w69_
	);
	LUT3 #(
		.INIT('h7f)
	) name8 (
		\59GAT(10)_pad ,
		\75GAT(15)_pad ,
		\80GAT(16)_pad ,
		_w70_
	);
	LUT3 #(
		.INIT('h7f)
	) name9 (
		\36GAT(6)_pad ,
		\59GAT(10)_pad ,
		\80GAT(16)_pad ,
		_w71_
	);
	LUT3 #(
		.INIT('h7f)
	) name10 (
		\36GAT(6)_pad ,
		\42GAT(7)_pad ,
		\59GAT(10)_pad ,
		_w72_
	);
	LUT3 #(
		.INIT('he0)
	) name11 (
		\87GAT(19)_pad ,
		\88GAT(20)_pad ,
		\90GAT(22)_pad ,
		_w73_
	);
	LUT2 #(
		.INIT('h7)
	) name12 (
		_w62_,
		_w68_,
		_w74_
	);
	LUT4 #(
		.INIT('h8000)
	) name13 (
		\13GAT(2)_pad ,
		\1GAT(0)_pad ,
		\55GAT(9)_pad ,
		\8GAT(1)_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\29GAT(5)_pad ,
		\68GAT(11)_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\59GAT(10)_pad ,
		\68GAT(11)_pad ,
		_w78_
	);
	LUT3 #(
		.INIT('h80)
	) name17 (
		\74GAT(14)_pad ,
		_w75_,
		_w78_,
		_w79_
	);
	LUT3 #(
		.INIT('he0)
	) name18 (
		\87GAT(19)_pad ,
		\88GAT(20)_pad ,
		\89GAT(21)_pad ,
		_w80_
	);
	LUT4 #(
		.INIT('h6996)
	) name19 (
		\111GAT(27)_pad ,
		\126GAT(30)_pad ,
		\91GAT(23)_pad ,
		\96GAT(24)_pad ,
		_w81_
	);
	LUT4 #(
		.INIT('h9669)
	) name20 (
		\101GAT(25)_pad ,
		\116GAT(28)_pad ,
		\121GAT(29)_pad ,
		\135GAT(32)_pad ,
		_w82_
	);
	LUT2 #(
		.INIT('h9)
	) name21 (
		\106GAT(26)_pad ,
		\130GAT(31)_pad ,
		_w83_
	);
	LUT3 #(
		.INIT('h96)
	) name22 (
		_w81_,
		_w82_,
		_w83_,
		_w84_
	);
	LUT4 #(
		.INIT('h6996)
	) name23 (
		\130GAT(31)_pad ,
		\171GAT(42)_pad ,
		\177GAT(43)_pad ,
		\183GAT(44)_pad ,
		_w85_
	);
	LUT4 #(
		.INIT('h9669)
	) name24 (
		\159GAT(40)_pad ,
		\189GAT(45)_pad ,
		\195GAT(46)_pad ,
		\207GAT(48)_pad ,
		_w86_
	);
	LUT2 #(
		.INIT('h9)
	) name25 (
		\165GAT(41)_pad ,
		\201GAT(47)_pad ,
		_w87_
	);
	LUT3 #(
		.INIT('h96)
	) name26 (
		_w85_,
		_w86_,
		_w87_,
		_w88_
	);
	LUT3 #(
		.INIT('h80)
	) name27 (
		\42GAT(7)_pad ,
		\59GAT(10)_pad ,
		\75GAT(15)_pad ,
		_w89_
	);
	LUT4 #(
		.INIT('h8000)
	) name28 (
		\17GAT(3)_pad ,
		\1GAT(0)_pad ,
		\51GAT(8)_pad ,
		\8GAT(1)_pad ,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		_w89_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h9)
	) name30 (
		\17GAT(3)_pad ,
		\42GAT(7)_pad ,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\156GAT(39)_pad ,
		\59GAT(10)_pad ,
		_w93_
	);
	LUT3 #(
		.INIT('h08)
	) name32 (
		_w66_,
		_w93_,
		_w92_,
		_w94_
	);
	LUT3 #(
		.INIT('ha8)
	) name33 (
		\126GAT(30)_pad ,
		_w91_,
		_w94_,
		_w95_
	);
	LUT4 #(
		.INIT('h8000)
	) name34 (
		\1GAT(0)_pad ,
		\26GAT(4)_pad ,
		\51GAT(8)_pad ,
		\55GAT(9)_pad ,
		_w96_
	);
	LUT4 #(
		.INIT('h4000)
	) name35 (
		\268GAT(59)_pad ,
		\29GAT(5)_pad ,
		\75GAT(15)_pad ,
		\80GAT(16)_pad ,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h8000)
	) name37 (
		\17GAT(3)_pad ,
		\1GAT(0)_pad ,
		\26GAT(4)_pad ,
		\51GAT(8)_pad ,
		_w99_
	);
	LUT4 #(
		.INIT('h2a22)
	) name38 (
		\153GAT(38)_pad ,
		\1GAT(0)_pad ,
		_w93_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w98_,
		_w100_,
		_w101_
	);
	LUT4 #(
		.INIT('h4844)
	) name40 (
		\201GAT(47)_pad ,
		\261GAT(57)_pad ,
		_w95_,
		_w101_,
		_w102_
	);
	LUT4 #(
		.INIT('h2122)
	) name41 (
		\201GAT(47)_pad ,
		\261GAT(57)_pad ,
		_w95_,
		_w101_,
		_w103_
	);
	LUT3 #(
		.INIT('h02)
	) name42 (
		\219GAT(50)_pad ,
		_w103_,
		_w102_,
		_w104_
	);
	LUT4 #(
		.INIT('h4844)
	) name43 (
		\201GAT(47)_pad ,
		\228GAT(51)_pad ,
		_w95_,
		_w101_,
		_w105_
	);
	LUT3 #(
		.INIT('h07)
	) name44 (
		\201GAT(47)_pad ,
		\237GAT(52)_pad ,
		\246GAT(53)_pad ,
		_w106_
	);
	LUT3 #(
		.INIT('h80)
	) name45 (
		\42GAT(7)_pad ,
		\72GAT(12)_pad ,
		\73GAT(13)_pad ,
		_w107_
	);
	LUT4 #(
		.INIT('h8000)
	) name46 (
		\201GAT(47)_pad ,
		_w75_,
		_w78_,
		_w107_,
		_w108_
	);
	LUT4 #(
		.INIT('h0777)
	) name47 (
		\121GAT(29)_pad ,
		\210GAT(49)_pad ,
		\255GAT(54)_pad ,
		\267GAT(58)_pad ,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w108_,
		_w109_,
		_w110_
	);
	LUT4 #(
		.INIT('hf400)
	) name49 (
		_w95_,
		_w101_,
		_w106_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w105_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('hb)
	) name51 (
		_w104_,
		_w112_,
		_w113_
	);
	LUT3 #(
		.INIT('ha8)
	) name52 (
		\111GAT(27)_pad ,
		_w91_,
		_w94_,
		_w114_
	);
	LUT4 #(
		.INIT('h2a22)
	) name53 (
		\143GAT(34)_pad ,
		\1GAT(0)_pad ,
		_w93_,
		_w99_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w98_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w114_,
		_w116_,
		_w117_
	);
	LUT3 #(
		.INIT('h65)
	) name56 (
		\183GAT(44)_pad ,
		_w114_,
		_w116_,
		_w118_
	);
	LUT3 #(
		.INIT('ha8)
	) name57 (
		\121GAT(29)_pad ,
		_w91_,
		_w94_,
		_w119_
	);
	LUT4 #(
		.INIT('h2a22)
	) name58 (
		\149GAT(36)_pad ,
		\1GAT(0)_pad ,
		_w93_,
		_w99_,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w98_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w119_,
		_w121_,
		_w122_
	);
	LUT4 #(
		.INIT('h1711)
	) name61 (
		\201GAT(47)_pad ,
		\261GAT(57)_pad ,
		_w95_,
		_w101_,
		_w123_
	);
	LUT3 #(
		.INIT('ha8)
	) name62 (
		\116GAT(28)_pad ,
		_w91_,
		_w94_,
		_w124_
	);
	LUT4 #(
		.INIT('h2a22)
	) name63 (
		\146GAT(35)_pad ,
		\1GAT(0)_pad ,
		_w93_,
		_w99_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w98_,
		_w125_,
		_w126_
	);
	LUT3 #(
		.INIT('h10)
	) name65 (
		\189GAT(45)_pad ,
		_w124_,
		_w126_,
		_w127_
	);
	LUT4 #(
		.INIT('h002b)
	) name66 (
		\195GAT(46)_pad ,
		_w122_,
		_w123_,
		_w127_,
		_w128_
	);
	LUT3 #(
		.INIT('h8a)
	) name67 (
		\189GAT(45)_pad ,
		_w124_,
		_w126_,
		_w129_
	);
	LUT4 #(
		.INIT('h2228)
	) name68 (
		\219GAT(50)_pad ,
		_w118_,
		_w128_,
		_w129_,
		_w130_
	);
	LUT4 #(
		.INIT('h4844)
	) name69 (
		\183GAT(44)_pad ,
		\228GAT(51)_pad ,
		_w114_,
		_w116_,
		_w131_
	);
	LUT3 #(
		.INIT('h07)
	) name70 (
		\183GAT(44)_pad ,
		\237GAT(52)_pad ,
		\246GAT(53)_pad ,
		_w132_
	);
	LUT4 #(
		.INIT('h8000)
	) name71 (
		\183GAT(44)_pad ,
		_w75_,
		_w78_,
		_w107_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\106GAT(26)_pad ,
		\210GAT(49)_pad ,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w133_,
		_w134_,
		_w135_
	);
	LUT4 #(
		.INIT('hf400)
	) name74 (
		_w114_,
		_w116_,
		_w132_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		_w131_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('hb)
	) name76 (
		_w130_,
		_w137_,
		_w138_
	);
	LUT3 #(
		.INIT('h65)
	) name77 (
		\189GAT(45)_pad ,
		_w124_,
		_w126_,
		_w139_
	);
	LUT3 #(
		.INIT('hd4)
	) name78 (
		\195GAT(46)_pad ,
		_w122_,
		_w123_,
		_w140_
	);
	LUT4 #(
		.INIT('h4844)
	) name79 (
		\189GAT(45)_pad ,
		\228GAT(51)_pad ,
		_w124_,
		_w126_,
		_w141_
	);
	LUT3 #(
		.INIT('h07)
	) name80 (
		\189GAT(45)_pad ,
		\237GAT(52)_pad ,
		\246GAT(53)_pad ,
		_w142_
	);
	LUT4 #(
		.INIT('h8000)
	) name81 (
		\189GAT(45)_pad ,
		_w75_,
		_w78_,
		_w107_,
		_w143_
	);
	LUT4 #(
		.INIT('h0777)
	) name82 (
		\111GAT(27)_pad ,
		\210GAT(49)_pad ,
		\255GAT(54)_pad ,
		\259GAT(55)_pad ,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w143_,
		_w144_,
		_w145_
	);
	LUT4 #(
		.INIT('hf400)
	) name84 (
		_w124_,
		_w126_,
		_w142_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w141_,
		_w146_,
		_w147_
	);
	LUT4 #(
		.INIT('h82ff)
	) name86 (
		\219GAT(50)_pad ,
		_w139_,
		_w140_,
		_w147_,
		_w148_
	);
	LUT3 #(
		.INIT('h65)
	) name87 (
		\195GAT(46)_pad ,
		_w119_,
		_w121_,
		_w149_
	);
	LUT3 #(
		.INIT('h82)
	) name88 (
		\219GAT(50)_pad ,
		_w123_,
		_w149_,
		_w150_
	);
	LUT4 #(
		.INIT('h4844)
	) name89 (
		\195GAT(46)_pad ,
		\228GAT(51)_pad ,
		_w119_,
		_w121_,
		_w151_
	);
	LUT3 #(
		.INIT('h07)
	) name90 (
		\195GAT(46)_pad ,
		\237GAT(52)_pad ,
		\246GAT(53)_pad ,
		_w152_
	);
	LUT4 #(
		.INIT('h8000)
	) name91 (
		\195GAT(46)_pad ,
		_w75_,
		_w78_,
		_w107_,
		_w153_
	);
	LUT4 #(
		.INIT('h0777)
	) name92 (
		\116GAT(28)_pad ,
		\210GAT(49)_pad ,
		\255GAT(54)_pad ,
		\260GAT(56)_pad ,
		_w154_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT4 #(
		.INIT('hf400)
	) name94 (
		_w119_,
		_w121_,
		_w152_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w151_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('hb)
	) name96 (
		_w150_,
		_w157_,
		_w158_
	);
	LUT3 #(
		.INIT('ha8)
	) name97 (
		\106GAT(26)_pad ,
		_w91_,
		_w94_,
		_w159_
	);
	LUT3 #(
		.INIT('h20)
	) name98 (
		\153GAT(38)_pad ,
		_w93_,
		_w96_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\138GAT(33)_pad ,
		\152GAT(37)_pad ,
		_w161_
	);
	LUT3 #(
		.INIT('h07)
	) name100 (
		_w97_,
		_w99_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w160_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w159_,
		_w163_,
		_w164_
	);
	LUT3 #(
		.INIT('h65)
	) name103 (
		\177GAT(43)_pad ,
		_w159_,
		_w163_,
		_w165_
	);
	LUT4 #(
		.INIT('h444d)
	) name104 (
		\183GAT(44)_pad ,
		_w117_,
		_w128_,
		_w129_,
		_w166_
	);
	LUT4 #(
		.INIT('h4844)
	) name105 (
		\177GAT(43)_pad ,
		\228GAT(51)_pad ,
		_w159_,
		_w163_,
		_w167_
	);
	LUT3 #(
		.INIT('h07)
	) name106 (
		\177GAT(43)_pad ,
		\237GAT(52)_pad ,
		\246GAT(53)_pad ,
		_w168_
	);
	LUT4 #(
		.INIT('h8000)
	) name107 (
		\177GAT(43)_pad ,
		_w75_,
		_w78_,
		_w107_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\101GAT(25)_pad ,
		\210GAT(49)_pad ,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w169_,
		_w170_,
		_w171_
	);
	LUT4 #(
		.INIT('hf400)
	) name110 (
		_w159_,
		_w163_,
		_w168_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w167_,
		_w172_,
		_w173_
	);
	LUT4 #(
		.INIT('h82ff)
	) name112 (
		\219GAT(50)_pad ,
		_w165_,
		_w166_,
		_w173_,
		_w174_
	);
	LUT3 #(
		.INIT('ha8)
	) name113 (
		\91GAT(23)_pad ,
		_w91_,
		_w94_,
		_w175_
	);
	LUT3 #(
		.INIT('h20)
	) name114 (
		\143GAT(34)_pad ,
		_w93_,
		_w96_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\138GAT(33)_pad ,
		\8GAT(1)_pad ,
		_w177_
	);
	LUT3 #(
		.INIT('h07)
	) name116 (
		_w97_,
		_w99_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w176_,
		_w178_,
		_w179_
	);
	LUT3 #(
		.INIT('h8a)
	) name118 (
		\159GAT(40)_pad ,
		_w175_,
		_w179_,
		_w180_
	);
	LUT3 #(
		.INIT('h10)
	) name119 (
		\159GAT(40)_pad ,
		_w175_,
		_w179_,
		_w181_
	);
	LUT3 #(
		.INIT('ha8)
	) name120 (
		\101GAT(25)_pad ,
		_w91_,
		_w94_,
		_w182_
	);
	LUT3 #(
		.INIT('h20)
	) name121 (
		\149GAT(36)_pad ,
		_w93_,
		_w96_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\138GAT(33)_pad ,
		\17GAT(3)_pad ,
		_w184_
	);
	LUT3 #(
		.INIT('h07)
	) name123 (
		_w97_,
		_w99_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		_w183_,
		_w185_,
		_w186_
	);
	LUT3 #(
		.INIT('h8a)
	) name125 (
		\171GAT(42)_pad ,
		_w182_,
		_w186_,
		_w187_
	);
	LUT3 #(
		.INIT('hd4)
	) name126 (
		\177GAT(43)_pad ,
		_w164_,
		_w166_,
		_w188_
	);
	LUT4 #(
		.INIT('h00d4)
	) name127 (
		\177GAT(43)_pad ,
		_w164_,
		_w166_,
		_w187_,
		_w189_
	);
	LUT3 #(
		.INIT('h10)
	) name128 (
		\171GAT(42)_pad ,
		_w182_,
		_w186_,
		_w190_
	);
	LUT3 #(
		.INIT('ha8)
	) name129 (
		\96GAT(24)_pad ,
		_w91_,
		_w94_,
		_w191_
	);
	LUT3 #(
		.INIT('h20)
	) name130 (
		\146GAT(35)_pad ,
		_w93_,
		_w96_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\138GAT(33)_pad ,
		\51GAT(8)_pad ,
		_w193_
	);
	LUT3 #(
		.INIT('h07)
	) name132 (
		_w97_,
		_w99_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		_w192_,
		_w194_,
		_w195_
	);
	LUT3 #(
		.INIT('h10)
	) name134 (
		\165GAT(41)_pad ,
		_w191_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w190_,
		_w196_,
		_w197_
	);
	LUT3 #(
		.INIT('h8a)
	) name136 (
		\165GAT(41)_pad ,
		_w191_,
		_w195_,
		_w198_
	);
	LUT3 #(
		.INIT('h0b)
	) name137 (
		_w189_,
		_w197_,
		_w198_,
		_w199_
	);
	LUT4 #(
		.INIT('h5510)
	) name138 (
		_w181_,
		_w189_,
		_w197_,
		_w198_,
		_w200_
	);
	LUT2 #(
		.INIT('he)
	) name139 (
		_w180_,
		_w200_,
		_w201_
	);
	LUT3 #(
		.INIT('h65)
	) name140 (
		\159GAT(40)_pad ,
		_w175_,
		_w179_,
		_w202_
	);
	LUT4 #(
		.INIT('h4844)
	) name141 (
		\159GAT(40)_pad ,
		\228GAT(51)_pad ,
		_w175_,
		_w179_,
		_w203_
	);
	LUT3 #(
		.INIT('h07)
	) name142 (
		\159GAT(40)_pad ,
		\237GAT(52)_pad ,
		\246GAT(53)_pad ,
		_w204_
	);
	LUT4 #(
		.INIT('h8000)
	) name143 (
		\159GAT(40)_pad ,
		_w75_,
		_w78_,
		_w107_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\210GAT(49)_pad ,
		\268GAT(59)_pad ,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w205_,
		_w206_,
		_w207_
	);
	LUT4 #(
		.INIT('hf400)
	) name146 (
		_w175_,
		_w179_,
		_w204_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		_w203_,
		_w208_,
		_w209_
	);
	LUT4 #(
		.INIT('h82ff)
	) name148 (
		\219GAT(50)_pad ,
		_w199_,
		_w202_,
		_w209_,
		_w210_
	);
	LUT3 #(
		.INIT('h65)
	) name149 (
		\165GAT(41)_pad ,
		_w191_,
		_w195_,
		_w211_
	);
	LUT4 #(
		.INIT('h002b)
	) name150 (
		\177GAT(43)_pad ,
		_w164_,
		_w166_,
		_w190_,
		_w212_
	);
	LUT4 #(
		.INIT('h0a28)
	) name151 (
		\219GAT(50)_pad ,
		_w187_,
		_w211_,
		_w212_,
		_w213_
	);
	LUT4 #(
		.INIT('h4844)
	) name152 (
		\165GAT(41)_pad ,
		\228GAT(51)_pad ,
		_w191_,
		_w195_,
		_w214_
	);
	LUT3 #(
		.INIT('h07)
	) name153 (
		\165GAT(41)_pad ,
		\237GAT(52)_pad ,
		\246GAT(53)_pad ,
		_w215_
	);
	LUT4 #(
		.INIT('h8000)
	) name154 (
		\165GAT(41)_pad ,
		_w75_,
		_w78_,
		_w107_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\210GAT(49)_pad ,
		\91GAT(23)_pad ,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w216_,
		_w217_,
		_w218_
	);
	LUT4 #(
		.INIT('hf400)
	) name157 (
		_w191_,
		_w195_,
		_w215_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		_w214_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('hb)
	) name159 (
		_w213_,
		_w220_,
		_w221_
	);
	LUT3 #(
		.INIT('h65)
	) name160 (
		\171GAT(42)_pad ,
		_w182_,
		_w186_,
		_w222_
	);
	LUT4 #(
		.INIT('h4844)
	) name161 (
		\171GAT(42)_pad ,
		\228GAT(51)_pad ,
		_w182_,
		_w186_,
		_w223_
	);
	LUT3 #(
		.INIT('h07)
	) name162 (
		\171GAT(42)_pad ,
		\237GAT(52)_pad ,
		\246GAT(53)_pad ,
		_w224_
	);
	LUT4 #(
		.INIT('h8000)
	) name163 (
		\171GAT(42)_pad ,
		_w75_,
		_w78_,
		_w107_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\210GAT(49)_pad ,
		\96GAT(24)_pad ,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w225_,
		_w226_,
		_w227_
	);
	LUT4 #(
		.INIT('hf400)
	) name166 (
		_w182_,
		_w186_,
		_w224_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		_w223_,
		_w228_,
		_w229_
	);
	LUT4 #(
		.INIT('h82ff)
	) name168 (
		\219GAT(50)_pad ,
		_w188_,
		_w222_,
		_w229_,
		_w230_
	);
	assign \273GAT(103)  = _w62_ ;
	assign \388GAT(133)_pad  = _w63_ ;
	assign \389GAT(132)_pad  = _w64_ ;
	assign \391GAT(124)_pad  = _w65_ ;
	assign \393GAT(165)  = _w66_ ;
	assign \418GAT(168)_pad  = _w67_ ;
	assign \419GAT(164)_pad  = _w69_ ;
	assign \420GAT(158)_pad  = _w70_ ;
	assign \421GAT(162)_pad  = _w71_ ;
	assign \422GAT(161)_pad  = _w72_ ;
	assign \423GAT(155)_pad  = _w73_ ;
	assign \446GAT(183)_pad  = _w74_ ;
	assign \448GAT(179)_pad  = _w77_ ;
	assign \449GAT(176)_pad  = _w79_ ;
	assign \450GAT(173)_pad  = _w80_ ;
	assign \767GAT(349)_pad  = _w84_ ;
	assign \768GAT(334)_pad  = _w88_ ;
	assign \811GAT(378)  = _w113_ ;
	assign \837GAT(396)  = _w138_ ;
	assign \838GAT(395)  = _w148_ ;
	assign \839GAT(394)  = _w158_ ;
	assign \854GAT(419)  = _w174_ ;
	assign \866GAT(426)_pad  = _w201_ ;
	assign \867GAT(432)  = _w210_ ;
	assign \868GAT(431)  = _w221_ ;
	assign \869GAT(430)  = _w230_ ;
endmodule;