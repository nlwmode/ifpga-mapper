module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	output v_pad ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		j_pad,
		q_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		i_pad,
		q_pad,
		_w23_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		r_pad,
		_w22_,
		_w24_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		_w23_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		l_pad,
		q_pad,
		_w26_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		k_pad,
		q_pad,
		_w27_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		r_pad,
		_w26_,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w27_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w25_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		s_pad,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		p_pad,
		q_pad,
		_w32_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		o_pad,
		q_pad,
		_w33_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		r_pad,
		_w32_,
		_w34_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w33_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		n_pad,
		q_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		m_pad,
		q_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		r_pad,
		_w36_,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w37_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w35_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		s_pad,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		t_pad,
		_w31_,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w41_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		b_pad,
		q_pad,
		_w44_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		a_pad,
		q_pad,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		r_pad,
		_w44_,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		d_pad,
		q_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		c_pad,
		q_pad,
		_w49_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		r_pad,
		_w48_,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w47_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		s_pad,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		h_pad,
		q_pad,
		_w54_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		g_pad,
		q_pad,
		_w55_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		r_pad,
		_w54_,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		f_pad,
		q_pad,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		e_pad,
		q_pad,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		r_pad,
		_w58_,
		_w60_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		_w59_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w57_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		s_pad,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		t_pad,
		_w53_,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w63_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w43_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		u_pad,
		_w66_,
		_w67_
	);
	assign v_pad = _w67_ ;
endmodule;