module top( \G10_pad  , \G11_pad  , \G12_pad  , \G13_pad  , \G14_pad  , \G15_pad  , \G16_pad  , \G18_pad  , \G19_pad  , \G20_pad  , \G22_pad  , \G23_pad  , \G24_pad  , \G25_pad  , \G26_pad  , \G28_pad  , \G2_pad  , \G30_pad  , \G31_pad  , \G32_pad  , \G33_pad  , \G34_pad  , \G35_pad  , \G3_pad  , \G4_pad  , \G5_pad  , \G64_reg/NET0131  , \G65_reg/NET0131  , \G66_reg/NET0131  , \G69_reg/NET0131  , \G6_pad  , \G70_reg/NET0131  , \G71_reg/NET0131  , \G72_reg/NET0131  , \G73_reg/NET0131  , \G74_reg/NET0131  , \G75_reg/NET0131  , \G76_reg/NET0131  , \G77_reg/NET0131  , \G79_reg/NET0131  , \G81_reg/NET0131  , \G8_pad  , \G9_pad  , \G100BF_pad  , \G103BF_pad  , \G104BF_pad  , \G105BF_pad  , \G107_pad  , \G83_pad  , \G84_pad  , \G86BF_pad  , \G87BF_pad  , \G88BF_pad  , \G89BF_pad  , \G90_pad  , \G95BF_pad  , \G96BF_pad  , \G97BF_pad  , \G98BF_pad  , \G99BF_pad  , \_al_n0  , \_al_n1  , \g1049/_0_  , \g1081/_0_  , \g1115/_0_  , \g13/_1_  , \g809/_0_  , \g810/_0_  , \g814/_0_  , \g825/_2_  , \g834/_0_  , \g863/_0_  , \g870/_0_  , \g871/_0_  , \g916/_0_  , \g917/_0_  , \g940/_3_  );
  input \G10_pad  ;
  input \G11_pad  ;
  input \G12_pad  ;
  input \G13_pad  ;
  input \G14_pad  ;
  input \G15_pad  ;
  input \G16_pad  ;
  input \G18_pad  ;
  input \G19_pad  ;
  input \G20_pad  ;
  input \G22_pad  ;
  input \G23_pad  ;
  input \G24_pad  ;
  input \G25_pad  ;
  input \G26_pad  ;
  input \G28_pad  ;
  input \G2_pad  ;
  input \G30_pad  ;
  input \G31_pad  ;
  input \G32_pad  ;
  input \G33_pad  ;
  input \G34_pad  ;
  input \G35_pad  ;
  input \G3_pad  ;
  input \G4_pad  ;
  input \G5_pad  ;
  input \G64_reg/NET0131  ;
  input \G65_reg/NET0131  ;
  input \G66_reg/NET0131  ;
  input \G69_reg/NET0131  ;
  input \G6_pad  ;
  input \G70_reg/NET0131  ;
  input \G71_reg/NET0131  ;
  input \G72_reg/NET0131  ;
  input \G73_reg/NET0131  ;
  input \G74_reg/NET0131  ;
  input \G75_reg/NET0131  ;
  input \G76_reg/NET0131  ;
  input \G77_reg/NET0131  ;
  input \G79_reg/NET0131  ;
  input \G81_reg/NET0131  ;
  input \G8_pad  ;
  input \G9_pad  ;
  output \G100BF_pad  ;
  output \G103BF_pad  ;
  output \G104BF_pad  ;
  output \G105BF_pad  ;
  output \G107_pad  ;
  output \G83_pad  ;
  output \G84_pad  ;
  output \G86BF_pad  ;
  output \G87BF_pad  ;
  output \G88BF_pad  ;
  output \G89BF_pad  ;
  output \G90_pad  ;
  output \G95BF_pad  ;
  output \G96BF_pad  ;
  output \G97BF_pad  ;
  output \G98BF_pad  ;
  output \G99BF_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1049/_0_  ;
  output \g1081/_0_  ;
  output \g1115/_0_  ;
  output \g13/_1_  ;
  output \g809/_0_  ;
  output \g810/_0_  ;
  output \g814/_0_  ;
  output \g825/_2_  ;
  output \g834/_0_  ;
  output \g863/_0_  ;
  output \g870/_0_  ;
  output \g871/_0_  ;
  output \g916/_0_  ;
  output \g917/_0_  ;
  output \g940/_3_  ;
  wire n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 ;
  assign n44 = ~\G4_pad  & \G69_reg/NET0131  ;
  assign n45 = \G35_pad  & n44 ;
  assign n47 = ~\G10_pad  & ~\G13_pad  ;
  assign n48 = ~\G3_pad  & \G9_pad  ;
  assign n49 = n47 & n48 ;
  assign n50 = ~\G11_pad  & ~\G3_pad  ;
  assign n46 = ~\G2_pad  & \G66_reg/NET0131  ;
  assign n51 = \G24_pad  & ~n46 ;
  assign n52 = ~n50 & n51 ;
  assign n53 = ~n49 & n52 ;
  assign n54 = ~\G3_pad  & ~n53 ;
  assign n55 = \G77_reg/NET0131  & ~n54 ;
  assign n56 = \G10_pad  & ~\G13_pad  ;
  assign n57 = ~\G3_pad  & ~\G9_pad  ;
  assign n58 = n56 & n57 ;
  assign n59 = \G23_pad  & ~\G65_reg/NET0131  ;
  assign n60 = ~n50 & n59 ;
  assign n61 = ~n58 & n60 ;
  assign n62 = ~\G3_pad  & ~n61 ;
  assign n63 = \G76_reg/NET0131  & ~n62 ;
  assign n64 = ~\G2_pad  & \G64_reg/NET0131  ;
  assign n65 = ~n63 & n64 ;
  assign n66 = ~n55 & n65 ;
  assign n67 = ~\G9_pad  & n47 ;
  assign n68 = \G11_pad  & ~n67 ;
  assign n69 = ~\G3_pad  & ~n68 ;
  assign n70 = \G22_pad  & ~n69 ;
  assign n71 = ~n66 & n70 ;
  assign n72 = ~\G3_pad  & ~n71 ;
  assign n73 = \G75_reg/NET0131  & ~n72 ;
  assign n74 = \G14_pad  & n73 ;
  assign n75 = \G15_pad  & n63 ;
  assign n76 = \G16_pad  & n55 ;
  assign n77 = \G18_pad  & ~\G4_pad  ;
  assign n78 = \G79_reg/NET0131  & n77 ;
  assign n79 = \G19_pad  & ~\G4_pad  ;
  assign n80 = \G65_reg/NET0131  & n79 ;
  assign n81 = \G20_pad  & ~\G4_pad  ;
  assign n82 = \G81_reg/NET0131  & n81 ;
  assign n83 = n48 & n56 ;
  assign n84 = \G25_pad  & ~n50 ;
  assign n85 = ~n83 & n84 ;
  assign n95 = \G74_reg/NET0131  & n71 ;
  assign n96 = ~\G4_pad  & \G73_reg/NET0131  ;
  assign n97 = n67 & n96 ;
  assign n98 = n95 & n97 ;
  assign n91 = \G70_reg/NET0131  & n53 ;
  assign n92 = \G9_pad  & n44 ;
  assign n93 = n47 & n92 ;
  assign n94 = n91 & n93 ;
  assign n87 = \G72_reg/NET0131  & n61 ;
  assign n86 = ~\G4_pad  & \G71_reg/NET0131  ;
  assign n88 = ~\G9_pad  & n56 ;
  assign n89 = n86 & n88 ;
  assign n90 = n87 & n89 ;
  assign n99 = \G12_pad  & \G26_pad  ;
  assign n100 = ~n90 & n99 ;
  assign n101 = ~n94 & n100 ;
  assign n102 = ~n98 & n101 ;
  assign n103 = \G30_pad  & n95 ;
  assign n104 = \G31_pad  & n96 ;
  assign n105 = \G32_pad  & n87 ;
  assign n106 = \G33_pad  & n86 ;
  assign n107 = \G34_pad  & n91 ;
  assign n108 = ~\G2_pad  & ~n55 ;
  assign n109 = n63 & n108 ;
  assign n110 = ~n71 & n96 ;
  assign n111 = ~n95 & ~n110 ;
  assign n112 = \G2_pad  & ~\G5_pad  ;
  assign n113 = n63 & ~n112 ;
  assign n114 = \G5_pad  & n86 ;
  assign n115 = n87 & n114 ;
  assign n116 = ~n55 & n115 ;
  assign n117 = ~n73 & n116 ;
  assign n118 = ~n113 & ~n117 ;
  assign n119 = \G2_pad  & ~\G6_pad  ;
  assign n120 = n55 & ~n119 ;
  assign n121 = \G6_pad  & n44 ;
  assign n122 = ~n63 & n121 ;
  assign n123 = n91 & n122 ;
  assign n124 = ~n73 & n123 ;
  assign n125 = ~n120 & ~n124 ;
  assign n126 = \G2_pad  & ~\G8_pad  ;
  assign n127 = n73 & ~n126 ;
  assign n128 = \G8_pad  & n96 ;
  assign n129 = ~n63 & n128 ;
  assign n130 = ~n55 & n129 ;
  assign n131 = n95 & n130 ;
  assign n132 = ~n127 & ~n131 ;
  assign n133 = ~n63 & n108 ;
  assign n134 = n73 & n133 ;
  assign n135 = ~n95 & n96 ;
  assign n136 = ~\G2_pad  & n55 ;
  assign n137 = n44 & ~n53 ;
  assign n138 = ~n91 & ~n137 ;
  assign n139 = n44 & ~n91 ;
  assign n140 = n86 & ~n87 ;
  assign n141 = ~n61 & n86 ;
  assign n142 = ~n87 & ~n141 ;
  assign n143 = \G11_pad  & \G12_pad  ;
  assign n144 = \G13_pad  & \G28_pad  ;
  assign n145 = n143 & n144 ;
  assign \G100BF_pad  = ~n45 ;
  assign \G103BF_pad  = ~n74 ;
  assign \G104BF_pad  = ~n75 ;
  assign \G105BF_pad  = ~n76 ;
  assign \G107_pad  = n78 ;
  assign \G83_pad  = n80 ;
  assign \G84_pad  = n82 ;
  assign \G86BF_pad  = ~n71 ;
  assign \G87BF_pad  = ~n61 ;
  assign \G88BF_pad  = ~n53 ;
  assign \G89BF_pad  = ~n85 ;
  assign \G90_pad  = n102 ;
  assign \G95BF_pad  = ~n103 ;
  assign \G96BF_pad  = ~n104 ;
  assign \G97BF_pad  = ~n105 ;
  assign \G98BF_pad  = ~n106 ;
  assign \G99BF_pad  = ~n107 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1049/_0_  = n109 ;
  assign \g1081/_0_  = n73 ;
  assign \g1115/_0_  = ~n111 ;
  assign \g13/_1_  = n55 ;
  assign \g809/_0_  = ~n118 ;
  assign \g810/_0_  = ~n125 ;
  assign \g814/_0_  = ~n132 ;
  assign \g825/_2_  = n134 ;
  assign \g834/_0_  = ~n135 ;
  assign \g863/_0_  = n136 ;
  assign \g870/_0_  = ~n138 ;
  assign \g871/_0_  = ~n139 ;
  assign \g916/_0_  = ~n140 ;
  assign \g917/_0_  = ~n142 ;
  assign \g940/_3_  = n145 ;
endmodule
