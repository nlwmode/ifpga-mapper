module top (\G0_pad , \G11_reg/NET0131 , \G12_reg/NET0131 , \G13_reg/NET0131 , \G14_reg/NET0131 , \G15_reg/NET0131 , \G16_reg/NET0131 , \G17_reg/NET0131 , \G18_reg/NET0131 , \G19_reg/NET0131 , \G1_pad , \G20_reg/NET0131 , \G21_reg/NET0131 , \G22_reg/NET0131 , \G23_reg/NET0131 , \G24_reg/NET0131 , \G28_reg/NET0131 , \G29_reg/NET0131 , \G2_pad , \G31_reg/NET0131 , \G119_pad , \G167_pad , \_al_n0 , \_al_n1 , \g43/_3_ , \g754/_0_ , \g757/_0_ , \g760/_0_ , \g768/_2_ , \g770/_2_ , \g773/_0_ , \g786/_2_ , \g792/_0_ , \g793/_0_ , \g796/_0_ , \g804/_0_ , \g808/_0_ , \g817/_0_ , \g825/_0_ , \g834/_0_ , \g837/_0_ , \g838/_0_ , \g839/_0_ , \g840/_0_ , \g843/_0_ );
	input \G0_pad  ;
	input \G11_reg/NET0131  ;
	input \G12_reg/NET0131  ;
	input \G13_reg/NET0131  ;
	input \G14_reg/NET0131  ;
	input \G15_reg/NET0131  ;
	input \G16_reg/NET0131  ;
	input \G17_reg/NET0131  ;
	input \G18_reg/NET0131  ;
	input \G19_reg/NET0131  ;
	input \G1_pad  ;
	input \G20_reg/NET0131  ;
	input \G21_reg/NET0131  ;
	input \G22_reg/NET0131  ;
	input \G23_reg/NET0131  ;
	input \G24_reg/NET0131  ;
	input \G28_reg/NET0131  ;
	input \G29_reg/NET0131  ;
	input \G2_pad  ;
	input \G31_reg/NET0131  ;
	output \G119_pad  ;
	output \G167_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g43/_3_  ;
	output \g754/_0_  ;
	output \g757/_0_  ;
	output \g760/_0_  ;
	output \g768/_2_  ;
	output \g770/_2_  ;
	output \g773/_0_  ;
	output \g786/_2_  ;
	output \g792/_0_  ;
	output \g793/_0_  ;
	output \g796/_0_  ;
	output \g804/_0_  ;
	output \g808/_0_  ;
	output \g817/_0_  ;
	output \g825/_0_  ;
	output \g834/_0_  ;
	output \g837/_0_  ;
	output \g838/_0_  ;
	output \g839/_0_  ;
	output \g840/_0_  ;
	output \g843/_0_  ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\G11_reg/NET0131 ,
		\G12_reg/NET0131 ,
		_w21_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\G13_reg/NET0131 ,
		_w21_,
		_w22_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\G14_reg/NET0131 ,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\G31_reg/NET0131 ,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\G15_reg/NET0131 ,
		\G16_reg/NET0131 ,
		_w25_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		\G17_reg/NET0131 ,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\G18_reg/NET0131 ,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w24_,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\G19_reg/NET0131 ,
		\G20_reg/NET0131 ,
		_w29_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\G21_reg/NET0131 ,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		_w28_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\G22_reg/NET0131 ,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\G0_pad ,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\G19_reg/NET0131 ,
		\G20_reg/NET0131 ,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w28_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\G19_reg/NET0131 ,
		_w28_,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\G20_reg/NET0131 ,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w35_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w33_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\G15_reg/NET0131 ,
		_w24_,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\G16_reg/NET0131 ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\G17_reg/NET0131 ,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\G0_pad ,
		_w28_,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\G18_reg/NET0131 ,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		_w42_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\G0_pad ,
		\G18_reg/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w42_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w45_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\G22_reg/NET0131 ,
		_w31_,
		_w49_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\G21_reg/NET0131 ,
		\G22_reg/NET0131 ,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w35_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w49_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\G0_pad ,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\G17_reg/NET0131 ,
		_w41_,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w42_,
		_w43_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\G21_reg/NET0131 ,
		_w35_,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\G21_reg/NET0131 ,
		_w35_,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w57_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w33_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		\G19_reg/NET0131 ,
		_w28_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w36_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w33_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\G16_reg/NET0131 ,
		_w40_,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		_w41_,
		_w43_,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		_w64_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\G11_reg/NET0131 ,
		\G12_reg/NET0131 ,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\G13_reg/NET0131 ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\G14_reg/NET0131 ,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\G0_pad ,
		_w23_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w69_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		\G21_reg/NET0131 ,
		\G24_reg/NET0131 ,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\G22_reg/NET0131 ,
		_w29_,
		_w73_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		_w72_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\G19_reg/NET0131 ,
		\G20_reg/NET0131 ,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		\G23_reg/NET0131 ,
		_w50_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\G24_reg/NET0131 ,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\G0_pad ,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		\G0_pad ,
		\G21_reg/NET0131 ,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\G23_reg/NET0131 ,
		_w29_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w80_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w79_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		\G17_reg/NET0131 ,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\G0_pad ,
		_w74_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\G15_reg/NET0131 ,
		_w24_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w40_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w43_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		\G21_reg/NET0131 ,
		\G22_reg/NET0131 ,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\G23_reg/NET0131 ,
		_w50_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w90_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		\G0_pad ,
		_w29_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w92_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w79_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w84_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\G13_reg/NET0131 ,
		_w67_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w68_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w70_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\G22_reg/NET0131 ,
		_w29_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\G23_reg/NET0131 ,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		_w80_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w78_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w21_,
		_w67_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w70_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\G19_reg/NET0131 ,
		\G22_reg/NET0131 ,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w34_,
		_w72_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\G0_pad ,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\G22_reg/NET0131 ,
		_w75_,
		_w110_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		_w72_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\G0_pad ,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\G11_reg/NET0131 ,
		_w70_,
		_w113_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\G1_pad ,
		\G31_reg/NET0131 ,
		_w114_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		\G1_pad ,
		\G31_reg/NET0131 ,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w114_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\G0_pad ,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\G23_reg/NET0131 ,
		\G2_pad ,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		\G23_reg/NET0131 ,
		\G2_pad ,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w118_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		\G0_pad ,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		\G0_pad ,
		_w34_,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w72_,
		_w122_,
		_w123_
	);
	assign \G119_pad  = \G28_reg/NET0131 ;
	assign \G167_pad  = \G29_reg/NET0131 ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g43/_3_  = _w39_ ;
	assign \g754/_0_  = _w48_ ;
	assign \g757/_0_  = _w53_ ;
	assign \g760/_0_  = _w56_ ;
	assign \g768/_2_  = _w60_ ;
	assign \g770/_2_  = _w63_ ;
	assign \g773/_0_  = _w66_ ;
	assign \g786/_2_  = _w71_ ;
	assign \g792/_0_  = _w86_ ;
	assign \g793/_0_  = _w89_ ;
	assign \g796/_0_  = _w96_ ;
	assign \g804/_0_  = _w99_ ;
	assign \g808/_0_  = _w103_ ;
	assign \g817/_0_  = _w83_ ;
	assign \g825/_0_  = _w105_ ;
	assign \g834/_0_  = _w109_ ;
	assign \g837/_0_  = _w112_ ;
	assign \g838/_0_  = _w113_ ;
	assign \g839/_0_  = _w117_ ;
	assign \g840/_0_  = _w121_ ;
	assign \g843/_0_  = _w123_ ;
endmodule;