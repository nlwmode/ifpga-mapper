module top( \1(0)_pad  , \100(77)_pad  , \101(78)_pad  , \102(79)_pad  , \103(80)_pad  , \104(81)_pad  , \105(82)_pad  , \106(83)_pad  , \107(84)_pad  , \108(85)_pad  , \11(8)_pad  , \111(86)_pad  , \112(87)_pad  , \113(88)_pad  , \114(89)_pad  , \115(90)_pad  , \116(91)_pad  , \117(92)_pad  , \118(93)_pad  , \119(94)_pad  , \120(95)_pad  , \123(96)_pad  , \124(97)_pad  , \125(98)_pad  , \126(99)_pad  , \127(100)_pad  , \128(101)_pad  , \129(102)_pad  , \130(103)_pad  , \131(104)_pad  , \132(105)_pad  , \1341(200)_pad  , \1348(201)_pad  , \135(106)_pad  , \136(107)_pad  , \137(108)_pad  , \138(109)_pad  , \1384(202)_pad  , \139(110)_pad  , \14(9)_pad  , \140(111)_pad  , \141(112)_pad  , \142(113)_pad  , \15(10)_pad  , \16(11)_pad  , \19(12)_pad  , \1956(203)_pad  , \1961(204)_pad  , \1966(205)_pad  , \1971(206)_pad  , \1976(207)_pad  , \1981(208)_pad  , \1986(209)_pad  , \1991(210)_pad  , \1996(211)_pad  , \2(1)_pad  , \20(13)_pad  , \2067(213)_pad  , \2072(214)_pad  , \2078(215)_pad  , \2084(216)_pad  , \2090(217)_pad  , \2096(218)_pad  , \21(14)_pad  , \2100(219)_pad  , \2104(220)_pad  , \2105(221)_pad  , \2106(222)_pad  , \22(15)_pad  , \23(16)_pad  , \24(17)_pad  , \2427(223)_pad  , \2430(224)_pad  , \2435(225)_pad  , \2438(226)_pad  , \2443(227)_pad  , \2446(228)_pad  , \2451(229)_pad  , \2454(230)_pad  , \2474(231)_pad  , \25(18)_pad  , \26(19)_pad  , \2678(232)_pad  , \27(20)_pad  , \28(21)_pad  , \29(22)_pad  , \3(2)_pad  , \32(23)_pad  , \33(24)_pad  , \34(25)_pad  , \35(26)_pad  , \36(27)_pad  , \37(28)_pad  , \4(3)_pad  , \40(29)_pad  , \409(298)_pad  , \43(30)_pad  , \44(31)_pad  , \47(32)_pad  , \48(33)_pad  , \483(191)_pad  , \49(34)_pad  , \5(4)_pad  , \50(35)_pad  , \51(36)_pad  , \52(37)_pad  , \53(38)_pad  , \54(39)_pad  , \543(192)_pad  , \55(40)_pad  , \559(193)_pad  , \56(41)_pad  , \567(194)_pad  , \57(42)_pad  , \6(5)_pad  , \60(43)_pad  , \61(44)_pad  , \62(45)_pad  , \63(46)_pad  , \64(47)_pad  , \65(48)_pad  , \651(195)_pad  , \66(49)_pad  , \661(196)_pad  , \67(50)_pad  , \68(51)_pad  , \69(52)_pad  , \7(6)_pad  , \72(53)_pad  , \73(54)_pad  , \74(55)_pad  , \75(56)_pad  , \76(57)_pad  , \77(58)_pad  , \78(59)_pad  , \79(60)_pad  , \8(7)_pad  , \80(61)_pad  , \81(62)_pad  , \82(63)_pad  , \85(64)_pad  , \86(65)_pad  , \860(197)_pad  , \868(198)_pad  , \87(66)_pad  , \88(67)_pad  , \89(68)_pad  , \90(69)_pad  , \91(70)_pad  , \92(71)_pad  , \93(72)_pad  , \94(73)_pad  , \95(74)_pad  , \96(75)_pad  , \99(76)_pad  , \145(1358)_pad  , \148(851)_pad  , \150(1277)_pad  , \153(671)_pad  , \156(1046)_pad  , \158(349)_pad  , \160(609)_pad  , \162(612)_pad  , \164(607)_pad  , \166(625)_pad  , \168(623)_pad  , \171(621)_pad  , \173(389)_pad  , \176(803)_pad  , \188(761)_pad  , \217(423)_pad  , \218(311)_pad  , \219(302)_pad  , \220(306)_pad  , \221(305)_pad  , \223(413)_pad  , \225(1424)_pad  , \227(1179)_pad  , \229(1180)_pad  , \234(376)_pad  , \235(307)_pad  , \236(303)_pad  , \237(309)_pad  , \238(304)_pad  , \259(414)_pad  , \261(506)_pad  , \282(922)_pad  , \284(847)_pad  , \286(696)_pad  , \288(700)_pad  , \290(704)_pad  , \295(1400)_pad  , \297(849)_pad  , \299(692)_pad  , \301(694)_pad  , \303(698)_pad  , \305(702)_pad  , \325(507)_pad  , \329(1414)_pad  , \_al_n0  , \u1082_syn_3  , \u1396_syn_3  , \u1414_syn_3  , \u1447_syn_3  , \u538_syn_3  , \u539_syn_3  );
  input \1(0)_pad  ;
  input \100(77)_pad  ;
  input \101(78)_pad  ;
  input \102(79)_pad  ;
  input \103(80)_pad  ;
  input \104(81)_pad  ;
  input \105(82)_pad  ;
  input \106(83)_pad  ;
  input \107(84)_pad  ;
  input \108(85)_pad  ;
  input \11(8)_pad  ;
  input \111(86)_pad  ;
  input \112(87)_pad  ;
  input \113(88)_pad  ;
  input \114(89)_pad  ;
  input \115(90)_pad  ;
  input \116(91)_pad  ;
  input \117(92)_pad  ;
  input \118(93)_pad  ;
  input \119(94)_pad  ;
  input \120(95)_pad  ;
  input \123(96)_pad  ;
  input \124(97)_pad  ;
  input \125(98)_pad  ;
  input \126(99)_pad  ;
  input \127(100)_pad  ;
  input \128(101)_pad  ;
  input \129(102)_pad  ;
  input \130(103)_pad  ;
  input \131(104)_pad  ;
  input \132(105)_pad  ;
  input \1341(200)_pad  ;
  input \1348(201)_pad  ;
  input \135(106)_pad  ;
  input \136(107)_pad  ;
  input \137(108)_pad  ;
  input \138(109)_pad  ;
  input \1384(202)_pad  ;
  input \139(110)_pad  ;
  input \14(9)_pad  ;
  input \140(111)_pad  ;
  input \141(112)_pad  ;
  input \142(113)_pad  ;
  input \15(10)_pad  ;
  input \16(11)_pad  ;
  input \19(12)_pad  ;
  input \1956(203)_pad  ;
  input \1961(204)_pad  ;
  input \1966(205)_pad  ;
  input \1971(206)_pad  ;
  input \1976(207)_pad  ;
  input \1981(208)_pad  ;
  input \1986(209)_pad  ;
  input \1991(210)_pad  ;
  input \1996(211)_pad  ;
  input \2(1)_pad  ;
  input \20(13)_pad  ;
  input \2067(213)_pad  ;
  input \2072(214)_pad  ;
  input \2078(215)_pad  ;
  input \2084(216)_pad  ;
  input \2090(217)_pad  ;
  input \2096(218)_pad  ;
  input \21(14)_pad  ;
  input \2100(219)_pad  ;
  input \2104(220)_pad  ;
  input \2105(221)_pad  ;
  input \2106(222)_pad  ;
  input \22(15)_pad  ;
  input \23(16)_pad  ;
  input \24(17)_pad  ;
  input \2427(223)_pad  ;
  input \2430(224)_pad  ;
  input \2435(225)_pad  ;
  input \2438(226)_pad  ;
  input \2443(227)_pad  ;
  input \2446(228)_pad  ;
  input \2451(229)_pad  ;
  input \2454(230)_pad  ;
  input \2474(231)_pad  ;
  input \25(18)_pad  ;
  input \26(19)_pad  ;
  input \2678(232)_pad  ;
  input \27(20)_pad  ;
  input \28(21)_pad  ;
  input \29(22)_pad  ;
  input \3(2)_pad  ;
  input \32(23)_pad  ;
  input \33(24)_pad  ;
  input \34(25)_pad  ;
  input \35(26)_pad  ;
  input \36(27)_pad  ;
  input \37(28)_pad  ;
  input \4(3)_pad  ;
  input \40(29)_pad  ;
  input \409(298)_pad  ;
  input \43(30)_pad  ;
  input \44(31)_pad  ;
  input \47(32)_pad  ;
  input \48(33)_pad  ;
  input \483(191)_pad  ;
  input \49(34)_pad  ;
  input \5(4)_pad  ;
  input \50(35)_pad  ;
  input \51(36)_pad  ;
  input \52(37)_pad  ;
  input \53(38)_pad  ;
  input \54(39)_pad  ;
  input \543(192)_pad  ;
  input \55(40)_pad  ;
  input \559(193)_pad  ;
  input \56(41)_pad  ;
  input \567(194)_pad  ;
  input \57(42)_pad  ;
  input \6(5)_pad  ;
  input \60(43)_pad  ;
  input \61(44)_pad  ;
  input \62(45)_pad  ;
  input \63(46)_pad  ;
  input \64(47)_pad  ;
  input \65(48)_pad  ;
  input \651(195)_pad  ;
  input \66(49)_pad  ;
  input \661(196)_pad  ;
  input \67(50)_pad  ;
  input \68(51)_pad  ;
  input \69(52)_pad  ;
  input \7(6)_pad  ;
  input \72(53)_pad  ;
  input \73(54)_pad  ;
  input \74(55)_pad  ;
  input \75(56)_pad  ;
  input \76(57)_pad  ;
  input \77(58)_pad  ;
  input \78(59)_pad  ;
  input \79(60)_pad  ;
  input \8(7)_pad  ;
  input \80(61)_pad  ;
  input \81(62)_pad  ;
  input \82(63)_pad  ;
  input \85(64)_pad  ;
  input \86(65)_pad  ;
  input \860(197)_pad  ;
  input \868(198)_pad  ;
  input \87(66)_pad  ;
  input \88(67)_pad  ;
  input \89(68)_pad  ;
  input \90(69)_pad  ;
  input \91(70)_pad  ;
  input \92(71)_pad  ;
  input \93(72)_pad  ;
  input \94(73)_pad  ;
  input \95(74)_pad  ;
  input \96(75)_pad  ;
  input \99(76)_pad  ;
  output \145(1358)_pad  ;
  output \148(851)_pad  ;
  output \150(1277)_pad  ;
  output \153(671)_pad  ;
  output \156(1046)_pad  ;
  output \158(349)_pad  ;
  output \160(609)_pad  ;
  output \162(612)_pad  ;
  output \164(607)_pad  ;
  output \166(625)_pad  ;
  output \168(623)_pad  ;
  output \171(621)_pad  ;
  output \173(389)_pad  ;
  output \176(803)_pad  ;
  output \188(761)_pad  ;
  output \217(423)_pad  ;
  output \218(311)_pad  ;
  output \219(302)_pad  ;
  output \220(306)_pad  ;
  output \221(305)_pad  ;
  output \223(413)_pad  ;
  output \225(1424)_pad  ;
  output \227(1179)_pad  ;
  output \229(1180)_pad  ;
  output \234(376)_pad  ;
  output \235(307)_pad  ;
  output \236(303)_pad  ;
  output \237(309)_pad  ;
  output \238(304)_pad  ;
  output \259(414)_pad  ;
  output \261(506)_pad  ;
  output \282(922)_pad  ;
  output \284(847)_pad  ;
  output \286(696)_pad  ;
  output \288(700)_pad  ;
  output \290(704)_pad  ;
  output \295(1400)_pad  ;
  output \297(849)_pad  ;
  output \299(692)_pad  ;
  output \301(694)_pad  ;
  output \303(698)_pad  ;
  output \305(702)_pad  ;
  output \325(507)_pad  ;
  output \329(1414)_pad  ;
  output \_al_n0  ;
  output \u1082_syn_3  ;
  output \u1396_syn_3  ;
  output \u1414_syn_3  ;
  output \u1447_syn_3  ;
  output \u538_syn_3  ;
  output \u539_syn_3  ;
  wire n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 ;
  assign n156 = \543(192)_pad  & ~\651(195)_pad  ;
  assign n157 = \54(39)_pad  & n156 ;
  assign n158 = \543(192)_pad  & \651(195)_pad  ;
  assign n159 = \79(60)_pad  & n158 ;
  assign n164 = ~n157 & ~n159 ;
  assign n160 = ~\543(192)_pad  & \651(195)_pad  ;
  assign n161 = \66(49)_pad  & n160 ;
  assign n162 = ~\543(192)_pad  & ~\651(195)_pad  ;
  assign n163 = \92(71)_pad  & n162 ;
  assign n165 = ~n161 & ~n163 ;
  assign n166 = n164 & n165 ;
  assign n167 = \559(193)_pad  & n166 ;
  assign n168 = ~\860(197)_pad  & n167 ;
  assign n169 = \43(30)_pad  & n156 ;
  assign n170 = \68(51)_pad  & n158 ;
  assign n173 = ~n169 & ~n170 ;
  assign n171 = \56(41)_pad  & n160 ;
  assign n172 = \81(62)_pad  & n162 ;
  assign n174 = ~n171 & ~n172 ;
  assign n175 = n173 & n174 ;
  assign n176 = \860(197)_pad  & n175 ;
  assign n177 = ~n168 & ~n176 ;
  assign n178 = \55(40)_pad  & n156 ;
  assign n179 = \80(61)_pad  & n158 ;
  assign n182 = ~n178 & ~n179 ;
  assign n180 = \67(50)_pad  & n160 ;
  assign n181 = \93(72)_pad  & n162 ;
  assign n183 = ~n180 & ~n181 ;
  assign n184 = n182 & n183 ;
  assign n185 = n175 & ~n184 ;
  assign n186 = ~n175 & n184 ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = n177 & ~n187 ;
  assign n189 = ~n177 & n187 ;
  assign n190 = ~n188 & ~n189 ;
  assign n191 = n166 & ~n168 ;
  assign n379 = \16(11)_pad  & ~n175 ;
  assign n380 = ~\16(11)_pad  & \19(12)_pad  ;
  assign n381 = ~n379 & ~n380 ;
  assign n383 = ~\1341(200)_pad  & n381 ;
  assign n339 = ~\16(11)_pad  & ~\23(16)_pad  ;
  assign n340 = \87(66)_pad  & n162 ;
  assign n343 = ~n160 & ~n340 ;
  assign n341 = \74(55)_pad  & n158 ;
  assign n342 = \49(34)_pad  & n156 ;
  assign n344 = ~n341 & ~n342 ;
  assign n345 = n343 & n344 ;
  assign n346 = \16(11)_pad  & n345 ;
  assign n347 = ~n339 & ~n346 ;
  assign n378 = ~\1976(207)_pad  & ~n347 ;
  assign n382 = \1341(200)_pad  & ~n381 ;
  assign n399 = ~n378 & ~n382 ;
  assign n400 = ~n383 & n399 ;
  assign n350 = ~\16(11)_pad  & ~\22(15)_pad  ;
  assign n351 = \50(35)_pad  & n156 ;
  assign n352 = \75(56)_pad  & n158 ;
  assign n355 = ~n351 & ~n352 ;
  assign n353 = \62(45)_pad  & n160 ;
  assign n354 = \88(67)_pad  & n162 ;
  assign n356 = ~n353 & ~n354 ;
  assign n357 = n355 & n356 ;
  assign n358 = \16(11)_pad  & n357 ;
  assign n359 = ~n350 & ~n358 ;
  assign n364 = ~\1971(206)_pad  & ~n359 ;
  assign n231 = ~\16(11)_pad  & \21(14)_pad  ;
  assign n232 = \51(36)_pad  & n156 ;
  assign n233 = \76(57)_pad  & n158 ;
  assign n236 = ~n232 & ~n233 ;
  assign n234 = \63(46)_pad  & n160 ;
  assign n235 = \89(68)_pad  & n162 ;
  assign n237 = ~n234 & ~n235 ;
  assign n238 = n236 & n237 ;
  assign n239 = \16(11)_pad  & ~n238 ;
  assign n240 = ~n231 & ~n239 ;
  assign n365 = \1966(205)_pad  & ~n240 ;
  assign n397 = ~n364 & ~n365 ;
  assign n366 = ~\16(11)_pad  & \5(4)_pad  ;
  assign n367 = \52(37)_pad  & n156 ;
  assign n368 = \77(58)_pad  & n158 ;
  assign n371 = ~n367 & ~n368 ;
  assign n369 = \64(47)_pad  & n160 ;
  assign n370 = \90(69)_pad  & n162 ;
  assign n372 = ~n369 & ~n370 ;
  assign n373 = n371 & n372 ;
  assign n374 = \16(11)_pad  & ~n373 ;
  assign n375 = ~n366 & ~n374 ;
  assign n376 = ~\1961(204)_pad  & n375 ;
  assign n377 = \1961(204)_pad  & ~n375 ;
  assign n398 = ~n376 & ~n377 ;
  assign n401 = n397 & n398 ;
  assign n360 = \1971(206)_pad  & n359 ;
  assign n328 = ~\29(22)_pad  & ~\32(23)_pad  ;
  assign n192 = \2104(220)_pad  & ~\2105(221)_pad  ;
  assign n329 = \105(82)_pad  & n192 ;
  assign n194 = \2104(220)_pad  & \2105(221)_pad  ;
  assign n330 = \117(92)_pad  & n194 ;
  assign n333 = ~n329 & ~n330 ;
  assign n196 = ~\2104(220)_pad  & \2105(221)_pad  ;
  assign n331 = \129(102)_pad  & n196 ;
  assign n198 = ~\2104(220)_pad  & ~\2105(221)_pad  ;
  assign n332 = \141(112)_pad  & n198 ;
  assign n334 = ~n331 & ~n332 ;
  assign n335 = n333 & n334 ;
  assign n336 = \29(22)_pad  & n335 ;
  assign n337 = ~n328 & ~n336 ;
  assign n361 = \1996(211)_pad  & n337 ;
  assign n395 = ~n360 & ~n361 ;
  assign n209 = ~\29(22)_pad  & ~\33(24)_pad  ;
  assign n210 = \103(80)_pad  & n192 ;
  assign n211 = \115(90)_pad  & n194 ;
  assign n214 = ~n210 & ~n211 ;
  assign n212 = \127(100)_pad  & n196 ;
  assign n213 = \139(110)_pad  & n198 ;
  assign n215 = ~n212 & ~n213 ;
  assign n216 = n214 & n215 ;
  assign n217 = \29(22)_pad  & n216 ;
  assign n218 = ~n209 & ~n217 ;
  assign n362 = \2072(214)_pad  & n218 ;
  assign n316 = ~\26(19)_pad  & ~\29(22)_pad  ;
  assign n317 = \104(81)_pad  & n192 ;
  assign n318 = \116(91)_pad  & n194 ;
  assign n321 = ~n317 & ~n318 ;
  assign n319 = \128(101)_pad  & n196 ;
  assign n320 = \140(111)_pad  & n198 ;
  assign n322 = ~n319 & ~n320 ;
  assign n323 = n321 & n322 ;
  assign n324 = \29(22)_pad  & n323 ;
  assign n325 = ~n316 & ~n324 ;
  assign n363 = ~\2067(213)_pad  & ~n325 ;
  assign n396 = ~n362 & ~n363 ;
  assign n402 = n395 & n396 ;
  assign n411 = n401 & n402 ;
  assign n412 = n400 & n411 ;
  assign n246 = \48(33)_pad  & n156 ;
  assign n247 = \73(54)_pad  & n158 ;
  assign n250 = ~n246 & ~n247 ;
  assign n248 = \61(44)_pad  & n160 ;
  assign n249 = \86(65)_pad  & n162 ;
  assign n251 = ~n248 & ~n249 ;
  assign n252 = n250 & n251 ;
  assign n253 = \16(11)_pad  & ~n252 ;
  assign n254 = ~\16(11)_pad  & \6(5)_pad  ;
  assign n255 = ~n253 & ~n254 ;
  assign n256 = ~\1981(208)_pad  & ~n255 ;
  assign n257 = \1981(208)_pad  & n255 ;
  assign n258 = ~n256 & ~n257 ;
  assign n193 = \100(77)_pad  & n192 ;
  assign n195 = \112(87)_pad  & n194 ;
  assign n200 = ~n193 & ~n195 ;
  assign n197 = \124(97)_pad  & n196 ;
  assign n199 = \136(107)_pad  & n198 ;
  assign n201 = ~n197 & ~n199 ;
  assign n202 = n200 & n201 ;
  assign n203 = \29(22)_pad  & ~n202 ;
  assign n204 = ~\29(22)_pad  & \35(26)_pad  ;
  assign n205 = ~n203 & ~n204 ;
  assign n206 = ~\2090(217)_pad  & ~n205 ;
  assign n207 = \2090(217)_pad  & n205 ;
  assign n208 = ~n206 & ~n207 ;
  assign n219 = ~\2072(214)_pad  & ~n218 ;
  assign n259 = \99(76)_pad  & n192 ;
  assign n260 = \111(86)_pad  & n194 ;
  assign n263 = ~n259 & ~n260 ;
  assign n261 = \123(96)_pad  & n196 ;
  assign n262 = \135(106)_pad  & n198 ;
  assign n264 = ~n261 & ~n262 ;
  assign n265 = n263 & n264 ;
  assign n266 = \29(22)_pad  & n265 ;
  assign n278 = ~\28(21)_pad  & ~\29(22)_pad  ;
  assign n384 = \11(8)_pad  & ~n278 ;
  assign n385 = ~n266 & n384 ;
  assign n386 = ~n219 & n385 ;
  assign n407 = ~n208 & n386 ;
  assign n408 = ~n258 & n407 ;
  assign n242 = ~\16(11)_pad  & \4(3)_pad  ;
  assign n243 = \16(11)_pad  & ~n166 ;
  assign n244 = ~n242 & ~n243 ;
  assign n279 = ~\1348(201)_pad  & n244 ;
  assign n267 = ~\16(11)_pad  & \24(17)_pad  ;
  assign n268 = \47(32)_pad  & n156 ;
  assign n269 = \72(53)_pad  & n158 ;
  assign n272 = ~n268 & ~n269 ;
  assign n270 = \60(43)_pad  & n160 ;
  assign n271 = \85(64)_pad  & n162 ;
  assign n273 = ~n270 & ~n271 ;
  assign n274 = n272 & n273 ;
  assign n275 = \16(11)_pad  & ~n274 ;
  assign n276 = ~n267 & ~n275 ;
  assign n280 = \1986(209)_pad  & ~n276 ;
  assign n389 = ~n279 & ~n280 ;
  assign n281 = \25(18)_pad  & ~\29(22)_pad  ;
  assign n282 = \95(74)_pad  & n192 ;
  assign n283 = \107(84)_pad  & n194 ;
  assign n286 = ~n282 & ~n283 ;
  assign n284 = \119(94)_pad  & n196 ;
  assign n285 = \131(104)_pad  & n198 ;
  assign n287 = ~n284 & ~n285 ;
  assign n288 = n286 & n287 ;
  assign n289 = \29(22)_pad  & ~n288 ;
  assign n290 = ~n281 & ~n289 ;
  assign n291 = \1991(210)_pad  & ~n290 ;
  assign n292 = ~\29(22)_pad  & ~\34(25)_pad  ;
  assign n293 = \101(78)_pad  & n192 ;
  assign n294 = \113(88)_pad  & n194 ;
  assign n297 = ~n293 & ~n294 ;
  assign n295 = \125(98)_pad  & n196 ;
  assign n296 = \137(108)_pad  & n198 ;
  assign n298 = ~n295 & ~n296 ;
  assign n299 = n297 & n298 ;
  assign n300 = \29(22)_pad  & n299 ;
  assign n301 = ~n292 & ~n300 ;
  assign n302 = \2084(216)_pad  & n301 ;
  assign n390 = ~n291 & ~n302 ;
  assign n405 = n389 & n390 ;
  assign n220 = \27(20)_pad  & ~\29(22)_pad  ;
  assign n221 = \102(79)_pad  & n192 ;
  assign n222 = \114(89)_pad  & n194 ;
  assign n225 = ~n221 & ~n222 ;
  assign n223 = \126(99)_pad  & n196 ;
  assign n224 = \138(109)_pad  & n198 ;
  assign n226 = ~n223 & ~n224 ;
  assign n227 = n225 & n226 ;
  assign n228 = \29(22)_pad  & ~n227 ;
  assign n229 = ~n220 & ~n228 ;
  assign n230 = ~\2078(215)_pad  & n229 ;
  assign n241 = ~\1966(205)_pad  & n240 ;
  assign n387 = ~n230 & ~n241 ;
  assign n245 = \1348(201)_pad  & ~n244 ;
  assign n277 = ~\1986(209)_pad  & n276 ;
  assign n388 = ~n245 & ~n277 ;
  assign n406 = n387 & n388 ;
  assign n409 = n405 & n406 ;
  assign n327 = ~\1991(210)_pad  & n290 ;
  assign n338 = ~\1996(211)_pad  & ~n337 ;
  assign n393 = ~n327 & ~n338 ;
  assign n348 = \1976(207)_pad  & n347 ;
  assign n349 = \2078(215)_pad  & ~n229 ;
  assign n394 = ~n348 & ~n349 ;
  assign n403 = n393 & n394 ;
  assign n303 = ~\16(11)_pad  & \20(13)_pad  ;
  assign n304 = \53(38)_pad  & n156 ;
  assign n305 = \78(59)_pad  & n158 ;
  assign n308 = ~n304 & ~n305 ;
  assign n306 = \65(48)_pad  & n160 ;
  assign n307 = \91(70)_pad  & n162 ;
  assign n309 = ~n306 & ~n307 ;
  assign n310 = n308 & n309 ;
  assign n311 = \16(11)_pad  & ~n310 ;
  assign n312 = ~n303 & ~n311 ;
  assign n313 = ~\1956(203)_pad  & n312 ;
  assign n314 = \1956(203)_pad  & ~n312 ;
  assign n391 = ~n313 & ~n314 ;
  assign n315 = ~\2084(216)_pad  & ~n301 ;
  assign n326 = \2067(213)_pad  & n325 ;
  assign n392 = ~n315 & ~n326 ;
  assign n404 = n391 & n392 ;
  assign n410 = n403 & n404 ;
  assign n413 = n409 & n410 ;
  assign n414 = n408 & n413 ;
  assign n415 = n412 & n414 ;
  assign n417 = ~\2096(218)_pad  & n265 ;
  assign n416 = \2096(218)_pad  & ~n265 ;
  assign n418 = ~\2100(219)_pad  & ~n416 ;
  assign n419 = ~n417 & n418 ;
  assign n420 = \2072(214)_pad  & \2078(215)_pad  ;
  assign n421 = \2084(216)_pad  & \2090(217)_pad  ;
  assign n422 = n420 & n421 ;
  assign n423 = \409(298)_pad  & \94(73)_pad  ;
  assign n424 = \108(85)_pad  & \120(95)_pad  ;
  assign n425 = \57(42)_pad  & \69(52)_pad  ;
  assign n426 = n424 & n425 ;
  assign n427 = \567(194)_pad  & ~n426 ;
  assign n428 = \132(105)_pad  & \44(31)_pad  ;
  assign n429 = \82(63)_pad  & \96(75)_pad  ;
  assign n430 = n428 & n429 ;
  assign n431 = \2106(222)_pad  & ~n430 ;
  assign n432 = ~n427 & ~n431 ;
  assign n433 = \483(191)_pad  & \661(196)_pad  ;
  assign n434 = \36(27)_pad  & n433 ;
  assign n435 = n432 & n434 ;
  assign n436 = \1(0)_pad  & \3(2)_pad  ;
  assign n437 = n433 & ~n436 ;
  assign n438 = n432 & n437 ;
  assign n439 = \661(196)_pad  & \7(6)_pad  ;
  assign n440 = \2106(222)_pad  & n439 ;
  assign n441 = n310 & ~n357 ;
  assign n442 = ~n310 & n357 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = n187 & ~n252 ;
  assign n445 = ~n187 & n252 ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = n274 & n446 ;
  assign n448 = ~n274 & ~n446 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = n345 & ~n449 ;
  assign n451 = ~n345 & n449 ;
  assign n452 = ~n450 & ~n451 ;
  assign n453 = n443 & n452 ;
  assign n454 = ~n443 & ~n452 ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = n166 & ~n373 ;
  assign n457 = ~n166 & n373 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = n238 & n458 ;
  assign n460 = ~n238 & ~n458 ;
  assign n461 = ~n459 & ~n460 ;
  assign n463 = ~n455 & ~n461 ;
  assign n462 = n455 & n461 ;
  assign n464 = ~\37(28)_pad  & ~n462 ;
  assign n465 = ~n463 & n464 ;
  assign n494 = ~n202 & n265 ;
  assign n495 = n202 & ~n265 ;
  assign n496 = ~n494 & ~n495 ;
  assign n497 = n299 & n496 ;
  assign n498 = ~n299 & ~n496 ;
  assign n499 = ~n497 & ~n498 ;
  assign n500 = \106(83)_pad  & n192 ;
  assign n501 = \118(93)_pad  & n194 ;
  assign n504 = ~n500 & ~n501 ;
  assign n502 = \130(103)_pad  & n196 ;
  assign n503 = \142(113)_pad  & n198 ;
  assign n505 = ~n502 & ~n503 ;
  assign n506 = n504 & n505 ;
  assign n507 = n227 & ~n506 ;
  assign n508 = ~n227 & n506 ;
  assign n509 = ~n507 & ~n508 ;
  assign n510 = n323 & ~n335 ;
  assign n511 = ~n323 & n335 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = n216 & n512 ;
  assign n514 = ~n216 & ~n512 ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = n288 & ~n515 ;
  assign n517 = ~n288 & n515 ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = n509 & n518 ;
  assign n520 = ~n509 & ~n518 ;
  assign n521 = ~n519 & ~n520 ;
  assign n523 = n499 & ~n521 ;
  assign n522 = ~n499 & n521 ;
  assign n524 = ~\37(28)_pad  & ~n522 ;
  assign n525 = ~n523 & n524 ;
  assign n466 = \1341(200)_pad  & ~\1348(201)_pad  ;
  assign n467 = ~\1341(200)_pad  & \1348(201)_pad  ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = ~\2435(225)_pad  & ~\2438(226)_pad  ;
  assign n470 = \2435(225)_pad  & \2438(226)_pad  ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = n468 & ~n471 ;
  assign n473 = ~n468 & n471 ;
  assign n474 = ~n472 & ~n473 ;
  assign n475 = ~\2446(228)_pad  & ~\2454(230)_pad  ;
  assign n476 = \2446(228)_pad  & \2454(230)_pad  ;
  assign n477 = ~n475 & ~n476 ;
  assign n478 = ~\2427(223)_pad  & ~\2430(224)_pad  ;
  assign n479 = \2427(223)_pad  & \2430(224)_pad  ;
  assign n480 = ~n478 & ~n479 ;
  assign n481 = \2443(227)_pad  & ~\2451(229)_pad  ;
  assign n482 = ~\2443(227)_pad  & \2451(229)_pad  ;
  assign n483 = ~n481 & ~n482 ;
  assign n484 = n480 & ~n483 ;
  assign n485 = ~n480 & n483 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = ~n477 & n486 ;
  assign n488 = n477 & ~n486 ;
  assign n489 = ~n487 & ~n488 ;
  assign n491 = ~n474 & ~n489 ;
  assign n490 = n474 & n489 ;
  assign n492 = \14(9)_pad  & ~n490 ;
  assign n493 = ~n491 & n492 ;
  assign n546 = \1971(206)_pad  & ~\1981(208)_pad  ;
  assign n547 = ~\1971(206)_pad  & \1981(208)_pad  ;
  assign n548 = ~n546 & ~n547 ;
  assign n549 = ~\1976(207)_pad  & ~\2474(231)_pad  ;
  assign n550 = \1976(207)_pad  & \2474(231)_pad  ;
  assign n551 = ~n549 & ~n550 ;
  assign n552 = n548 & ~n551 ;
  assign n553 = ~n548 & n551 ;
  assign n554 = ~n552 & ~n553 ;
  assign n555 = ~\1961(204)_pad  & ~\1986(209)_pad  ;
  assign n556 = \1961(204)_pad  & \1986(209)_pad  ;
  assign n557 = ~n555 & ~n556 ;
  assign n558 = \1966(205)_pad  & ~\1991(210)_pad  ;
  assign n559 = ~\1966(205)_pad  & \1991(210)_pad  ;
  assign n560 = ~n558 & ~n559 ;
  assign n561 = n557 & n560 ;
  assign n562 = ~n557 & ~n560 ;
  assign n563 = ~n561 & ~n562 ;
  assign n564 = \1956(203)_pad  & ~\1996(211)_pad  ;
  assign n565 = ~\1956(203)_pad  & \1996(211)_pad  ;
  assign n566 = ~n564 & ~n565 ;
  assign n567 = n563 & ~n566 ;
  assign n568 = ~n563 & n566 ;
  assign n569 = ~n567 & ~n568 ;
  assign n570 = n554 & n569 ;
  assign n571 = ~n554 & ~n569 ;
  assign n572 = ~n570 & ~n571 ;
  assign n526 = ~\2072(214)_pad  & ~\2078(215)_pad  ;
  assign n527 = ~n420 & ~n526 ;
  assign n528 = \2096(218)_pad  & ~n527 ;
  assign n529 = ~\2096(218)_pad  & n527 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = \2084(216)_pad  & ~n530 ;
  assign n532 = ~\2084(216)_pad  & n530 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = ~\2090(217)_pad  & ~\2678(232)_pad  ;
  assign n535 = \2090(217)_pad  & \2678(232)_pad  ;
  assign n536 = ~n534 & ~n535 ;
  assign n537 = \2067(213)_pad  & n536 ;
  assign n538 = ~\2067(213)_pad  & ~n536 ;
  assign n539 = ~n537 & ~n538 ;
  assign n540 = \2100(219)_pad  & ~n539 ;
  assign n541 = ~\2100(219)_pad  & n539 ;
  assign n542 = ~n540 & ~n541 ;
  assign n543 = n533 & n542 ;
  assign n544 = ~n533 & ~n542 ;
  assign n545 = ~n543 & ~n544 ;
  assign n573 = n432 & ~n545 ;
  assign n574 = ~n572 & n573 ;
  assign n575 = ~n493 & n574 ;
  assign n576 = ~n525 & n575 ;
  assign n577 = ~n465 & n576 ;
  assign n578 = \567(194)_pad  & n439 ;
  assign n579 = \15(10)_pad  & \2(1)_pad  ;
  assign n580 = \661(196)_pad  & n579 ;
  assign n581 = n426 & n430 ;
  assign n582 = ~\868(198)_pad  & n175 ;
  assign n583 = ~\559(193)_pad  & \868(198)_pad  ;
  assign n584 = n166 & n583 ;
  assign n585 = ~n582 & ~n584 ;
  assign n586 = \868(198)_pad  & ~n373 ;
  assign n587 = ~\868(198)_pad  & ~n166 ;
  assign n588 = ~n586 & ~n587 ;
  assign n589 = n167 & n455 ;
  assign n590 = ~n167 & ~n455 ;
  assign n591 = ~n589 & ~n590 ;
  assign n592 = \868(198)_pad  & ~n591 ;
  assign n593 = ~\868(198)_pad  & ~n184 ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = \868(198)_pad  & ~n238 ;
  assign n596 = ~\868(198)_pad  & ~n310 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = ~\1384(202)_pad  & ~n227 ;
  assign n599 = \40(29)_pad  & n299 ;
  assign n600 = n598 & n599 ;
  assign n605 = \1348(201)_pad  & ~n600 ;
  assign n606 = \2067(213)_pad  & n600 ;
  assign n607 = ~n605 & ~n606 ;
  assign n610 = ~n166 & ~n607 ;
  assign n611 = \1341(200)_pad  & ~n600 ;
  assign n609 = \1996(211)_pad  & n600 ;
  assign n612 = n175 & ~n609 ;
  assign n613 = ~n611 & n612 ;
  assign n614 = ~n610 & n613 ;
  assign n601 = \1956(203)_pad  & ~n600 ;
  assign n602 = \2072(214)_pad  & n600 ;
  assign n603 = ~n601 & ~n602 ;
  assign n604 = n310 & n603 ;
  assign n608 = n166 & n607 ;
  assign n615 = ~n604 & ~n608 ;
  assign n616 = ~n614 & n615 ;
  assign n624 = \1961(204)_pad  & ~n600 ;
  assign n625 = \2078(215)_pad  & n600 ;
  assign n626 = ~n624 & ~n625 ;
  assign n628 = ~n373 & ~n626 ;
  assign n623 = ~n310 & ~n603 ;
  assign n627 = n373 & n626 ;
  assign n630 = ~n623 & ~n627 ;
  assign n631 = ~n628 & n630 ;
  assign n618 = \1966(205)_pad  & ~n600 ;
  assign n617 = \2084(216)_pad  & n600 ;
  assign n619 = \8(7)_pad  & ~n617 ;
  assign n620 = ~n618 & n619 ;
  assign n621 = \8(7)_pad  & ~n238 ;
  assign n622 = ~n620 & n621 ;
  assign n629 = n238 & n620 ;
  assign n632 = ~n622 & ~n629 ;
  assign n633 = n631 & n632 ;
  assign n634 = ~n616 & n633 ;
  assign n635 = ~n622 & n627 ;
  assign n636 = ~n629 & ~n635 ;
  assign n637 = ~n634 & n636 ;
  assign n648 = \1971(206)_pad  & ~n600 ;
  assign n647 = \2090(217)_pad  & n600 ;
  assign n649 = \8(7)_pad  & ~n647 ;
  assign n650 = ~n648 & n649 ;
  assign n652 = \8(7)_pad  & ~n357 ;
  assign n653 = ~n650 & n652 ;
  assign n651 = n357 & n650 ;
  assign n638 = \8(7)_pad  & ~n600 ;
  assign n639 = ~\1976(207)_pad  & n345 ;
  assign n640 = n638 & n639 ;
  assign n641 = \1981(208)_pad  & ~n252 ;
  assign n642 = n638 & n641 ;
  assign n654 = ~n640 & ~n642 ;
  assign n643 = \1976(207)_pad  & ~n345 ;
  assign n644 = n638 & n643 ;
  assign n645 = ~\1981(208)_pad  & n252 ;
  assign n646 = n638 & n645 ;
  assign n655 = ~n644 & ~n646 ;
  assign n656 = n654 & n655 ;
  assign n657 = ~n651 & n656 ;
  assign n658 = ~n653 & n657 ;
  assign n659 = ~n637 & n658 ;
  assign n660 = ~n644 & n651 ;
  assign n661 = ~n640 & ~n660 ;
  assign n662 = ~n642 & ~n661 ;
  assign n663 = ~n646 & ~n662 ;
  assign n664 = ~n659 & n663 ;
  assign n665 = ~n598 & n599 ;
  assign n666 = ~\2067(213)_pad  & n323 ;
  assign n667 = \1986(209)_pad  & ~n274 ;
  assign n676 = ~n666 & ~n667 ;
  assign n668 = \1991(210)_pad  & ~n288 ;
  assign n669 = ~\1986(209)_pad  & n274 ;
  assign n677 = ~n668 & ~n669 ;
  assign n678 = n676 & n677 ;
  assign n670 = \2067(213)_pad  & ~n323 ;
  assign n671 = \1996(211)_pad  & ~n335 ;
  assign n672 = ~n670 & ~n671 ;
  assign n673 = ~\1991(210)_pad  & n288 ;
  assign n674 = ~\1996(211)_pad  & n335 ;
  assign n675 = ~n673 & ~n674 ;
  assign n679 = n672 & n675 ;
  assign n680 = n678 & n679 ;
  assign n681 = n665 & ~n680 ;
  assign n682 = ~n664 & ~n681 ;
  assign n683 = ~n668 & n669 ;
  assign n684 = n675 & ~n683 ;
  assign n685 = n672 & ~n684 ;
  assign n686 = ~n666 & ~n685 ;
  assign n687 = n665 & ~n686 ;
  assign n688 = ~n682 & ~n687 ;
  assign \145(1358)_pad  = n190 ;
  assign \148(851)_pad  = ~n191 ;
  assign \150(1277)_pad  = ~n415 ;
  assign \153(671)_pad  = ~n176 ;
  assign \156(1046)_pad  = ~n419 ;
  assign \158(349)_pad  = ~n422 ;
  assign \160(609)_pad  = n299 ;
  assign \162(612)_pad  = n202 ;
  assign \164(607)_pad  = n227 ;
  assign \166(625)_pad  = n357 ;
  assign \168(623)_pad  = n238 ;
  assign \171(621)_pad  = n373 ;
  assign \173(389)_pad  = n423 ;
  assign \176(803)_pad  = ~n435 ;
  assign \188(761)_pad  = ~n438 ;
  assign \217(423)_pad  = ~n440 ;
  assign \218(311)_pad  = ~\44(31)_pad  ;
  assign \219(302)_pad  = ~\132(105)_pad  ;
  assign \220(306)_pad  = ~\82(63)_pad  ;
  assign \221(305)_pad  = ~\96(75)_pad  ;
  assign \223(413)_pad  = ~n439 ;
  assign \225(1424)_pad  = ~n577 ;
  assign \227(1179)_pad  = n545 ;
  assign \229(1180)_pad  = n572 ;
  assign \234(376)_pad  = ~n578 ;
  assign \235(307)_pad  = ~\69(52)_pad  ;
  assign \236(303)_pad  = ~\120(95)_pad  ;
  assign \237(309)_pad  = ~\57(42)_pad  ;
  assign \238(304)_pad  = ~\108(85)_pad  ;
  assign \259(414)_pad  = ~n580 ;
  assign \261(506)_pad  = ~n581 ;
  assign \282(922)_pad  = n585 ;
  assign \284(847)_pad  = ~n588 ;
  assign \286(696)_pad  = ~n238 ;
  assign \288(700)_pad  = ~n345 ;
  assign \290(704)_pad  = ~n274 ;
  assign \295(1400)_pad  = ~n594 ;
  assign \297(849)_pad  = ~n597 ;
  assign \299(692)_pad  = ~n310 ;
  assign \301(694)_pad  = ~n373 ;
  assign \303(698)_pad  = ~n357 ;
  assign \305(702)_pad  = ~n252 ;
  assign \325(507)_pad  = n581 ;
  assign \329(1414)_pad  = ~n688 ;
  assign \_al_n0  = 1'b0 ;
  assign \u1082_syn_3  = n432 ;
  assign \u1396_syn_3  = n577 ;
  assign \u1414_syn_3  = n465 ;
  assign \u1447_syn_3  = n525 ;
  assign \u538_syn_3  = n415 ;
  assign \u539_syn_3  = n493 ;
endmodule
