module top( \n1035gat_reg/NET0131  , \n1045gat_reg/NET0131  , \n1068gat_reg/NET0131  , \n1072gat_reg/NET0131  , \n1080gat_reg/NET0131  , \n1121gat_reg/NET0131  , \n1135gat_reg/NET0131  , \n1148gat_reg/NET0131  , \n1197gat_reg/NET0131  , \n1226gat_reg/NET0131  , \n1241gat_reg/NET0131  , \n1282gat_reg/NET0131  , \n1294gat_reg/NET0131  , \n1312gat_reg/NET0131  , \n1316gat_reg/NET0131  , \n1332gat_reg/NET0131  , \n1336gat_reg/NET0131  , \n1340gat_reg/NET0131  , \n1363gat_reg/NET0131  , \n1389gat_reg/NET0131  , \n1394gat_reg/NET0131  , \n1433gat_reg/NET0131  , \n1456gat_reg/NET0131  , \n1462gat_reg/NET0131  , \n148gat_reg/NET0131  , \n1496gat_reg/NET0131  , \n1508gat_reg/NET0131  , \n1525gat_reg/NET0131  , \n152gat_reg/NET0131  , \n156gat_reg/NET0131  , \n1588gat_reg/NET0131  , \n1596gat_reg/NET0131  , \n160gat_reg/NET0131  , \n1675gat_reg/NET0131  , \n1678gat_reg/NET0131  , \n1740gat_reg/NET0131  , \n1748gat_reg/NET0131  , \n1763gat_reg/NET0131  , \n1767gat_reg/NET0131  , \n1771gat_reg/NET0131  , \n1775gat_reg/NET0131  , \n1807gat_reg/NET0131  , \n1821gat_reg/NET0131  , \n1829gat_reg/NET0131  , \n1834gat_reg/NET0131  , \n1850gat_reg/NET0131  , \n1871gat_reg/NET0131  , \n1880gat_reg/NET0131  , \n1899gat_reg/NET0131  , \n1975gat_reg/NET0131  , \n2021gat_reg/NET0131  , \n2025gat_reg/NET0131  , \n2029gat_reg/NET0131  , \n2033gat_reg/NET0131  , \n2037gat_reg/NET0131  , \n2040gat_reg/NET0131  , \n2044gat_reg/NET0131  , \n2061gat_reg/NET0131  , \n2084gat_reg/NET0131  , \n2091gat_reg/NET0131  , \n2095gat_reg/NET0131  , \n2099gat_reg/NET0131  , \n2102gat_reg/NET0131  , \n2110gat_reg/NET0131  , \n2117gat_reg/NET0131  , \n2121gat_reg/NET0131  , \n2125gat_reg/NET0131  , \n2135gat_reg/NET0131  , \n2139gat_reg/NET0131  , \n2143gat_reg/NET0131  , \n2155gat_reg/NET0131  , \n2169gat_reg/NET0131  , \n2176gat_reg/NET0131  , \n2179gat_reg/NET0131  , \n2182gat_reg/NET0131  , \n2190gat_reg/NET0131  , \n2203gat_reg/NET0131  , \n2207gat_reg/NET0131  , \n2262gat_reg/NET0131  , \n2266gat_reg/NET0131  , \n2270gat_reg/NET0131  , \n2319gat_reg/NET0131  , \n2339gat_reg/NET0131  , \n2343gat_reg/NET0131  , \n2347gat_reg/NET0131  , \n2390gat_reg/NET0131  , \n2394gat_reg/NET0131  , \n2399gat_reg/NET0131  , \n2403gat_reg/NET0131  , \n2407gat_reg/NET0131  , \n2440gat_reg/NET0131  , \n2446gat_reg/NET0131  , \n2450gat_reg/NET0131  , \n2454gat_reg/NET0131  , \n2458gat_reg/NET0131  , \n2464gat_reg/NET0131  , \n2468gat_reg/NET0131  , \n2472gat_reg/NET0131  , \n2476gat_reg/NET0131  , \n2490gat_reg/NET0131  , \n2495gat_reg/NET0131  , \n2502gat_reg/NET0131  , \n2506gat_reg/NET0131  , \n2510gat_reg/NET0131  , \n2514gat_reg/NET0131  , \n2518gat_reg/NET0131  , \n2526gat_reg/NET0131  , \n2543gat_reg/NET0131  , \n2562gat_reg/NET0131  , \n256gat_reg/NET0131  , \n2588gat_reg/NET0131  , \n2592gat_reg/NET0131  , \n2599gat_reg/NET0131  , \n2622gat_reg/NET0131  , \n2626gat_reg/NET0131  , \n2630gat_reg/NET0131  , \n2634gat_reg/NET0131  , \n2640gat_reg/NET0131  , \n2644gat_reg/NET0131  , \n2658gat_reg/NET0131  , \n271gat_reg/NET0131  , \n3065gat_pad  , \n3066gat_pad  , \n3067gat_pad  , \n3068gat_pad  , \n3069gat_pad  , \n3070gat_pad  , \n3071gat_pad  , \n3072gat_pad  , \n3073gat_pad  , \n3074gat_pad  , \n3075gat_pad  , \n3076gat_pad  , \n3077gat_pad  , \n3078gat_pad  , \n3079gat_pad  , \n3080gat_pad  , \n3081gat_pad  , \n3082gat_pad  , \n3083gat_pad  , \n3084gat_pad  , \n3085gat_pad  , \n3086gat_pad  , \n3087gat_pad  , \n3088gat_pad  , \n3089gat_pad  , \n3090gat_pad  , \n3091gat_pad  , \n3092gat_pad  , \n3093gat_pad  , \n3094gat_pad  , \n3095gat_pad  , \n3097gat_pad  , \n3098gat_pad  , \n3099gat_pad  , \n3100gat_pad  , \n314gat_reg/NET0131  , \n318gat_reg/NET0131  , \n322gat_reg/NET0131  , \n327gat_reg/NET0131  , \n331gat_reg/NET0131  , \n337gat_reg/NET0131  , \n341gat_reg/NET0131  , \n366gat_reg/NET0131  , \n384gat_reg/NET0131  , \n388gat_reg/NET0131  , \n398gat_reg/NET0131  , \n402gat_reg/NET0131  , \n463gat_reg/NET0131  , \n470gat_reg/NET0131  , \n553gat_reg/NET0131  , \n561gat_reg/NET0131  , \n580gat_reg/NET0131  , \n584gat_reg/NET0131  , \n614gat_reg/NET0131  , \n659gat_reg/NET0131  , \n667gat_reg/NET0131  , \n673gat_reg/NET0131  , \n680gat_reg/NET0131  , \n684gat_reg/NET0131  , \n699gat_reg/NET0131  , \n707gat_reg/NET0131  , \n777gat_reg/NET0131  , \n816gat_reg/NET0131  , \n820gat_reg/NET0131  , \n824gat_reg/NET0131  , \n830gat_reg/NET0131  , \n834gat_reg/NET0131  , \n838gat_reg/NET0131  , \n842gat_reg/NET0131  , \n846gat_reg/NET0131  , \n861gat_reg/NET0131  , \n865gat_reg/NET0131  , \n883gat_reg/NET0131  , \n919gat_reg/NET0131  , \n931gat_reg/NET0131  , \n957gat_reg/NET0131  , \_al_n0  , \g17_dup/_0_  , \g6952/_2_  , \g6953/_2_  , \g6961/_0_  , \g7076/_0_  , \g7077/_0_  , \g7079/_0_  , \g7081/_0_  , \g7082/_0_  , \g7083/_0_  , \g7146/_0_  , \g7147/_0_  , \g7148/_0_  , \g7149/_0_  , \g7150/_0_  , \g7151/_0_  , \g7152/_0_  , \g7153/_0_  , \g7154/_0_  , \g7156/_2_  , \g7161/_2_  , \g7165/_2_  , \g7174/_0_  , \g7180/_00_  , \g7182/_3_  , \g7191/_0_  , \g7204/_0_  , \g7209/_3_  , \g7220/_0_  , \g7229/_0_  , \g7233/_0_  , \g7234/_0_  , \g7235/_0_  , \g7236/_0_  , \g7237/_0_  , \g7238/_0_  , \g7241/_3_  , \g7264/_0_  , \g7265/_0_  , \g7266/_0_  , \g7267/_0_  , \g7268/_0_  , \g7301/_0_  , \g7326/_3_  , \g7350/_2_  , \g7352/_0_  , \g7356/_0_  , \g7359/_0_  , \g7389/_3_  , \g7417/_0_  , \g7418/_0_  , \g7419/_0_  , \g7444/_0_  , \g7445/_0_  , \g7449/_3_  , \g7451/_3_  , \g7454/_0_  , \g7467/_3_  , \g7476/_0_  , \g7480/_0_  , \g7494/_0_  , \g7509/_0_  , \g7514/_0_  , \g7517/_3_  , \g7524/_0_  , \g7558/_0_  , \g7560/_0_  , \g7561/_0_  , \g7563/_0_  , \g7567/_0_  , \g7572/_0_  , \g7579/_0_  , \g7605/_0_  , \g7625/_0_  , \g7627/_0_  , \g7671/_0_  , \g7675/_0_  , \g7689/_0_  , \g7697/_0_  , \g7743/_1_  , \g7764/_1_  , \g7769/_0_  , \g7771/_2_  , \g7779/_0_  , \g7852/_0_  , \g7873/_0_  , \g7884/_3_  , \g7889/_0_  , \g7902/_1_  , \g7992/_3_  , \g7994/_3_  , \g7996/_3_  , \g7998/_3_  , \g8000/_3_  , \g8002/_3_  , \g8004/_3_  , \g8006/_3_  , \g8008/_3_  , \g8150/_0_  , \g8151/_0_  , \g8157/_0_  , \g8163/_0_  , \g8172/_0_  , \g8197/_0_  , \g8211/_0_  , \g8223/_0_  , \g8237/_0_  , \g8251/_0_  , \g8261/_0_  , \g8272/_0_  , \g8287/_0_  , \g8647/_0_  , \g8671/_0_  , \g8672/_0_  , \g8735/_0_  , \g8766/_0_  , \g8811/_0_  , \g8821/_0_  , \g8856/_0_  , \g8858/_3_  , \g8868/_0_  , \g8880/_2_  , \g8886/_0_  , \g8900/_0_  , \g8932/_0_  , \g8991/_3_  , \g9014/_3_  , \g9074/_0_  , \g9091/_0_  , \g9105/_0_  , \g9107/_1_  , \g9111/_0_  , \n1332gat_reg/P0001  , \n1363gat_reg/P0001  , \n1394gat_reg/P0001  , \n1433gat_reg/P0001  , \n1775gat_reg/P0001  , \n2025gat_reg/P0001  , \n2029gat_reg/P0001  , \n2033gat_reg/P0001  , \n2044gat_reg/P0001  , \n2121gat_reg/P0001  , \n2125gat_reg/P0001  , \n2458gat_reg/P0001  , \n2472gat_reg/P0001  , \n2592gat_reg/P0001  , \n3104gat_pad  , \n3105gat_pad  , \n3106gat_pad  , \n3107gat_pad  , \n3108gat_pad  , \n3109gat_pad  , \n3110gat_pad  , \n3111gat_pad  , \n3112gat_pad  , \n3113gat_pad  , \n3114gat_pad  , \n3116gat_pad  , \n3117gat_pad  , \n3118gat_pad  , \n3119gat_pad  , \n3120gat_pad  , \n3121gat_pad  , \n3122gat_pad  , \n3123gat_pad  , \n3124gat_pad  , \n3125gat_pad  , \n3126gat_pad  , \n3127gat_pad  , \n3128gat_pad  , \n3130gat_pad  , \n3131gat_pad  , \n3132gat_pad  , \n3133gat_pad  , \n3134gat_pad  , \n3135gat_pad  , \n3136gat_pad  , \n3137gat_pad  , \n3138gat_pad  , \n3140gat_pad  , \n3142gat_pad  , \n3143gat_pad  , \n3144gat_pad  , \n3145gat_pad  , \n3146gat_pad  , \n3147gat_pad  , \n3148gat_pad  , \n3149gat_pad  , \n3150gat_pad  , \n3151gat_pad  , \n684gat_reg/P0001  , \n824gat_reg/P0001  , \n883gat_reg/P0001  );
  input \n1035gat_reg/NET0131  ;
  input \n1045gat_reg/NET0131  ;
  input \n1068gat_reg/NET0131  ;
  input \n1072gat_reg/NET0131  ;
  input \n1080gat_reg/NET0131  ;
  input \n1121gat_reg/NET0131  ;
  input \n1135gat_reg/NET0131  ;
  input \n1148gat_reg/NET0131  ;
  input \n1197gat_reg/NET0131  ;
  input \n1226gat_reg/NET0131  ;
  input \n1241gat_reg/NET0131  ;
  input \n1282gat_reg/NET0131  ;
  input \n1294gat_reg/NET0131  ;
  input \n1312gat_reg/NET0131  ;
  input \n1316gat_reg/NET0131  ;
  input \n1332gat_reg/NET0131  ;
  input \n1336gat_reg/NET0131  ;
  input \n1340gat_reg/NET0131  ;
  input \n1363gat_reg/NET0131  ;
  input \n1389gat_reg/NET0131  ;
  input \n1394gat_reg/NET0131  ;
  input \n1433gat_reg/NET0131  ;
  input \n1456gat_reg/NET0131  ;
  input \n1462gat_reg/NET0131  ;
  input \n148gat_reg/NET0131  ;
  input \n1496gat_reg/NET0131  ;
  input \n1508gat_reg/NET0131  ;
  input \n1525gat_reg/NET0131  ;
  input \n152gat_reg/NET0131  ;
  input \n156gat_reg/NET0131  ;
  input \n1588gat_reg/NET0131  ;
  input \n1596gat_reg/NET0131  ;
  input \n160gat_reg/NET0131  ;
  input \n1675gat_reg/NET0131  ;
  input \n1678gat_reg/NET0131  ;
  input \n1740gat_reg/NET0131  ;
  input \n1748gat_reg/NET0131  ;
  input \n1763gat_reg/NET0131  ;
  input \n1767gat_reg/NET0131  ;
  input \n1771gat_reg/NET0131  ;
  input \n1775gat_reg/NET0131  ;
  input \n1807gat_reg/NET0131  ;
  input \n1821gat_reg/NET0131  ;
  input \n1829gat_reg/NET0131  ;
  input \n1834gat_reg/NET0131  ;
  input \n1850gat_reg/NET0131  ;
  input \n1871gat_reg/NET0131  ;
  input \n1880gat_reg/NET0131  ;
  input \n1899gat_reg/NET0131  ;
  input \n1975gat_reg/NET0131  ;
  input \n2021gat_reg/NET0131  ;
  input \n2025gat_reg/NET0131  ;
  input \n2029gat_reg/NET0131  ;
  input \n2033gat_reg/NET0131  ;
  input \n2037gat_reg/NET0131  ;
  input \n2040gat_reg/NET0131  ;
  input \n2044gat_reg/NET0131  ;
  input \n2061gat_reg/NET0131  ;
  input \n2084gat_reg/NET0131  ;
  input \n2091gat_reg/NET0131  ;
  input \n2095gat_reg/NET0131  ;
  input \n2099gat_reg/NET0131  ;
  input \n2102gat_reg/NET0131  ;
  input \n2110gat_reg/NET0131  ;
  input \n2117gat_reg/NET0131  ;
  input \n2121gat_reg/NET0131  ;
  input \n2125gat_reg/NET0131  ;
  input \n2135gat_reg/NET0131  ;
  input \n2139gat_reg/NET0131  ;
  input \n2143gat_reg/NET0131  ;
  input \n2155gat_reg/NET0131  ;
  input \n2169gat_reg/NET0131  ;
  input \n2176gat_reg/NET0131  ;
  input \n2179gat_reg/NET0131  ;
  input \n2182gat_reg/NET0131  ;
  input \n2190gat_reg/NET0131  ;
  input \n2203gat_reg/NET0131  ;
  input \n2207gat_reg/NET0131  ;
  input \n2262gat_reg/NET0131  ;
  input \n2266gat_reg/NET0131  ;
  input \n2270gat_reg/NET0131  ;
  input \n2319gat_reg/NET0131  ;
  input \n2339gat_reg/NET0131  ;
  input \n2343gat_reg/NET0131  ;
  input \n2347gat_reg/NET0131  ;
  input \n2390gat_reg/NET0131  ;
  input \n2394gat_reg/NET0131  ;
  input \n2399gat_reg/NET0131  ;
  input \n2403gat_reg/NET0131  ;
  input \n2407gat_reg/NET0131  ;
  input \n2440gat_reg/NET0131  ;
  input \n2446gat_reg/NET0131  ;
  input \n2450gat_reg/NET0131  ;
  input \n2454gat_reg/NET0131  ;
  input \n2458gat_reg/NET0131  ;
  input \n2464gat_reg/NET0131  ;
  input \n2468gat_reg/NET0131  ;
  input \n2472gat_reg/NET0131  ;
  input \n2476gat_reg/NET0131  ;
  input \n2490gat_reg/NET0131  ;
  input \n2495gat_reg/NET0131  ;
  input \n2502gat_reg/NET0131  ;
  input \n2506gat_reg/NET0131  ;
  input \n2510gat_reg/NET0131  ;
  input \n2514gat_reg/NET0131  ;
  input \n2518gat_reg/NET0131  ;
  input \n2526gat_reg/NET0131  ;
  input \n2543gat_reg/NET0131  ;
  input \n2562gat_reg/NET0131  ;
  input \n256gat_reg/NET0131  ;
  input \n2588gat_reg/NET0131  ;
  input \n2592gat_reg/NET0131  ;
  input \n2599gat_reg/NET0131  ;
  input \n2622gat_reg/NET0131  ;
  input \n2626gat_reg/NET0131  ;
  input \n2630gat_reg/NET0131  ;
  input \n2634gat_reg/NET0131  ;
  input \n2640gat_reg/NET0131  ;
  input \n2644gat_reg/NET0131  ;
  input \n2658gat_reg/NET0131  ;
  input \n271gat_reg/NET0131  ;
  input \n3065gat_pad  ;
  input \n3066gat_pad  ;
  input \n3067gat_pad  ;
  input \n3068gat_pad  ;
  input \n3069gat_pad  ;
  input \n3070gat_pad  ;
  input \n3071gat_pad  ;
  input \n3072gat_pad  ;
  input \n3073gat_pad  ;
  input \n3074gat_pad  ;
  input \n3075gat_pad  ;
  input \n3076gat_pad  ;
  input \n3077gat_pad  ;
  input \n3078gat_pad  ;
  input \n3079gat_pad  ;
  input \n3080gat_pad  ;
  input \n3081gat_pad  ;
  input \n3082gat_pad  ;
  input \n3083gat_pad  ;
  input \n3084gat_pad  ;
  input \n3085gat_pad  ;
  input \n3086gat_pad  ;
  input \n3087gat_pad  ;
  input \n3088gat_pad  ;
  input \n3089gat_pad  ;
  input \n3090gat_pad  ;
  input \n3091gat_pad  ;
  input \n3092gat_pad  ;
  input \n3093gat_pad  ;
  input \n3094gat_pad  ;
  input \n3095gat_pad  ;
  input \n3097gat_pad  ;
  input \n3098gat_pad  ;
  input \n3099gat_pad  ;
  input \n3100gat_pad  ;
  input \n314gat_reg/NET0131  ;
  input \n318gat_reg/NET0131  ;
  input \n322gat_reg/NET0131  ;
  input \n327gat_reg/NET0131  ;
  input \n331gat_reg/NET0131  ;
  input \n337gat_reg/NET0131  ;
  input \n341gat_reg/NET0131  ;
  input \n366gat_reg/NET0131  ;
  input \n384gat_reg/NET0131  ;
  input \n388gat_reg/NET0131  ;
  input \n398gat_reg/NET0131  ;
  input \n402gat_reg/NET0131  ;
  input \n463gat_reg/NET0131  ;
  input \n470gat_reg/NET0131  ;
  input \n553gat_reg/NET0131  ;
  input \n561gat_reg/NET0131  ;
  input \n580gat_reg/NET0131  ;
  input \n584gat_reg/NET0131  ;
  input \n614gat_reg/NET0131  ;
  input \n659gat_reg/NET0131  ;
  input \n667gat_reg/NET0131  ;
  input \n673gat_reg/NET0131  ;
  input \n680gat_reg/NET0131  ;
  input \n684gat_reg/NET0131  ;
  input \n699gat_reg/NET0131  ;
  input \n707gat_reg/NET0131  ;
  input \n777gat_reg/NET0131  ;
  input \n816gat_reg/NET0131  ;
  input \n820gat_reg/NET0131  ;
  input \n824gat_reg/NET0131  ;
  input \n830gat_reg/NET0131  ;
  input \n834gat_reg/NET0131  ;
  input \n838gat_reg/NET0131  ;
  input \n842gat_reg/NET0131  ;
  input \n846gat_reg/NET0131  ;
  input \n861gat_reg/NET0131  ;
  input \n865gat_reg/NET0131  ;
  input \n883gat_reg/NET0131  ;
  input \n919gat_reg/NET0131  ;
  input \n931gat_reg/NET0131  ;
  input \n957gat_reg/NET0131  ;
  output \_al_n0  ;
  output \g17_dup/_0_  ;
  output \g6952/_2_  ;
  output \g6953/_2_  ;
  output \g6961/_0_  ;
  output \g7076/_0_  ;
  output \g7077/_0_  ;
  output \g7079/_0_  ;
  output \g7081/_0_  ;
  output \g7082/_0_  ;
  output \g7083/_0_  ;
  output \g7146/_0_  ;
  output \g7147/_0_  ;
  output \g7148/_0_  ;
  output \g7149/_0_  ;
  output \g7150/_0_  ;
  output \g7151/_0_  ;
  output \g7152/_0_  ;
  output \g7153/_0_  ;
  output \g7154/_0_  ;
  output \g7156/_2_  ;
  output \g7161/_2_  ;
  output \g7165/_2_  ;
  output \g7174/_0_  ;
  output \g7180/_00_  ;
  output \g7182/_3_  ;
  output \g7191/_0_  ;
  output \g7204/_0_  ;
  output \g7209/_3_  ;
  output \g7220/_0_  ;
  output \g7229/_0_  ;
  output \g7233/_0_  ;
  output \g7234/_0_  ;
  output \g7235/_0_  ;
  output \g7236/_0_  ;
  output \g7237/_0_  ;
  output \g7238/_0_  ;
  output \g7241/_3_  ;
  output \g7264/_0_  ;
  output \g7265/_0_  ;
  output \g7266/_0_  ;
  output \g7267/_0_  ;
  output \g7268/_0_  ;
  output \g7301/_0_  ;
  output \g7326/_3_  ;
  output \g7350/_2_  ;
  output \g7352/_0_  ;
  output \g7356/_0_  ;
  output \g7359/_0_  ;
  output \g7389/_3_  ;
  output \g7417/_0_  ;
  output \g7418/_0_  ;
  output \g7419/_0_  ;
  output \g7444/_0_  ;
  output \g7445/_0_  ;
  output \g7449/_3_  ;
  output \g7451/_3_  ;
  output \g7454/_0_  ;
  output \g7467/_3_  ;
  output \g7476/_0_  ;
  output \g7480/_0_  ;
  output \g7494/_0_  ;
  output \g7509/_0_  ;
  output \g7514/_0_  ;
  output \g7517/_3_  ;
  output \g7524/_0_  ;
  output \g7558/_0_  ;
  output \g7560/_0_  ;
  output \g7561/_0_  ;
  output \g7563/_0_  ;
  output \g7567/_0_  ;
  output \g7572/_0_  ;
  output \g7579/_0_  ;
  output \g7605/_0_  ;
  output \g7625/_0_  ;
  output \g7627/_0_  ;
  output \g7671/_0_  ;
  output \g7675/_0_  ;
  output \g7689/_0_  ;
  output \g7697/_0_  ;
  output \g7743/_1_  ;
  output \g7764/_1_  ;
  output \g7769/_0_  ;
  output \g7771/_2_  ;
  output \g7779/_0_  ;
  output \g7852/_0_  ;
  output \g7873/_0_  ;
  output \g7884/_3_  ;
  output \g7889/_0_  ;
  output \g7902/_1_  ;
  output \g7992/_3_  ;
  output \g7994/_3_  ;
  output \g7996/_3_  ;
  output \g7998/_3_  ;
  output \g8000/_3_  ;
  output \g8002/_3_  ;
  output \g8004/_3_  ;
  output \g8006/_3_  ;
  output \g8008/_3_  ;
  output \g8150/_0_  ;
  output \g8151/_0_  ;
  output \g8157/_0_  ;
  output \g8163/_0_  ;
  output \g8172/_0_  ;
  output \g8197/_0_  ;
  output \g8211/_0_  ;
  output \g8223/_0_  ;
  output \g8237/_0_  ;
  output \g8251/_0_  ;
  output \g8261/_0_  ;
  output \g8272/_0_  ;
  output \g8287/_0_  ;
  output \g8647/_0_  ;
  output \g8671/_0_  ;
  output \g8672/_0_  ;
  output \g8735/_0_  ;
  output \g8766/_0_  ;
  output \g8811/_0_  ;
  output \g8821/_0_  ;
  output \g8856/_0_  ;
  output \g8858/_3_  ;
  output \g8868/_0_  ;
  output \g8880/_2_  ;
  output \g8886/_0_  ;
  output \g8900/_0_  ;
  output \g8932/_0_  ;
  output \g8991/_3_  ;
  output \g9014/_3_  ;
  output \g9074/_0_  ;
  output \g9091/_0_  ;
  output \g9105/_0_  ;
  output \g9107/_1_  ;
  output \g9111/_0_  ;
  output \n1332gat_reg/P0001  ;
  output \n1363gat_reg/P0001  ;
  output \n1394gat_reg/P0001  ;
  output \n1433gat_reg/P0001  ;
  output \n1775gat_reg/P0001  ;
  output \n2025gat_reg/P0001  ;
  output \n2029gat_reg/P0001  ;
  output \n2033gat_reg/P0001  ;
  output \n2044gat_reg/P0001  ;
  output \n2121gat_reg/P0001  ;
  output \n2125gat_reg/P0001  ;
  output \n2458gat_reg/P0001  ;
  output \n2472gat_reg/P0001  ;
  output \n2592gat_reg/P0001  ;
  output \n3104gat_pad  ;
  output \n3105gat_pad  ;
  output \n3106gat_pad  ;
  output \n3107gat_pad  ;
  output \n3108gat_pad  ;
  output \n3109gat_pad  ;
  output \n3110gat_pad  ;
  output \n3111gat_pad  ;
  output \n3112gat_pad  ;
  output \n3113gat_pad  ;
  output \n3114gat_pad  ;
  output \n3116gat_pad  ;
  output \n3117gat_pad  ;
  output \n3118gat_pad  ;
  output \n3119gat_pad  ;
  output \n3120gat_pad  ;
  output \n3121gat_pad  ;
  output \n3122gat_pad  ;
  output \n3123gat_pad  ;
  output \n3124gat_pad  ;
  output \n3125gat_pad  ;
  output \n3126gat_pad  ;
  output \n3127gat_pad  ;
  output \n3128gat_pad  ;
  output \n3130gat_pad  ;
  output \n3131gat_pad  ;
  output \n3132gat_pad  ;
  output \n3133gat_pad  ;
  output \n3134gat_pad  ;
  output \n3135gat_pad  ;
  output \n3136gat_pad  ;
  output \n3137gat_pad  ;
  output \n3138gat_pad  ;
  output \n3140gat_pad  ;
  output \n3142gat_pad  ;
  output \n3143gat_pad  ;
  output \n3144gat_pad  ;
  output \n3145gat_pad  ;
  output \n3146gat_pad  ;
  output \n3147gat_pad  ;
  output \n3148gat_pad  ;
  output \n3149gat_pad  ;
  output \n3150gat_pad  ;
  output \n3151gat_pad  ;
  output \n684gat_reg/P0001  ;
  output \n824gat_reg/P0001  ;
  output \n883gat_reg/P0001  ;
  wire n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 ;
  assign n198 = \n398gat_reg/NET0131  & ~\n402gat_reg/NET0131  ;
  assign n199 = ~\n2454gat_reg/NET0131  & \n846gat_reg/NET0131  ;
  assign n200 = n198 & n199 ;
  assign n201 = ~\n553gat_reg/NET0131  & ~\n777gat_reg/NET0131  ;
  assign n202 = \n553gat_reg/NET0131  & \n777gat_reg/NET0131  ;
  assign n203 = ~n201 & ~n202 ;
  assign n204 = ~\n366gat_reg/NET0131  & ~\n561gat_reg/NET0131  ;
  assign n205 = \n366gat_reg/NET0131  & \n561gat_reg/NET0131  ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = ~\n314gat_reg/NET0131  & n206 ;
  assign n208 = \n314gat_reg/NET0131  & ~n206 ;
  assign n209 = ~n207 & ~n208 ;
  assign n210 = ~n203 & ~n209 ;
  assign n211 = n203 & n209 ;
  assign n212 = ~n210 & ~n211 ;
  assign n213 = \n3088gat_pad  & \n3095gat_pad  ;
  assign n214 = \n3087gat_pad  & \n3093gat_pad  ;
  assign n215 = ~n213 & ~n214 ;
  assign n216 = \n3087gat_pad  & \n3095gat_pad  ;
  assign n217 = \n3086gat_pad  & \n3093gat_pad  ;
  assign n218 = ~n216 & ~n217 ;
  assign n219 = n215 & ~n218 ;
  assign n220 = \n3086gat_pad  & \n3095gat_pad  ;
  assign n221 = \n3085gat_pad  & \n3093gat_pad  ;
  assign n222 = ~n220 & ~n221 ;
  assign n223 = n219 & ~n222 ;
  assign n224 = ~\n318gat_reg/NET0131  & ~\n322gat_reg/NET0131  ;
  assign n225 = \n318gat_reg/NET0131  & \n322gat_reg/NET0131  ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = \n659gat_reg/NET0131  & ~n226 ;
  assign n228 = ~\n659gat_reg/NET0131  & n226 ;
  assign n229 = ~n227 & ~n228 ;
  assign n230 = n223 & ~n229 ;
  assign n231 = ~n212 & n230 ;
  assign n232 = n223 & n229 ;
  assign n233 = n212 & n232 ;
  assign n234 = ~n231 & ~n233 ;
  assign n235 = \n820gat_reg/NET0131  & ~n215 ;
  assign n236 = n218 & ~n235 ;
  assign n237 = ~n215 & ~n218 ;
  assign n238 = ~\n842gat_reg/NET0131  & n237 ;
  assign n239 = ~n236 & ~n238 ;
  assign n240 = ~n222 & ~n239 ;
  assign n241 = ~\n1241gat_reg/NET0131  & n222 ;
  assign n242 = n237 & n241 ;
  assign n243 = \n673gat_reg/NET0131  & n222 ;
  assign n244 = n219 & n243 ;
  assign n245 = ~n242 & ~n244 ;
  assign n246 = ~n240 & n245 ;
  assign n247 = n234 & n246 ;
  assign n248 = ~\n3083gat_pad  & ~\n3084gat_pad  ;
  assign n249 = \n3093gat_pad  & n248 ;
  assign n250 = ~\n3085gat_pad  & ~\n3086gat_pad  ;
  assign n251 = ~\n3088gat_pad  & ~n250 ;
  assign n252 = n249 & n251 ;
  assign n253 = ~\n3085gat_pad  & n248 ;
  assign n254 = \n3086gat_pad  & \n3087gat_pad  ;
  assign n255 = n213 & n254 ;
  assign n256 = n253 & n255 ;
  assign n257 = ~n252 & ~n256 ;
  assign n258 = ~n247 & ~n257 ;
  assign n259 = ~\n3086gat_pad  & ~\n3087gat_pad  ;
  assign n260 = \n3095gat_pad  & ~n259 ;
  assign n261 = n253 & n260 ;
  assign n262 = n249 & ~n250 ;
  assign n263 = n221 & n254 ;
  assign n264 = \n3088gat_pad  & ~n263 ;
  assign n265 = n262 & n264 ;
  assign n266 = ~n261 & ~n265 ;
  assign n267 = ~\n1035gat_reg/NET0131  & ~\n1121gat_reg/NET0131  ;
  assign n268 = \n1035gat_reg/NET0131  & \n1121gat_reg/NET0131  ;
  assign n269 = ~n267 & ~n268 ;
  assign n270 = \n1226gat_reg/NET0131  & ~\n1282gat_reg/NET0131  ;
  assign n271 = ~n269 & n270 ;
  assign n272 = \n1226gat_reg/NET0131  & \n1282gat_reg/NET0131  ;
  assign n273 = n269 & n272 ;
  assign n274 = ~n271 & ~n273 ;
  assign n275 = ~\n1226gat_reg/NET0131  & \n1282gat_reg/NET0131  ;
  assign n276 = ~n269 & n275 ;
  assign n277 = ~\n1226gat_reg/NET0131  & ~\n1282gat_reg/NET0131  ;
  assign n278 = n269 & n277 ;
  assign n279 = ~n276 & ~n278 ;
  assign n280 = n274 & n279 ;
  assign n281 = \n1135gat_reg/NET0131  & ~\n931gat_reg/NET0131  ;
  assign n282 = ~\n1135gat_reg/NET0131  & \n931gat_reg/NET0131  ;
  assign n283 = ~n281 & ~n282 ;
  assign n284 = \n1045gat_reg/NET0131  & ~\n1072gat_reg/NET0131  ;
  assign n285 = ~\n1045gat_reg/NET0131  & \n1072gat_reg/NET0131  ;
  assign n286 = ~n284 & ~n285 ;
  assign n287 = ~n222 & n286 ;
  assign n288 = n219 & n287 ;
  assign n289 = ~n283 & n288 ;
  assign n290 = ~n280 & n289 ;
  assign n291 = n283 & n288 ;
  assign n292 = n280 & n291 ;
  assign n293 = ~n290 & ~n292 ;
  assign n294 = n283 & ~n286 ;
  assign n295 = n223 & n294 ;
  assign n296 = ~n280 & n295 ;
  assign n297 = ~n283 & ~n286 ;
  assign n298 = n223 & n297 ;
  assign n299 = n280 & n298 ;
  assign n300 = ~n296 & ~n299 ;
  assign n301 = n293 & n300 ;
  assign n302 = ~\n842gat_reg/NET0131  & n222 ;
  assign n303 = n237 & n302 ;
  assign n304 = ~n215 & n218 ;
  assign n305 = ~\n830gat_reg/NET0131  & ~n222 ;
  assign n306 = n304 & n305 ;
  assign n307 = ~n303 & ~n306 ;
  assign n308 = n301 & n307 ;
  assign n309 = ~n266 & ~n308 ;
  assign n310 = ~n258 & ~n309 ;
  assign n311 = \n2476gat_reg/NET0131  & \n2518gat_reg/NET0131  ;
  assign n312 = \n2464gat_reg/NET0131  & n311 ;
  assign n313 = \n2526gat_reg/NET0131  & \n2599gat_reg/NET0131  ;
  assign n314 = \n2468gat_reg/NET0131  & ~\n3090gat_pad  ;
  assign n315 = n313 & n314 ;
  assign n316 = n312 & n315 ;
  assign n317 = ~\n659gat_reg/NET0131  & \n667gat_reg/NET0131  ;
  assign n318 = ~n226 & n317 ;
  assign n319 = \n659gat_reg/NET0131  & \n667gat_reg/NET0131  ;
  assign n320 = n226 & n319 ;
  assign n321 = ~n318 & ~n320 ;
  assign n322 = ~n212 & ~n321 ;
  assign n323 = \n667gat_reg/NET0131  & ~n229 ;
  assign n324 = n212 & n323 ;
  assign n325 = ~n322 & ~n324 ;
  assign n326 = ~\n667gat_reg/NET0131  & ~n229 ;
  assign n327 = ~n212 & n326 ;
  assign n328 = ~\n659gat_reg/NET0131  & ~\n667gat_reg/NET0131  ;
  assign n329 = ~n226 & n328 ;
  assign n330 = \n659gat_reg/NET0131  & ~\n667gat_reg/NET0131  ;
  assign n331 = n226 & n330 ;
  assign n332 = ~n329 & ~n331 ;
  assign n333 = n212 & ~n332 ;
  assign n334 = ~n327 & ~n333 ;
  assign n335 = n325 & n334 ;
  assign n336 = \n3069gat_pad  & \n3093gat_pad  ;
  assign n337 = \n3078gat_pad  & \n3095gat_pad  ;
  assign n338 = ~n336 & ~n337 ;
  assign n339 = \n2155gat_reg/NET0131  & ~\n2622gat_reg/NET0131  ;
  assign n340 = \n2490gat_reg/NET0131  & \n2543gat_reg/NET0131  ;
  assign n341 = ~\n2626gat_reg/NET0131  & \n2630gat_reg/NET0131  ;
  assign n342 = n340 & n341 ;
  assign n343 = n339 & n342 ;
  assign n344 = ~\n2543gat_reg/NET0131  & \n2630gat_reg/NET0131  ;
  assign n345 = ~\n2622gat_reg/NET0131  & \n2626gat_reg/NET0131  ;
  assign n346 = ~\n2155gat_reg/NET0131  & ~\n2490gat_reg/NET0131  ;
  assign n347 = n345 & n346 ;
  assign n348 = n344 & n347 ;
  assign n349 = ~n343 & ~n348 ;
  assign n350 = ~\n2203gat_reg/NET0131  & ~\n2207gat_reg/NET0131  ;
  assign n351 = ~\n2343gat_reg/NET0131  & \n2399gat_reg/NET0131  ;
  assign n352 = \n2562gat_reg/NET0131  & n351 ;
  assign n353 = n350 & n352 ;
  assign n354 = ~n349 & ~n353 ;
  assign n355 = \n398gat_reg/NET0131  & \n402gat_reg/NET0131  ;
  assign n356 = ~\n919gat_reg/NET0131  & n199 ;
  assign n357 = n355 & n356 ;
  assign n358 = ~\n398gat_reg/NET0131  & ~\n402gat_reg/NET0131  ;
  assign n359 = n199 & ~n358 ;
  assign n360 = ~\n398gat_reg/NET0131  & ~\n919gat_reg/NET0131  ;
  assign n361 = ~n355 & ~n360 ;
  assign n362 = n359 & n361 ;
  assign n363 = ~n357 & ~n362 ;
  assign n364 = \n2343gat_reg/NET0131  & \n2399gat_reg/NET0131  ;
  assign n365 = ~\n2207gat_reg/NET0131  & ~n364 ;
  assign n366 = \n2203gat_reg/NET0131  & ~\n2207gat_reg/NET0131  ;
  assign n367 = ~\n2207gat_reg/NET0131  & \n2562gat_reg/NET0131  ;
  assign n368 = ~n366 & ~n367 ;
  assign n369 = ~n365 & n368 ;
  assign n370 = ~n363 & ~n369 ;
  assign n371 = n354 & n370 ;
  assign n372 = n338 & ~n371 ;
  assign n373 = \n3070gat_pad  & \n3093gat_pad  ;
  assign n374 = \n3079gat_pad  & \n3095gat_pad  ;
  assign n375 = ~n373 & ~n374 ;
  assign n376 = ~n371 & n375 ;
  assign n377 = \n3072gat_pad  & \n3093gat_pad  ;
  assign n378 = \n3081gat_pad  & \n3095gat_pad  ;
  assign n379 = ~n377 & ~n378 ;
  assign n380 = ~n371 & n379 ;
  assign n381 = \n3071gat_pad  & \n3093gat_pad  ;
  assign n382 = \n3080gat_pad  & \n3095gat_pad  ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = ~n371 & n383 ;
  assign n385 = \n3065gat_pad  & \n3093gat_pad  ;
  assign n386 = \n3074gat_pad  & \n3095gat_pad  ;
  assign n387 = ~n385 & ~n386 ;
  assign n388 = ~n371 & n387 ;
  assign n389 = \n3073gat_pad  & \n3093gat_pad  ;
  assign n390 = \n3082gat_pad  & \n3095gat_pad  ;
  assign n391 = ~n389 & ~n390 ;
  assign n392 = ~n371 & n391 ;
  assign n393 = \n1871gat_reg/NET0131  & ~\n3085gat_pad  ;
  assign n394 = n248 & n393 ;
  assign n395 = \n3094gat_pad  & n216 ;
  assign n396 = n394 & n395 ;
  assign n397 = ~\n3088gat_pad  & n220 ;
  assign n398 = n394 & n397 ;
  assign n399 = n396 & n398 ;
  assign n400 = \n1871gat_reg/NET0131  & \n3093gat_pad  ;
  assign n401 = n248 & n400 ;
  assign n402 = ~\n3087gat_pad  & \n3088gat_pad  ;
  assign n403 = n401 & n402 ;
  assign n404 = ~\n3091gat_pad  & ~\n3092gat_pad  ;
  assign n405 = \n3085gat_pad  & \n3086gat_pad  ;
  assign n406 = ~n404 & n405 ;
  assign n407 = n403 & n406 ;
  assign n408 = ~n399 & ~n407 ;
  assign n409 = \n3068gat_pad  & ~n408 ;
  assign n410 = ~n371 & ~n409 ;
  assign n411 = \n3065gat_pad  & ~n408 ;
  assign n412 = ~n371 & ~n411 ;
  assign n413 = \n3069gat_pad  & ~n408 ;
  assign n414 = ~n371 & ~n413 ;
  assign n415 = \n3066gat_pad  & ~n408 ;
  assign n416 = ~n371 & ~n415 ;
  assign n417 = \n3067gat_pad  & ~n408 ;
  assign n418 = ~n371 & ~n417 ;
  assign n419 = \n3070gat_pad  & ~n408 ;
  assign n420 = ~n371 & ~n419 ;
  assign n421 = \n3073gat_pad  & ~n408 ;
  assign n422 = ~n371 & ~n421 ;
  assign n423 = \n3072gat_pad  & ~n408 ;
  assign n424 = ~n371 & ~n423 ;
  assign n425 = \n3071gat_pad  & ~n408 ;
  assign n426 = ~n371 & ~n425 ;
  assign n427 = ~\n2403gat_reg/NET0131  & ~\n402gat_reg/NET0131  ;
  assign n428 = \n2403gat_reg/NET0131  & \n402gat_reg/NET0131  ;
  assign n429 = ~n427 & ~n428 ;
  assign n430 = \n2347gat_reg/NET0131  & ~\n2407gat_reg/NET0131  ;
  assign n431 = \n398gat_reg/NET0131  & n430 ;
  assign n432 = ~n429 & n431 ;
  assign n433 = ~\n2394gat_reg/NET0131  & ~\n2440gat_reg/NET0131  ;
  assign n434 = ~\n846gat_reg/NET0131  & ~\n919gat_reg/NET0131  ;
  assign n435 = n433 & n434 ;
  assign n436 = ~\n846gat_reg/NET0131  & \n919gat_reg/NET0131  ;
  assign n437 = ~\n2394gat_reg/NET0131  & \n2440gat_reg/NET0131  ;
  assign n438 = n436 & n437 ;
  assign n439 = \n2394gat_reg/NET0131  & ~\n2440gat_reg/NET0131  ;
  assign n440 = \n846gat_reg/NET0131  & ~\n919gat_reg/NET0131  ;
  assign n441 = n439 & n440 ;
  assign n442 = ~n438 & ~n441 ;
  assign n443 = ~n435 & n442 ;
  assign n444 = n432 & ~n443 ;
  assign n445 = \n846gat_reg/NET0131  & \n919gat_reg/NET0131  ;
  assign n446 = \n2394gat_reg/NET0131  & \n2440gat_reg/NET0131  ;
  assign n447 = n445 & n446 ;
  assign n448 = n432 & n447 ;
  assign n449 = ~\n2347gat_reg/NET0131  & \n2403gat_reg/NET0131  ;
  assign n450 = ~\n2407gat_reg/NET0131  & n449 ;
  assign n451 = n446 & n450 ;
  assign n452 = ~n448 & ~n451 ;
  assign n453 = ~n444 & n452 ;
  assign n454 = ~\n1763gat_reg/NET0131  & ~\n1880gat_reg/NET0131  ;
  assign n455 = \n2102gat_reg/NET0131  & ~n454 ;
  assign n456 = \n1850gat_reg/NET0131  & \n2143gat_reg/NET0131  ;
  assign n457 = ~\n1899gat_reg/NET0131  & ~\n2061gat_reg/NET0131  ;
  assign n458 = ~\n2139gat_reg/NET0131  & n457 ;
  assign n459 = n456 & n458 ;
  assign n460 = n455 & n459 ;
  assign n461 = \n2061gat_reg/NET0131  & ~n455 ;
  assign n462 = ~\n1899gat_reg/NET0131  & \n2139gat_reg/NET0131  ;
  assign n463 = ~\n1850gat_reg/NET0131  & \n2143gat_reg/NET0131  ;
  assign n464 = n462 & n463 ;
  assign n465 = n461 & n464 ;
  assign n466 = ~n460 & ~n465 ;
  assign n467 = \n1767gat_reg/NET0131  & \n1834gat_reg/NET0131  ;
  assign n468 = \n1880gat_reg/NET0131  & n467 ;
  assign n469 = ~n466 & ~n468 ;
  assign n470 = ~n453 & n469 ;
  assign n471 = \n1880gat_reg/NET0131  & \n2021gat_reg/NET0131  ;
  assign n472 = ~\n1312gat_reg/NET0131  & \n1775gat_reg/NET0131  ;
  assign n473 = \n3100gat_pad  & ~n472 ;
  assign n474 = \n2510gat_reg/NET0131  & \n2588gat_reg/NET0131  ;
  assign n475 = \n2658gat_reg/NET0131  & n474 ;
  assign n476 = \n2502gat_reg/NET0131  & \n2506gat_reg/NET0131  ;
  assign n477 = ~n472 & n476 ;
  assign n478 = n475 & n477 ;
  assign n479 = ~n473 & ~n478 ;
  assign n480 = ~n471 & ~n479 ;
  assign n481 = ~n470 & n480 ;
  assign n482 = n437 & n450 ;
  assign n483 = n465 & ~n482 ;
  assign n484 = ~n470 & n483 ;
  assign n485 = ~\n2490gat_reg/NET0131  & ~\n2634gat_reg/NET0131  ;
  assign n486 = \n2490gat_reg/NET0131  & \n2634gat_reg/NET0131  ;
  assign n487 = ~n485 & ~n486 ;
  assign n488 = \n2622gat_reg/NET0131  & ~\n2626gat_reg/NET0131  ;
  assign n489 = ~n345 & ~n488 ;
  assign n490 = \n2543gat_reg/NET0131  & ~\n2630gat_reg/NET0131  ;
  assign n491 = ~n344 & ~n490 ;
  assign n492 = n489 & n491 ;
  assign n493 = ~n489 & ~n491 ;
  assign n494 = ~n492 & ~n493 ;
  assign n495 = n487 & n494 ;
  assign n496 = ~n487 & ~n494 ;
  assign n497 = ~n495 & ~n496 ;
  assign n498 = n459 & ~n470 ;
  assign n499 = ~\n1740gat_reg/NET0131  & n464 ;
  assign n500 = n461 & n499 ;
  assign n501 = ~\n1496gat_reg/NET0131  & ~\n2091gat_reg/NET0131  ;
  assign n502 = n455 & ~n501 ;
  assign n503 = n459 & n502 ;
  assign n504 = ~n500 & ~n503 ;
  assign n505 = ~\n2061gat_reg/NET0131  & n456 ;
  assign n506 = n462 & n505 ;
  assign n507 = n455 & n501 ;
  assign n508 = n506 & n507 ;
  assign n509 = ~\n2139gat_reg/NET0131  & ~\n2143gat_reg/NET0131  ;
  assign n510 = n457 & n509 ;
  assign n511 = \n1850gat_reg/NET0131  & n510 ;
  assign n512 = \n1740gat_reg/NET0131  & ~n455 ;
  assign n513 = n511 & n512 ;
  assign n514 = ~n508 & ~n513 ;
  assign n515 = n504 & n514 ;
  assign n516 = ~n437 & ~n455 ;
  assign n517 = n450 & ~n516 ;
  assign n518 = ~\n2190gat_reg/NET0131  & ~\n2262gat_reg/NET0131  ;
  assign n519 = ~\n2135gat_reg/NET0131  & ~\n2179gat_reg/NET0131  ;
  assign n520 = n518 & n519 ;
  assign n521 = \n2182gat_reg/NET0131  & ~n520 ;
  assign n522 = n517 & ~n521 ;
  assign n523 = ~n439 & n455 ;
  assign n524 = n522 & ~n523 ;
  assign n525 = ~n515 & n524 ;
  assign n526 = \n2630gat_reg/NET0131  & n340 ;
  assign n527 = n488 & n526 ;
  assign n528 = \n2562gat_reg/NET0131  & n364 ;
  assign n529 = n366 & n528 ;
  assign n530 = n527 & n529 ;
  assign n531 = n475 & n476 ;
  assign n532 = ~\n3100gat_pad  & ~n531 ;
  assign n533 = ~\n2135gat_reg/NET0131  & n518 ;
  assign n534 = \n2135gat_reg/NET0131  & ~n518 ;
  assign n535 = ~n533 & ~n534 ;
  assign n536 = \n2099gat_reg/NET0131  & ~n471 ;
  assign n537 = \n2037gat_reg/NET0131  & \n2095gat_reg/NET0131  ;
  assign n538 = ~n536 & n537 ;
  assign n539 = n535 & n538 ;
  assign n540 = ~n532 & n539 ;
  assign n541 = \n2190gat_reg/NET0131  & ~\n2262gat_reg/NET0131  ;
  assign n542 = \n2266gat_reg/NET0131  & ~n541 ;
  assign n543 = ~\n2266gat_reg/NET0131  & n541 ;
  assign n544 = ~n542 & ~n543 ;
  assign n545 = n538 & n544 ;
  assign n546 = ~n532 & n545 ;
  assign n547 = \n684gat_reg/NET0131  & ~\n816gat_reg/NET0131  ;
  assign n548 = ~\n684gat_reg/NET0131  & \n816gat_reg/NET0131  ;
  assign n549 = ~n547 & ~n548 ;
  assign n550 = \n699gat_reg/NET0131  & ~\n824gat_reg/NET0131  ;
  assign n551 = ~\n699gat_reg/NET0131  & \n824gat_reg/NET0131  ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = ~\n680gat_reg/NET0131  & ~\n883gat_reg/NET0131  ;
  assign n554 = \n680gat_reg/NET0131  & \n883gat_reg/NET0131  ;
  assign n555 = ~n553 & ~n554 ;
  assign n556 = ~n552 & ~n555 ;
  assign n557 = n552 & n555 ;
  assign n558 = ~n556 & ~n557 ;
  assign n559 = ~\n580gat_reg/NET0131  & ~\n820gat_reg/NET0131  ;
  assign n560 = \n580gat_reg/NET0131  & \n820gat_reg/NET0131  ;
  assign n561 = ~n559 & ~n560 ;
  assign n562 = \n584gat_reg/NET0131  & n561 ;
  assign n563 = ~\n584gat_reg/NET0131  & ~n561 ;
  assign n564 = ~n562 & ~n563 ;
  assign n565 = ~n558 & ~n564 ;
  assign n566 = n558 & n564 ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = ~n549 & ~n567 ;
  assign n569 = n549 & n567 ;
  assign n570 = ~n568 & ~n569 ;
  assign n571 = ~\n2390gat_reg/NET0131  & ~\n2495gat_reg/NET0131  ;
  assign n572 = \n2390gat_reg/NET0131  & \n2495gat_reg/NET0131  ;
  assign n573 = ~n571 & ~n572 ;
  assign n574 = \n2270gat_reg/NET0131  & ~\n2339gat_reg/NET0131  ;
  assign n575 = ~\n2270gat_reg/NET0131  & \n2339gat_reg/NET0131  ;
  assign n576 = ~n574 & ~n575 ;
  assign n577 = n573 & n576 ;
  assign n578 = ~n573 & ~n576 ;
  assign n579 = ~n577 & ~n578 ;
  assign n580 = \n2190gat_reg/NET0131  & \n2262gat_reg/NET0131  ;
  assign n581 = n538 & ~n580 ;
  assign n582 = ~n532 & n581 ;
  assign n583 = ~n532 & n538 ;
  assign n584 = \n1899gat_reg/NET0131  & \n2139gat_reg/NET0131  ;
  assign n585 = n583 & ~n584 ;
  assign n586 = n515 & n585 ;
  assign n587 = \n2143gat_reg/NET0131  & ~n458 ;
  assign n588 = ~n510 & ~n587 ;
  assign n589 = n583 & n588 ;
  assign n590 = n515 & n589 ;
  assign n591 = ~\n1899gat_reg/NET0131  & ~\n2139gat_reg/NET0131  ;
  assign n592 = \n2061gat_reg/NET0131  & n591 ;
  assign n593 = ~\n2061gat_reg/NET0131  & ~n591 ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = n583 & ~n594 ;
  assign n596 = n515 & n595 ;
  assign n597 = ~\n1850gat_reg/NET0131  & ~n510 ;
  assign n598 = ~n511 & ~n597 ;
  assign n599 = n583 & ~n598 ;
  assign n600 = n515 & n599 ;
  assign n601 = ~n457 & ~n462 ;
  assign n602 = ~n510 & ~n601 ;
  assign n603 = \n1975gat_reg/NET0131  & n602 ;
  assign n604 = ~\n1975gat_reg/NET0131  & ~n602 ;
  assign n605 = ~n603 & ~n604 ;
  assign n606 = n583 & ~n605 ;
  assign n607 = n515 & n606 ;
  assign n608 = ~n434 & ~n445 ;
  assign n609 = ~\n398gat_reg/NET0131  & \n402gat_reg/NET0131  ;
  assign n610 = ~n198 & ~n609 ;
  assign n611 = ~n608 & ~n610 ;
  assign n612 = n608 & n610 ;
  assign n613 = ~n611 & ~n612 ;
  assign n614 = ~\n830gat_reg/NET0131  & ~\n834gat_reg/NET0131  ;
  assign n615 = \n830gat_reg/NET0131  & \n834gat_reg/NET0131  ;
  assign n616 = ~n614 & ~n615 ;
  assign n617 = \n614gat_reg/NET0131  & ~\n838gat_reg/NET0131  ;
  assign n618 = ~\n614gat_reg/NET0131  & \n838gat_reg/NET0131  ;
  assign n619 = ~n617 & ~n618 ;
  assign n620 = \n707gat_reg/NET0131  & n619 ;
  assign n621 = ~n616 & n620 ;
  assign n622 = ~n613 & n621 ;
  assign n623 = ~\n707gat_reg/NET0131  & n619 ;
  assign n624 = n616 & n623 ;
  assign n625 = ~n613 & n624 ;
  assign n626 = ~n622 & ~n625 ;
  assign n627 = ~n616 & n623 ;
  assign n628 = n616 & n620 ;
  assign n629 = ~n627 & ~n628 ;
  assign n630 = n613 & ~n629 ;
  assign n631 = n626 & ~n630 ;
  assign n632 = \n707gat_reg/NET0131  & ~n619 ;
  assign n633 = ~n616 & n632 ;
  assign n634 = n613 & n633 ;
  assign n635 = ~\n707gat_reg/NET0131  & ~n619 ;
  assign n636 = n616 & n635 ;
  assign n637 = n613 & n636 ;
  assign n638 = ~n634 & ~n637 ;
  assign n639 = ~n616 & n635 ;
  assign n640 = ~n613 & n639 ;
  assign n641 = n616 & n632 ;
  assign n642 = ~n613 & n641 ;
  assign n643 = ~n640 & ~n642 ;
  assign n644 = n638 & n643 ;
  assign n645 = n631 & n644 ;
  assign n646 = n517 & ~n523 ;
  assign n647 = n583 & ~n646 ;
  assign n648 = ~\n2403gat_reg/NET0131  & n433 ;
  assign n649 = ~\n2347gat_reg/NET0131  & ~n648 ;
  assign n650 = \n2347gat_reg/NET0131  & ~\n2403gat_reg/NET0131  ;
  assign n651 = n433 & n650 ;
  assign n652 = ~n649 & ~n651 ;
  assign n653 = n647 & ~n652 ;
  assign n654 = ~\n2347gat_reg/NET0131  & ~\n2407gat_reg/NET0131  ;
  assign n655 = n648 & n654 ;
  assign n656 = ~\n2347gat_reg/NET0131  & ~\n2403gat_reg/NET0131  ;
  assign n657 = n433 & n656 ;
  assign n658 = \n2407gat_reg/NET0131  & ~n657 ;
  assign n659 = ~n655 & ~n658 ;
  assign n660 = n647 & n659 ;
  assign n661 = ~\n2644gat_reg/NET0131  & n439 ;
  assign n662 = ~\n2440gat_reg/NET0131  & ~\n2644gat_reg/NET0131  ;
  assign n663 = n650 & n662 ;
  assign n664 = ~n661 & ~n663 ;
  assign n665 = ~\n2440gat_reg/NET0131  & n650 ;
  assign n666 = \n2644gat_reg/NET0131  & ~n439 ;
  assign n667 = ~n665 & n666 ;
  assign n668 = n538 & ~n667 ;
  assign n669 = ~n532 & n668 ;
  assign n670 = ~n646 & n669 ;
  assign n671 = n664 & n670 ;
  assign n672 = \n2403gat_reg/NET0131  & ~n433 ;
  assign n673 = ~n648 & ~n672 ;
  assign n674 = n538 & n673 ;
  assign n675 = ~n532 & n674 ;
  assign n676 = ~n646 & n675 ;
  assign n677 = ~\n2440gat_reg/NET0131  & ~n455 ;
  assign n678 = ~\n2440gat_reg/NET0131  & ~n450 ;
  assign n679 = ~n677 & ~n678 ;
  assign n680 = ~\n2394gat_reg/NET0131  & n455 ;
  assign n681 = ~\n2394gat_reg/NET0131  & ~n450 ;
  assign n682 = ~n680 & ~n681 ;
  assign n683 = n679 & n682 ;
  assign n684 = n583 & ~n683 ;
  assign n685 = ~\n2347gat_reg/NET0131  & \n2407gat_reg/NET0131  ;
  assign n686 = ~\n2403gat_reg/NET0131  & n685 ;
  assign n687 = n437 & n686 ;
  assign n688 = ~n466 & n687 ;
  assign n689 = \n1850gat_reg/NET0131  & ~\n2143gat_reg/NET0131  ;
  assign n690 = \n2061gat_reg/NET0131  & n462 ;
  assign n691 = ~n455 & n690 ;
  assign n692 = n689 & n691 ;
  assign n693 = ~\n2454gat_reg/NET0131  & ~\n846gat_reg/NET0131  ;
  assign n694 = n355 & n693 ;
  assign n695 = n363 & ~n694 ;
  assign n696 = ~\n1316gat_reg/NET0131  & ~\n1775gat_reg/NET0131  ;
  assign n697 = ~\n2040gat_reg/NET0131  & n696 ;
  assign n698 = \n1241gat_reg/NET0131  & ~\n957gat_reg/NET0131  ;
  assign n699 = ~\n1241gat_reg/NET0131  & \n957gat_reg/NET0131  ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = \n1294gat_reg/NET0131  & ~\n673gat_reg/NET0131  ;
  assign n702 = ~\n1294gat_reg/NET0131  & \n673gat_reg/NET0131  ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = ~\n1068gat_reg/NET0131  & ~\n861gat_reg/NET0131  ;
  assign n705 = \n1068gat_reg/NET0131  & \n861gat_reg/NET0131  ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = ~n703 & ~n706 ;
  assign n708 = n703 & n706 ;
  assign n709 = ~n707 & ~n708 ;
  assign n710 = ~\n1148gat_reg/NET0131  & ~\n865gat_reg/NET0131  ;
  assign n711 = \n1148gat_reg/NET0131  & \n865gat_reg/NET0131  ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = \n1080gat_reg/NET0131  & n712 ;
  assign n714 = ~\n1080gat_reg/NET0131  & ~n712 ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = ~n709 & ~n715 ;
  assign n717 = n709 & n715 ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = ~n700 & ~n718 ;
  assign n720 = n700 & n718 ;
  assign n721 = ~n719 & ~n720 ;
  assign n722 = ~\n2454gat_reg/NET0131  & n198 ;
  assign n723 = n436 & n722 ;
  assign n724 = \n2446gat_reg/NET0131  & \n2450gat_reg/NET0131  ;
  assign n725 = ~\n3100gat_pad  & ~n724 ;
  assign n726 = \n1821gat_reg/NET0131  & ~\n1829gat_reg/NET0131  ;
  assign n727 = \n2472gat_reg/NET0131  & ~n726 ;
  assign n728 = ~n725 & n727 ;
  assign n729 = n723 & n728 ;
  assign n730 = ~\n2454gat_reg/NET0131  & ~\n271gat_reg/NET0131  ;
  assign n731 = n728 & n730 ;
  assign n732 = n434 & n722 ;
  assign n733 = n728 & n732 ;
  assign n734 = ~\n2454gat_reg/NET0131  & ~\n388gat_reg/NET0131  ;
  assign n735 = n198 & n734 ;
  assign n736 = n445 & n735 ;
  assign n737 = \n331gat_reg/NET0131  & ~n736 ;
  assign n738 = n216 & n394 ;
  assign n739 = \n3094gat_pad  & ~n738 ;
  assign n740 = \n3088gat_pad  & n220 ;
  assign n741 = n394 & n740 ;
  assign n742 = n739 & n741 ;
  assign n743 = ~\n3088gat_pad  & n401 ;
  assign n744 = \n3085gat_pad  & ~\n3086gat_pad  ;
  assign n745 = ~n404 & n744 ;
  assign n746 = \n3087gat_pad  & n745 ;
  assign n747 = n743 & n746 ;
  assign n748 = ~\n331gat_reg/NET0131  & ~\n388gat_reg/NET0131  ;
  assign n749 = n445 & n748 ;
  assign n750 = n722 & n749 ;
  assign n751 = ~n747 & ~n750 ;
  assign n752 = ~n742 & n751 ;
  assign n753 = ~n737 & n752 ;
  assign n754 = \n3080gat_pad  & n741 ;
  assign n755 = n739 & n754 ;
  assign n756 = \n3071gat_pad  & ~\n3088gat_pad  ;
  assign n757 = n401 & n756 ;
  assign n758 = n746 & n757 ;
  assign n759 = ~n755 & ~n758 ;
  assign n760 = ~n753 & n759 ;
  assign n761 = \n3087gat_pad  & \n3088gat_pad  ;
  assign n762 = n745 & n761 ;
  assign n763 = n401 & n762 ;
  assign n764 = \n3065gat_pad  & n763 ;
  assign n765 = \n3065gat_pad  & n741 ;
  assign n766 = n739 & n765 ;
  assign n767 = ~n764 & ~n766 ;
  assign n768 = ~n742 & ~n763 ;
  assign n769 = ~\n152gat_reg/NET0131  & ~\n156gat_reg/NET0131  ;
  assign n770 = n198 & n769 ;
  assign n771 = ~\n256gat_reg/NET0131  & ~\n919gat_reg/NET0131  ;
  assign n772 = n199 & n771 ;
  assign n773 = n770 & n772 ;
  assign n774 = ~\n148gat_reg/NET0131  & ~n773 ;
  assign n775 = \n148gat_reg/NET0131  & n773 ;
  assign n776 = ~n774 & ~n775 ;
  assign n777 = n768 & ~n776 ;
  assign n778 = n767 & ~n777 ;
  assign n779 = n198 & n356 ;
  assign n780 = ~\n152gat_reg/NET0131  & \n256gat_reg/NET0131  ;
  assign n781 = ~\n156gat_reg/NET0131  & ~n780 ;
  assign n782 = n779 & ~n781 ;
  assign n783 = ~\n470gat_reg/NET0131  & ~n782 ;
  assign n784 = \n470gat_reg/NET0131  & ~n781 ;
  assign n785 = n779 & n784 ;
  assign n786 = ~n783 & ~n785 ;
  assign n787 = n768 & ~n786 ;
  assign n788 = \n3073gat_pad  & n763 ;
  assign n789 = \n3073gat_pad  & n741 ;
  assign n790 = n739 & n789 ;
  assign n791 = ~n788 & ~n790 ;
  assign n792 = ~n787 & n791 ;
  assign n793 = ~\n3084gat_pad  & ~\n3085gat_pad  ;
  assign n794 = \n3084gat_pad  & \n3085gat_pad  ;
  assign n795 = ~n793 & ~n794 ;
  assign n796 = \n3089gat_pad  & n795 ;
  assign n797 = ~\n3089gat_pad  & ~n795 ;
  assign n798 = ~n796 & ~n797 ;
  assign n799 = ~\n3083gat_pad  & ~\n3088gat_pad  ;
  assign n800 = \n3083gat_pad  & \n3088gat_pad  ;
  assign n801 = ~n799 & ~n800 ;
  assign n802 = ~n254 & ~n259 ;
  assign n803 = n801 & ~n802 ;
  assign n804 = ~n798 & n803 ;
  assign n805 = n801 & n802 ;
  assign n806 = n798 & n805 ;
  assign n807 = ~n804 & ~n806 ;
  assign n808 = ~n801 & ~n802 ;
  assign n809 = n798 & n808 ;
  assign n810 = ~n801 & n802 ;
  assign n811 = ~n798 & n810 ;
  assign n812 = ~n809 & ~n811 ;
  assign n813 = n807 & n812 ;
  assign n814 = n356 & n770 ;
  assign n815 = \n256gat_reg/NET0131  & ~n814 ;
  assign n816 = ~n773 & ~n815 ;
  assign n817 = n768 & n816 ;
  assign n818 = \n3066gat_pad  & n763 ;
  assign n819 = \n3066gat_pad  & n741 ;
  assign n820 = n739 & n819 ;
  assign n821 = ~n818 & ~n820 ;
  assign n822 = ~n817 & n821 ;
  assign n823 = ~n742 & ~n747 ;
  assign n824 = \n327gat_reg/NET0131  & ~n750 ;
  assign n825 = ~\n2454gat_reg/NET0131  & ~\n327gat_reg/NET0131  ;
  assign n826 = n198 & n825 ;
  assign n827 = n749 & n826 ;
  assign n828 = ~n824 & ~n827 ;
  assign n829 = n823 & n828 ;
  assign n830 = \n3079gat_pad  & n741 ;
  assign n831 = n739 & n830 ;
  assign n832 = \n3070gat_pad  & \n3087gat_pad  ;
  assign n833 = n745 & n832 ;
  assign n834 = n743 & n833 ;
  assign n835 = ~n831 & ~n834 ;
  assign n836 = ~n829 & n835 ;
  assign n837 = ~\n156gat_reg/NET0131  & n198 ;
  assign n838 = n356 & n837 ;
  assign n839 = \n152gat_reg/NET0131  & ~n838 ;
  assign n840 = ~n763 & ~n814 ;
  assign n841 = ~n742 & n840 ;
  assign n842 = ~n839 & n841 ;
  assign n843 = \n3067gat_pad  & n763 ;
  assign n844 = \n3067gat_pad  & n741 ;
  assign n845 = n739 & n844 ;
  assign n846 = ~n843 & ~n845 ;
  assign n847 = ~n842 & n846 ;
  assign n848 = \n919gat_reg/NET0131  & n609 ;
  assign n849 = n199 & n848 ;
  assign n850 = ~n694 & ~n849 ;
  assign n851 = ~n357 & ~n722 ;
  assign n852 = n850 & n851 ;
  assign n853 = \n156gat_reg/NET0131  & ~n779 ;
  assign n854 = ~n838 & ~n853 ;
  assign n855 = n768 & n854 ;
  assign n856 = \n3068gat_pad  & n763 ;
  assign n857 = \n3068gat_pad  & n741 ;
  assign n858 = n739 & n857 ;
  assign n859 = ~n856 & ~n858 ;
  assign n860 = ~n855 & n859 ;
  assign n861 = \n3067gat_pad  & \n3087gat_pad  ;
  assign n862 = n745 & n861 ;
  assign n863 = n743 & n862 ;
  assign n864 = \n3076gat_pad  & n741 ;
  assign n865 = n739 & n864 ;
  assign n866 = ~n863 & ~n865 ;
  assign n867 = \n3068gat_pad  & \n3087gat_pad  ;
  assign n868 = n745 & n867 ;
  assign n869 = n743 & n868 ;
  assign n870 = \n3077gat_pad  & n741 ;
  assign n871 = n739 & n870 ;
  assign n872 = ~n869 & ~n871 ;
  assign n873 = \n3065gat_pad  & \n3087gat_pad  ;
  assign n874 = n745 & n873 ;
  assign n875 = n743 & n874 ;
  assign n876 = \n3074gat_pad  & n741 ;
  assign n877 = n739 & n876 ;
  assign n878 = ~n875 & ~n877 ;
  assign n879 = \n3066gat_pad  & \n3087gat_pad  ;
  assign n880 = n745 & n879 ;
  assign n881 = n743 & n880 ;
  assign n882 = \n3075gat_pad  & n741 ;
  assign n883 = n739 & n882 ;
  assign n884 = ~n881 & ~n883 ;
  assign n885 = \n2203gat_reg/NET0131  & \n2207gat_reg/NET0131  ;
  assign n886 = ~n350 & ~n885 ;
  assign n887 = ~\n2562gat_reg/NET0131  & ~\n2640gat_reg/NET0131  ;
  assign n888 = \n2562gat_reg/NET0131  & \n2640gat_reg/NET0131  ;
  assign n889 = ~n887 & ~n888 ;
  assign n890 = \n2343gat_reg/NET0131  & ~\n2399gat_reg/NET0131  ;
  assign n891 = ~n351 & ~n890 ;
  assign n892 = n889 & n891 ;
  assign n893 = ~n889 & ~n891 ;
  assign n894 = ~n892 & ~n893 ;
  assign n895 = n886 & n894 ;
  assign n896 = ~n886 & ~n894 ;
  assign n897 = ~n895 & ~n896 ;
  assign n898 = \n2117gat_reg/NET0131  & ~\n2125gat_reg/NET0131  ;
  assign n899 = ~n725 & n898 ;
  assign n900 = n396 & n741 ;
  assign n901 = \n3087gat_pad  & ~\n3088gat_pad  ;
  assign n902 = n401 & n901 ;
  assign n903 = n406 & n902 ;
  assign n904 = ~n900 & ~n903 ;
  assign n905 = \n2319gat_reg/NET0131  & ~\n3099gat_pad  ;
  assign n906 = ~n357 & n850 ;
  assign n907 = n439 & n686 ;
  assign n908 = n511 & n907 ;
  assign n909 = \n2403gat_reg/NET0131  & n446 ;
  assign n910 = \n2061gat_reg/NET0131  & n456 ;
  assign n911 = n430 & n462 ;
  assign n912 = n910 & n911 ;
  assign n913 = n909 & n912 ;
  assign n914 = n459 & n907 ;
  assign n915 = n505 & n584 ;
  assign n916 = n687 & n915 ;
  assign n917 = n456 & n592 ;
  assign n918 = n687 & n917 ;
  assign n919 = \n1312gat_reg/NET0131  & n462 ;
  assign n920 = n910 & n919 ;
  assign n921 = \n1899gat_reg/NET0131  & ~\n2139gat_reg/NET0131  ;
  assign n922 = n910 & n921 ;
  assign n923 = n355 & n445 ;
  assign n924 = \n3066gat_pad  & \n3093gat_pad  ;
  assign n925 = \n3075gat_pad  & \n3095gat_pad  ;
  assign n926 = ~n924 & ~n925 ;
  assign n927 = \n3068gat_pad  & \n3093gat_pad  ;
  assign n928 = \n3077gat_pad  & \n3095gat_pad  ;
  assign n929 = ~n927 & ~n928 ;
  assign n930 = \n3067gat_pad  & \n3093gat_pad  ;
  assign n931 = \n3076gat_pad  & \n3095gat_pad  ;
  assign n932 = ~n930 & ~n931 ;
  assign n933 = ~\n271gat_reg/NET0131  & ~\n842gat_reg/NET0131  ;
  assign n934 = \n271gat_reg/NET0131  & \n842gat_reg/NET0131  ;
  assign n935 = ~n933 & ~n934 ;
  assign n936 = \n337gat_reg/NET0131  & ~\n341gat_reg/NET0131  ;
  assign n937 = ~\n337gat_reg/NET0131  & \n341gat_reg/NET0131  ;
  assign n938 = ~n936 & ~n937 ;
  assign n939 = ~\n160gat_reg/NET0131  & n938 ;
  assign n940 = ~n935 & n939 ;
  assign n941 = n613 & n940 ;
  assign n942 = \n160gat_reg/NET0131  & n938 ;
  assign n943 = n935 & n942 ;
  assign n944 = n613 & n943 ;
  assign n945 = ~n941 & ~n944 ;
  assign n946 = ~n935 & n942 ;
  assign n947 = ~n613 & n946 ;
  assign n948 = n935 & n939 ;
  assign n949 = ~n613 & n948 ;
  assign n950 = ~n947 & ~n949 ;
  assign n951 = n945 & n950 ;
  assign n952 = \n160gat_reg/NET0131  & ~n938 ;
  assign n953 = ~n935 & n952 ;
  assign n954 = n613 & n953 ;
  assign n955 = ~\n160gat_reg/NET0131  & ~n938 ;
  assign n956 = n935 & n955 ;
  assign n957 = n613 & n956 ;
  assign n958 = ~n954 & ~n957 ;
  assign n959 = ~n935 & n955 ;
  assign n960 = ~n613 & n959 ;
  assign n961 = n935 & n952 ;
  assign n962 = ~n613 & n961 ;
  assign n963 = ~n960 & ~n962 ;
  assign n964 = n958 & n963 ;
  assign n965 = n951 & n964 ;
  assign n966 = ~n371 & n932 ;
  assign n967 = ~n371 & n929 ;
  assign n968 = \n384gat_reg/NET0131  & ~n827 ;
  assign n969 = ~\n327gat_reg/NET0131  & ~\n384gat_reg/NET0131  ;
  assign n970 = n750 & n969 ;
  assign n971 = ~n968 & ~n970 ;
  assign n972 = n823 & n971 ;
  assign n973 = \n3078gat_pad  & n741 ;
  assign n974 = n739 & n973 ;
  assign n975 = \n3069gat_pad  & \n3087gat_pad  ;
  assign n976 = n745 & n975 ;
  assign n977 = n743 & n976 ;
  assign n978 = ~n974 & ~n977 ;
  assign n979 = ~n972 & n978 ;
  assign n980 = n515 & n583 ;
  assign n981 = n445 & n722 ;
  assign n982 = \n327gat_reg/NET0131  & ~\n331gat_reg/NET0131  ;
  assign n983 = ~\n388gat_reg/NET0131  & ~n982 ;
  assign n984 = \n463gat_reg/NET0131  & ~n983 ;
  assign n985 = n981 & n984 ;
  assign n986 = n981 & ~n983 ;
  assign n987 = ~\n463gat_reg/NET0131  & ~n986 ;
  assign n988 = ~n985 & ~n987 ;
  assign n989 = n823 & ~n988 ;
  assign n990 = \n3082gat_pad  & n741 ;
  assign n991 = n739 & n990 ;
  assign n992 = \n3073gat_pad  & \n3087gat_pad  ;
  assign n993 = n745 & n992 ;
  assign n994 = n743 & n993 ;
  assign n995 = ~n991 & ~n994 ;
  assign n996 = ~n989 & n995 ;
  assign n997 = ~n371 & n926 ;
  assign n998 = \n388gat_reg/NET0131  & ~n981 ;
  assign n999 = ~n736 & ~n998 ;
  assign n1000 = n823 & n999 ;
  assign n1001 = \n3081gat_pad  & n741 ;
  assign n1002 = n739 & n1001 ;
  assign n1003 = \n3072gat_pad  & \n3087gat_pad  ;
  assign n1004 = n745 & n1003 ;
  assign n1005 = n743 & n1004 ;
  assign n1006 = ~n1002 & ~n1005 ;
  assign n1007 = ~n1000 & n1006 ;
  assign n1008 = ~n470 & ~n471 ;
  assign n1009 = \n1312gat_reg/NET0131  & ~\n2169gat_reg/NET0131  ;
  assign n1010 = \n3100gat_pad  & n1009 ;
  assign n1011 = n476 & n1009 ;
  assign n1012 = n475 & n1011 ;
  assign n1013 = ~n1010 & ~n1012 ;
  assign n1014 = ~n470 & ~n1013 ;
  assign n1015 = \n1197gat_reg/NET0131  & n286 ;
  assign n1016 = ~n283 & n1015 ;
  assign n1017 = ~n280 & n1016 ;
  assign n1018 = n283 & n1015 ;
  assign n1019 = n280 & n1018 ;
  assign n1020 = ~n1017 & ~n1019 ;
  assign n1021 = \n1197gat_reg/NET0131  & ~n286 ;
  assign n1022 = n283 & n1021 ;
  assign n1023 = ~n280 & n1022 ;
  assign n1024 = ~n283 & n1021 ;
  assign n1025 = n280 & n1024 ;
  assign n1026 = ~n1023 & ~n1025 ;
  assign n1027 = n1020 & n1026 ;
  assign n1028 = ~\n1197gat_reg/NET0131  & ~n286 ;
  assign n1029 = ~n283 & n1028 ;
  assign n1030 = ~n280 & n1029 ;
  assign n1031 = n283 & n1028 ;
  assign n1032 = n280 & n1031 ;
  assign n1033 = ~n1030 & ~n1032 ;
  assign n1034 = ~\n1197gat_reg/NET0131  & n286 ;
  assign n1035 = n283 & n1034 ;
  assign n1036 = ~n280 & n1035 ;
  assign n1037 = ~n283 & n1034 ;
  assign n1038 = n280 & n1037 ;
  assign n1039 = ~n1036 & ~n1038 ;
  assign n1040 = n1033 & n1039 ;
  assign n1041 = n1027 & n1040 ;
  assign n1042 = ~\n3085gat_pad  & \n3086gat_pad  ;
  assign n1043 = n402 & n1042 ;
  assign n1044 = n401 & n1043 ;
  assign n1045 = ~n404 & n1044 ;
  assign n1046 = ~\n3086gat_pad  & ~n213 ;
  assign n1047 = n396 & n1046 ;
  assign n1048 = ~n1045 & ~n1047 ;
  assign n1049 = n598 & n1048 ;
  assign n1050 = n398 & n739 ;
  assign n1051 = n403 & n745 ;
  assign n1052 = ~n588 & ~n1051 ;
  assign n1053 = ~n1050 & n1052 ;
  assign n1054 = \n1771gat_reg/NET0131  & \n1775gat_reg/NET0131  ;
  assign n1055 = \n1871gat_reg/NET0131  & ~n1054 ;
  assign n1056 = \n1035gat_reg/NET0131  & ~n659 ;
  assign n1057 = \n1072gat_reg/NET0131  & ~n651 ;
  assign n1058 = ~n649 & n1057 ;
  assign n1059 = \n1121gat_reg/NET0131  & \n2403gat_reg/NET0131  ;
  assign n1060 = ~n433 & n1059 ;
  assign n1061 = \n1121gat_reg/NET0131  & ~\n2403gat_reg/NET0131  ;
  assign n1062 = n433 & n1061 ;
  assign n1063 = ~n1060 & ~n1062 ;
  assign n1064 = \n931gat_reg/NET0131  & n446 ;
  assign n1065 = \n1135gat_reg/NET0131  & \n2135gat_reg/NET0131  ;
  assign n1066 = ~n518 & n1065 ;
  assign n1067 = \n1135gat_reg/NET0131  & ~\n2135gat_reg/NET0131  ;
  assign n1068 = n518 & n1067 ;
  assign n1069 = ~n1066 & ~n1068 ;
  assign n1070 = \n1282gat_reg/NET0131  & n580 ;
  assign n1071 = n283 & n286 ;
  assign n1072 = ~n280 & n1071 ;
  assign n1073 = ~n283 & n286 ;
  assign n1074 = n280 & n1073 ;
  assign n1075 = ~n1072 & ~n1074 ;
  assign n1076 = ~n280 & n297 ;
  assign n1077 = n280 & n294 ;
  assign n1078 = ~n1076 & ~n1077 ;
  assign n1079 = n1075 & n1078 ;
  assign n1080 = ~\n659gat_reg/NET0131  & ~n222 ;
  assign n1081 = n219 & n1080 ;
  assign n1082 = ~\n1068gat_reg/NET0131  & n222 ;
  assign n1083 = n237 & n1082 ;
  assign n1084 = ~n1081 & ~n1083 ;
  assign n1085 = ~\n680gat_reg/NET0131  & ~n222 ;
  assign n1086 = n304 & n1085 ;
  assign n1087 = ~\n271gat_reg/NET0131  & ~n222 ;
  assign n1088 = n237 & n1087 ;
  assign n1089 = ~n1086 & ~n1088 ;
  assign n1090 = n1084 & n1089 ;
  assign n1091 = n261 & ~n1090 ;
  assign n1092 = n813 & ~n1091 ;
  assign n1093 = ~\n580gat_reg/NET0131  & ~n222 ;
  assign n1094 = n304 & n1093 ;
  assign n1095 = ~\n337gat_reg/NET0131  & ~n222 ;
  assign n1096 = n237 & n1095 ;
  assign n1097 = ~n1094 & ~n1096 ;
  assign n1098 = ~\n861gat_reg/NET0131  & n222 ;
  assign n1099 = n237 & n1098 ;
  assign n1100 = ~\n777gat_reg/NET0131  & ~n222 ;
  assign n1101 = n219 & n1100 ;
  assign n1102 = ~n1099 & ~n1101 ;
  assign n1103 = n1097 & n1102 ;
  assign n1104 = n261 & ~n1103 ;
  assign n1105 = n965 & ~n1104 ;
  assign n1106 = ~\n816gat_reg/NET0131  & ~n222 ;
  assign n1107 = n304 & n1106 ;
  assign n1108 = ~\n160gat_reg/NET0131  & ~n222 ;
  assign n1109 = n237 & n1108 ;
  assign n1110 = ~n1107 & ~n1109 ;
  assign n1111 = ~\n957gat_reg/NET0131  & n222 ;
  assign n1112 = n237 & n1111 ;
  assign n1113 = ~\n553gat_reg/NET0131  & ~n222 ;
  assign n1114 = n219 & n1113 ;
  assign n1115 = ~n1112 & ~n1114 ;
  assign n1116 = n1110 & n1115 ;
  assign n1117 = n261 & ~n1116 ;
  assign n1118 = n721 & ~n1117 ;
  assign n1119 = ~\n322gat_reg/NET0131  & ~n222 ;
  assign n1120 = n219 & n1119 ;
  assign n1121 = ~\n865gat_reg/NET0131  & n222 ;
  assign n1122 = n237 & n1121 ;
  assign n1123 = ~n1120 & ~n1122 ;
  assign n1124 = ~\n584gat_reg/NET0131  & ~n222 ;
  assign n1125 = n304 & n1124 ;
  assign n1126 = ~\n341gat_reg/NET0131  & ~n222 ;
  assign n1127 = n237 & n1126 ;
  assign n1128 = ~n1125 & ~n1127 ;
  assign n1129 = n1123 & n1128 ;
  assign n1130 = n261 & ~n1129 ;
  assign n1131 = n965 & ~n1130 ;
  assign n1132 = ~\n314gat_reg/NET0131  & ~n222 ;
  assign n1133 = n219 & n1132 ;
  assign n1134 = ~\n1148gat_reg/NET0131  & n222 ;
  assign n1135 = n237 & n1134 ;
  assign n1136 = ~n1133 & ~n1135 ;
  assign n1137 = ~\n398gat_reg/NET0131  & ~n222 ;
  assign n1138 = n237 & n1137 ;
  assign n1139 = ~\n699gat_reg/NET0131  & ~n222 ;
  assign n1140 = n304 & n1139 ;
  assign n1141 = ~n1138 & ~n1140 ;
  assign n1142 = n1136 & n1141 ;
  assign n1143 = n261 & ~n1142 ;
  assign n1144 = n570 & ~n1143 ;
  assign n1145 = ~\n318gat_reg/NET0131  & ~n222 ;
  assign n1146 = n219 & n1145 ;
  assign n1147 = ~\n1080gat_reg/NET0131  & n222 ;
  assign n1148 = n237 & n1147 ;
  assign n1149 = ~n1146 & ~n1148 ;
  assign n1150 = ~\n402gat_reg/NET0131  & ~n222 ;
  assign n1151 = n237 & n1150 ;
  assign n1152 = ~\n684gat_reg/NET0131  & ~n222 ;
  assign n1153 = n304 & n1152 ;
  assign n1154 = ~n1151 & ~n1153 ;
  assign n1155 = n1149 & n1154 ;
  assign n1156 = n261 & ~n1155 ;
  assign n1157 = n645 & ~n1156 ;
  assign n1158 = ~\n561gat_reg/NET0131  & ~n222 ;
  assign n1159 = n219 & n1158 ;
  assign n1160 = ~\n1294gat_reg/NET0131  & n222 ;
  assign n1161 = n237 & n1160 ;
  assign n1162 = ~n1159 & ~n1161 ;
  assign n1163 = ~\n824gat_reg/NET0131  & ~n222 ;
  assign n1164 = n304 & n1163 ;
  assign n1165 = ~\n846gat_reg/NET0131  & ~n222 ;
  assign n1166 = n237 & n1165 ;
  assign n1167 = ~n1164 & ~n1166 ;
  assign n1168 = n1162 & n1167 ;
  assign n1169 = n261 & ~n1168 ;
  assign n1170 = n335 & ~n1169 ;
  assign n1171 = ~\n919gat_reg/NET0131  & ~n215 ;
  assign n1172 = ~n222 & ~n1171 ;
  assign n1173 = ~n218 & ~n243 ;
  assign n1174 = ~n1172 & n1173 ;
  assign n1175 = ~\n366gat_reg/NET0131  & ~n222 ;
  assign n1176 = n219 & n1175 ;
  assign n1177 = ~\n883gat_reg/NET0131  & ~n222 ;
  assign n1178 = n304 & n1177 ;
  assign n1179 = ~n1176 & ~n1178 ;
  assign n1180 = ~n1174 & n1179 ;
  assign n1181 = n261 & ~n1180 ;
  assign n1182 = ~n1041 & ~n1181 ;
  assign n1183 = ~n261 & n579 ;
  assign n1184 = n246 & n579 ;
  assign n1185 = n234 & n1184 ;
  assign n1186 = ~n1183 & ~n1185 ;
  assign n1187 = ~n257 & ~n1090 ;
  assign n1188 = ~\n271gat_reg/NET0131  & n222 ;
  assign n1189 = n237 & n1188 ;
  assign n1190 = ~\n1035gat_reg/NET0131  & ~n222 ;
  assign n1191 = n219 & n1190 ;
  assign n1192 = ~\n834gat_reg/NET0131  & ~n222 ;
  assign n1193 = n304 & n1192 ;
  assign n1194 = ~n1191 & ~n1193 ;
  assign n1195 = ~n1189 & n1194 ;
  assign n1196 = ~n266 & ~n1195 ;
  assign n1197 = ~n1187 & ~n1196 ;
  assign n1198 = ~n257 & ~n1103 ;
  assign n1199 = ~\n1072gat_reg/NET0131  & ~n222 ;
  assign n1200 = n219 & n1199 ;
  assign n1201 = ~\n337gat_reg/NET0131  & n222 ;
  assign n1202 = n237 & n1201 ;
  assign n1203 = ~\n838gat_reg/NET0131  & ~n222 ;
  assign n1204 = n304 & n1203 ;
  assign n1205 = ~n1202 & ~n1204 ;
  assign n1206 = ~n1200 & n1205 ;
  assign n1207 = ~n266 & ~n1206 ;
  assign n1208 = ~n1198 & ~n1207 ;
  assign n1209 = ~n257 & ~n1116 ;
  assign n1210 = ~\n1121gat_reg/NET0131  & ~n222 ;
  assign n1211 = n219 & n1210 ;
  assign n1212 = ~\n160gat_reg/NET0131  & n222 ;
  assign n1213 = n237 & n1212 ;
  assign n1214 = ~\n707gat_reg/NET0131  & ~n222 ;
  assign n1215 = n304 & n1214 ;
  assign n1216 = ~n1213 & ~n1215 ;
  assign n1217 = ~n1211 & n1216 ;
  assign n1218 = ~n266 & ~n1217 ;
  assign n1219 = ~n1209 & ~n1218 ;
  assign n1220 = ~n257 & ~n1129 ;
  assign n1221 = ~\n931gat_reg/NET0131  & ~n222 ;
  assign n1222 = n219 & n1221 ;
  assign n1223 = ~\n341gat_reg/NET0131  & n222 ;
  assign n1224 = n237 & n1223 ;
  assign n1225 = ~\n614gat_reg/NET0131  & ~n222 ;
  assign n1226 = n304 & n1225 ;
  assign n1227 = ~n1224 & ~n1226 ;
  assign n1228 = ~n1222 & n1227 ;
  assign n1229 = ~n266 & ~n1228 ;
  assign n1230 = ~n1220 & ~n1229 ;
  assign n1231 = ~\n1045gat_reg/NET0131  & ~n222 ;
  assign n1232 = n219 & n1231 ;
  assign n1233 = n304 & n1137 ;
  assign n1234 = ~\n398gat_reg/NET0131  & n222 ;
  assign n1235 = n237 & n1234 ;
  assign n1236 = ~n1233 & ~n1235 ;
  assign n1237 = ~n1232 & n1236 ;
  assign n1238 = ~n266 & ~n1237 ;
  assign n1239 = ~n257 & ~n1142 ;
  assign n1240 = ~n1238 & ~n1239 ;
  assign n1241 = ~\n1135gat_reg/NET0131  & ~n222 ;
  assign n1242 = n219 & n1241 ;
  assign n1243 = n304 & n1150 ;
  assign n1244 = ~\n402gat_reg/NET0131  & n222 ;
  assign n1245 = n237 & n1244 ;
  assign n1246 = ~n1243 & ~n1245 ;
  assign n1247 = ~n1242 & n1246 ;
  assign n1248 = ~n266 & ~n1247 ;
  assign n1249 = ~n257 & ~n1155 ;
  assign n1250 = ~n1248 & ~n1249 ;
  assign n1251 = ~\n1282gat_reg/NET0131  & ~n222 ;
  assign n1252 = n219 & n1251 ;
  assign n1253 = n304 & n1165 ;
  assign n1254 = ~\n846gat_reg/NET0131  & n222 ;
  assign n1255 = n237 & n1254 ;
  assign n1256 = ~n1253 & ~n1255 ;
  assign n1257 = ~n1252 & n1256 ;
  assign n1258 = ~n266 & ~n1257 ;
  assign n1259 = ~n257 & ~n1168 ;
  assign n1260 = ~n1258 & ~n1259 ;
  assign n1261 = ~\n1226gat_reg/NET0131  & ~n222 ;
  assign n1262 = n219 & n1261 ;
  assign n1263 = ~\n919gat_reg/NET0131  & ~n222 ;
  assign n1264 = n304 & n1263 ;
  assign n1265 = ~\n919gat_reg/NET0131  & n222 ;
  assign n1266 = n237 & n1265 ;
  assign n1267 = ~n1264 & ~n1266 ;
  assign n1268 = ~n1262 & n1267 ;
  assign n1269 = ~n266 & ~n1268 ;
  assign n1270 = ~n257 & ~n1180 ;
  assign n1271 = ~n1269 & ~n1270 ;
  assign n1272 = ~\n2562gat_reg/NET0131  & n364 ;
  assign n1273 = n350 & n1272 ;
  assign n1274 = n200 & n1273 ;
  assign n1275 = n527 & n1274 ;
  assign n1276 = ~\n1462gat_reg/NET0131  & ~n455 ;
  assign n1277 = \n1394gat_reg/NET0131  & ~n468 ;
  assign n1278 = n1276 & n1277 ;
  assign n1279 = ~\n1508gat_reg/NET0131  & n1278 ;
  assign n1280 = ~\n1340gat_reg/NET0131  & ~n455 ;
  assign n1281 = ~n353 & n1280 ;
  assign n1282 = ~\n1508gat_reg/NET0131  & n1281 ;
  assign n1283 = ~n695 & n1282 ;
  assign n1284 = ~n1279 & ~n1283 ;
  assign n1285 = ~\n1394gat_reg/NET0131  & ~n694 ;
  assign n1286 = ~\n1596gat_reg/NET0131  & ~n1285 ;
  assign n1287 = n455 & ~n1286 ;
  assign n1288 = \n1462gat_reg/NET0131  & ~\n1678gat_reg/NET0131  ;
  assign n1289 = ~\n1678gat_reg/NET0131  & \n2102gat_reg/NET0131  ;
  assign n1290 = ~n454 & n1289 ;
  assign n1291 = ~n1288 & ~n1290 ;
  assign n1292 = ~n1287 & ~n1291 ;
  assign n1293 = ~\n1394gat_reg/NET0131  & \n2102gat_reg/NET0131  ;
  assign n1294 = ~n454 & n1293 ;
  assign n1295 = ~\n1525gat_reg/NET0131  & n1294 ;
  assign n1296 = ~n363 & n1295 ;
  assign n1297 = \n1829gat_reg/NET0131  & \n3097gat_pad  ;
  assign n1298 = n471 & n1297 ;
  assign n1299 = \n1821gat_reg/NET0131  & ~n1298 ;
  assign n1300 = ~\n1775gat_reg/NET0131  & \n1871gat_reg/NET0131  ;
  assign n1301 = ~\n3098gat_pad  & n1300 ;
  assign n1302 = ~n1299 & n1301 ;
  assign n1303 = ~\n1588gat_reg/NET0131  & \n2102gat_reg/NET0131  ;
  assign n1304 = ~n454 & n1303 ;
  assign n1305 = \n1596gat_reg/NET0131  & n1304 ;
  assign n1306 = ~n1302 & ~n1305 ;
  assign n1307 = ~n1296 & n1306 ;
  assign n1308 = ~n1292 & n1307 ;
  assign n1309 = n1284 & n1308 ;
  assign n1310 = n468 & ~n694 ;
  assign n1311 = ~\n1748gat_reg/NET0131  & ~n1310 ;
  assign n1312 = \n1336gat_reg/NET0131  & ~\n1748gat_reg/NET0131  ;
  assign n1313 = ~n363 & n1312 ;
  assign n1314 = ~n1311 & ~n1313 ;
  assign n1315 = n455 & ~n1314 ;
  assign n1316 = ~\n1675gat_reg/NET0131  & n1294 ;
  assign n1317 = ~n363 & n1316 ;
  assign n1318 = n455 & ~n1317 ;
  assign n1319 = ~\n1456gat_reg/NET0131  & ~n468 ;
  assign n1320 = ~\n1340gat_reg/NET0131  & ~\n1456gat_reg/NET0131  ;
  assign n1321 = ~n1319 & ~n1320 ;
  assign n1322 = ~n694 & ~n1319 ;
  assign n1323 = n363 & n1322 ;
  assign n1324 = ~n1321 & ~n1323 ;
  assign n1325 = \n1340gat_reg/NET0131  & ~\n1807gat_reg/NET0131  ;
  assign n1326 = ~n1317 & ~n1325 ;
  assign n1327 = ~n1324 & n1326 ;
  assign n1328 = ~n1318 & ~n1327 ;
  assign n1329 = ~n1315 & ~n1328 ;
  assign n1330 = \n1678gat_reg/NET0131  & \n2102gat_reg/NET0131  ;
  assign n1331 = ~n454 & n1330 ;
  assign n1332 = \n1508gat_reg/NET0131  & ~n455 ;
  assign n1333 = ~\n1394gat_reg/NET0131  & ~n468 ;
  assign n1334 = ~n1332 & n1333 ;
  assign n1335 = ~n1331 & n1334 ;
  assign n1336 = \n1871gat_reg/NET0131  & ~\n2592gat_reg/NET0131  ;
  assign n1337 = ~\n673gat_reg/NET0131  & n1336 ;
  assign n1338 = ~\n1389gat_reg/NET0131  & ~n1337 ;
  assign n1339 = ~n1335 & n1338 ;
  assign n1340 = ~n850 & n1272 ;
  assign n1341 = \n2084gat_reg/NET0131  & ~n849 ;
  assign n1342 = n528 & ~n1341 ;
  assign n1343 = ~n1340 & ~n1342 ;
  assign n1344 = ~\n1068gat_reg/NET0131  & \n2562gat_reg/NET0131  ;
  assign n1345 = n351 & n1344 ;
  assign n1346 = ~\n2562gat_reg/NET0131  & ~\n865gat_reg/NET0131  ;
  assign n1347 = n890 & n1346 ;
  assign n1348 = ~n1345 & ~n1347 ;
  assign n1349 = \n2562gat_reg/NET0131  & ~\n957gat_reg/NET0131  ;
  assign n1350 = n890 & n1349 ;
  assign n1351 = ~\n2562gat_reg/NET0131  & ~\n861gat_reg/NET0131  ;
  assign n1352 = n351 & n1351 ;
  assign n1353 = ~n1350 & ~n1352 ;
  assign n1354 = n1348 & n1353 ;
  assign n1355 = ~n468 & ~n1354 ;
  assign n1356 = \n2562gat_reg/NET0131  & ~\n816gat_reg/NET0131  ;
  assign n1357 = n890 & n1356 ;
  assign n1358 = \n2562gat_reg/NET0131  & ~\n680gat_reg/NET0131  ;
  assign n1359 = n351 & n1358 ;
  assign n1360 = ~n1357 & ~n1359 ;
  assign n1361 = ~\n2562gat_reg/NET0131  & ~\n580gat_reg/NET0131  ;
  assign n1362 = n351 & n1361 ;
  assign n1363 = ~\n2562gat_reg/NET0131  & ~\n584gat_reg/NET0131  ;
  assign n1364 = n890 & n1363 ;
  assign n1365 = ~n1362 & ~n1364 ;
  assign n1366 = n1360 & n1365 ;
  assign n1367 = n468 & ~n1366 ;
  assign n1368 = ~n1355 & ~n1367 ;
  assign n1369 = n1343 & n1368 ;
  assign n1370 = n885 & ~n1369 ;
  assign n1371 = \n1880gat_reg/NET0131  & \n699gat_reg/NET0131  ;
  assign n1372 = n467 & n1371 ;
  assign n1373 = \n1148gat_reg/NET0131  & ~n468 ;
  assign n1374 = ~\n2343gat_reg/NET0131  & ~\n2399gat_reg/NET0131  ;
  assign n1375 = \n2562gat_reg/NET0131  & n885 ;
  assign n1376 = n1374 & n1375 ;
  assign n1377 = ~n1373 & n1376 ;
  assign n1378 = ~n1372 & n1377 ;
  assign n1379 = \n1880gat_reg/NET0131  & \n684gat_reg/NET0131  ;
  assign n1380 = n467 & n1379 ;
  assign n1381 = \n1080gat_reg/NET0131  & ~n468 ;
  assign n1382 = ~\n2562gat_reg/NET0131  & n885 ;
  assign n1383 = n1374 & n1382 ;
  assign n1384 = ~n1381 & n1383 ;
  assign n1385 = ~n1380 & n1384 ;
  assign n1386 = ~n1378 & ~n1385 ;
  assign n1387 = ~n1370 & n1386 ;
  assign n1388 = ~n1335 & ~n1337 ;
  assign n1389 = ~\n160gat_reg/NET0131  & \n2562gat_reg/NET0131  ;
  assign n1390 = n890 & n1389 ;
  assign n1391 = \n2562gat_reg/NET0131  & ~\n271gat_reg/NET0131  ;
  assign n1392 = n351 & n1391 ;
  assign n1393 = ~n1390 & ~n1392 ;
  assign n1394 = ~\n2562gat_reg/NET0131  & ~\n337gat_reg/NET0131  ;
  assign n1395 = n351 & n1394 ;
  assign n1396 = ~n468 & ~n1395 ;
  assign n1397 = ~\n2562gat_reg/NET0131  & ~\n341gat_reg/NET0131  ;
  assign n1398 = n890 & n1397 ;
  assign n1399 = n1396 & ~n1398 ;
  assign n1400 = n1393 & n1399 ;
  assign n1401 = ~\n2562gat_reg/NET0131  & ~\n614gat_reg/NET0131  ;
  assign n1402 = n890 & n1401 ;
  assign n1403 = n468 & ~n1402 ;
  assign n1404 = \n2562gat_reg/NET0131  & ~\n707gat_reg/NET0131  ;
  assign n1405 = n890 & n1404 ;
  assign n1406 = ~\n2562gat_reg/NET0131  & ~\n838gat_reg/NET0131  ;
  assign n1407 = n351 & n1406 ;
  assign n1408 = \n2562gat_reg/NET0131  & ~\n834gat_reg/NET0131  ;
  assign n1409 = n351 & n1408 ;
  assign n1410 = ~n1407 & ~n1409 ;
  assign n1411 = ~n1405 & n1410 ;
  assign n1412 = n1403 & n1411 ;
  assign n1413 = ~n1400 & ~n1412 ;
  assign n1414 = \n1294gat_reg/NET0131  & ~n468 ;
  assign n1415 = \n1880gat_reg/NET0131  & \n824gat_reg/NET0131  ;
  assign n1416 = n467 & n1415 ;
  assign n1417 = n528 & ~n1416 ;
  assign n1418 = ~n1414 & n1417 ;
  assign n1419 = \n673gat_reg/NET0131  & ~n468 ;
  assign n1420 = \n1880gat_reg/NET0131  & \n883gat_reg/NET0131  ;
  assign n1421 = n467 & n1420 ;
  assign n1422 = n1272 & ~n1421 ;
  assign n1423 = ~n1419 & n1422 ;
  assign n1424 = ~n1418 & ~n1423 ;
  assign n1425 = ~n1413 & n1424 ;
  assign n1426 = ~\n2203gat_reg/NET0131  & \n2207gat_reg/NET0131  ;
  assign n1427 = ~n1425 & n1426 ;
  assign n1428 = n1388 & ~n1427 ;
  assign n1429 = n1387 & n1428 ;
  assign n1430 = ~n1339 & ~n1429 ;
  assign n1431 = ~\n919gat_reg/NET0131  & ~n229 ;
  assign n1432 = ~n212 & n1431 ;
  assign n1433 = ~\n659gat_reg/NET0131  & ~\n919gat_reg/NET0131  ;
  assign n1434 = ~n226 & n1433 ;
  assign n1435 = \n659gat_reg/NET0131  & ~\n919gat_reg/NET0131  ;
  assign n1436 = n226 & n1435 ;
  assign n1437 = ~n1434 & ~n1436 ;
  assign n1438 = n212 & ~n1437 ;
  assign n1439 = ~n1432 & ~n1438 ;
  assign n1440 = n350 & n528 ;
  assign n1441 = \n919gat_reg/NET0131  & ~n229 ;
  assign n1442 = n212 & n1441 ;
  assign n1443 = ~n203 & n694 ;
  assign n1444 = n209 & n1443 ;
  assign n1445 = ~\n659gat_reg/NET0131  & \n919gat_reg/NET0131  ;
  assign n1446 = ~n226 & n1445 ;
  assign n1447 = \n659gat_reg/NET0131  & \n919gat_reg/NET0131  ;
  assign n1448 = n226 & n1447 ;
  assign n1449 = ~n1446 & ~n1448 ;
  assign n1450 = n694 & n1449 ;
  assign n1451 = n203 & n694 ;
  assign n1452 = ~n209 & n1451 ;
  assign n1453 = ~n1450 & ~n1452 ;
  assign n1454 = ~n1444 & n1453 ;
  assign n1455 = ~n1442 & ~n1454 ;
  assign n1456 = n1440 & n1455 ;
  assign n1457 = n1439 & n1456 ;
  assign n1458 = \n2562gat_reg/NET0131  & ~\n561gat_reg/NET0131  ;
  assign n1459 = n1374 & n1458 ;
  assign n1460 = \n2562gat_reg/NET0131  & ~\n659gat_reg/NET0131  ;
  assign n1461 = n364 & n1460 ;
  assign n1462 = ~n1459 & ~n1461 ;
  assign n1463 = ~\n2562gat_reg/NET0131  & ~\n318gat_reg/NET0131  ;
  assign n1464 = n890 & n1463 ;
  assign n1465 = ~\n2562gat_reg/NET0131  & ~\n777gat_reg/NET0131  ;
  assign n1466 = n364 & n1465 ;
  assign n1467 = ~n1464 & ~n1466 ;
  assign n1468 = n1462 & n1467 ;
  assign n1469 = ~\n2562gat_reg/NET0131  & ~\n322gat_reg/NET0131  ;
  assign n1470 = n351 & n1469 ;
  assign n1471 = \n2562gat_reg/NET0131  & ~\n314gat_reg/NET0131  ;
  assign n1472 = n890 & n1471 ;
  assign n1473 = ~n1470 & ~n1472 ;
  assign n1474 = \n2562gat_reg/NET0131  & ~\n553gat_reg/NET0131  ;
  assign n1475 = n351 & n1474 ;
  assign n1476 = ~\n2562gat_reg/NET0131  & ~\n366gat_reg/NET0131  ;
  assign n1477 = n1374 & n1476 ;
  assign n1478 = ~n1475 & ~n1477 ;
  assign n1479 = n1473 & n1478 ;
  assign n1480 = n1468 & n1479 ;
  assign n1481 = n366 & n694 ;
  assign n1482 = ~n1480 & n1481 ;
  assign n1483 = ~n497 & ~n1482 ;
  assign n1484 = ~n1457 & n1483 ;
  assign n1485 = ~n1430 & n1484 ;
  assign n1486 = n897 & ~n1482 ;
  assign n1487 = ~n1457 & n1486 ;
  assign n1488 = ~n1430 & n1487 ;
  assign n1489 = \n2514gat_reg/NET0131  & n1054 ;
  assign n1490 = ~n694 & ~n1489 ;
  assign n1491 = n363 & n1490 ;
  assign n1492 = \n1871gat_reg/NET0131  & \n2514gat_reg/NET0131  ;
  assign n1493 = n1054 & n1492 ;
  assign n1494 = \n2169gat_reg/NET0131  & \n2176gat_reg/NET0131  ;
  assign n1495 = \n2033gat_reg/NET0131  & n1494 ;
  assign n1496 = \n2110gat_reg/NET0131  & n537 ;
  assign n1497 = n1495 & n1496 ;
  assign n1498 = ~n1493 & n1497 ;
  assign n1499 = ~\n2454gat_reg/NET0131  & ~\n337gat_reg/NET0131  ;
  assign n1500 = n594 & ~n1499 ;
  assign n1501 = n738 & n1046 ;
  assign n1502 = n584 & ~n1044 ;
  assign n1503 = ~n1501 & n1502 ;
  assign \_al_n0  = 1'b0 ;
  assign \g17_dup/_0_  = n200 ;
  assign \g6952/_2_  = ~n310 ;
  assign \g6953/_2_  = ~n316 ;
  assign \g6961/_0_  = n335 ;
  assign \g7076/_0_  = ~n372 ;
  assign \g7077/_0_  = ~n376 ;
  assign \g7079/_0_  = ~n380 ;
  assign \g7081/_0_  = ~n384 ;
  assign \g7082/_0_  = ~n388 ;
  assign \g7083/_0_  = ~n392 ;
  assign \g7146/_0_  = ~n410 ;
  assign \g7147/_0_  = ~n412 ;
  assign \g7148/_0_  = ~n414 ;
  assign \g7149/_0_  = ~n416 ;
  assign \g7150/_0_  = ~n418 ;
  assign \g7151/_0_  = ~n420 ;
  assign \g7152/_0_  = ~n422 ;
  assign \g7153/_0_  = ~n424 ;
  assign \g7154/_0_  = ~n426 ;
  assign \g7156/_2_  = n481 ;
  assign \g7161/_2_  = n484 ;
  assign \g7165/_2_  = ~n497 ;
  assign \g7174/_0_  = n498 ;
  assign \g7180/_00_  = n525 ;
  assign \g7182/_3_  = n530 ;
  assign \g7191/_0_  = n540 ;
  assign \g7204/_0_  = ~n546 ;
  assign \g7209/_3_  = n570 ;
  assign \g7220/_0_  = ~\n2543gat_reg/NET0131  ;
  assign \g7229/_0_  = n579 ;
  assign \g7233/_0_  = n582 ;
  assign \g7234/_0_  = n586 ;
  assign \g7235/_0_  = n590 ;
  assign \g7236/_0_  = n596 ;
  assign \g7237/_0_  = n600 ;
  assign \g7238/_0_  = ~n607 ;
  assign \g7241/_3_  = n645 ;
  assign \g7264/_0_  = n653 ;
  assign \g7265/_0_  = n660 ;
  assign \g7266/_0_  = ~n671 ;
  assign \g7267/_0_  = n676 ;
  assign \g7268/_0_  = n684 ;
  assign \g7301/_0_  = n688 ;
  assign \g7326/_3_  = n692 ;
  assign \g7350/_2_  = ~n695 ;
  assign \g7352/_0_  = ~\n838gat_reg/NET0131  ;
  assign \g7356/_0_  = n697 ;
  assign \g7359/_0_  = ~n531 ;
  assign \g7389/_3_  = n721 ;
  assign \g7417/_0_  = n729 ;
  assign \g7418/_0_  = n731 ;
  assign \g7419/_0_  = n733 ;
  assign \g7444/_0_  = ~n760 ;
  assign \g7445/_0_  = ~n778 ;
  assign \g7449/_3_  = ~n792 ;
  assign \g7451/_3_  = n813 ;
  assign \g7454/_0_  = ~\n707gat_reg/NET0131  ;
  assign \g7467/_3_  = ~n822 ;
  assign \g7476/_0_  = ~\n614gat_reg/NET0131  ;
  assign \g7480/_0_  = ~n836 ;
  assign \g7494/_0_  = ~n847 ;
  assign \g7509/_0_  = ~\n2176gat_reg/NET0131  ;
  assign \g7514/_0_  = ~n852 ;
  assign \g7517/_3_  = ~n860 ;
  assign \g7524/_0_  = ~\n2095gat_reg/NET0131  ;
  assign \g7558/_0_  = ~n866 ;
  assign \g7560/_0_  = ~n872 ;
  assign \g7561/_0_  = ~n878 ;
  assign \g7563/_0_  = ~n884 ;
  assign \g7567/_0_  = n897 ;
  assign \g7572/_0_  = ~\n1821gat_reg/NET0131  ;
  assign \g7579/_0_  = n899 ;
  assign \g7605/_0_  = ~n904 ;
  assign \g7625/_0_  = n905 ;
  assign \g7627/_0_  = ~n906 ;
  assign \g7671/_0_  = n908 ;
  assign \g7675/_0_  = n913 ;
  assign \g7689/_0_  = n914 ;
  assign \g7697/_0_  = n916 ;
  assign \g7743/_1_  = n723 ;
  assign \g7764/_1_  = n732 ;
  assign \g7769/_0_  = n918 ;
  assign \g7771/_2_  = n915 ;
  assign \g7779/_0_  = n920 ;
  assign \g7852/_0_  = n922 ;
  assign \g7873/_0_  = n923 ;
  assign \g7884/_3_  = n506 ;
  assign \g7889/_0_  = ~\n2110gat_reg/NET0131  ;
  assign \g7902/_1_  = n730 ;
  assign \g7992/_3_  = ~n926 ;
  assign \g7994/_3_  = ~n375 ;
  assign \g7996/_3_  = ~n383 ;
  assign \g7998/_3_  = ~n929 ;
  assign \g8000/_3_  = ~n932 ;
  assign \g8002/_3_  = ~n338 ;
  assign \g8004/_3_  = ~n391 ;
  assign \g8006/_3_  = ~n387 ;
  assign \g8008/_3_  = ~n379 ;
  assign \g8150/_0_  = ~\n2626gat_reg/NET0131  ;
  assign \g8151/_0_  = ~\n2495gat_reg/NET0131  ;
  assign \g8157/_0_  = ~\n2037gat_reg/NET0131  ;
  assign \g8163/_0_  = ~\n830gat_reg/NET0131  ;
  assign \g8172/_0_  = ~\n2490gat_reg/NET0131  ;
  assign \g8197/_0_  = ~\n834gat_reg/NET0131  ;
  assign \g8211/_0_  = ~\n2562gat_reg/NET0131  ;
  assign \g8223/_0_  = ~\n2634gat_reg/NET0131  ;
  assign \g8237/_0_  = ~\n2203gat_reg/NET0131  ;
  assign \g8251/_0_  = ~\n2640gat_reg/NET0131  ;
  assign \g8261/_0_  = ~\n820gat_reg/NET0131  ;
  assign \g8272/_0_  = ~\n1316gat_reg/NET0131  ;
  assign \g8287/_0_  = ~\n699gat_reg/NET0131  ;
  assign \g8647/_0_  = ~\n2207gat_reg/NET0131  ;
  assign \g8671/_0_  = ~\n2343gat_reg/NET0131  ;
  assign \g8672/_0_  = ~\n2399gat_reg/NET0131  ;
  assign \g8735/_0_  = n965 ;
  assign \g8766/_0_  = ~n966 ;
  assign \g8811/_0_  = ~n967 ;
  assign \g8821/_0_  = ~n979 ;
  assign \g8856/_0_  = n647 ;
  assign \g8858/_3_  = n583 ;
  assign \g8868/_0_  = ~n455 ;
  assign \g8880/_2_  = n980 ;
  assign \g8886/_0_  = ~n996 ;
  assign \g8900/_0_  = ~n997 ;
  assign \g8932/_0_  = ~n1007 ;
  assign \g8991/_3_  = n1008 ;
  assign \g9014/_3_  = n1014 ;
  assign \g9074/_0_  = n511 ;
  assign \g9091/_0_  = ~\n2622gat_reg/NET0131  ;
  assign \g9105/_0_  = ~\n2630gat_reg/NET0131  ;
  assign \g9107/_1_  = ~n363 ;
  assign \g9111/_0_  = ~n1041 ;
  assign \n1332gat_reg/P0001  = ~\n1332gat_reg/NET0131  ;
  assign \n1363gat_reg/P0001  = ~\n1363gat_reg/NET0131  ;
  assign \n1394gat_reg/P0001  = ~\n1394gat_reg/NET0131  ;
  assign \n1433gat_reg/P0001  = ~\n1433gat_reg/NET0131  ;
  assign \n1775gat_reg/P0001  = ~\n1775gat_reg/NET0131  ;
  assign \n2025gat_reg/P0001  = ~\n2025gat_reg/NET0131  ;
  assign \n2029gat_reg/P0001  = ~\n2029gat_reg/NET0131  ;
  assign \n2033gat_reg/P0001  = ~\n2033gat_reg/NET0131  ;
  assign \n2044gat_reg/P0001  = ~\n2044gat_reg/NET0131  ;
  assign \n2121gat_reg/P0001  = ~\n2121gat_reg/NET0131  ;
  assign \n2125gat_reg/P0001  = ~\n2125gat_reg/NET0131  ;
  assign \n2458gat_reg/P0001  = ~\n2458gat_reg/NET0131  ;
  assign \n2472gat_reg/P0001  = ~\n2472gat_reg/NET0131  ;
  assign \n2592gat_reg/P0001  = ~\n2592gat_reg/NET0131  ;
  assign \n3104gat_pad  = ~n1049 ;
  assign \n3105gat_pad  = ~n1053 ;
  assign \n3106gat_pad  = ~\n1871gat_reg/NET0131  ;
  assign \n3107gat_pad  = n1055 ;
  assign \n3108gat_pad  = ~n1056 ;
  assign \n3109gat_pad  = ~n1058 ;
  assign \n3110gat_pad  = n1063 ;
  assign \n3111gat_pad  = ~n1064 ;
  assign \n3112gat_pad  = ~1'b0 ;
  assign \n3113gat_pad  = n1069 ;
  assign \n3114gat_pad  = ~n1070 ;
  assign \n3116gat_pad  = n1079 ;
  assign \n3117gat_pad  = ~n1092 ;
  assign \n3118gat_pad  = ~n1105 ;
  assign \n3119gat_pad  = ~n1118 ;
  assign \n3120gat_pad  = ~n1131 ;
  assign \n3121gat_pad  = ~n1144 ;
  assign \n3122gat_pad  = ~n1157 ;
  assign \n3123gat_pad  = ~n1170 ;
  assign \n3124gat_pad  = ~n1182 ;
  assign \n3125gat_pad  = n1186 ;
  assign \n3126gat_pad  = ~\n2339gat_reg/NET0131  ;
  assign \n3127gat_pad  = ~\n2270gat_reg/NET0131  ;
  assign \n3128gat_pad  = ~\n2390gat_reg/NET0131  ;
  assign \n3130gat_pad  = ~n1197 ;
  assign \n3131gat_pad  = ~n1208 ;
  assign \n3132gat_pad  = ~n1219 ;
  assign \n3133gat_pad  = ~n1230 ;
  assign \n3134gat_pad  = ~n1240 ;
  assign \n3135gat_pad  = ~n1250 ;
  assign \n3136gat_pad  = ~n1260 ;
  assign \n3137gat_pad  = ~n1271 ;
  assign \n3138gat_pad  = n1275 ;
  assign \n3140gat_pad  = ~n1309 ;
  assign \n3142gat_pad  = ~n1329 ;
  assign \n3143gat_pad  = ~n1485 ;
  assign \n3144gat_pad  = ~n1488 ;
  assign \n3145gat_pad  = n1491 ;
  assign \n3146gat_pad  = n1498 ;
  assign \n3147gat_pad  = ~n724 ;
  assign \n3148gat_pad  = ~\n2450gat_reg/NET0131  ;
  assign \n3149gat_pad  = ~n468 ;
  assign \n3150gat_pad  = ~n1500 ;
  assign \n3151gat_pad  = ~n1503 ;
  assign \n684gat_reg/P0001  = ~\n684gat_reg/NET0131  ;
  assign \n824gat_reg/P0001  = ~\n824gat_reg/NET0131  ;
  assign \n883gat_reg/P0001  = ~\n883gat_reg/NET0131  ;
endmodule
