module top (mc_cke_pad_o__pad, mc_vpen_pad_o_pad, \mem_ack_r_reg/P0001 , \poc_o[0]_pad , \poc_o[10]_pad , \poc_o[11]_pad , \poc_o[12]_pad , \poc_o[13]_pad , \poc_o[14]_pad , \poc_o[15]_pad , \poc_o[16]_pad , \poc_o[17]_pad , \poc_o[18]_pad , \poc_o[19]_pad , \poc_o[1]_pad , \poc_o[20]_pad , \poc_o[21]_pad , \poc_o[22]_pad , \poc_o[23]_pad , \poc_o[24]_pad , \poc_o[25]_pad , \poc_o[26]_pad , \poc_o[27]_pad , \poc_o[28]_pad , \poc_o[29]_pad , \poc_o[2]_pad , \poc_o[30]_pad , \poc_o[31]_pad , \poc_o[3]_pad , \poc_o[4]_pad , \poc_o[5]_pad , \poc_o[6]_pad , \poc_o[7]_pad , \poc_o[8]_pad , \poc_o[9]_pad , suspended_o_pad, \u0_cs_reg[0]/NET0131 , \u0_cs_reg[1]/NET0131 , \u0_csc_mask_r_reg[0]/NET0131 , \u0_csc_mask_r_reg[10]/NET0131 , \u0_csc_mask_r_reg[1]/NET0131 , \u0_csc_mask_r_reg[2]/NET0131 , \u0_csc_mask_r_reg[3]/NET0131 , \u0_csc_mask_r_reg[4]/NET0131 , \u0_csc_mask_r_reg[5]/NET0131 , \u0_csc_mask_r_reg[6]/NET0131 , \u0_csc_mask_r_reg[7]/NET0131 , \u0_csc_mask_r_reg[8]/NET0131 , \u0_csc_mask_r_reg[9]/NET0131 , \u0_csc_reg[10]/NET0131 , \u0_csc_reg[11]/NET0131 , \u0_csc_reg[1]/NET0131 , \u0_csc_reg[2]/NET0131 , \u0_csc_reg[3]/NET0131 , \u0_csc_reg[4]/NET0131 , \u0_csc_reg[5]/NET0131 , \u0_csc_reg[6]/NET0131 , \u0_csc_reg[7]/NET0131 , \u0_csc_reg[9]/NET0131 , \u0_csr_r2_reg[0]/NET0131 , \u0_csr_r2_reg[1]/NET0131 , \u0_csr_r2_reg[2]/NET0131 , \u0_csr_r2_reg[3]/NET0131 , \u0_csr_r2_reg[4]/NET0131 , \u0_csr_r2_reg[5]/NET0131 , \u0_csr_r2_reg[6]/NET0131 , \u0_csr_r2_reg[7]/NET0131 , \u0_csr_r_reg[0]/P0001 , \u0_csr_r_reg[10]/NET0131 , \u0_csr_r_reg[2]/NET0131 , \u0_csr_r_reg[3]/NET0131 , \u0_csr_r_reg[4]/NET0131 , \u0_csr_r_reg[5]/NET0131 , \u0_csr_r_reg[6]/NET0131 , \u0_csr_r_reg[7]/NET0131 , \u0_csr_r_reg[8]/NET0131 , \u0_csr_r_reg[9]/NET0131 , \u0_init_ack_r_reg/P0001 , \u0_init_req_reg/NET0131 , \u0_lmr_ack_r_reg/P0001 , \u0_lmr_req_reg/NET0131 , \u0_rf_we_reg/NET0131 , \u0_rst_r2_reg/NET0131 , \u0_sp_csc_reg[10]/NET0131 , \u0_sp_csc_reg[1]/NET0131 , \u0_sp_csc_reg[2]/NET0131 , \u0_sp_csc_reg[3]/NET0131 , \u0_sp_csc_reg[4]/NET0131 , \u0_sp_csc_reg[5]/NET0131 , \u0_sp_csc_reg[6]/NET0131 , \u0_sp_csc_reg[7]/NET0131 , \u0_sp_csc_reg[9]/NET0131 , \u0_sp_tms_reg[0]/NET0131 , \u0_sp_tms_reg[10]/NET0131 , \u0_sp_tms_reg[11]/NET0131 , \u0_sp_tms_reg[12]/NET0131 , \u0_sp_tms_reg[13]/NET0131 , \u0_sp_tms_reg[14]/NET0131 , \u0_sp_tms_reg[15]/NET0131 , \u0_sp_tms_reg[16]/NET0131 , \u0_sp_tms_reg[17]/NET0131 , \u0_sp_tms_reg[18]/NET0131 , \u0_sp_tms_reg[19]/NET0131 , \u0_sp_tms_reg[1]/NET0131 , \u0_sp_tms_reg[20]/NET0131 , \u0_sp_tms_reg[21]/NET0131 , \u0_sp_tms_reg[22]/NET0131 , \u0_sp_tms_reg[23]/NET0131 , \u0_sp_tms_reg[24]/NET0131 , \u0_sp_tms_reg[25]/NET0131 , \u0_sp_tms_reg[26]/NET0131 , \u0_sp_tms_reg[27]/NET0131 , \u0_sp_tms_reg[2]/NET0131 , \u0_sp_tms_reg[3]/NET0131 , \u0_sp_tms_reg[4]/NET0131 , \u0_sp_tms_reg[5]/NET0131 , \u0_sp_tms_reg[6]/NET0131 , \u0_sp_tms_reg[7]/NET0131 , \u0_sp_tms_reg[8]/NET0131 , \u0_sp_tms_reg[9]/NET0131 , \u0_spec_req_cs_reg[0]/NET0131 , \u0_spec_req_cs_reg[1]/NET0131 , \u0_sreq_cs_le_reg/NET0131 , \u0_tms_reg[0]/NET0131 , \u0_tms_reg[10]/NET0131 , \u0_tms_reg[11]/NET0131 , \u0_tms_reg[12]/NET0131 , \u0_tms_reg[13]/NET0131 , \u0_tms_reg[14]/NET0131 , \u0_tms_reg[15]/NET0131 , \u0_tms_reg[16]/NET0131 , \u0_tms_reg[17]/NET0131 , \u0_tms_reg[18]/NET0131 , \u0_tms_reg[19]/NET0131 , \u0_tms_reg[1]/NET0131 , \u0_tms_reg[20]/NET0131 , \u0_tms_reg[21]/NET0131 , \u0_tms_reg[22]/NET0131 , \u0_tms_reg[23]/NET0131 , \u0_tms_reg[24]/NET0131 , \u0_tms_reg[25]/NET0131 , \u0_tms_reg[26]/NET0131 , \u0_tms_reg[27]/NET0131 , \u0_tms_reg[2]/NET0131 , \u0_tms_reg[3]/NET0131 , \u0_tms_reg[4]/NET0131 , \u0_tms_reg[5]/NET0131 , \u0_tms_reg[6]/NET0131 , \u0_tms_reg[7]/NET0131 , \u0_tms_reg[8]/NET0131 , \u0_tms_reg[9]/NET0131 , \u0_u0_addr_r_reg[2]/P0001 , \u0_u0_addr_r_reg[3]/P0001 , \u0_u0_addr_r_reg[4]/P0001 , \u0_u0_addr_r_reg[5]/P0001 , \u0_u0_addr_r_reg[6]/P0001 , \u0_u0_csc_reg[0]/NET0131 , \u0_u0_csc_reg[10]/P0001 , \u0_u0_csc_reg[11]/P0001 , \u0_u0_csc_reg[12]/P0001 , \u0_u0_csc_reg[13]/P0001 , \u0_u0_csc_reg[14]/P0001 , \u0_u0_csc_reg[15]/P0001 , \u0_u0_csc_reg[16]/P0001 , \u0_u0_csc_reg[17]/P0001 , \u0_u0_csc_reg[18]/P0001 , \u0_u0_csc_reg[19]/P0001 , \u0_u0_csc_reg[1]/NET0131 , \u0_u0_csc_reg[20]/P0001 , \u0_u0_csc_reg[21]/P0001 , \u0_u0_csc_reg[22]/P0001 , \u0_u0_csc_reg[23]/P0001 , \u0_u0_csc_reg[24]/P0001 , \u0_u0_csc_reg[25]/P0001 , \u0_u0_csc_reg[26]/P0001 , \u0_u0_csc_reg[27]/P0001 , \u0_u0_csc_reg[28]/P0001 , \u0_u0_csc_reg[29]/P0001 , \u0_u0_csc_reg[2]/NET0131 , \u0_u0_csc_reg[30]/P0001 , \u0_u0_csc_reg[31]/P0001 , \u0_u0_csc_reg[3]/NET0131 , \u0_u0_csc_reg[4]/P0001 , \u0_u0_csc_reg[5]/P0001 , \u0_u0_csc_reg[6]/P0001 , \u0_u0_csc_reg[7]/P0001 , \u0_u0_csc_reg[8]/P0001 , \u0_u0_csc_reg[9]/P0001 , \u0_u0_init_req_reg/NET0131 , \u0_u0_init_req_we_reg/NET0131 , \u0_u0_inited_reg/NET0131 , \u0_u0_lmr_req_reg/NET0131 , \u0_u0_lmr_req_we_reg/NET0131 , \u0_u0_tms_reg[0]/P0001 , \u0_u0_tms_reg[10]/P0001 , \u0_u0_tms_reg[11]/P0001 , \u0_u0_tms_reg[12]/P0001 , \u0_u0_tms_reg[13]/P0001 , \u0_u0_tms_reg[14]/P0001 , \u0_u0_tms_reg[15]/P0001 , \u0_u0_tms_reg[16]/P0001 , \u0_u0_tms_reg[17]/P0001 , \u0_u0_tms_reg[18]/P0001 , \u0_u0_tms_reg[19]/P0001 , \u0_u0_tms_reg[1]/P0001 , \u0_u0_tms_reg[20]/P0001 , \u0_u0_tms_reg[21]/P0001 , \u0_u0_tms_reg[22]/P0001 , \u0_u0_tms_reg[23]/P0001 , \u0_u0_tms_reg[24]/P0001 , \u0_u0_tms_reg[25]/P0001 , \u0_u0_tms_reg[26]/P0001 , \u0_u0_tms_reg[27]/P0001 , \u0_u0_tms_reg[28]/P0001 , \u0_u0_tms_reg[29]/P0001 , \u0_u0_tms_reg[2]/P0001 , \u0_u0_tms_reg[30]/P0001 , \u0_u0_tms_reg[31]/P0001 , \u0_u0_tms_reg[3]/P0001 , \u0_u0_tms_reg[4]/P0001 , \u0_u0_tms_reg[5]/P0001 , \u0_u0_tms_reg[6]/P0001 , \u0_u0_tms_reg[7]/P0001 , \u0_u0_tms_reg[8]/P0001 , \u0_u0_tms_reg[9]/P0001 , \u0_u1_csc_reg[0]/NET0131 , \u0_u1_csc_reg[10]/P0001 , \u0_u1_csc_reg[11]/P0001 , \u0_u1_csc_reg[12]/P0001 , \u0_u1_csc_reg[13]/P0001 , \u0_u1_csc_reg[14]/P0001 , \u0_u1_csc_reg[15]/P0001 , \u0_u1_csc_reg[16]/P0001 , \u0_u1_csc_reg[17]/P0001 , \u0_u1_csc_reg[18]/P0001 , \u0_u1_csc_reg[19]/P0001 , \u0_u1_csc_reg[1]/NET0131 , \u0_u1_csc_reg[20]/P0001 , \u0_u1_csc_reg[21]/P0001 , \u0_u1_csc_reg[22]/P0001 , \u0_u1_csc_reg[23]/P0001 , \u0_u1_csc_reg[24]/P0001 , \u0_u1_csc_reg[25]/P0001 , \u0_u1_csc_reg[26]/P0001 , \u0_u1_csc_reg[27]/P0001 , \u0_u1_csc_reg[28]/P0001 , \u0_u1_csc_reg[29]/P0001 , \u0_u1_csc_reg[2]/NET0131 , \u0_u1_csc_reg[30]/P0001 , \u0_u1_csc_reg[31]/P0001 , \u0_u1_csc_reg[3]/NET0131 , \u0_u1_csc_reg[4]/P0001 , \u0_u1_csc_reg[5]/P0001 , \u0_u1_csc_reg[6]/P0001 , \u0_u1_csc_reg[7]/P0001 , \u0_u1_csc_reg[8]/P0001 , \u0_u1_csc_reg[9]/P0001 , \u0_u1_init_req_reg/NET0131 , \u0_u1_init_req_we_reg/NET0131 , \u0_u1_inited_reg/NET0131 , \u0_u1_lmr_req_reg/NET0131 , \u0_u1_lmr_req_we_reg/NET0131 , \u0_u1_tms_reg[0]/P0001 , \u0_u1_tms_reg[10]/P0001 , \u0_u1_tms_reg[11]/P0001 , \u0_u1_tms_reg[12]/P0001 , \u0_u1_tms_reg[13]/P0001 , \u0_u1_tms_reg[14]/P0001 , \u0_u1_tms_reg[15]/P0001 , \u0_u1_tms_reg[16]/P0001 , \u0_u1_tms_reg[17]/P0001 , \u0_u1_tms_reg[18]/P0001 , \u0_u1_tms_reg[19]/P0001 , \u0_u1_tms_reg[1]/P0001 , \u0_u1_tms_reg[20]/P0001 , \u0_u1_tms_reg[21]/P0001 , \u0_u1_tms_reg[22]/P0001 , \u0_u1_tms_reg[23]/P0001 , \u0_u1_tms_reg[24]/P0001 , \u0_u1_tms_reg[25]/P0001 , \u0_u1_tms_reg[26]/P0001 , \u0_u1_tms_reg[27]/P0001 , \u0_u1_tms_reg[28]/P0001 , \u0_u1_tms_reg[29]/P0001 , \u0_u1_tms_reg[2]/P0001 , \u0_u1_tms_reg[30]/P0001 , \u0_u1_tms_reg[31]/P0001 , \u0_u1_tms_reg[3]/P0001 , \u0_u1_tms_reg[4]/P0001 , \u0_u1_tms_reg[5]/P0001 , \u0_u1_tms_reg[6]/P0001 , \u0_u1_tms_reg[7]/P0001 , \u0_u1_tms_reg[8]/P0001 , \u0_u1_tms_reg[9]/P0001 , \u0_wp_err_reg/NET0131 , \u1_acs_addr_reg[0]/P0001 , \u1_acs_addr_reg[10]/P0001 , \u1_acs_addr_reg[11]/P0001 , \u1_acs_addr_reg[12]/P0001 , \u1_acs_addr_reg[13]/P0001 , \u1_acs_addr_reg[14]/P0001 , \u1_acs_addr_reg[15]/P0001 , \u1_acs_addr_reg[16]/P0001 , \u1_acs_addr_reg[17]/P0001 , \u1_acs_addr_reg[18]/P0001 , \u1_acs_addr_reg[19]/P0001 , \u1_acs_addr_reg[1]/P0001 , \u1_acs_addr_reg[20]/P0001 , \u1_acs_addr_reg[21]/P0001 , \u1_acs_addr_reg[22]/P0001 , \u1_acs_addr_reg[23]/P0001 , \u1_acs_addr_reg[2]/P0001 , \u1_acs_addr_reg[3]/P0001 , \u1_acs_addr_reg[4]/P0001 , \u1_acs_addr_reg[5]/P0001 , \u1_acs_addr_reg[6]/P0001 , \u1_acs_addr_reg[7]/P0001 , \u1_acs_addr_reg[8]/P0001 , \u1_acs_addr_reg[9]/P0001 , \u1_bank_adr_reg[0]/P0001 , \u1_bank_adr_reg[1]/P0001 , \u1_col_adr_reg[0]/P0001 , \u1_col_adr_reg[1]/P0001 , \u1_col_adr_reg[2]/P0001 , \u1_col_adr_reg[3]/P0001 , \u1_col_adr_reg[4]/P0001 , \u1_col_adr_reg[5]/P0001 , \u1_col_adr_reg[6]/P0001 , \u1_col_adr_reg[7]/P0001 , \u1_col_adr_reg[8]/P0001 , \u1_col_adr_reg[9]/P0001 , \u1_row_adr_reg[0]/P0001 , \u1_row_adr_reg[10]/P0001 , \u1_row_adr_reg[11]/P0001 , \u1_row_adr_reg[12]/P0001 , \u1_row_adr_reg[1]/P0001 , \u1_row_adr_reg[2]/P0001 , \u1_row_adr_reg[3]/P0001 , \u1_row_adr_reg[4]/P0001 , \u1_row_adr_reg[5]/P0001 , \u1_row_adr_reg[6]/P0001 , \u1_row_adr_reg[7]/P0001 , \u1_row_adr_reg[8]/P0001 , \u1_row_adr_reg[9]/P0001 , \u1_sram_addr_reg[0]/P0001 , \u1_sram_addr_reg[10]/P0001 , \u1_sram_addr_reg[11]/P0001 , \u1_sram_addr_reg[12]/P0001 , \u1_sram_addr_reg[13]/P0001 , \u1_sram_addr_reg[14]/P0001 , \u1_sram_addr_reg[15]/P0001 , \u1_sram_addr_reg[16]/P0001 , \u1_sram_addr_reg[17]/P0001 , \u1_sram_addr_reg[18]/P0001 , \u1_sram_addr_reg[19]/P0001 , \u1_sram_addr_reg[1]/P0001 , \u1_sram_addr_reg[20]/P0001 , \u1_sram_addr_reg[21]/P0001 , \u1_sram_addr_reg[22]/P0001 , \u1_sram_addr_reg[23]/P0001 , \u1_sram_addr_reg[2]/P0001 , \u1_sram_addr_reg[3]/P0001 , \u1_sram_addr_reg[4]/P0001 , \u1_sram_addr_reg[5]/P0001 , \u1_sram_addr_reg[6]/P0001 , \u1_sram_addr_reg[7]/P0001 , \u1_sram_addr_reg[8]/P0001 , \u1_sram_addr_reg[9]/P0001 , \u1_u0_out_r_reg[0]/P0001 , \u1_u0_out_r_reg[10]/P0001 , \u1_u0_out_r_reg[11]/P0001 , \u1_u0_out_r_reg[12]/P0001 , \u1_u0_out_r_reg[1]/P0001 , \u1_u0_out_r_reg[2]/P0001 , \u1_u0_out_r_reg[3]/P0001 , \u1_u0_out_r_reg[4]/P0001 , \u1_u0_out_r_reg[5]/P0001 , \u1_u0_out_r_reg[6]/P0001 , \u1_u0_out_r_reg[7]/P0001 , \u1_u0_out_r_reg[8]/P0001 , \u1_u0_out_r_reg[9]/P0001 , \u2_bank_open_reg/P0001 , \u2_row_same_reg/P0001 , \u2_u0_b0_last_row_reg[0]/P0001 , \u2_u0_b0_last_row_reg[10]/P0001 , \u2_u0_b0_last_row_reg[11]/P0001 , \u2_u0_b0_last_row_reg[12]/P0001 , \u2_u0_b0_last_row_reg[1]/P0001 , \u2_u0_b0_last_row_reg[2]/P0001 , \u2_u0_b0_last_row_reg[3]/P0001 , \u2_u0_b0_last_row_reg[4]/P0001 , \u2_u0_b0_last_row_reg[5]/P0001 , \u2_u0_b0_last_row_reg[6]/P0001 , \u2_u0_b0_last_row_reg[7]/P0001 , \u2_u0_b0_last_row_reg[8]/P0001 , \u2_u0_b0_last_row_reg[9]/P0001 , \u2_u0_b1_last_row_reg[0]/P0001 , \u2_u0_b1_last_row_reg[10]/P0001 , \u2_u0_b1_last_row_reg[11]/P0001 , \u2_u0_b1_last_row_reg[12]/P0001 , \u2_u0_b1_last_row_reg[1]/P0001 , \u2_u0_b1_last_row_reg[2]/P0001 , \u2_u0_b1_last_row_reg[3]/P0001 , \u2_u0_b1_last_row_reg[4]/P0001 , \u2_u0_b1_last_row_reg[5]/P0001 , \u2_u0_b1_last_row_reg[6]/P0001 , \u2_u0_b1_last_row_reg[7]/P0001 , \u2_u0_b1_last_row_reg[8]/P0001 , \u2_u0_b1_last_row_reg[9]/P0001 , \u2_u0_b2_last_row_reg[0]/P0001 , \u2_u0_b2_last_row_reg[10]/P0001 , \u2_u0_b2_last_row_reg[11]/P0001 , \u2_u0_b2_last_row_reg[12]/P0001 , \u2_u0_b2_last_row_reg[1]/P0001 , \u2_u0_b2_last_row_reg[2]/P0001 , \u2_u0_b2_last_row_reg[3]/P0001 , \u2_u0_b2_last_row_reg[4]/P0001 , \u2_u0_b2_last_row_reg[5]/P0001 , \u2_u0_b2_last_row_reg[6]/P0001 , \u2_u0_b2_last_row_reg[7]/P0001 , \u2_u0_b2_last_row_reg[8]/P0001 , \u2_u0_b2_last_row_reg[9]/P0001 , \u2_u0_b3_last_row_reg[0]/P0001 , \u2_u0_b3_last_row_reg[10]/P0001 , \u2_u0_b3_last_row_reg[11]/P0001 , \u2_u0_b3_last_row_reg[12]/P0001 , \u2_u0_b3_last_row_reg[1]/P0001 , \u2_u0_b3_last_row_reg[2]/P0001 , \u2_u0_b3_last_row_reg[3]/P0001 , \u2_u0_b3_last_row_reg[4]/P0001 , \u2_u0_b3_last_row_reg[5]/P0001 , \u2_u0_b3_last_row_reg[6]/P0001 , \u2_u0_b3_last_row_reg[7]/P0001 , \u2_u0_b3_last_row_reg[8]/P0001 , \u2_u0_b3_last_row_reg[9]/P0001 , \u2_u0_bank0_open_reg/NET0131 , \u2_u0_bank1_open_reg/NET0131 , \u2_u0_bank2_open_reg/NET0131 , \u2_u0_bank3_open_reg/NET0131 , \u2_u1_b0_last_row_reg[0]/P0001 , \u2_u1_b0_last_row_reg[10]/P0001 , \u2_u1_b0_last_row_reg[11]/P0001 , \u2_u1_b0_last_row_reg[12]/P0001 , \u2_u1_b0_last_row_reg[1]/P0001 , \u2_u1_b0_last_row_reg[2]/P0001 , \u2_u1_b0_last_row_reg[3]/P0001 , \u2_u1_b0_last_row_reg[4]/P0001 , \u2_u1_b0_last_row_reg[5]/P0001 , \u2_u1_b0_last_row_reg[6]/P0001 , \u2_u1_b0_last_row_reg[7]/P0001 , \u2_u1_b0_last_row_reg[8]/P0001 , \u2_u1_b0_last_row_reg[9]/P0001 , \u2_u1_b1_last_row_reg[0]/P0001 , \u2_u1_b1_last_row_reg[10]/P0001 , \u2_u1_b1_last_row_reg[11]/P0001 , \u2_u1_b1_last_row_reg[12]/P0001 , \u2_u1_b1_last_row_reg[1]/P0001 , \u2_u1_b1_last_row_reg[2]/P0001 , \u2_u1_b1_last_row_reg[3]/P0001 , \u2_u1_b1_last_row_reg[4]/P0001 , \u2_u1_b1_last_row_reg[5]/P0001 , \u2_u1_b1_last_row_reg[6]/P0001 , \u2_u1_b1_last_row_reg[7]/P0001 , \u2_u1_b1_last_row_reg[8]/P0001 , \u2_u1_b1_last_row_reg[9]/P0001 , \u2_u1_b2_last_row_reg[0]/P0001 , \u2_u1_b2_last_row_reg[10]/P0001 , \u2_u1_b2_last_row_reg[11]/P0001 , \u2_u1_b2_last_row_reg[12]/P0001 , \u2_u1_b2_last_row_reg[1]/P0001 , \u2_u1_b2_last_row_reg[2]/P0001 , \u2_u1_b2_last_row_reg[3]/P0001 , \u2_u1_b2_last_row_reg[4]/P0001 , \u2_u1_b2_last_row_reg[5]/P0001 , \u2_u1_b2_last_row_reg[6]/P0001 , \u2_u1_b2_last_row_reg[7]/P0001 , \u2_u1_b2_last_row_reg[8]/P0001 , \u2_u1_b2_last_row_reg[9]/P0001 , \u2_u1_b3_last_row_reg[0]/P0001 , \u2_u1_b3_last_row_reg[10]/P0001 , \u2_u1_b3_last_row_reg[11]/P0001 , \u2_u1_b3_last_row_reg[12]/P0001 , \u2_u1_b3_last_row_reg[1]/P0001 , \u2_u1_b3_last_row_reg[2]/P0001 , \u2_u1_b3_last_row_reg[3]/P0001 , \u2_u1_b3_last_row_reg[4]/P0001 , \u2_u1_b3_last_row_reg[5]/P0001 , \u2_u1_b3_last_row_reg[6]/P0001 , \u2_u1_b3_last_row_reg[7]/P0001 , \u2_u1_b3_last_row_reg[8]/P0001 , \u2_u1_b3_last_row_reg[9]/P0001 , \u2_u1_bank0_open_reg/NET0131 , \u2_u1_bank1_open_reg/NET0131 , \u2_u1_bank2_open_reg/NET0131 , \u2_u1_bank3_open_reg/NET0131 , \u3_byte0_reg[0]/P0001 , \u3_byte0_reg[1]/P0001 , \u3_byte0_reg[2]/P0001 , \u3_byte0_reg[3]/P0001 , \u3_byte0_reg[4]/P0001 , \u3_byte0_reg[5]/P0001 , \u3_byte0_reg[6]/P0001 , \u3_byte0_reg[7]/P0001 , \u3_byte1_reg[0]/P0001 , \u3_byte1_reg[1]/P0001 , \u3_byte1_reg[2]/P0001 , \u3_byte1_reg[3]/P0001 , \u3_byte1_reg[4]/P0001 , \u3_byte1_reg[5]/P0001 , \u3_byte1_reg[6]/P0001 , \u3_byte1_reg[7]/P0001 , \u3_byte2_reg[0]/P0001 , \u3_byte2_reg[1]/P0001 , \u3_byte2_reg[2]/P0001 , \u3_byte2_reg[3]/P0001 , \u3_byte2_reg[4]/P0001 , \u3_byte2_reg[5]/P0001 , \u3_byte2_reg[6]/P0001 , \u3_byte2_reg[7]/P0001 , \u3_u0_r0_reg[0]/P0001 , \u3_u0_r0_reg[10]/P0001 , \u3_u0_r0_reg[11]/P0001 , \u3_u0_r0_reg[12]/P0001 , \u3_u0_r0_reg[13]/P0001 , \u3_u0_r0_reg[14]/P0001 , \u3_u0_r0_reg[15]/P0001 , \u3_u0_r0_reg[16]/P0001 , \u3_u0_r0_reg[17]/P0001 , \u3_u0_r0_reg[18]/P0001 , \u3_u0_r0_reg[19]/P0001 , \u3_u0_r0_reg[1]/P0001 , \u3_u0_r0_reg[20]/P0001 , \u3_u0_r0_reg[21]/P0001 , \u3_u0_r0_reg[22]/P0001 , \u3_u0_r0_reg[23]/P0001 , \u3_u0_r0_reg[24]/P0001 , \u3_u0_r0_reg[25]/P0001 , \u3_u0_r0_reg[26]/P0001 , \u3_u0_r0_reg[27]/P0001 , \u3_u0_r0_reg[28]/P0001 , \u3_u0_r0_reg[29]/P0001 , \u3_u0_r0_reg[2]/P0001 , \u3_u0_r0_reg[30]/P0001 , \u3_u0_r0_reg[31]/P0001 , \u3_u0_r0_reg[32]/P0001 , \u3_u0_r0_reg[33]/P0001 , \u3_u0_r0_reg[34]/P0001 , \u3_u0_r0_reg[35]/P0001 , \u3_u0_r0_reg[3]/P0001 , \u3_u0_r0_reg[4]/P0001 , \u3_u0_r0_reg[5]/P0001 , \u3_u0_r0_reg[6]/P0001 , \u3_u0_r0_reg[7]/P0001 , \u3_u0_r0_reg[8]/P0001 , \u3_u0_r0_reg[9]/P0001 , \u3_u0_r1_reg[0]/P0001 , \u3_u0_r1_reg[10]/P0001 , \u3_u0_r1_reg[11]/P0001 , \u3_u0_r1_reg[12]/P0001 , \u3_u0_r1_reg[13]/P0001 , \u3_u0_r1_reg[14]/P0001 , \u3_u0_r1_reg[15]/P0001 , \u3_u0_r1_reg[16]/P0001 , \u3_u0_r1_reg[17]/P0001 , \u3_u0_r1_reg[18]/P0001 , \u3_u0_r1_reg[19]/P0001 , \u3_u0_r1_reg[1]/P0001 , \u3_u0_r1_reg[20]/P0001 , \u3_u0_r1_reg[21]/P0001 , \u3_u0_r1_reg[22]/P0001 , \u3_u0_r1_reg[23]/P0001 , \u3_u0_r1_reg[24]/P0001 , \u3_u0_r1_reg[25]/P0001 , \u3_u0_r1_reg[26]/P0001 , \u3_u0_r1_reg[27]/P0001 , \u3_u0_r1_reg[28]/P0001 , \u3_u0_r1_reg[29]/P0001 , \u3_u0_r1_reg[2]/P0001 , \u3_u0_r1_reg[30]/P0001 , \u3_u0_r1_reg[31]/P0001 , \u3_u0_r1_reg[32]/P0001 , \u3_u0_r1_reg[33]/P0001 , \u3_u0_r1_reg[34]/P0001 , \u3_u0_r1_reg[35]/P0001 , \u3_u0_r1_reg[3]/P0001 , \u3_u0_r1_reg[4]/P0001 , \u3_u0_r1_reg[5]/P0001 , \u3_u0_r1_reg[6]/P0001 , \u3_u0_r1_reg[7]/P0001 , \u3_u0_r1_reg[8]/P0001 , \u3_u0_r1_reg[9]/P0001 , \u3_u0_r2_reg[0]/P0001 , \u3_u0_r2_reg[10]/P0001 , \u3_u0_r2_reg[11]/P0001 , \u3_u0_r2_reg[12]/P0001 , \u3_u0_r2_reg[13]/P0001 , \u3_u0_r2_reg[14]/P0001 , \u3_u0_r2_reg[15]/P0001 , \u3_u0_r2_reg[16]/P0001 , \u3_u0_r2_reg[17]/P0001 , \u3_u0_r2_reg[18]/P0001 , \u3_u0_r2_reg[19]/P0001 , \u3_u0_r2_reg[1]/P0001 , \u3_u0_r2_reg[20]/P0001 , \u3_u0_r2_reg[21]/P0001 , \u3_u0_r2_reg[22]/P0001 , \u3_u0_r2_reg[23]/P0001 , \u3_u0_r2_reg[24]/P0001 , \u3_u0_r2_reg[25]/P0001 , \u3_u0_r2_reg[26]/P0001 , \u3_u0_r2_reg[27]/P0001 , \u3_u0_r2_reg[28]/P0001 , \u3_u0_r2_reg[29]/P0001 , \u3_u0_r2_reg[2]/P0001 , \u3_u0_r2_reg[30]/P0001 , \u3_u0_r2_reg[31]/P0001 , \u3_u0_r2_reg[32]/P0001 , \u3_u0_r2_reg[33]/P0001 , \u3_u0_r2_reg[34]/P0001 , \u3_u0_r2_reg[35]/P0001 , \u3_u0_r2_reg[3]/P0001 , \u3_u0_r2_reg[4]/P0001 , \u3_u0_r2_reg[5]/P0001 , \u3_u0_r2_reg[6]/P0001 , \u3_u0_r2_reg[7]/P0001 , \u3_u0_r2_reg[8]/P0001 , \u3_u0_r2_reg[9]/P0001 , \u3_u0_r3_reg[0]/P0001 , \u3_u0_r3_reg[10]/P0001 , \u3_u0_r3_reg[11]/P0001 , \u3_u0_r3_reg[12]/P0001 , \u3_u0_r3_reg[13]/P0001 , \u3_u0_r3_reg[14]/P0001 , \u3_u0_r3_reg[15]/P0001 , \u3_u0_r3_reg[16]/P0001 , \u3_u0_r3_reg[17]/P0001 , \u3_u0_r3_reg[18]/P0001 , \u3_u0_r3_reg[19]/P0001 , \u3_u0_r3_reg[1]/P0001 , \u3_u0_r3_reg[20]/P0001 , \u3_u0_r3_reg[21]/P0001 , \u3_u0_r3_reg[22]/P0001 , \u3_u0_r3_reg[23]/P0001 , \u3_u0_r3_reg[24]/P0001 , \u3_u0_r3_reg[25]/P0001 , \u3_u0_r3_reg[26]/P0001 , \u3_u0_r3_reg[27]/P0001 , \u3_u0_r3_reg[28]/P0001 , \u3_u0_r3_reg[29]/P0001 , \u3_u0_r3_reg[2]/P0001 , \u3_u0_r3_reg[30]/P0001 , \u3_u0_r3_reg[31]/P0001 , \u3_u0_r3_reg[32]/P0001 , \u3_u0_r3_reg[33]/P0001 , \u3_u0_r3_reg[34]/P0001 , \u3_u0_r3_reg[35]/P0001 , \u3_u0_r3_reg[3]/P0001 , \u3_u0_r3_reg[4]/P0001 , \u3_u0_r3_reg[5]/P0001 , \u3_u0_r3_reg[6]/P0001 , \u3_u0_r3_reg[7]/P0001 , \u3_u0_r3_reg[8]/P0001 , \u3_u0_r3_reg[9]/P0001 , \u3_u0_rd_adr_reg[0]/NET0131 , \u3_u0_rd_adr_reg[1]/NET0131 , \u3_u0_rd_adr_reg[2]/NET0131 , \u3_u0_rd_adr_reg[3]/NET0131 , \u3_u0_wr_adr_reg[0]/NET0131 , \u3_u0_wr_adr_reg[1]/NET0131 , \u3_u0_wr_adr_reg[2]/NET0131 , \u3_u0_wr_adr_reg[3]/NET0131 , \u4_ps_cnt_reg[0]/NET0131 , \u4_ps_cnt_reg[1]/NET0131 , \u4_ps_cnt_reg[2]/NET0131 , \u4_ps_cnt_reg[3]/NET0131 , \u4_ps_cnt_reg[4]/NET0131 , \u4_ps_cnt_reg[5]/NET0131 , \u4_ps_cnt_reg[6]/NET0131 , \u4_ps_cnt_reg[7]/NET0131 , \u4_rfr_ce_reg/NET0131 , \u4_rfr_clr_reg/P0001 , \u4_rfr_cnt_reg[0]/NET0131 , \u4_rfr_cnt_reg[1]/NET0131 , \u4_rfr_cnt_reg[2]/NET0131 , \u4_rfr_cnt_reg[3]/NET0131 , \u4_rfr_cnt_reg[4]/NET0131 , \u4_rfr_cnt_reg[5]/NET0131 , \u4_rfr_cnt_reg[6]/NET0131 , \u4_rfr_cnt_reg[7]/NET0131 , \u4_rfr_early_reg/NET0131 , \u4_rfr_en_reg/NET0131 , \u4_rfr_req_reg/NET0131 , \u5_ack_cnt_reg[0]/NET0131 , \u5_ack_cnt_reg[1]/NET0131 , \u5_ack_cnt_reg[2]/NET0131 , \u5_ack_cnt_reg[3]/NET0131 , \u5_ap_en_reg/NET0131 , \u5_burst_act_rd_reg/P0001 , \u5_burst_cnt_reg[0]/NET0131 , \u5_burst_cnt_reg[10]/NET0131 , \u5_burst_cnt_reg[1]/NET0131 , \u5_burst_cnt_reg[2]/NET0131 , \u5_burst_cnt_reg[3]/NET0131 , \u5_burst_cnt_reg[4]/NET0131 , \u5_burst_cnt_reg[5]/NET0131 , \u5_burst_cnt_reg[6]/NET0131 , \u5_burst_cnt_reg[7]/NET0131 , \u5_burst_cnt_reg[8]/NET0131 , \u5_burst_cnt_reg[9]/NET0131 , \u5_cke_o_del_reg/P0001 , \u5_cke_r_reg/NET0131 , \u5_cmd_a10_r_reg/P0001 , \u5_cmd_asserted2_reg/NET0131 , \u5_cmd_asserted_reg/NET0131 , \u5_cmd_del_reg[0]/NET0131 , \u5_cmd_del_reg[1]/NET0131 , \u5_cmd_del_reg[2]/NET0131 , \u5_cmd_del_reg[3]/NET0131 , \u5_cnt_reg/NET0131 , \u5_cs_le_r_reg/P0001 , \u5_cs_le_reg/P0001 , \u5_data_oe_r2_reg/NET0131 , \u5_data_oe_reg/NET0131 , \u5_dv_r_reg/NET0131 , \u5_ir_cnt_done_reg/P0001 , \u5_ir_cnt_reg[0]/P0001 , \u5_ir_cnt_reg[1]/P0001 , \u5_ir_cnt_reg[2]/P0001 , \u5_ir_cnt_reg[3]/P0001 , \u5_lmr_ack_reg/NET0131 , \u5_lookup_ready1_reg/NET0131 , \u5_lookup_ready2_reg/NET0131 , \u5_mc_adv_r1_reg/NET0131 , \u5_mc_adv_r_reg/NET0131 , \u5_mc_c_oe_reg/NET0131 , \u5_mc_le_reg/NET0131 , \u5_mem_ack_r_reg/NET0131 , \u5_no_wb_cycle_reg/NET0131 , \u5_oe__reg/NET0131 , \u5_pack_le0_reg/P0001 , \u5_pack_le1_reg/P0001 , \u5_resume_req_r_reg/NET0131 , \u5_rfr_ack_r_reg/NET0131 , \u5_state_reg[0]/NET0131 , \u5_state_reg[10]/NET0131 , \u5_state_reg[11]/NET0131 , \u5_state_reg[12]/NET0131 , \u5_state_reg[13]/NET0131 , \u5_state_reg[14]/NET0131 , \u5_state_reg[15]/NET0131 , \u5_state_reg[16]/NET0131 , \u5_state_reg[17]/NET0131 , \u5_state_reg[18]/NET0131 , \u5_state_reg[19]/NET0131 , \u5_state_reg[1]/NET0131 , \u5_state_reg[20]/NET0131 , \u5_state_reg[21]/NET0131 , \u5_state_reg[22]/NET0131 , \u5_state_reg[23]/NET0131 , \u5_state_reg[24]/NET0131 , \u5_state_reg[25]/NET0131 , \u5_state_reg[26]/NET0131 , \u5_state_reg[27]/NET0131 , \u5_state_reg[28]/NET0131 , \u5_state_reg[29]/NET0131 , \u5_state_reg[2]/NET0131 , \u5_state_reg[30]/NET0131 , \u5_state_reg[31]/NET0131 , \u5_state_reg[32]/NET0131 , \u5_state_reg[33]/NET0131 , \u5_state_reg[34]/NET0131 , \u5_state_reg[35]/NET0131 , \u5_state_reg[36]/NET0131 , \u5_state_reg[37]/NET0131 , \u5_state_reg[38]/NET0131 , \u5_state_reg[39]/NET0131 , \u5_state_reg[3]/NET0131 , \u5_state_reg[40]/NET0131 , \u5_state_reg[41]/NET0131 , \u5_state_reg[42]/NET0131 , \u5_state_reg[43]/NET0131 , \u5_state_reg[44]/NET0131 , \u5_state_reg[45]/NET0131 , \u5_state_reg[46]/NET0131 , \u5_state_reg[47]/NET0131 , \u5_state_reg[48]/NET0131 , \u5_state_reg[49]/NET0131 , \u5_state_reg[4]/NET0131 , \u5_state_reg[50]/NET0131 , \u5_state_reg[51]/NET0131 , \u5_state_reg[52]/NET0131 , \u5_state_reg[53]/NET0131 , \u5_state_reg[54]/NET0131 , \u5_state_reg[55]/NET0131 , \u5_state_reg[56]/NET0131 , \u5_state_reg[57]/NET0131 , \u5_state_reg[58]/NET0131 , \u5_state_reg[59]/NET0131 , \u5_state_reg[5]/NET0131 , \u5_state_reg[60]/NET0131 , \u5_state_reg[61]/NET0131 , \u5_state_reg[62]/NET0131 , \u5_state_reg[63]/NET0131 , \u5_state_reg[64]/NET0131 , \u5_state_reg[65]/NET0131 , \u5_state_reg[6]/NET0131 , \u5_state_reg[7]/NET0131 , \u5_state_reg[8]/NET0131 , \u5_state_reg[9]/NET0131 , \u5_susp_req_r_reg/NET0131 , \u5_susp_sel_r_reg/NET0131 , \u5_timer2_reg[0]/P0001 , \u5_timer2_reg[1]/P0001 , \u5_timer2_reg[2]/P0001 , \u5_timer2_reg[3]/P0001 , \u5_timer2_reg[4]/P0001 , \u5_timer2_reg[5]/P0001 , \u5_timer2_reg[6]/P0001 , \u5_timer2_reg[7]/P0001 , \u5_timer2_reg[8]/P0001 , \u5_timer_reg[0]/NET0131 , \u5_timer_reg[1]/NET0131 , \u5_timer_reg[2]/NET0131 , \u5_timer_reg[3]/NET0131 , \u5_timer_reg[4]/NET0131 , \u5_timer_reg[5]/NET0131 , \u5_timer_reg[6]/NET0131 , \u5_timer_reg[7]/NET0131 , \u5_tmr2_done_reg/NET0131 , \u5_tmr_done_reg/NET0131 , \u5_wb_cycle_reg/NET0131 , \u5_wb_stb_first_reg/NET0131 , \u5_wb_wait_r_reg/P0001 , \u5_wb_write_go_r_reg/NET0131 , \u5_wr_cycle_reg/NET0131 , \u6_read_go_r1_reg/NET0131 , \u6_read_go_r_reg/NET0131 , \u6_rmw_en_reg/NET0131 , \u6_rmw_r_reg/NET0131 , \u6_wb_first_r_reg/NET0131 , \u6_wr_hold_reg/NET0131 , \u6_write_go_r1_reg/NET0131 , \u6_write_go_r_reg/NET0131 , \u7_mc_ack_r_reg/NET0131 , \u7_mc_br_r_reg/P0001 , \u7_mc_data_ir_reg[0]/P0001 , \u7_mc_data_ir_reg[10]/P0001 , \u7_mc_data_ir_reg[11]/P0001 , \u7_mc_data_ir_reg[12]/P0001 , \u7_mc_data_ir_reg[13]/P0001 , \u7_mc_data_ir_reg[14]/P0001 , \u7_mc_data_ir_reg[15]/P0001 , \u7_mc_data_ir_reg[16]/P0001 , \u7_mc_data_ir_reg[17]/P0001 , \u7_mc_data_ir_reg[18]/P0001 , \u7_mc_data_ir_reg[19]/P0001 , \u7_mc_data_ir_reg[1]/P0001 , \u7_mc_data_ir_reg[20]/P0001 , \u7_mc_data_ir_reg[21]/P0001 , \u7_mc_data_ir_reg[22]/P0001 , \u7_mc_data_ir_reg[23]/P0001 , \u7_mc_data_ir_reg[24]/P0001 , \u7_mc_data_ir_reg[25]/P0001 , \u7_mc_data_ir_reg[26]/P0001 , \u7_mc_data_ir_reg[27]/P0001 , \u7_mc_data_ir_reg[28]/P0001 , \u7_mc_data_ir_reg[29]/P0001 , \u7_mc_data_ir_reg[2]/P0001 , \u7_mc_data_ir_reg[30]/P0001 , \u7_mc_data_ir_reg[31]/P0001 , \u7_mc_data_ir_reg[3]/P0001 , \u7_mc_data_ir_reg[4]/P0001 , \u7_mc_data_ir_reg[5]/P0001 , \u7_mc_data_ir_reg[6]/P0001 , \u7_mc_data_ir_reg[7]/P0001 , \u7_mc_data_ir_reg[8]/P0001 , \u7_mc_data_ir_reg[9]/P0001 , \u7_mc_dqm_r2_reg[0]/P0001 , \u7_mc_dqm_r2_reg[1]/P0001 , \u7_mc_dqm_r2_reg[2]/P0001 , \u7_mc_dqm_r2_reg[3]/P0001 , \u7_mc_dqm_r_reg[0]/P0001 , \u7_mc_dqm_r_reg[1]/P0001 , \u7_mc_dqm_r_reg[2]/P0001 , \u7_mc_dqm_r_reg[3]/P0001 , wb_ack_o_pad, \wb_addr_i[0]_pad , \wb_addr_i[10]_pad , \wb_addr_i[11]_pad , \wb_addr_i[12]_pad , \wb_addr_i[13]_pad , \wb_addr_i[14]_pad , \wb_addr_i[15]_pad , \wb_addr_i[16]_pad , \wb_addr_i[17]_pad , \wb_addr_i[18]_pad , \wb_addr_i[19]_pad , \wb_addr_i[1]_pad , \wb_addr_i[20]_pad , \wb_addr_i[21]_pad , \wb_addr_i[22]_pad , \wb_addr_i[23]_pad , \wb_addr_i[24]_pad , \wb_addr_i[25]_pad , \wb_addr_i[26]_pad , \wb_addr_i[27]_pad , \wb_addr_i[28]_pad , \wb_addr_i[29]_pad , \wb_addr_i[2]_pad , \wb_addr_i[30]_pad , \wb_addr_i[31]_pad , \wb_addr_i[3]_pad , \wb_addr_i[4]_pad , \wb_addr_i[5]_pad , \wb_addr_i[6]_pad , \wb_addr_i[7]_pad , \wb_addr_i[8]_pad , \wb_addr_i[9]_pad , wb_cyc_i_pad, \wb_data_i[0]_pad , \wb_data_i[10]_pad , \wb_data_i[11]_pad , \wb_data_i[12]_pad , \wb_data_i[13]_pad , \wb_data_i[14]_pad , \wb_data_i[15]_pad , \wb_data_i[16]_pad , \wb_data_i[17]_pad , \wb_data_i[18]_pad , \wb_data_i[19]_pad , \wb_data_i[1]_pad , \wb_data_i[20]_pad , \wb_data_i[21]_pad , \wb_data_i[22]_pad , \wb_data_i[23]_pad , \wb_data_i[24]_pad , \wb_data_i[25]_pad , \wb_data_i[26]_pad , \wb_data_i[27]_pad , \wb_data_i[28]_pad , \wb_data_i[29]_pad , \wb_data_i[2]_pad , \wb_data_i[30]_pad , \wb_data_i[31]_pad , \wb_data_i[3]_pad , \wb_data_i[4]_pad , \wb_data_i[5]_pad , \wb_data_i[6]_pad , \wb_data_i[7]_pad , \wb_data_i[8]_pad , \wb_data_i[9]_pad , wb_err_o_pad, \wb_sel_i[0]_pad , \wb_sel_i[1]_pad , \wb_sel_i[2]_pad , \wb_sel_i[3]_pad , wb_stb_i_pad, wb_we_i_pad, \_al_n0 , \_al_n1 , \g22/_0_ , \g23/_0_ , \g25_dup61718/_2_ , \g43466/_0_ , \g43467/_0_ , \g43468/_0_ , \g43469/_0_ , \g43470/_0_ , \g43471/_0_ , \g43472/_0_ , \g43473/_0_ , \g43474/_0_ , \g43475/_0_ , \g43476/_0_ , \g43477/_0_ , \g43478/_0_ , \g43512/_0_ , \g43513/_0_ , \g43544/_3_ , \g43545/_0_ , \g43554/_0_ , \g43555/_0_ , \g43557/_0_ , \g43558/_0_ , \g43571/_2_ , \g43632/_0_ , \g43633/_0_ , \g43635/_0_ , \g43636/_0_ , \g43637/_0_ , \g43638/_0_ , \g43639/_0_ , \g43640/_0_ , \g43642/_0_ , \g43662/_0_ , \g43663/_0_ , \g43664/_0_ , \g43665/_0_ , \g43668/_0_ , \g43670/_0_ , \g43671/_0_ , \g43673/_0_ , \g43674/_0_ , \g43692/_0_ , \g43695/_0_ , \g43696/_0_ , \g43697/_0_ , \g43698/_0_ , \g43700/_0_ , \g43701/_0_ , \g43703/_0_ , \g43705/_0_ , \g43707/_0_ , \g43708/_0_ , \g43710/_0_ , \g43717/_0_ , \g43719/_0_ , \g43720/_0_ , \g43721/_0_ , \g43722/_1_ , \g43723/_0_ , \g43725/_0_ , \g43729/_0_ , \g43731/_0_ , \g43734/_0_ , \g43735/_0_ , \g43737/_0_ , \g43744/_0_ , \g43747/_0_ , \g43760/_2_ , \g43770/_1_ , \g43775/_2_ , \g43780/_2_ , \g43786/_0_ , \g43787/_1_ , \g43847/_0_ , \g43848/_1_ , \g43858/_1_ , \g43891/_3_ , \g43895/_0_ , \g43934/_0_ , \g43936/_3_ , \g43954/_3_ , \g43961/_0_ , \g44016/_1_ , \g44067/_0_ , \g44094/_0_ , \g44096/_0_ , \g44104/_0_ , \g44122/_0_ , \g44172/_0_ , \g44209/_0_ , \g44219/_0_ , \g44220/_0_ , \g44222/_0_ , \g44223/_0_ , \g44241/_2_ , \g44252/_0_ , \g44253/_0_ , \g44255/_2_ , \g44263/_2_ , \g44470/_0_ , \g44538/_0_ , \g44539/_0_ , \g44540/_0_ , \g44541/_0_ , \g44542/_0_ , \g44543/_0_ , \g44544/_0_ , \g44545/_0_ , \g44546/_0_ , \g44547/_0_ , \g44548/_0_ , \g44549/_0_ , \g44550/_0_ , \g44551/_0_ , \g44552/_0_ , \g44553/_0_ , \g44554/_0_ , \g44555/_0_ , \g44556/_0_ , \g44557/_0_ , \g44558/_0_ , \g44559/_0_ , \g44560/_0_ , \g44561/_0_ , \g44562/_0_ , \g44563/_0_ , \g44564/_0_ , \g44565/_0_ , \g44566/_0_ , \g44567/_0_ , \g44568/_0_ , \g44569/_0_ , \g44570/_0_ , \g44571/_0_ , \g44572/_0_ , \g44573/_0_ , \g44574/_0_ , \g44575/_0_ , \g44576/_0_ , \g44577/_0_ , \g44578/_0_ , \g44579/_0_ , \g44580/_0_ , \g44581/_0_ , \g44582/_0_ , \g44583/_0_ , \g44584/_0_ , \g44585/_0_ , \g44586/_0_ , \g44588/_0_ , \g44589/_0_ , \g44590/_0_ , \g44591/_0_ , \g44592/_0_ , \g44593/_0_ , \g44594/_0_ , \g44595/_0_ , \g44596/_0_ , \g44636/_2_ , \g44646/_0_ , \g44647/_0_ , \g44648/_0_ , \g44649/_0_ , \g44650/_0_ , \g44651/_0_ , \g44652/_0_ , \g44653/_0_ , \g44654/_0_ , \g44655/_0_ , \g44656/_0_ , \g44657/_0_ , \g44665/_0_ , \g44666/_0_ , \g44667/_0_ , \g44668/_0_ , \g44752/_0_ , \g44753/_0_ , \g44873/_0_ , \g44939/_0_ , \g44942/_0_ , \g44945/_0_ , \g45023/_2_ , \g45090/_0_ , \g45141/_0_ , \g45147/_3_ , \g45155/_0_ , \g45190/_0_ , \g45195/_2_ , \g45199/_2_ , \g45201/_2_ , \g45324/_0_ , \g45334/_2_ , \g45336/_0_ , \g45388/_0_ , \g45391/_0_ , \g45413/_2_ , \g45530/_0_ , \g45532/_0_ , \g45533/_0_ , \g45534/_0_ , \g45739/_2_ , \g45743/_2_ , \g45767/_0_ , \g45782/_0_ , \g45830/_3_ , \g45834/_3_ , \g45835/_3_ , \g45836/_3_ , \g45837/_3_ , \g45839/_3_ , \g45840/_3_ , \g45841/_3_ , \g45842/_3_ , \g45843/_3_ , \g45844/_3_ , \g45845/_3_ , \g46191/_0_ , \g46193/_3_ , \g46256/_3_ , \g46257/_3_ , \g46258/_3_ , \g46259/_3_ , \g46260/_3_ , \g46261/_3_ , \g46262/_3_ , \g46263/_3_ , \g46278/_0_ , \g46292/_0_ , \g46293/_0_ , \g46312/_0_ , \g46367/_2_ , \g46370/_2_ , \g46380/_2_ , \g46386/_2_ , \g46388/_2_ , \g46392/_2_ , \g46395/_2_ , \g46399/_2_ , \g46420/_0_ , \g46446/_0_ , \g46493/_0_ , \g46510/_0_ , \g46669/_2_ , \g46691/_0_ , \g46708/_0_ , \g46721/_00_ , \g46776/_0_ , \g46777/_0_ , \g46778/_0_ , \g46779/_0_ , \g46780/_0_ , \g46782/_0_ , \g46784/_0_ , \g46932/_0_ , \g47112/_0_ , \g47124/_0_ , \g47265/_0_ , \g47270/_0_ , \g47275/_0_ , \g47300/_1_ , \g47305/_1_ , \g47338/_0_ , \g47339/_0_ , \g47352/_0_ , \g47699/_3_ , \g47711/_0_ , \g47719/_3_ , \g47721/_3_ , \g47723/_3_ , \g47853/_0_ , \g48094/_0_ , \g48095/_0_ , \g48177/_2_ , \g48194/_0_ , \g48369/_2_ , \g48371/_2_ , \g48373/_2_ , \g48375/_2_ , \g48377/_2_ , \g48379/_2_ , \g48381/_2_ , \g48383/_2_ , \g48385/_2_ , \g48535/_0_ , \g48569/_0_ , \g48570/_0_ , \g48571/_0_ , \g48836/_0_ , \g48843/_0_ , \g49187/_3_ , \g49375/_2_ , \g49633/_0_ , \g49788/_1_ , \g49800/_1_ , \g49802/_1_ , \g49806/_1_ , \g49853/_1_ , \g49883/_0_ , \g49884/_0_ , \g49885/_0_ , \g49886/_0_ , \g49976/_1_ , \g50038/_0_ , \g50082/_0_ , \g50083/_0_ , \g50167/_3_ , \g50168/_3_ , \g50169/_3_ , \g50170/_3_ , \g50171/_3_ , \g50177/_0_ , \g50190/_0_ , \g50236/_0_ , \g50251/_3_ , \g50256/_0_ , \g50318/_3_ , \g50319/_3_ , \g50350/_3_ , \g50351/_3_ , \g50352/_3_ , \g50353/_3_ , \g50354/_3_ , \g50355/_3_ , \g50361/_2_ , \g50366/_0_ , \g50393/_0_ , \g50552/_1_ , \g51108/_0_ , \g51160/_0_ , \g51290/_1_ , \g51327/_3_ , \g51328/_3_ , \g51329/_3_ , \g51330/_3_ , \g51331/_3_ , \g51332/_3_ , \g51333/_3_ , \g51334/_3_ , \g51339/_3_ , \g51340/_3_ , \g51341/_3_ , \g51342/_3_ , \g51343/_3_ , \g51346/_0_ , \g51347/_0_ , \g51348/_0_ , \g51381/_3_ , \g51382/_3_ , \g51383/_3_ , \g51386/_3_ , \g51387/_3_ , \g51405/_3_ , \g51410/_3_ , \g51883/_0_ , \g51916/_0_ , \g51947/_0_ , \g51948/_0_ , \g51949/_0_ , \g51950/_0_ , \g51951/_0_ , \g51952/_0_ , \g51953/_0_ , \g51954/_0_ , \g51955/_0_ , \g51956/_0_ , \g51957/_0_ , \g51958/_0_ , \g51959/_0_ , \g51960/_0_ , \g51961/_0_ , \g51962/_0_ , \g51963/_0_ , \g51964/_0_ , \g51965/_0_ , \g51967/_0_ , \g51968/_0_ , \g51969/_0_ , \g51970/_0_ , \g51971/_0_ , \g51972/_0_ , \g51973/_0_ , \g51974/_0_ , \g51975/_0_ , \g51976/_0_ , \g51977/_0_ , \g51978/_0_ , \g51979/_0_ , \g51980/_0_ , \g51981/_0_ , \g51982/_0_ , \g51983/_0_ , \g51984/_0_ , \g51985/_0_ , \g51986/_0_ , \g51987/_0_ , \g51988/_0_ , \g51989/_0_ , \g51990/_0_ , \g51991/_0_ , \g51992/_0_ , \g51993/_0_ , \g51994/_0_ , \g51995/_0_ , \g51996/_0_ , \g51997/_0_ , \g51998/_0_ , \g51999/_0_ , \g52000/_0_ , \g52001/_0_ , \g52002/_0_ , \g52003/_0_ , \g52004/_0_ , \g52005/_0_ , \g52006/_0_ , \g52007/_0_ , \g52008/_0_ , \g52009/_0_ , \g52010/_0_ , \g52011/_0_ , \g52012/_0_ , \g52013/_0_ , \g52014/_0_ , \g52015/_0_ , \g52016/_0_ , \g52017/_0_ , \g52018/_0_ , \g52019/_0_ , \g52020/_0_ , \g52021/_0_ , \g52022/_0_ , \g52023/_0_ , \g52024/_0_ , \g52025/_0_ , \g52026/_0_ , \g52027/_0_ , \g52028/_0_ , \g52029/_0_ , \g52030/_0_ , \g52031/_0_ , \g52032/_0_ , \g52033/_0_ , \g52034/_0_ , \g52035/_0_ , \g52036/_0_ , \g52037/_0_ , \g52038/_0_ , \g52039/_0_ , \g52040/_0_ , \g52041/_0_ , \g52042/_0_ , \g52043/_0_ , \g52044/_0_ , \g52045/_0_ , \g52046/_0_ , \g52047/_0_ , \g52049/_0_ , \g52050/_0_ , \g52051/_0_ , \g52052/_0_ , \g52053/_0_ , \g52054/_0_ , \g52055/_0_ , \g52056/_0_ , \g52057/_0_ , \g52058/_0_ , \g52061/_0_ , \g52065/_0_ , \g52066/_0_ , \g52067/_0_ , \g52068/_0_ , \g52069/_0_ , \g52070/_0_ , \g52071/_0_ , \g52073/_0_ , \g52074/_0_ , \g52075/_0_ , \g52082/_0_ , \g52083/_0_ , \g52158/_0_ , \g52201/_0_ , \g52202/_0_ , \g52346/_0_ , \g52351/_0_ , \g52390/_0_ , \g52847/_0_ , \g52854/_0_ , \g52968/_0_ , \g52969/_0_ , \g52970/_0_ , \g52971/_0_ , \g52984/_0_ , \g52994/_0_ , \g53019/_0_ , \g53030/_0_ , \g53094/_1_ , \g53106/_0_ , \g53150/_0_ , \g53256/_0_ , \g53297/_0_ , \g53345/_0_ , \g53359/_0_ , \g53375/_0_ , \g53474/_1__syn_2 , \g53475/_2_ , \g53593/_0_ , \g53643/_1_ , \g53655/_0_ , \g53710/_0_ , \g53786/_0_ , \g53837/_0_ , \g53888/_1_ , \g53909/_0_ , \g54253/_2_ , \g54394/_3_ , \g54413/_0_ , \g55420/_0_ , \g55587/_0_ , \g55852/_0_ , \g57020/_0_ , \g59450/_0_ , \g59488/_2_ , \g59752/_0_ , \g59786/_0_ , \g59854/_0_ , \g59878/_0_ , \g59902/_0_ , \g59924/_0_ , \g59947/_0_ , \g59972/_0_ , \g59996/_0_ , \g60017/_0_ , \g60040/_0_ , \g60064/_0_ , \g60095/_0_ , \g60119/_0_ , \g60145/_1_ , \g60165/_0_ , \g60407/_2_ , \g60408/_0_ , \g60613/_2_ , \g60649/_0_ , \g60771/_0_ , \g60908/_1_ , \g60911/_0_ , \g60977/_0_ , \g61/_0_ , \g61002/_0_ , \g61308/_0_ , \g61312/_1_ , \g61314/_0_ , \g61319/_1_ , \g61342/_1_ , \g61360/_0_ , \g61377/_0_ , \g61423/_1_ , \g61426/_0_ , \g61479/_1_ , \g61523/_1_ , \g61558/_1_ , \g61652/_0_ , \g61866/_0_ , \g61868/_1_ , \g61887/_0_ , \u7_mc_dqm_r_reg[0]/P0001_reg_syn_3 , \u7_mc_dqm_r_reg[1]/P0001_reg_syn_3 , \u7_mc_dqm_r_reg[2]/P0001_reg_syn_3 , \u7_mc_dqm_r_reg[3]/P0001_reg_syn_3 , \u7_mc_we__reg/_05_ );
	input mc_cke_pad_o__pad ;
	input mc_vpen_pad_o_pad ;
	input \mem_ack_r_reg/P0001  ;
	input \poc_o[0]_pad  ;
	input \poc_o[10]_pad  ;
	input \poc_o[11]_pad  ;
	input \poc_o[12]_pad  ;
	input \poc_o[13]_pad  ;
	input \poc_o[14]_pad  ;
	input \poc_o[15]_pad  ;
	input \poc_o[16]_pad  ;
	input \poc_o[17]_pad  ;
	input \poc_o[18]_pad  ;
	input \poc_o[19]_pad  ;
	input \poc_o[1]_pad  ;
	input \poc_o[20]_pad  ;
	input \poc_o[21]_pad  ;
	input \poc_o[22]_pad  ;
	input \poc_o[23]_pad  ;
	input \poc_o[24]_pad  ;
	input \poc_o[25]_pad  ;
	input \poc_o[26]_pad  ;
	input \poc_o[27]_pad  ;
	input \poc_o[28]_pad  ;
	input \poc_o[29]_pad  ;
	input \poc_o[2]_pad  ;
	input \poc_o[30]_pad  ;
	input \poc_o[31]_pad  ;
	input \poc_o[3]_pad  ;
	input \poc_o[4]_pad  ;
	input \poc_o[5]_pad  ;
	input \poc_o[6]_pad  ;
	input \poc_o[7]_pad  ;
	input \poc_o[8]_pad  ;
	input \poc_o[9]_pad  ;
	input suspended_o_pad ;
	input \u0_cs_reg[0]/NET0131  ;
	input \u0_cs_reg[1]/NET0131  ;
	input \u0_csc_mask_r_reg[0]/NET0131  ;
	input \u0_csc_mask_r_reg[10]/NET0131  ;
	input \u0_csc_mask_r_reg[1]/NET0131  ;
	input \u0_csc_mask_r_reg[2]/NET0131  ;
	input \u0_csc_mask_r_reg[3]/NET0131  ;
	input \u0_csc_mask_r_reg[4]/NET0131  ;
	input \u0_csc_mask_r_reg[5]/NET0131  ;
	input \u0_csc_mask_r_reg[6]/NET0131  ;
	input \u0_csc_mask_r_reg[7]/NET0131  ;
	input \u0_csc_mask_r_reg[8]/NET0131  ;
	input \u0_csc_mask_r_reg[9]/NET0131  ;
	input \u0_csc_reg[10]/NET0131  ;
	input \u0_csc_reg[11]/NET0131  ;
	input \u0_csc_reg[1]/NET0131  ;
	input \u0_csc_reg[2]/NET0131  ;
	input \u0_csc_reg[3]/NET0131  ;
	input \u0_csc_reg[4]/NET0131  ;
	input \u0_csc_reg[5]/NET0131  ;
	input \u0_csc_reg[6]/NET0131  ;
	input \u0_csc_reg[7]/NET0131  ;
	input \u0_csc_reg[9]/NET0131  ;
	input \u0_csr_r2_reg[0]/NET0131  ;
	input \u0_csr_r2_reg[1]/NET0131  ;
	input \u0_csr_r2_reg[2]/NET0131  ;
	input \u0_csr_r2_reg[3]/NET0131  ;
	input \u0_csr_r2_reg[4]/NET0131  ;
	input \u0_csr_r2_reg[5]/NET0131  ;
	input \u0_csr_r2_reg[6]/NET0131  ;
	input \u0_csr_r2_reg[7]/NET0131  ;
	input \u0_csr_r_reg[0]/P0001  ;
	input \u0_csr_r_reg[10]/NET0131  ;
	input \u0_csr_r_reg[2]/NET0131  ;
	input \u0_csr_r_reg[3]/NET0131  ;
	input \u0_csr_r_reg[4]/NET0131  ;
	input \u0_csr_r_reg[5]/NET0131  ;
	input \u0_csr_r_reg[6]/NET0131  ;
	input \u0_csr_r_reg[7]/NET0131  ;
	input \u0_csr_r_reg[8]/NET0131  ;
	input \u0_csr_r_reg[9]/NET0131  ;
	input \u0_init_ack_r_reg/P0001  ;
	input \u0_init_req_reg/NET0131  ;
	input \u0_lmr_ack_r_reg/P0001  ;
	input \u0_lmr_req_reg/NET0131  ;
	input \u0_rf_we_reg/NET0131  ;
	input \u0_rst_r2_reg/NET0131  ;
	input \u0_sp_csc_reg[10]/NET0131  ;
	input \u0_sp_csc_reg[1]/NET0131  ;
	input \u0_sp_csc_reg[2]/NET0131  ;
	input \u0_sp_csc_reg[3]/NET0131  ;
	input \u0_sp_csc_reg[4]/NET0131  ;
	input \u0_sp_csc_reg[5]/NET0131  ;
	input \u0_sp_csc_reg[6]/NET0131  ;
	input \u0_sp_csc_reg[7]/NET0131  ;
	input \u0_sp_csc_reg[9]/NET0131  ;
	input \u0_sp_tms_reg[0]/NET0131  ;
	input \u0_sp_tms_reg[10]/NET0131  ;
	input \u0_sp_tms_reg[11]/NET0131  ;
	input \u0_sp_tms_reg[12]/NET0131  ;
	input \u0_sp_tms_reg[13]/NET0131  ;
	input \u0_sp_tms_reg[14]/NET0131  ;
	input \u0_sp_tms_reg[15]/NET0131  ;
	input \u0_sp_tms_reg[16]/NET0131  ;
	input \u0_sp_tms_reg[17]/NET0131  ;
	input \u0_sp_tms_reg[18]/NET0131  ;
	input \u0_sp_tms_reg[19]/NET0131  ;
	input \u0_sp_tms_reg[1]/NET0131  ;
	input \u0_sp_tms_reg[20]/NET0131  ;
	input \u0_sp_tms_reg[21]/NET0131  ;
	input \u0_sp_tms_reg[22]/NET0131  ;
	input \u0_sp_tms_reg[23]/NET0131  ;
	input \u0_sp_tms_reg[24]/NET0131  ;
	input \u0_sp_tms_reg[25]/NET0131  ;
	input \u0_sp_tms_reg[26]/NET0131  ;
	input \u0_sp_tms_reg[27]/NET0131  ;
	input \u0_sp_tms_reg[2]/NET0131  ;
	input \u0_sp_tms_reg[3]/NET0131  ;
	input \u0_sp_tms_reg[4]/NET0131  ;
	input \u0_sp_tms_reg[5]/NET0131  ;
	input \u0_sp_tms_reg[6]/NET0131  ;
	input \u0_sp_tms_reg[7]/NET0131  ;
	input \u0_sp_tms_reg[8]/NET0131  ;
	input \u0_sp_tms_reg[9]/NET0131  ;
	input \u0_spec_req_cs_reg[0]/NET0131  ;
	input \u0_spec_req_cs_reg[1]/NET0131  ;
	input \u0_sreq_cs_le_reg/NET0131  ;
	input \u0_tms_reg[0]/NET0131  ;
	input \u0_tms_reg[10]/NET0131  ;
	input \u0_tms_reg[11]/NET0131  ;
	input \u0_tms_reg[12]/NET0131  ;
	input \u0_tms_reg[13]/NET0131  ;
	input \u0_tms_reg[14]/NET0131  ;
	input \u0_tms_reg[15]/NET0131  ;
	input \u0_tms_reg[16]/NET0131  ;
	input \u0_tms_reg[17]/NET0131  ;
	input \u0_tms_reg[18]/NET0131  ;
	input \u0_tms_reg[19]/NET0131  ;
	input \u0_tms_reg[1]/NET0131  ;
	input \u0_tms_reg[20]/NET0131  ;
	input \u0_tms_reg[21]/NET0131  ;
	input \u0_tms_reg[22]/NET0131  ;
	input \u0_tms_reg[23]/NET0131  ;
	input \u0_tms_reg[24]/NET0131  ;
	input \u0_tms_reg[25]/NET0131  ;
	input \u0_tms_reg[26]/NET0131  ;
	input \u0_tms_reg[27]/NET0131  ;
	input \u0_tms_reg[2]/NET0131  ;
	input \u0_tms_reg[3]/NET0131  ;
	input \u0_tms_reg[4]/NET0131  ;
	input \u0_tms_reg[5]/NET0131  ;
	input \u0_tms_reg[6]/NET0131  ;
	input \u0_tms_reg[7]/NET0131  ;
	input \u0_tms_reg[8]/NET0131  ;
	input \u0_tms_reg[9]/NET0131  ;
	input \u0_u0_addr_r_reg[2]/P0001  ;
	input \u0_u0_addr_r_reg[3]/P0001  ;
	input \u0_u0_addr_r_reg[4]/P0001  ;
	input \u0_u0_addr_r_reg[5]/P0001  ;
	input \u0_u0_addr_r_reg[6]/P0001  ;
	input \u0_u0_csc_reg[0]/NET0131  ;
	input \u0_u0_csc_reg[10]/P0001  ;
	input \u0_u0_csc_reg[11]/P0001  ;
	input \u0_u0_csc_reg[12]/P0001  ;
	input \u0_u0_csc_reg[13]/P0001  ;
	input \u0_u0_csc_reg[14]/P0001  ;
	input \u0_u0_csc_reg[15]/P0001  ;
	input \u0_u0_csc_reg[16]/P0001  ;
	input \u0_u0_csc_reg[17]/P0001  ;
	input \u0_u0_csc_reg[18]/P0001  ;
	input \u0_u0_csc_reg[19]/P0001  ;
	input \u0_u0_csc_reg[1]/NET0131  ;
	input \u0_u0_csc_reg[20]/P0001  ;
	input \u0_u0_csc_reg[21]/P0001  ;
	input \u0_u0_csc_reg[22]/P0001  ;
	input \u0_u0_csc_reg[23]/P0001  ;
	input \u0_u0_csc_reg[24]/P0001  ;
	input \u0_u0_csc_reg[25]/P0001  ;
	input \u0_u0_csc_reg[26]/P0001  ;
	input \u0_u0_csc_reg[27]/P0001  ;
	input \u0_u0_csc_reg[28]/P0001  ;
	input \u0_u0_csc_reg[29]/P0001  ;
	input \u0_u0_csc_reg[2]/NET0131  ;
	input \u0_u0_csc_reg[30]/P0001  ;
	input \u0_u0_csc_reg[31]/P0001  ;
	input \u0_u0_csc_reg[3]/NET0131  ;
	input \u0_u0_csc_reg[4]/P0001  ;
	input \u0_u0_csc_reg[5]/P0001  ;
	input \u0_u0_csc_reg[6]/P0001  ;
	input \u0_u0_csc_reg[7]/P0001  ;
	input \u0_u0_csc_reg[8]/P0001  ;
	input \u0_u0_csc_reg[9]/P0001  ;
	input \u0_u0_init_req_reg/NET0131  ;
	input \u0_u0_init_req_we_reg/NET0131  ;
	input \u0_u0_inited_reg/NET0131  ;
	input \u0_u0_lmr_req_reg/NET0131  ;
	input \u0_u0_lmr_req_we_reg/NET0131  ;
	input \u0_u0_tms_reg[0]/P0001  ;
	input \u0_u0_tms_reg[10]/P0001  ;
	input \u0_u0_tms_reg[11]/P0001  ;
	input \u0_u0_tms_reg[12]/P0001  ;
	input \u0_u0_tms_reg[13]/P0001  ;
	input \u0_u0_tms_reg[14]/P0001  ;
	input \u0_u0_tms_reg[15]/P0001  ;
	input \u0_u0_tms_reg[16]/P0001  ;
	input \u0_u0_tms_reg[17]/P0001  ;
	input \u0_u0_tms_reg[18]/P0001  ;
	input \u0_u0_tms_reg[19]/P0001  ;
	input \u0_u0_tms_reg[1]/P0001  ;
	input \u0_u0_tms_reg[20]/P0001  ;
	input \u0_u0_tms_reg[21]/P0001  ;
	input \u0_u0_tms_reg[22]/P0001  ;
	input \u0_u0_tms_reg[23]/P0001  ;
	input \u0_u0_tms_reg[24]/P0001  ;
	input \u0_u0_tms_reg[25]/P0001  ;
	input \u0_u0_tms_reg[26]/P0001  ;
	input \u0_u0_tms_reg[27]/P0001  ;
	input \u0_u0_tms_reg[28]/P0001  ;
	input \u0_u0_tms_reg[29]/P0001  ;
	input \u0_u0_tms_reg[2]/P0001  ;
	input \u0_u0_tms_reg[30]/P0001  ;
	input \u0_u0_tms_reg[31]/P0001  ;
	input \u0_u0_tms_reg[3]/P0001  ;
	input \u0_u0_tms_reg[4]/P0001  ;
	input \u0_u0_tms_reg[5]/P0001  ;
	input \u0_u0_tms_reg[6]/P0001  ;
	input \u0_u0_tms_reg[7]/P0001  ;
	input \u0_u0_tms_reg[8]/P0001  ;
	input \u0_u0_tms_reg[9]/P0001  ;
	input \u0_u1_csc_reg[0]/NET0131  ;
	input \u0_u1_csc_reg[10]/P0001  ;
	input \u0_u1_csc_reg[11]/P0001  ;
	input \u0_u1_csc_reg[12]/P0001  ;
	input \u0_u1_csc_reg[13]/P0001  ;
	input \u0_u1_csc_reg[14]/P0001  ;
	input \u0_u1_csc_reg[15]/P0001  ;
	input \u0_u1_csc_reg[16]/P0001  ;
	input \u0_u1_csc_reg[17]/P0001  ;
	input \u0_u1_csc_reg[18]/P0001  ;
	input \u0_u1_csc_reg[19]/P0001  ;
	input \u0_u1_csc_reg[1]/NET0131  ;
	input \u0_u1_csc_reg[20]/P0001  ;
	input \u0_u1_csc_reg[21]/P0001  ;
	input \u0_u1_csc_reg[22]/P0001  ;
	input \u0_u1_csc_reg[23]/P0001  ;
	input \u0_u1_csc_reg[24]/P0001  ;
	input \u0_u1_csc_reg[25]/P0001  ;
	input \u0_u1_csc_reg[26]/P0001  ;
	input \u0_u1_csc_reg[27]/P0001  ;
	input \u0_u1_csc_reg[28]/P0001  ;
	input \u0_u1_csc_reg[29]/P0001  ;
	input \u0_u1_csc_reg[2]/NET0131  ;
	input \u0_u1_csc_reg[30]/P0001  ;
	input \u0_u1_csc_reg[31]/P0001  ;
	input \u0_u1_csc_reg[3]/NET0131  ;
	input \u0_u1_csc_reg[4]/P0001  ;
	input \u0_u1_csc_reg[5]/P0001  ;
	input \u0_u1_csc_reg[6]/P0001  ;
	input \u0_u1_csc_reg[7]/P0001  ;
	input \u0_u1_csc_reg[8]/P0001  ;
	input \u0_u1_csc_reg[9]/P0001  ;
	input \u0_u1_init_req_reg/NET0131  ;
	input \u0_u1_init_req_we_reg/NET0131  ;
	input \u0_u1_inited_reg/NET0131  ;
	input \u0_u1_lmr_req_reg/NET0131  ;
	input \u0_u1_lmr_req_we_reg/NET0131  ;
	input \u0_u1_tms_reg[0]/P0001  ;
	input \u0_u1_tms_reg[10]/P0001  ;
	input \u0_u1_tms_reg[11]/P0001  ;
	input \u0_u1_tms_reg[12]/P0001  ;
	input \u0_u1_tms_reg[13]/P0001  ;
	input \u0_u1_tms_reg[14]/P0001  ;
	input \u0_u1_tms_reg[15]/P0001  ;
	input \u0_u1_tms_reg[16]/P0001  ;
	input \u0_u1_tms_reg[17]/P0001  ;
	input \u0_u1_tms_reg[18]/P0001  ;
	input \u0_u1_tms_reg[19]/P0001  ;
	input \u0_u1_tms_reg[1]/P0001  ;
	input \u0_u1_tms_reg[20]/P0001  ;
	input \u0_u1_tms_reg[21]/P0001  ;
	input \u0_u1_tms_reg[22]/P0001  ;
	input \u0_u1_tms_reg[23]/P0001  ;
	input \u0_u1_tms_reg[24]/P0001  ;
	input \u0_u1_tms_reg[25]/P0001  ;
	input \u0_u1_tms_reg[26]/P0001  ;
	input \u0_u1_tms_reg[27]/P0001  ;
	input \u0_u1_tms_reg[28]/P0001  ;
	input \u0_u1_tms_reg[29]/P0001  ;
	input \u0_u1_tms_reg[2]/P0001  ;
	input \u0_u1_tms_reg[30]/P0001  ;
	input \u0_u1_tms_reg[31]/P0001  ;
	input \u0_u1_tms_reg[3]/P0001  ;
	input \u0_u1_tms_reg[4]/P0001  ;
	input \u0_u1_tms_reg[5]/P0001  ;
	input \u0_u1_tms_reg[6]/P0001  ;
	input \u0_u1_tms_reg[7]/P0001  ;
	input \u0_u1_tms_reg[8]/P0001  ;
	input \u0_u1_tms_reg[9]/P0001  ;
	input \u0_wp_err_reg/NET0131  ;
	input \u1_acs_addr_reg[0]/P0001  ;
	input \u1_acs_addr_reg[10]/P0001  ;
	input \u1_acs_addr_reg[11]/P0001  ;
	input \u1_acs_addr_reg[12]/P0001  ;
	input \u1_acs_addr_reg[13]/P0001  ;
	input \u1_acs_addr_reg[14]/P0001  ;
	input \u1_acs_addr_reg[15]/P0001  ;
	input \u1_acs_addr_reg[16]/P0001  ;
	input \u1_acs_addr_reg[17]/P0001  ;
	input \u1_acs_addr_reg[18]/P0001  ;
	input \u1_acs_addr_reg[19]/P0001  ;
	input \u1_acs_addr_reg[1]/P0001  ;
	input \u1_acs_addr_reg[20]/P0001  ;
	input \u1_acs_addr_reg[21]/P0001  ;
	input \u1_acs_addr_reg[22]/P0001  ;
	input \u1_acs_addr_reg[23]/P0001  ;
	input \u1_acs_addr_reg[2]/P0001  ;
	input \u1_acs_addr_reg[3]/P0001  ;
	input \u1_acs_addr_reg[4]/P0001  ;
	input \u1_acs_addr_reg[5]/P0001  ;
	input \u1_acs_addr_reg[6]/P0001  ;
	input \u1_acs_addr_reg[7]/P0001  ;
	input \u1_acs_addr_reg[8]/P0001  ;
	input \u1_acs_addr_reg[9]/P0001  ;
	input \u1_bank_adr_reg[0]/P0001  ;
	input \u1_bank_adr_reg[1]/P0001  ;
	input \u1_col_adr_reg[0]/P0001  ;
	input \u1_col_adr_reg[1]/P0001  ;
	input \u1_col_adr_reg[2]/P0001  ;
	input \u1_col_adr_reg[3]/P0001  ;
	input \u1_col_adr_reg[4]/P0001  ;
	input \u1_col_adr_reg[5]/P0001  ;
	input \u1_col_adr_reg[6]/P0001  ;
	input \u1_col_adr_reg[7]/P0001  ;
	input \u1_col_adr_reg[8]/P0001  ;
	input \u1_col_adr_reg[9]/P0001  ;
	input \u1_row_adr_reg[0]/P0001  ;
	input \u1_row_adr_reg[10]/P0001  ;
	input \u1_row_adr_reg[11]/P0001  ;
	input \u1_row_adr_reg[12]/P0001  ;
	input \u1_row_adr_reg[1]/P0001  ;
	input \u1_row_adr_reg[2]/P0001  ;
	input \u1_row_adr_reg[3]/P0001  ;
	input \u1_row_adr_reg[4]/P0001  ;
	input \u1_row_adr_reg[5]/P0001  ;
	input \u1_row_adr_reg[6]/P0001  ;
	input \u1_row_adr_reg[7]/P0001  ;
	input \u1_row_adr_reg[8]/P0001  ;
	input \u1_row_adr_reg[9]/P0001  ;
	input \u1_sram_addr_reg[0]/P0001  ;
	input \u1_sram_addr_reg[10]/P0001  ;
	input \u1_sram_addr_reg[11]/P0001  ;
	input \u1_sram_addr_reg[12]/P0001  ;
	input \u1_sram_addr_reg[13]/P0001  ;
	input \u1_sram_addr_reg[14]/P0001  ;
	input \u1_sram_addr_reg[15]/P0001  ;
	input \u1_sram_addr_reg[16]/P0001  ;
	input \u1_sram_addr_reg[17]/P0001  ;
	input \u1_sram_addr_reg[18]/P0001  ;
	input \u1_sram_addr_reg[19]/P0001  ;
	input \u1_sram_addr_reg[1]/P0001  ;
	input \u1_sram_addr_reg[20]/P0001  ;
	input \u1_sram_addr_reg[21]/P0001  ;
	input \u1_sram_addr_reg[22]/P0001  ;
	input \u1_sram_addr_reg[23]/P0001  ;
	input \u1_sram_addr_reg[2]/P0001  ;
	input \u1_sram_addr_reg[3]/P0001  ;
	input \u1_sram_addr_reg[4]/P0001  ;
	input \u1_sram_addr_reg[5]/P0001  ;
	input \u1_sram_addr_reg[6]/P0001  ;
	input \u1_sram_addr_reg[7]/P0001  ;
	input \u1_sram_addr_reg[8]/P0001  ;
	input \u1_sram_addr_reg[9]/P0001  ;
	input \u1_u0_out_r_reg[0]/P0001  ;
	input \u1_u0_out_r_reg[10]/P0001  ;
	input \u1_u0_out_r_reg[11]/P0001  ;
	input \u1_u0_out_r_reg[12]/P0001  ;
	input \u1_u0_out_r_reg[1]/P0001  ;
	input \u1_u0_out_r_reg[2]/P0001  ;
	input \u1_u0_out_r_reg[3]/P0001  ;
	input \u1_u0_out_r_reg[4]/P0001  ;
	input \u1_u0_out_r_reg[5]/P0001  ;
	input \u1_u0_out_r_reg[6]/P0001  ;
	input \u1_u0_out_r_reg[7]/P0001  ;
	input \u1_u0_out_r_reg[8]/P0001  ;
	input \u1_u0_out_r_reg[9]/P0001  ;
	input \u2_bank_open_reg/P0001  ;
	input \u2_row_same_reg/P0001  ;
	input \u2_u0_b0_last_row_reg[0]/P0001  ;
	input \u2_u0_b0_last_row_reg[10]/P0001  ;
	input \u2_u0_b0_last_row_reg[11]/P0001  ;
	input \u2_u0_b0_last_row_reg[12]/P0001  ;
	input \u2_u0_b0_last_row_reg[1]/P0001  ;
	input \u2_u0_b0_last_row_reg[2]/P0001  ;
	input \u2_u0_b0_last_row_reg[3]/P0001  ;
	input \u2_u0_b0_last_row_reg[4]/P0001  ;
	input \u2_u0_b0_last_row_reg[5]/P0001  ;
	input \u2_u0_b0_last_row_reg[6]/P0001  ;
	input \u2_u0_b0_last_row_reg[7]/P0001  ;
	input \u2_u0_b0_last_row_reg[8]/P0001  ;
	input \u2_u0_b0_last_row_reg[9]/P0001  ;
	input \u2_u0_b1_last_row_reg[0]/P0001  ;
	input \u2_u0_b1_last_row_reg[10]/P0001  ;
	input \u2_u0_b1_last_row_reg[11]/P0001  ;
	input \u2_u0_b1_last_row_reg[12]/P0001  ;
	input \u2_u0_b1_last_row_reg[1]/P0001  ;
	input \u2_u0_b1_last_row_reg[2]/P0001  ;
	input \u2_u0_b1_last_row_reg[3]/P0001  ;
	input \u2_u0_b1_last_row_reg[4]/P0001  ;
	input \u2_u0_b1_last_row_reg[5]/P0001  ;
	input \u2_u0_b1_last_row_reg[6]/P0001  ;
	input \u2_u0_b1_last_row_reg[7]/P0001  ;
	input \u2_u0_b1_last_row_reg[8]/P0001  ;
	input \u2_u0_b1_last_row_reg[9]/P0001  ;
	input \u2_u0_b2_last_row_reg[0]/P0001  ;
	input \u2_u0_b2_last_row_reg[10]/P0001  ;
	input \u2_u0_b2_last_row_reg[11]/P0001  ;
	input \u2_u0_b2_last_row_reg[12]/P0001  ;
	input \u2_u0_b2_last_row_reg[1]/P0001  ;
	input \u2_u0_b2_last_row_reg[2]/P0001  ;
	input \u2_u0_b2_last_row_reg[3]/P0001  ;
	input \u2_u0_b2_last_row_reg[4]/P0001  ;
	input \u2_u0_b2_last_row_reg[5]/P0001  ;
	input \u2_u0_b2_last_row_reg[6]/P0001  ;
	input \u2_u0_b2_last_row_reg[7]/P0001  ;
	input \u2_u0_b2_last_row_reg[8]/P0001  ;
	input \u2_u0_b2_last_row_reg[9]/P0001  ;
	input \u2_u0_b3_last_row_reg[0]/P0001  ;
	input \u2_u0_b3_last_row_reg[10]/P0001  ;
	input \u2_u0_b3_last_row_reg[11]/P0001  ;
	input \u2_u0_b3_last_row_reg[12]/P0001  ;
	input \u2_u0_b3_last_row_reg[1]/P0001  ;
	input \u2_u0_b3_last_row_reg[2]/P0001  ;
	input \u2_u0_b3_last_row_reg[3]/P0001  ;
	input \u2_u0_b3_last_row_reg[4]/P0001  ;
	input \u2_u0_b3_last_row_reg[5]/P0001  ;
	input \u2_u0_b3_last_row_reg[6]/P0001  ;
	input \u2_u0_b3_last_row_reg[7]/P0001  ;
	input \u2_u0_b3_last_row_reg[8]/P0001  ;
	input \u2_u0_b3_last_row_reg[9]/P0001  ;
	input \u2_u0_bank0_open_reg/NET0131  ;
	input \u2_u0_bank1_open_reg/NET0131  ;
	input \u2_u0_bank2_open_reg/NET0131  ;
	input \u2_u0_bank3_open_reg/NET0131  ;
	input \u2_u1_b0_last_row_reg[0]/P0001  ;
	input \u2_u1_b0_last_row_reg[10]/P0001  ;
	input \u2_u1_b0_last_row_reg[11]/P0001  ;
	input \u2_u1_b0_last_row_reg[12]/P0001  ;
	input \u2_u1_b0_last_row_reg[1]/P0001  ;
	input \u2_u1_b0_last_row_reg[2]/P0001  ;
	input \u2_u1_b0_last_row_reg[3]/P0001  ;
	input \u2_u1_b0_last_row_reg[4]/P0001  ;
	input \u2_u1_b0_last_row_reg[5]/P0001  ;
	input \u2_u1_b0_last_row_reg[6]/P0001  ;
	input \u2_u1_b0_last_row_reg[7]/P0001  ;
	input \u2_u1_b0_last_row_reg[8]/P0001  ;
	input \u2_u1_b0_last_row_reg[9]/P0001  ;
	input \u2_u1_b1_last_row_reg[0]/P0001  ;
	input \u2_u1_b1_last_row_reg[10]/P0001  ;
	input \u2_u1_b1_last_row_reg[11]/P0001  ;
	input \u2_u1_b1_last_row_reg[12]/P0001  ;
	input \u2_u1_b1_last_row_reg[1]/P0001  ;
	input \u2_u1_b1_last_row_reg[2]/P0001  ;
	input \u2_u1_b1_last_row_reg[3]/P0001  ;
	input \u2_u1_b1_last_row_reg[4]/P0001  ;
	input \u2_u1_b1_last_row_reg[5]/P0001  ;
	input \u2_u1_b1_last_row_reg[6]/P0001  ;
	input \u2_u1_b1_last_row_reg[7]/P0001  ;
	input \u2_u1_b1_last_row_reg[8]/P0001  ;
	input \u2_u1_b1_last_row_reg[9]/P0001  ;
	input \u2_u1_b2_last_row_reg[0]/P0001  ;
	input \u2_u1_b2_last_row_reg[10]/P0001  ;
	input \u2_u1_b2_last_row_reg[11]/P0001  ;
	input \u2_u1_b2_last_row_reg[12]/P0001  ;
	input \u2_u1_b2_last_row_reg[1]/P0001  ;
	input \u2_u1_b2_last_row_reg[2]/P0001  ;
	input \u2_u1_b2_last_row_reg[3]/P0001  ;
	input \u2_u1_b2_last_row_reg[4]/P0001  ;
	input \u2_u1_b2_last_row_reg[5]/P0001  ;
	input \u2_u1_b2_last_row_reg[6]/P0001  ;
	input \u2_u1_b2_last_row_reg[7]/P0001  ;
	input \u2_u1_b2_last_row_reg[8]/P0001  ;
	input \u2_u1_b2_last_row_reg[9]/P0001  ;
	input \u2_u1_b3_last_row_reg[0]/P0001  ;
	input \u2_u1_b3_last_row_reg[10]/P0001  ;
	input \u2_u1_b3_last_row_reg[11]/P0001  ;
	input \u2_u1_b3_last_row_reg[12]/P0001  ;
	input \u2_u1_b3_last_row_reg[1]/P0001  ;
	input \u2_u1_b3_last_row_reg[2]/P0001  ;
	input \u2_u1_b3_last_row_reg[3]/P0001  ;
	input \u2_u1_b3_last_row_reg[4]/P0001  ;
	input \u2_u1_b3_last_row_reg[5]/P0001  ;
	input \u2_u1_b3_last_row_reg[6]/P0001  ;
	input \u2_u1_b3_last_row_reg[7]/P0001  ;
	input \u2_u1_b3_last_row_reg[8]/P0001  ;
	input \u2_u1_b3_last_row_reg[9]/P0001  ;
	input \u2_u1_bank0_open_reg/NET0131  ;
	input \u2_u1_bank1_open_reg/NET0131  ;
	input \u2_u1_bank2_open_reg/NET0131  ;
	input \u2_u1_bank3_open_reg/NET0131  ;
	input \u3_byte0_reg[0]/P0001  ;
	input \u3_byte0_reg[1]/P0001  ;
	input \u3_byte0_reg[2]/P0001  ;
	input \u3_byte0_reg[3]/P0001  ;
	input \u3_byte0_reg[4]/P0001  ;
	input \u3_byte0_reg[5]/P0001  ;
	input \u3_byte0_reg[6]/P0001  ;
	input \u3_byte0_reg[7]/P0001  ;
	input \u3_byte1_reg[0]/P0001  ;
	input \u3_byte1_reg[1]/P0001  ;
	input \u3_byte1_reg[2]/P0001  ;
	input \u3_byte1_reg[3]/P0001  ;
	input \u3_byte1_reg[4]/P0001  ;
	input \u3_byte1_reg[5]/P0001  ;
	input \u3_byte1_reg[6]/P0001  ;
	input \u3_byte1_reg[7]/P0001  ;
	input \u3_byte2_reg[0]/P0001  ;
	input \u3_byte2_reg[1]/P0001  ;
	input \u3_byte2_reg[2]/P0001  ;
	input \u3_byte2_reg[3]/P0001  ;
	input \u3_byte2_reg[4]/P0001  ;
	input \u3_byte2_reg[5]/P0001  ;
	input \u3_byte2_reg[6]/P0001  ;
	input \u3_byte2_reg[7]/P0001  ;
	input \u3_u0_r0_reg[0]/P0001  ;
	input \u3_u0_r0_reg[10]/P0001  ;
	input \u3_u0_r0_reg[11]/P0001  ;
	input \u3_u0_r0_reg[12]/P0001  ;
	input \u3_u0_r0_reg[13]/P0001  ;
	input \u3_u0_r0_reg[14]/P0001  ;
	input \u3_u0_r0_reg[15]/P0001  ;
	input \u3_u0_r0_reg[16]/P0001  ;
	input \u3_u0_r0_reg[17]/P0001  ;
	input \u3_u0_r0_reg[18]/P0001  ;
	input \u3_u0_r0_reg[19]/P0001  ;
	input \u3_u0_r0_reg[1]/P0001  ;
	input \u3_u0_r0_reg[20]/P0001  ;
	input \u3_u0_r0_reg[21]/P0001  ;
	input \u3_u0_r0_reg[22]/P0001  ;
	input \u3_u0_r0_reg[23]/P0001  ;
	input \u3_u0_r0_reg[24]/P0001  ;
	input \u3_u0_r0_reg[25]/P0001  ;
	input \u3_u0_r0_reg[26]/P0001  ;
	input \u3_u0_r0_reg[27]/P0001  ;
	input \u3_u0_r0_reg[28]/P0001  ;
	input \u3_u0_r0_reg[29]/P0001  ;
	input \u3_u0_r0_reg[2]/P0001  ;
	input \u3_u0_r0_reg[30]/P0001  ;
	input \u3_u0_r0_reg[31]/P0001  ;
	input \u3_u0_r0_reg[32]/P0001  ;
	input \u3_u0_r0_reg[33]/P0001  ;
	input \u3_u0_r0_reg[34]/P0001  ;
	input \u3_u0_r0_reg[35]/P0001  ;
	input \u3_u0_r0_reg[3]/P0001  ;
	input \u3_u0_r0_reg[4]/P0001  ;
	input \u3_u0_r0_reg[5]/P0001  ;
	input \u3_u0_r0_reg[6]/P0001  ;
	input \u3_u0_r0_reg[7]/P0001  ;
	input \u3_u0_r0_reg[8]/P0001  ;
	input \u3_u0_r0_reg[9]/P0001  ;
	input \u3_u0_r1_reg[0]/P0001  ;
	input \u3_u0_r1_reg[10]/P0001  ;
	input \u3_u0_r1_reg[11]/P0001  ;
	input \u3_u0_r1_reg[12]/P0001  ;
	input \u3_u0_r1_reg[13]/P0001  ;
	input \u3_u0_r1_reg[14]/P0001  ;
	input \u3_u0_r1_reg[15]/P0001  ;
	input \u3_u0_r1_reg[16]/P0001  ;
	input \u3_u0_r1_reg[17]/P0001  ;
	input \u3_u0_r1_reg[18]/P0001  ;
	input \u3_u0_r1_reg[19]/P0001  ;
	input \u3_u0_r1_reg[1]/P0001  ;
	input \u3_u0_r1_reg[20]/P0001  ;
	input \u3_u0_r1_reg[21]/P0001  ;
	input \u3_u0_r1_reg[22]/P0001  ;
	input \u3_u0_r1_reg[23]/P0001  ;
	input \u3_u0_r1_reg[24]/P0001  ;
	input \u3_u0_r1_reg[25]/P0001  ;
	input \u3_u0_r1_reg[26]/P0001  ;
	input \u3_u0_r1_reg[27]/P0001  ;
	input \u3_u0_r1_reg[28]/P0001  ;
	input \u3_u0_r1_reg[29]/P0001  ;
	input \u3_u0_r1_reg[2]/P0001  ;
	input \u3_u0_r1_reg[30]/P0001  ;
	input \u3_u0_r1_reg[31]/P0001  ;
	input \u3_u0_r1_reg[32]/P0001  ;
	input \u3_u0_r1_reg[33]/P0001  ;
	input \u3_u0_r1_reg[34]/P0001  ;
	input \u3_u0_r1_reg[35]/P0001  ;
	input \u3_u0_r1_reg[3]/P0001  ;
	input \u3_u0_r1_reg[4]/P0001  ;
	input \u3_u0_r1_reg[5]/P0001  ;
	input \u3_u0_r1_reg[6]/P0001  ;
	input \u3_u0_r1_reg[7]/P0001  ;
	input \u3_u0_r1_reg[8]/P0001  ;
	input \u3_u0_r1_reg[9]/P0001  ;
	input \u3_u0_r2_reg[0]/P0001  ;
	input \u3_u0_r2_reg[10]/P0001  ;
	input \u3_u0_r2_reg[11]/P0001  ;
	input \u3_u0_r2_reg[12]/P0001  ;
	input \u3_u0_r2_reg[13]/P0001  ;
	input \u3_u0_r2_reg[14]/P0001  ;
	input \u3_u0_r2_reg[15]/P0001  ;
	input \u3_u0_r2_reg[16]/P0001  ;
	input \u3_u0_r2_reg[17]/P0001  ;
	input \u3_u0_r2_reg[18]/P0001  ;
	input \u3_u0_r2_reg[19]/P0001  ;
	input \u3_u0_r2_reg[1]/P0001  ;
	input \u3_u0_r2_reg[20]/P0001  ;
	input \u3_u0_r2_reg[21]/P0001  ;
	input \u3_u0_r2_reg[22]/P0001  ;
	input \u3_u0_r2_reg[23]/P0001  ;
	input \u3_u0_r2_reg[24]/P0001  ;
	input \u3_u0_r2_reg[25]/P0001  ;
	input \u3_u0_r2_reg[26]/P0001  ;
	input \u3_u0_r2_reg[27]/P0001  ;
	input \u3_u0_r2_reg[28]/P0001  ;
	input \u3_u0_r2_reg[29]/P0001  ;
	input \u3_u0_r2_reg[2]/P0001  ;
	input \u3_u0_r2_reg[30]/P0001  ;
	input \u3_u0_r2_reg[31]/P0001  ;
	input \u3_u0_r2_reg[32]/P0001  ;
	input \u3_u0_r2_reg[33]/P0001  ;
	input \u3_u0_r2_reg[34]/P0001  ;
	input \u3_u0_r2_reg[35]/P0001  ;
	input \u3_u0_r2_reg[3]/P0001  ;
	input \u3_u0_r2_reg[4]/P0001  ;
	input \u3_u0_r2_reg[5]/P0001  ;
	input \u3_u0_r2_reg[6]/P0001  ;
	input \u3_u0_r2_reg[7]/P0001  ;
	input \u3_u0_r2_reg[8]/P0001  ;
	input \u3_u0_r2_reg[9]/P0001  ;
	input \u3_u0_r3_reg[0]/P0001  ;
	input \u3_u0_r3_reg[10]/P0001  ;
	input \u3_u0_r3_reg[11]/P0001  ;
	input \u3_u0_r3_reg[12]/P0001  ;
	input \u3_u0_r3_reg[13]/P0001  ;
	input \u3_u0_r3_reg[14]/P0001  ;
	input \u3_u0_r3_reg[15]/P0001  ;
	input \u3_u0_r3_reg[16]/P0001  ;
	input \u3_u0_r3_reg[17]/P0001  ;
	input \u3_u0_r3_reg[18]/P0001  ;
	input \u3_u0_r3_reg[19]/P0001  ;
	input \u3_u0_r3_reg[1]/P0001  ;
	input \u3_u0_r3_reg[20]/P0001  ;
	input \u3_u0_r3_reg[21]/P0001  ;
	input \u3_u0_r3_reg[22]/P0001  ;
	input \u3_u0_r3_reg[23]/P0001  ;
	input \u3_u0_r3_reg[24]/P0001  ;
	input \u3_u0_r3_reg[25]/P0001  ;
	input \u3_u0_r3_reg[26]/P0001  ;
	input \u3_u0_r3_reg[27]/P0001  ;
	input \u3_u0_r3_reg[28]/P0001  ;
	input \u3_u0_r3_reg[29]/P0001  ;
	input \u3_u0_r3_reg[2]/P0001  ;
	input \u3_u0_r3_reg[30]/P0001  ;
	input \u3_u0_r3_reg[31]/P0001  ;
	input \u3_u0_r3_reg[32]/P0001  ;
	input \u3_u0_r3_reg[33]/P0001  ;
	input \u3_u0_r3_reg[34]/P0001  ;
	input \u3_u0_r3_reg[35]/P0001  ;
	input \u3_u0_r3_reg[3]/P0001  ;
	input \u3_u0_r3_reg[4]/P0001  ;
	input \u3_u0_r3_reg[5]/P0001  ;
	input \u3_u0_r3_reg[6]/P0001  ;
	input \u3_u0_r3_reg[7]/P0001  ;
	input \u3_u0_r3_reg[8]/P0001  ;
	input \u3_u0_r3_reg[9]/P0001  ;
	input \u3_u0_rd_adr_reg[0]/NET0131  ;
	input \u3_u0_rd_adr_reg[1]/NET0131  ;
	input \u3_u0_rd_adr_reg[2]/NET0131  ;
	input \u3_u0_rd_adr_reg[3]/NET0131  ;
	input \u3_u0_wr_adr_reg[0]/NET0131  ;
	input \u3_u0_wr_adr_reg[1]/NET0131  ;
	input \u3_u0_wr_adr_reg[2]/NET0131  ;
	input \u3_u0_wr_adr_reg[3]/NET0131  ;
	input \u4_ps_cnt_reg[0]/NET0131  ;
	input \u4_ps_cnt_reg[1]/NET0131  ;
	input \u4_ps_cnt_reg[2]/NET0131  ;
	input \u4_ps_cnt_reg[3]/NET0131  ;
	input \u4_ps_cnt_reg[4]/NET0131  ;
	input \u4_ps_cnt_reg[5]/NET0131  ;
	input \u4_ps_cnt_reg[6]/NET0131  ;
	input \u4_ps_cnt_reg[7]/NET0131  ;
	input \u4_rfr_ce_reg/NET0131  ;
	input \u4_rfr_clr_reg/P0001  ;
	input \u4_rfr_cnt_reg[0]/NET0131  ;
	input \u4_rfr_cnt_reg[1]/NET0131  ;
	input \u4_rfr_cnt_reg[2]/NET0131  ;
	input \u4_rfr_cnt_reg[3]/NET0131  ;
	input \u4_rfr_cnt_reg[4]/NET0131  ;
	input \u4_rfr_cnt_reg[5]/NET0131  ;
	input \u4_rfr_cnt_reg[6]/NET0131  ;
	input \u4_rfr_cnt_reg[7]/NET0131  ;
	input \u4_rfr_early_reg/NET0131  ;
	input \u4_rfr_en_reg/NET0131  ;
	input \u4_rfr_req_reg/NET0131  ;
	input \u5_ack_cnt_reg[0]/NET0131  ;
	input \u5_ack_cnt_reg[1]/NET0131  ;
	input \u5_ack_cnt_reg[2]/NET0131  ;
	input \u5_ack_cnt_reg[3]/NET0131  ;
	input \u5_ap_en_reg/NET0131  ;
	input \u5_burst_act_rd_reg/P0001  ;
	input \u5_burst_cnt_reg[0]/NET0131  ;
	input \u5_burst_cnt_reg[10]/NET0131  ;
	input \u5_burst_cnt_reg[1]/NET0131  ;
	input \u5_burst_cnt_reg[2]/NET0131  ;
	input \u5_burst_cnt_reg[3]/NET0131  ;
	input \u5_burst_cnt_reg[4]/NET0131  ;
	input \u5_burst_cnt_reg[5]/NET0131  ;
	input \u5_burst_cnt_reg[6]/NET0131  ;
	input \u5_burst_cnt_reg[7]/NET0131  ;
	input \u5_burst_cnt_reg[8]/NET0131  ;
	input \u5_burst_cnt_reg[9]/NET0131  ;
	input \u5_cke_o_del_reg/P0001  ;
	input \u5_cke_r_reg/NET0131  ;
	input \u5_cmd_a10_r_reg/P0001  ;
	input \u5_cmd_asserted2_reg/NET0131  ;
	input \u5_cmd_asserted_reg/NET0131  ;
	input \u5_cmd_del_reg[0]/NET0131  ;
	input \u5_cmd_del_reg[1]/NET0131  ;
	input \u5_cmd_del_reg[2]/NET0131  ;
	input \u5_cmd_del_reg[3]/NET0131  ;
	input \u5_cnt_reg/NET0131  ;
	input \u5_cs_le_r_reg/P0001  ;
	input \u5_cs_le_reg/P0001  ;
	input \u5_data_oe_r2_reg/NET0131  ;
	input \u5_data_oe_reg/NET0131  ;
	input \u5_dv_r_reg/NET0131  ;
	input \u5_ir_cnt_done_reg/P0001  ;
	input \u5_ir_cnt_reg[0]/P0001  ;
	input \u5_ir_cnt_reg[1]/P0001  ;
	input \u5_ir_cnt_reg[2]/P0001  ;
	input \u5_ir_cnt_reg[3]/P0001  ;
	input \u5_lmr_ack_reg/NET0131  ;
	input \u5_lookup_ready1_reg/NET0131  ;
	input \u5_lookup_ready2_reg/NET0131  ;
	input \u5_mc_adv_r1_reg/NET0131  ;
	input \u5_mc_adv_r_reg/NET0131  ;
	input \u5_mc_c_oe_reg/NET0131  ;
	input \u5_mc_le_reg/NET0131  ;
	input \u5_mem_ack_r_reg/NET0131  ;
	input \u5_no_wb_cycle_reg/NET0131  ;
	input \u5_oe__reg/NET0131  ;
	input \u5_pack_le0_reg/P0001  ;
	input \u5_pack_le1_reg/P0001  ;
	input \u5_resume_req_r_reg/NET0131  ;
	input \u5_rfr_ack_r_reg/NET0131  ;
	input \u5_state_reg[0]/NET0131  ;
	input \u5_state_reg[10]/NET0131  ;
	input \u5_state_reg[11]/NET0131  ;
	input \u5_state_reg[12]/NET0131  ;
	input \u5_state_reg[13]/NET0131  ;
	input \u5_state_reg[14]/NET0131  ;
	input \u5_state_reg[15]/NET0131  ;
	input \u5_state_reg[16]/NET0131  ;
	input \u5_state_reg[17]/NET0131  ;
	input \u5_state_reg[18]/NET0131  ;
	input \u5_state_reg[19]/NET0131  ;
	input \u5_state_reg[1]/NET0131  ;
	input \u5_state_reg[20]/NET0131  ;
	input \u5_state_reg[21]/NET0131  ;
	input \u5_state_reg[22]/NET0131  ;
	input \u5_state_reg[23]/NET0131  ;
	input \u5_state_reg[24]/NET0131  ;
	input \u5_state_reg[25]/NET0131  ;
	input \u5_state_reg[26]/NET0131  ;
	input \u5_state_reg[27]/NET0131  ;
	input \u5_state_reg[28]/NET0131  ;
	input \u5_state_reg[29]/NET0131  ;
	input \u5_state_reg[2]/NET0131  ;
	input \u5_state_reg[30]/NET0131  ;
	input \u5_state_reg[31]/NET0131  ;
	input \u5_state_reg[32]/NET0131  ;
	input \u5_state_reg[33]/NET0131  ;
	input \u5_state_reg[34]/NET0131  ;
	input \u5_state_reg[35]/NET0131  ;
	input \u5_state_reg[36]/NET0131  ;
	input \u5_state_reg[37]/NET0131  ;
	input \u5_state_reg[38]/NET0131  ;
	input \u5_state_reg[39]/NET0131  ;
	input \u5_state_reg[3]/NET0131  ;
	input \u5_state_reg[40]/NET0131  ;
	input \u5_state_reg[41]/NET0131  ;
	input \u5_state_reg[42]/NET0131  ;
	input \u5_state_reg[43]/NET0131  ;
	input \u5_state_reg[44]/NET0131  ;
	input \u5_state_reg[45]/NET0131  ;
	input \u5_state_reg[46]/NET0131  ;
	input \u5_state_reg[47]/NET0131  ;
	input \u5_state_reg[48]/NET0131  ;
	input \u5_state_reg[49]/NET0131  ;
	input \u5_state_reg[4]/NET0131  ;
	input \u5_state_reg[50]/NET0131  ;
	input \u5_state_reg[51]/NET0131  ;
	input \u5_state_reg[52]/NET0131  ;
	input \u5_state_reg[53]/NET0131  ;
	input \u5_state_reg[54]/NET0131  ;
	input \u5_state_reg[55]/NET0131  ;
	input \u5_state_reg[56]/NET0131  ;
	input \u5_state_reg[57]/NET0131  ;
	input \u5_state_reg[58]/NET0131  ;
	input \u5_state_reg[59]/NET0131  ;
	input \u5_state_reg[5]/NET0131  ;
	input \u5_state_reg[60]/NET0131  ;
	input \u5_state_reg[61]/NET0131  ;
	input \u5_state_reg[62]/NET0131  ;
	input \u5_state_reg[63]/NET0131  ;
	input \u5_state_reg[64]/NET0131  ;
	input \u5_state_reg[65]/NET0131  ;
	input \u5_state_reg[6]/NET0131  ;
	input \u5_state_reg[7]/NET0131  ;
	input \u5_state_reg[8]/NET0131  ;
	input \u5_state_reg[9]/NET0131  ;
	input \u5_susp_req_r_reg/NET0131  ;
	input \u5_susp_sel_r_reg/NET0131  ;
	input \u5_timer2_reg[0]/P0001  ;
	input \u5_timer2_reg[1]/P0001  ;
	input \u5_timer2_reg[2]/P0001  ;
	input \u5_timer2_reg[3]/P0001  ;
	input \u5_timer2_reg[4]/P0001  ;
	input \u5_timer2_reg[5]/P0001  ;
	input \u5_timer2_reg[6]/P0001  ;
	input \u5_timer2_reg[7]/P0001  ;
	input \u5_timer2_reg[8]/P0001  ;
	input \u5_timer_reg[0]/NET0131  ;
	input \u5_timer_reg[1]/NET0131  ;
	input \u5_timer_reg[2]/NET0131  ;
	input \u5_timer_reg[3]/NET0131  ;
	input \u5_timer_reg[4]/NET0131  ;
	input \u5_timer_reg[5]/NET0131  ;
	input \u5_timer_reg[6]/NET0131  ;
	input \u5_timer_reg[7]/NET0131  ;
	input \u5_tmr2_done_reg/NET0131  ;
	input \u5_tmr_done_reg/NET0131  ;
	input \u5_wb_cycle_reg/NET0131  ;
	input \u5_wb_stb_first_reg/NET0131  ;
	input \u5_wb_wait_r_reg/P0001  ;
	input \u5_wb_write_go_r_reg/NET0131  ;
	input \u5_wr_cycle_reg/NET0131  ;
	input \u6_read_go_r1_reg/NET0131  ;
	input \u6_read_go_r_reg/NET0131  ;
	input \u6_rmw_en_reg/NET0131  ;
	input \u6_rmw_r_reg/NET0131  ;
	input \u6_wb_first_r_reg/NET0131  ;
	input \u6_wr_hold_reg/NET0131  ;
	input \u6_write_go_r1_reg/NET0131  ;
	input \u6_write_go_r_reg/NET0131  ;
	input \u7_mc_ack_r_reg/NET0131  ;
	input \u7_mc_br_r_reg/P0001  ;
	input \u7_mc_data_ir_reg[0]/P0001  ;
	input \u7_mc_data_ir_reg[10]/P0001  ;
	input \u7_mc_data_ir_reg[11]/P0001  ;
	input \u7_mc_data_ir_reg[12]/P0001  ;
	input \u7_mc_data_ir_reg[13]/P0001  ;
	input \u7_mc_data_ir_reg[14]/P0001  ;
	input \u7_mc_data_ir_reg[15]/P0001  ;
	input \u7_mc_data_ir_reg[16]/P0001  ;
	input \u7_mc_data_ir_reg[17]/P0001  ;
	input \u7_mc_data_ir_reg[18]/P0001  ;
	input \u7_mc_data_ir_reg[19]/P0001  ;
	input \u7_mc_data_ir_reg[1]/P0001  ;
	input \u7_mc_data_ir_reg[20]/P0001  ;
	input \u7_mc_data_ir_reg[21]/P0001  ;
	input \u7_mc_data_ir_reg[22]/P0001  ;
	input \u7_mc_data_ir_reg[23]/P0001  ;
	input \u7_mc_data_ir_reg[24]/P0001  ;
	input \u7_mc_data_ir_reg[25]/P0001  ;
	input \u7_mc_data_ir_reg[26]/P0001  ;
	input \u7_mc_data_ir_reg[27]/P0001  ;
	input \u7_mc_data_ir_reg[28]/P0001  ;
	input \u7_mc_data_ir_reg[29]/P0001  ;
	input \u7_mc_data_ir_reg[2]/P0001  ;
	input \u7_mc_data_ir_reg[30]/P0001  ;
	input \u7_mc_data_ir_reg[31]/P0001  ;
	input \u7_mc_data_ir_reg[3]/P0001  ;
	input \u7_mc_data_ir_reg[4]/P0001  ;
	input \u7_mc_data_ir_reg[5]/P0001  ;
	input \u7_mc_data_ir_reg[6]/P0001  ;
	input \u7_mc_data_ir_reg[7]/P0001  ;
	input \u7_mc_data_ir_reg[8]/P0001  ;
	input \u7_mc_data_ir_reg[9]/P0001  ;
	input \u7_mc_dqm_r2_reg[0]/P0001  ;
	input \u7_mc_dqm_r2_reg[1]/P0001  ;
	input \u7_mc_dqm_r2_reg[2]/P0001  ;
	input \u7_mc_dqm_r2_reg[3]/P0001  ;
	input \u7_mc_dqm_r_reg[0]/P0001  ;
	input \u7_mc_dqm_r_reg[1]/P0001  ;
	input \u7_mc_dqm_r_reg[2]/P0001  ;
	input \u7_mc_dqm_r_reg[3]/P0001  ;
	input wb_ack_o_pad ;
	input \wb_addr_i[0]_pad  ;
	input \wb_addr_i[10]_pad  ;
	input \wb_addr_i[11]_pad  ;
	input \wb_addr_i[12]_pad  ;
	input \wb_addr_i[13]_pad  ;
	input \wb_addr_i[14]_pad  ;
	input \wb_addr_i[15]_pad  ;
	input \wb_addr_i[16]_pad  ;
	input \wb_addr_i[17]_pad  ;
	input \wb_addr_i[18]_pad  ;
	input \wb_addr_i[19]_pad  ;
	input \wb_addr_i[1]_pad  ;
	input \wb_addr_i[20]_pad  ;
	input \wb_addr_i[21]_pad  ;
	input \wb_addr_i[22]_pad  ;
	input \wb_addr_i[23]_pad  ;
	input \wb_addr_i[24]_pad  ;
	input \wb_addr_i[25]_pad  ;
	input \wb_addr_i[26]_pad  ;
	input \wb_addr_i[27]_pad  ;
	input \wb_addr_i[28]_pad  ;
	input \wb_addr_i[29]_pad  ;
	input \wb_addr_i[2]_pad  ;
	input \wb_addr_i[30]_pad  ;
	input \wb_addr_i[31]_pad  ;
	input \wb_addr_i[3]_pad  ;
	input \wb_addr_i[4]_pad  ;
	input \wb_addr_i[5]_pad  ;
	input \wb_addr_i[6]_pad  ;
	input \wb_addr_i[7]_pad  ;
	input \wb_addr_i[8]_pad  ;
	input \wb_addr_i[9]_pad  ;
	input wb_cyc_i_pad ;
	input \wb_data_i[0]_pad  ;
	input \wb_data_i[10]_pad  ;
	input \wb_data_i[11]_pad  ;
	input \wb_data_i[12]_pad  ;
	input \wb_data_i[13]_pad  ;
	input \wb_data_i[14]_pad  ;
	input \wb_data_i[15]_pad  ;
	input \wb_data_i[16]_pad  ;
	input \wb_data_i[17]_pad  ;
	input \wb_data_i[18]_pad  ;
	input \wb_data_i[19]_pad  ;
	input \wb_data_i[1]_pad  ;
	input \wb_data_i[20]_pad  ;
	input \wb_data_i[21]_pad  ;
	input \wb_data_i[22]_pad  ;
	input \wb_data_i[23]_pad  ;
	input \wb_data_i[24]_pad  ;
	input \wb_data_i[25]_pad  ;
	input \wb_data_i[26]_pad  ;
	input \wb_data_i[27]_pad  ;
	input \wb_data_i[28]_pad  ;
	input \wb_data_i[29]_pad  ;
	input \wb_data_i[2]_pad  ;
	input \wb_data_i[30]_pad  ;
	input \wb_data_i[31]_pad  ;
	input \wb_data_i[3]_pad  ;
	input \wb_data_i[4]_pad  ;
	input \wb_data_i[5]_pad  ;
	input \wb_data_i[6]_pad  ;
	input \wb_data_i[7]_pad  ;
	input \wb_data_i[8]_pad  ;
	input \wb_data_i[9]_pad  ;
	input wb_err_o_pad ;
	input \wb_sel_i[0]_pad  ;
	input \wb_sel_i[1]_pad  ;
	input \wb_sel_i[2]_pad  ;
	input \wb_sel_i[3]_pad  ;
	input wb_stb_i_pad ;
	input wb_we_i_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g22/_0_  ;
	output \g23/_0_  ;
	output \g25_dup61718/_2_  ;
	output \g43466/_0_  ;
	output \g43467/_0_  ;
	output \g43468/_0_  ;
	output \g43469/_0_  ;
	output \g43470/_0_  ;
	output \g43471/_0_  ;
	output \g43472/_0_  ;
	output \g43473/_0_  ;
	output \g43474/_0_  ;
	output \g43475/_0_  ;
	output \g43476/_0_  ;
	output \g43477/_0_  ;
	output \g43478/_0_  ;
	output \g43512/_0_  ;
	output \g43513/_0_  ;
	output \g43544/_3_  ;
	output \g43545/_0_  ;
	output \g43554/_0_  ;
	output \g43555/_0_  ;
	output \g43557/_0_  ;
	output \g43558/_0_  ;
	output \g43571/_2_  ;
	output \g43632/_0_  ;
	output \g43633/_0_  ;
	output \g43635/_0_  ;
	output \g43636/_0_  ;
	output \g43637/_0_  ;
	output \g43638/_0_  ;
	output \g43639/_0_  ;
	output \g43640/_0_  ;
	output \g43642/_0_  ;
	output \g43662/_0_  ;
	output \g43663/_0_  ;
	output \g43664/_0_  ;
	output \g43665/_0_  ;
	output \g43668/_0_  ;
	output \g43670/_0_  ;
	output \g43671/_0_  ;
	output \g43673/_0_  ;
	output \g43674/_0_  ;
	output \g43692/_0_  ;
	output \g43695/_0_  ;
	output \g43696/_0_  ;
	output \g43697/_0_  ;
	output \g43698/_0_  ;
	output \g43700/_0_  ;
	output \g43701/_0_  ;
	output \g43703/_0_  ;
	output \g43705/_0_  ;
	output \g43707/_0_  ;
	output \g43708/_0_  ;
	output \g43710/_0_  ;
	output \g43717/_0_  ;
	output \g43719/_0_  ;
	output \g43720/_0_  ;
	output \g43721/_0_  ;
	output \g43722/_1_  ;
	output \g43723/_0_  ;
	output \g43725/_0_  ;
	output \g43729/_0_  ;
	output \g43731/_0_  ;
	output \g43734/_0_  ;
	output \g43735/_0_  ;
	output \g43737/_0_  ;
	output \g43744/_0_  ;
	output \g43747/_0_  ;
	output \g43760/_2_  ;
	output \g43770/_1_  ;
	output \g43775/_2_  ;
	output \g43780/_2_  ;
	output \g43786/_0_  ;
	output \g43787/_1_  ;
	output \g43847/_0_  ;
	output \g43848/_1_  ;
	output \g43858/_1_  ;
	output \g43891/_3_  ;
	output \g43895/_0_  ;
	output \g43934/_0_  ;
	output \g43936/_3_  ;
	output \g43954/_3_  ;
	output \g43961/_0_  ;
	output \g44016/_1_  ;
	output \g44067/_0_  ;
	output \g44094/_0_  ;
	output \g44096/_0_  ;
	output \g44104/_0_  ;
	output \g44122/_0_  ;
	output \g44172/_0_  ;
	output \g44209/_0_  ;
	output \g44219/_0_  ;
	output \g44220/_0_  ;
	output \g44222/_0_  ;
	output \g44223/_0_  ;
	output \g44241/_2_  ;
	output \g44252/_0_  ;
	output \g44253/_0_  ;
	output \g44255/_2_  ;
	output \g44263/_2_  ;
	output \g44470/_0_  ;
	output \g44538/_0_  ;
	output \g44539/_0_  ;
	output \g44540/_0_  ;
	output \g44541/_0_  ;
	output \g44542/_0_  ;
	output \g44543/_0_  ;
	output \g44544/_0_  ;
	output \g44545/_0_  ;
	output \g44546/_0_  ;
	output \g44547/_0_  ;
	output \g44548/_0_  ;
	output \g44549/_0_  ;
	output \g44550/_0_  ;
	output \g44551/_0_  ;
	output \g44552/_0_  ;
	output \g44553/_0_  ;
	output \g44554/_0_  ;
	output \g44555/_0_  ;
	output \g44556/_0_  ;
	output \g44557/_0_  ;
	output \g44558/_0_  ;
	output \g44559/_0_  ;
	output \g44560/_0_  ;
	output \g44561/_0_  ;
	output \g44562/_0_  ;
	output \g44563/_0_  ;
	output \g44564/_0_  ;
	output \g44565/_0_  ;
	output \g44566/_0_  ;
	output \g44567/_0_  ;
	output \g44568/_0_  ;
	output \g44569/_0_  ;
	output \g44570/_0_  ;
	output \g44571/_0_  ;
	output \g44572/_0_  ;
	output \g44573/_0_  ;
	output \g44574/_0_  ;
	output \g44575/_0_  ;
	output \g44576/_0_  ;
	output \g44577/_0_  ;
	output \g44578/_0_  ;
	output \g44579/_0_  ;
	output \g44580/_0_  ;
	output \g44581/_0_  ;
	output \g44582/_0_  ;
	output \g44583/_0_  ;
	output \g44584/_0_  ;
	output \g44585/_0_  ;
	output \g44586/_0_  ;
	output \g44588/_0_  ;
	output \g44589/_0_  ;
	output \g44590/_0_  ;
	output \g44591/_0_  ;
	output \g44592/_0_  ;
	output \g44593/_0_  ;
	output \g44594/_0_  ;
	output \g44595/_0_  ;
	output \g44596/_0_  ;
	output \g44636/_2_  ;
	output \g44646/_0_  ;
	output \g44647/_0_  ;
	output \g44648/_0_  ;
	output \g44649/_0_  ;
	output \g44650/_0_  ;
	output \g44651/_0_  ;
	output \g44652/_0_  ;
	output \g44653/_0_  ;
	output \g44654/_0_  ;
	output \g44655/_0_  ;
	output \g44656/_0_  ;
	output \g44657/_0_  ;
	output \g44665/_0_  ;
	output \g44666/_0_  ;
	output \g44667/_0_  ;
	output \g44668/_0_  ;
	output \g44752/_0_  ;
	output \g44753/_0_  ;
	output \g44873/_0_  ;
	output \g44939/_0_  ;
	output \g44942/_0_  ;
	output \g44945/_0_  ;
	output \g45023/_2_  ;
	output \g45090/_0_  ;
	output \g45141/_0_  ;
	output \g45147/_3_  ;
	output \g45155/_0_  ;
	output \g45190/_0_  ;
	output \g45195/_2_  ;
	output \g45199/_2_  ;
	output \g45201/_2_  ;
	output \g45324/_0_  ;
	output \g45334/_2_  ;
	output \g45336/_0_  ;
	output \g45388/_0_  ;
	output \g45391/_0_  ;
	output \g45413/_2_  ;
	output \g45530/_0_  ;
	output \g45532/_0_  ;
	output \g45533/_0_  ;
	output \g45534/_0_  ;
	output \g45739/_2_  ;
	output \g45743/_2_  ;
	output \g45767/_0_  ;
	output \g45782/_0_  ;
	output \g45830/_3_  ;
	output \g45834/_3_  ;
	output \g45835/_3_  ;
	output \g45836/_3_  ;
	output \g45837/_3_  ;
	output \g45839/_3_  ;
	output \g45840/_3_  ;
	output \g45841/_3_  ;
	output \g45842/_3_  ;
	output \g45843/_3_  ;
	output \g45844/_3_  ;
	output \g45845/_3_  ;
	output \g46191/_0_  ;
	output \g46193/_3_  ;
	output \g46256/_3_  ;
	output \g46257/_3_  ;
	output \g46258/_3_  ;
	output \g46259/_3_  ;
	output \g46260/_3_  ;
	output \g46261/_3_  ;
	output \g46262/_3_  ;
	output \g46263/_3_  ;
	output \g46278/_0_  ;
	output \g46292/_0_  ;
	output \g46293/_0_  ;
	output \g46312/_0_  ;
	output \g46367/_2_  ;
	output \g46370/_2_  ;
	output \g46380/_2_  ;
	output \g46386/_2_  ;
	output \g46388/_2_  ;
	output \g46392/_2_  ;
	output \g46395/_2_  ;
	output \g46399/_2_  ;
	output \g46420/_0_  ;
	output \g46446/_0_  ;
	output \g46493/_0_  ;
	output \g46510/_0_  ;
	output \g46669/_2_  ;
	output \g46691/_0_  ;
	output \g46708/_0_  ;
	output \g46721/_00_  ;
	output \g46776/_0_  ;
	output \g46777/_0_  ;
	output \g46778/_0_  ;
	output \g46779/_0_  ;
	output \g46780/_0_  ;
	output \g46782/_0_  ;
	output \g46784/_0_  ;
	output \g46932/_0_  ;
	output \g47112/_0_  ;
	output \g47124/_0_  ;
	output \g47265/_0_  ;
	output \g47270/_0_  ;
	output \g47275/_0_  ;
	output \g47300/_1_  ;
	output \g47305/_1_  ;
	output \g47338/_0_  ;
	output \g47339/_0_  ;
	output \g47352/_0_  ;
	output \g47699/_3_  ;
	output \g47711/_0_  ;
	output \g47719/_3_  ;
	output \g47721/_3_  ;
	output \g47723/_3_  ;
	output \g47853/_0_  ;
	output \g48094/_0_  ;
	output \g48095/_0_  ;
	output \g48177/_2_  ;
	output \g48194/_0_  ;
	output \g48369/_2_  ;
	output \g48371/_2_  ;
	output \g48373/_2_  ;
	output \g48375/_2_  ;
	output \g48377/_2_  ;
	output \g48379/_2_  ;
	output \g48381/_2_  ;
	output \g48383/_2_  ;
	output \g48385/_2_  ;
	output \g48535/_0_  ;
	output \g48569/_0_  ;
	output \g48570/_0_  ;
	output \g48571/_0_  ;
	output \g48836/_0_  ;
	output \g48843/_0_  ;
	output \g49187/_3_  ;
	output \g49375/_2_  ;
	output \g49633/_0_  ;
	output \g49788/_1_  ;
	output \g49800/_1_  ;
	output \g49802/_1_  ;
	output \g49806/_1_  ;
	output \g49853/_1_  ;
	output \g49883/_0_  ;
	output \g49884/_0_  ;
	output \g49885/_0_  ;
	output \g49886/_0_  ;
	output \g49976/_1_  ;
	output \g50038/_0_  ;
	output \g50082/_0_  ;
	output \g50083/_0_  ;
	output \g50167/_3_  ;
	output \g50168/_3_  ;
	output \g50169/_3_  ;
	output \g50170/_3_  ;
	output \g50171/_3_  ;
	output \g50177/_0_  ;
	output \g50190/_0_  ;
	output \g50236/_0_  ;
	output \g50251/_3_  ;
	output \g50256/_0_  ;
	output \g50318/_3_  ;
	output \g50319/_3_  ;
	output \g50350/_3_  ;
	output \g50351/_3_  ;
	output \g50352/_3_  ;
	output \g50353/_3_  ;
	output \g50354/_3_  ;
	output \g50355/_3_  ;
	output \g50361/_2_  ;
	output \g50366/_0_  ;
	output \g50393/_0_  ;
	output \g50552/_1_  ;
	output \g51108/_0_  ;
	output \g51160/_0_  ;
	output \g51290/_1_  ;
	output \g51327/_3_  ;
	output \g51328/_3_  ;
	output \g51329/_3_  ;
	output \g51330/_3_  ;
	output \g51331/_3_  ;
	output \g51332/_3_  ;
	output \g51333/_3_  ;
	output \g51334/_3_  ;
	output \g51339/_3_  ;
	output \g51340/_3_  ;
	output \g51341/_3_  ;
	output \g51342/_3_  ;
	output \g51343/_3_  ;
	output \g51346/_0_  ;
	output \g51347/_0_  ;
	output \g51348/_0_  ;
	output \g51381/_3_  ;
	output \g51382/_3_  ;
	output \g51383/_3_  ;
	output \g51386/_3_  ;
	output \g51387/_3_  ;
	output \g51405/_3_  ;
	output \g51410/_3_  ;
	output \g51883/_0_  ;
	output \g51916/_0_  ;
	output \g51947/_0_  ;
	output \g51948/_0_  ;
	output \g51949/_0_  ;
	output \g51950/_0_  ;
	output \g51951/_0_  ;
	output \g51952/_0_  ;
	output \g51953/_0_  ;
	output \g51954/_0_  ;
	output \g51955/_0_  ;
	output \g51956/_0_  ;
	output \g51957/_0_  ;
	output \g51958/_0_  ;
	output \g51959/_0_  ;
	output \g51960/_0_  ;
	output \g51961/_0_  ;
	output \g51962/_0_  ;
	output \g51963/_0_  ;
	output \g51964/_0_  ;
	output \g51965/_0_  ;
	output \g51967/_0_  ;
	output \g51968/_0_  ;
	output \g51969/_0_  ;
	output \g51970/_0_  ;
	output \g51971/_0_  ;
	output \g51972/_0_  ;
	output \g51973/_0_  ;
	output \g51974/_0_  ;
	output \g51975/_0_  ;
	output \g51976/_0_  ;
	output \g51977/_0_  ;
	output \g51978/_0_  ;
	output \g51979/_0_  ;
	output \g51980/_0_  ;
	output \g51981/_0_  ;
	output \g51982/_0_  ;
	output \g51983/_0_  ;
	output \g51984/_0_  ;
	output \g51985/_0_  ;
	output \g51986/_0_  ;
	output \g51987/_0_  ;
	output \g51988/_0_  ;
	output \g51989/_0_  ;
	output \g51990/_0_  ;
	output \g51991/_0_  ;
	output \g51992/_0_  ;
	output \g51993/_0_  ;
	output \g51994/_0_  ;
	output \g51995/_0_  ;
	output \g51996/_0_  ;
	output \g51997/_0_  ;
	output \g51998/_0_  ;
	output \g51999/_0_  ;
	output \g52000/_0_  ;
	output \g52001/_0_  ;
	output \g52002/_0_  ;
	output \g52003/_0_  ;
	output \g52004/_0_  ;
	output \g52005/_0_  ;
	output \g52006/_0_  ;
	output \g52007/_0_  ;
	output \g52008/_0_  ;
	output \g52009/_0_  ;
	output \g52010/_0_  ;
	output \g52011/_0_  ;
	output \g52012/_0_  ;
	output \g52013/_0_  ;
	output \g52014/_0_  ;
	output \g52015/_0_  ;
	output \g52016/_0_  ;
	output \g52017/_0_  ;
	output \g52018/_0_  ;
	output \g52019/_0_  ;
	output \g52020/_0_  ;
	output \g52021/_0_  ;
	output \g52022/_0_  ;
	output \g52023/_0_  ;
	output \g52024/_0_  ;
	output \g52025/_0_  ;
	output \g52026/_0_  ;
	output \g52027/_0_  ;
	output \g52028/_0_  ;
	output \g52029/_0_  ;
	output \g52030/_0_  ;
	output \g52031/_0_  ;
	output \g52032/_0_  ;
	output \g52033/_0_  ;
	output \g52034/_0_  ;
	output \g52035/_0_  ;
	output \g52036/_0_  ;
	output \g52037/_0_  ;
	output \g52038/_0_  ;
	output \g52039/_0_  ;
	output \g52040/_0_  ;
	output \g52041/_0_  ;
	output \g52042/_0_  ;
	output \g52043/_0_  ;
	output \g52044/_0_  ;
	output \g52045/_0_  ;
	output \g52046/_0_  ;
	output \g52047/_0_  ;
	output \g52049/_0_  ;
	output \g52050/_0_  ;
	output \g52051/_0_  ;
	output \g52052/_0_  ;
	output \g52053/_0_  ;
	output \g52054/_0_  ;
	output \g52055/_0_  ;
	output \g52056/_0_  ;
	output \g52057/_0_  ;
	output \g52058/_0_  ;
	output \g52061/_0_  ;
	output \g52065/_0_  ;
	output \g52066/_0_  ;
	output \g52067/_0_  ;
	output \g52068/_0_  ;
	output \g52069/_0_  ;
	output \g52070/_0_  ;
	output \g52071/_0_  ;
	output \g52073/_0_  ;
	output \g52074/_0_  ;
	output \g52075/_0_  ;
	output \g52082/_0_  ;
	output \g52083/_0_  ;
	output \g52158/_0_  ;
	output \g52201/_0_  ;
	output \g52202/_0_  ;
	output \g52346/_0_  ;
	output \g52351/_0_  ;
	output \g52390/_0_  ;
	output \g52847/_0_  ;
	output \g52854/_0_  ;
	output \g52968/_0_  ;
	output \g52969/_0_  ;
	output \g52970/_0_  ;
	output \g52971/_0_  ;
	output \g52984/_0_  ;
	output \g52994/_0_  ;
	output \g53019/_0_  ;
	output \g53030/_0_  ;
	output \g53094/_1_  ;
	output \g53106/_0_  ;
	output \g53150/_0_  ;
	output \g53256/_0_  ;
	output \g53297/_0_  ;
	output \g53345/_0_  ;
	output \g53359/_0_  ;
	output \g53375/_0_  ;
	output \g53474/_1__syn_2  ;
	output \g53475/_2_  ;
	output \g53593/_0_  ;
	output \g53643/_1_  ;
	output \g53655/_0_  ;
	output \g53710/_0_  ;
	output \g53786/_0_  ;
	output \g53837/_0_  ;
	output \g53888/_1_  ;
	output \g53909/_0_  ;
	output \g54253/_2_  ;
	output \g54394/_3_  ;
	output \g54413/_0_  ;
	output \g55420/_0_  ;
	output \g55587/_0_  ;
	output \g55852/_0_  ;
	output \g57020/_0_  ;
	output \g59450/_0_  ;
	output \g59488/_2_  ;
	output \g59752/_0_  ;
	output \g59786/_0_  ;
	output \g59854/_0_  ;
	output \g59878/_0_  ;
	output \g59902/_0_  ;
	output \g59924/_0_  ;
	output \g59947/_0_  ;
	output \g59972/_0_  ;
	output \g59996/_0_  ;
	output \g60017/_0_  ;
	output \g60040/_0_  ;
	output \g60064/_0_  ;
	output \g60095/_0_  ;
	output \g60119/_0_  ;
	output \g60145/_1_  ;
	output \g60165/_0_  ;
	output \g60407/_2_  ;
	output \g60408/_0_  ;
	output \g60613/_2_  ;
	output \g60649/_0_  ;
	output \g60771/_0_  ;
	output \g60908/_1_  ;
	output \g60911/_0_  ;
	output \g60977/_0_  ;
	output \g61/_0_  ;
	output \g61002/_0_  ;
	output \g61308/_0_  ;
	output \g61312/_1_  ;
	output \g61314/_0_  ;
	output \g61319/_1_  ;
	output \g61342/_1_  ;
	output \g61360/_0_  ;
	output \g61377/_0_  ;
	output \g61423/_1_  ;
	output \g61426/_0_  ;
	output \g61479/_1_  ;
	output \g61523/_1_  ;
	output \g61558/_1_  ;
	output \g61652/_0_  ;
	output \g61866/_0_  ;
	output \g61868/_1_  ;
	output \g61887/_0_  ;
	output \u7_mc_dqm_r_reg[0]/P0001_reg_syn_3  ;
	output \u7_mc_dqm_r_reg[1]/P0001_reg_syn_3  ;
	output \u7_mc_dqm_r_reg[2]/P0001_reg_syn_3  ;
	output \u7_mc_dqm_r_reg[3]/P0001_reg_syn_3  ;
	output \u7_mc_we__reg/_05_  ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		_w959_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\u5_state_reg[50]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w960_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w959_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\u5_state_reg[63]/NET0131 ,
		\u5_state_reg[64]/NET0131 ,
		_w962_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\u5_state_reg[62]/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w963_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w962_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\u5_state_reg[60]/NET0131 ,
		\u5_state_reg[61]/NET0131 ,
		_w965_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w966_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w965_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w964_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\u5_state_reg[15]/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		_w969_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		_w970_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w969_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\u5_state_reg[6]/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\u5_state_reg[7]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w973_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w972_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		_w971_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		_w978_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w977_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\u5_state_reg[3]/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		_w980_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w979_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w976_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w975_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\u5_state_reg[38]/NET0131 ,
		\u5_state_reg[39]/NET0131 ,
		_w984_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w985_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w984_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\u5_state_reg[43]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w988_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w987_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w986_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w992_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w991_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		_w994_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\u5_state_reg[46]/NET0131 ,
		\u5_state_reg[49]/NET0131 ,
		_w995_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w994_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w993_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w990_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w999_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		_w1000_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w999_,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		_w1002_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\u5_state_reg[20]/NET0131 ,
		\u5_state_reg[21]/NET0131 ,
		_w1003_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w1002_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w1001_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		_w1006_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		_w1007_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w1006_,
		_w1007_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\u5_state_reg[32]/NET0131 ,
		\u5_state_reg[33]/NET0131 ,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		_w1010_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w1009_,
		_w1010_,
		_w1011_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w1008_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w1005_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w998_,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w983_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w1016_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w1015_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w968_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w961_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\u5_state_reg[56]/NET0131 ,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\u5_state_reg[54]/NET0131 ,
		\u5_state_reg[55]/NET0131 ,
		_w1021_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		\u5_state_reg[57]/NET0131 ,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w1020_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		\u5_dv_r_reg/NET0131 ,
		\u5_mc_adv_r_reg/NET0131 ,
		_w1024_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w1023_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\u5_state_reg[3]/NET0131 ,
		_w976_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\u5_state_reg[54]/NET0131 ,
		\u5_state_reg[55]/NET0131 ,
		_w1027_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		\u5_state_reg[56]/NET0131 ,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\u5_state_reg[57]/NET0131 ,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w961_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w968_,
		_w1016_,
		_w1031_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w1030_,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w1014_,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w975_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		\u5_state_reg[5]/NET0131 ,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w1026_,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w977_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w1037_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		\u5_cnt_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w1040_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\u5_burst_act_rd_reg/P0001 ,
		\u5_cke_o_del_reg/P0001 ,
		_w1041_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		_w1040_,
		_w1041_,
		_w1042_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w1039_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w1025_,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\u3_u0_wr_adr_reg[3]/NET0131 ,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w1046_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		wb_we_i_pad,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\u6_rmw_en_reg/NET0131 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1048_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		\u5_state_reg[26]/NET0131 ,
		_w1008_,
		_w1050_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\u5_lmr_ack_reg/NET0131 ,
		_w1050_,
		_w1051_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\u0_sp_csc_reg[1]/NET0131 ,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\u0_csc_reg[1]/NET0131 ,
		_w1051_,
		_w1053_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w1052_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		\u0_sp_csc_reg[3]/NET0131 ,
		_w1051_,
		_w1055_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\u0_csc_reg[3]/NET0131 ,
		_w1051_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w1055_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w1054_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		\u0_sp_csc_reg[2]/NET0131 ,
		_w1051_,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		\u0_csc_reg[2]/NET0131 ,
		_w1051_,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w1059_,
		_w1060_,
		_w1061_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w1058_,
		_w1061_,
		_w1062_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		_w998_,
		_w1032_,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w1001_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w983_,
		_w1012_,
		_w1065_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w1064_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		\u5_state_reg[21]/NET0131 ,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		_w1068_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\u5_state_reg[20]/NET0131 ,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w1067_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w983_,
		_w1004_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w1011_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w1064_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		\u5_state_reg[24]/NET0131 ,
		_w1006_,
		_w1074_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		\u5_state_reg[22]/NET0131 ,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		_w1073_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w1070_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\u5_state_reg[18]/NET0131 ,
		_w1067_,
		_w1078_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w1079_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		_w1078_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w983_,
		_w1013_,
		_w1081_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w1032_,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w990_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w993_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		\u5_state_reg[46]/NET0131 ,
		\u5_state_reg[49]/NET0131 ,
		_w1085_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w994_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w1084_,
		_w1086_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w1080_,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w982_,
		_w1033_,
		_w1089_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w971_,
		_w1089_,
		_w1090_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w973_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		\u5_state_reg[6]/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		_w1092_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w1091_,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		_w1088_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w995_,
		_w1084_,
		_w1095_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		_w1096_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w1017_,
		_w1030_,
		_w1098_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w967_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w963_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		\u5_state_reg[63]/NET0131 ,
		\u5_state_reg[64]/NET0131 ,
		_w1101_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w1100_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w1097_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\u5_state_reg[3]/NET0131 ,
		_w976_,
		_w1104_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		_w979_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w1035_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\u5_state_reg[57]/NET0131 ,
		_w1028_,
		_w1107_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w1019_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w1106_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		_w1110_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w960_,
		_w1029_,
		_w1111_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w1018_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		_w1110_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w1023_,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w962_,
		_w1099_,
		_w1115_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		\u5_state_reg[62]/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w1116_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w1115_,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w997_,
		_w1082_,
		_w1118_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w989_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		_w984_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		_w1119_,
		_w1121_,
		_w1122_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w1117_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w1114_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		_w1103_,
		_w1109_,
		_w1125_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		_w1094_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w1124_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w1077_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		_w1007_,
		_w1073_,
		_w1129_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w1129_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w1132_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		_w1133_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w986_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w1118_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		_w1132_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		\u5_state_reg[54]/NET0131 ,
		\u5_state_reg[55]/NET0131 ,
		_w1137_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		\u5_state_reg[57]/NET0131 ,
		_w1137_,
		_w1138_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w1020_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\u5_state_reg[62]/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w1140_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		_w1115_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w1142_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w986_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		_w1118_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		_w1145_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w1144_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w1147_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w1135_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		_w1149_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		_w1144_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w1148_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w959_,
		_w966_,
		_w1152_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w964_,
		_w965_,
		_w1153_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w1029_,
		_w1152_,
		_w1154_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w1153_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w1017_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		\u5_state_reg[50]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w1157_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w1156_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w1131_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w1136_,
		_w1146_,
		_w1160_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		_w1159_,
		_w1160_,
		_w1161_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w1139_,
		_w1141_,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w1151_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w1161_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w996_,
		_w1083_,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w992_,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		_w1167_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w1166_,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		_w1164_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\u0_sp_tms_reg[1]/NET0131 ,
		_w1051_,
		_w1170_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\u0_tms_reg[1]/NET0131 ,
		_w1051_,
		_w1171_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w1170_,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h2)
	) name214 (
		\u0_sp_tms_reg[2]/NET0131 ,
		_w1051_,
		_w1173_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		\u0_tms_reg[2]/NET0131 ,
		_w1051_,
		_w1174_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w1173_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w1172_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		\u0_sp_tms_reg[0]/NET0131 ,
		_w1051_,
		_w1177_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\u0_tms_reg[0]/NET0131 ,
		_w1051_,
		_w1178_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w1177_,
		_w1178_,
		_w1179_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		_w1176_,
		_w1179_,
		_w1180_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\u0_sp_tms_reg[9]/NET0131 ,
		_w1051_,
		_w1181_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\u0_tms_reg[9]/NET0131 ,
		_w1051_,
		_w1182_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w1181_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w1180_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1184_,
		_w1185_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w974_,
		_w1089_,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w969_,
		_w1186_,
		_w1187_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		_w1188_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w1187_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		_w1185_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		_w1008_,
		_w1071_,
		_w1191_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w1064_,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		\u5_state_reg[32]/NET0131 ,
		\u5_state_reg[33]/NET0131 ,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w1010_,
		_w1193_,
		_w1194_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w1192_,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		\u5_state_reg[32]/NET0131 ,
		_w1010_,
		_w1196_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\u5_state_reg[33]/NET0131 ,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w1192_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		_w1199_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w1166_,
		_w1199_,
		_w1200_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w1198_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h2)
	) name243 (
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		_w1202_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		_w1129_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w1009_,
		_w1192_,
		_w1204_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		_w1205_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w1204_,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		_w1203_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		_w1039_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		_w1201_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		_w1004_,
		_w1063_,
		_w1210_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		_w1065_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w999_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		_w1213_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w1212_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		_w1215_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w981_,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w1034_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w1214_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w970_,
		_w1186_,
		_w1219_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		\u5_state_reg[15]/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		_w1220_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		_w1219_,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w978_,
		_w1036_,
		_w1222_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		_w1223_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		_w1222_,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		\u5_state_reg[49]/NET0131 ,
		_w994_,
		_w1225_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		\u5_state_reg[46]/NET0131 ,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w1084_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w1224_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w1095_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w1221_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		_w1228_,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w966_,
		_w1098_,
		_w1233_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		\u5_state_reg[60]/NET0131 ,
		\u5_state_reg[61]/NET0131 ,
		_w1234_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w964_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w1233_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		\u5_state_reg[63]/NET0131 ,
		\u5_state_reg[64]/NET0131 ,
		_w1237_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w1100_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\u5_state_reg[56]/NET0131 ,
		\u5_state_reg[57]/NET0131 ,
		_w1239_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		_w1027_,
		_w1239_,
		_w1240_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w1019_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		_w991_,
		_w1165_,
		_w1242_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w1243_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w1242_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		_w1245_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		_w1037_,
		_w1245_,
		_w1246_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w1241_,
		_w1244_,
		_w1247_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w1246_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w1236_,
		_w1238_,
		_w1249_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w1248_,
		_w1249_,
		_w1250_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w972_,
		_w1090_,
		_w1251_
	);
	LUT2 #(
		.INIT('h2)
	) name293 (
		\u5_state_reg[7]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w1252_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		_w1251_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		\u5_state_reg[38]/NET0131 ,
		\u5_state_reg[39]/NET0131 ,
		_w1254_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		_w985_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w1256_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		_w984_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w1255_,
		_w1257_,
		_w1258_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		_w1119_,
		_w1258_,
		_w1259_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w1253_,
		_w1259_,
		_w1260_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		\u5_state_reg[20]/NET0131 ,
		_w1002_,
		_w1261_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		\u5_state_reg[21]/NET0131 ,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		_w1066_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		\u5_state_reg[60]/NET0131 ,
		\u5_state_reg[61]/NET0131 ,
		_w1264_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w964_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w1233_,
		_w1265_,
		_w1266_
	);
	LUT2 #(
		.INIT('h2)
	) name308 (
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		_w1267_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w981_,
		_w1267_,
		_w1268_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		_w1034_,
		_w1268_,
		_w1269_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w1266_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		\u5_state_reg[50]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w1271_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		_w1156_,
		_w1271_,
		_w1272_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w1263_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		_w1270_,
		_w1273_,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w1260_,
		_w1274_,
		_w1275_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		_w1250_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\u5_state_reg[5]/NET0131 ,
		_w979_,
		_w1277_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w1026_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w1034_,
		_w1278_,
		_w1279_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w968_,
		_w1030_,
		_w1280_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w1015_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w1282_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w1281_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w1279_,
		_w1283_,
		_w1284_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		_w1098_,
		_w1153_,
		_w1285_
	);
	LUT2 #(
		.INIT('h4)
	) name327 (
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w1286_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		_w1285_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		_w1284_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w1204_,
		_w1289_,
		_w1290_
	);
	LUT2 #(
		.INIT('h4)
	) name332 (
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w1291_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		_w1242_,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		_w1000_,
		_w1211_,
		_w1293_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w1294_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		_w1293_,
		_w1294_,
		_w1295_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w1290_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		_w1292_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w1288_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('h2)
	) name340 (
		\u5_state_reg[6]/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		_w1299_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w1091_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		\u5_state_reg[15]/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		_w1219_,
		_w1301_,
		_w1302_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w1300_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		_w1298_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		_w985_,
		_w1119_,
		_w1305_
	);
	LUT2 #(
		.INIT('h4)
	) name347 (
		\u5_state_reg[38]/NET0131 ,
		\u5_state_reg[39]/NET0131 ,
		_w1306_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w1308_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		_w1281_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w1307_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w1311_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		_w1285_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		_w1313_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		_w1112_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w1312_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		_w1310_,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		_w1190_,
		_w1195_,
		_w1317_
	);
	LUT2 #(
		.INIT('h8)
	) name359 (
		_w1218_,
		_w1317_,
		_w1318_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		_w1209_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		_w1232_,
		_w1316_,
		_w1320_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		_w1319_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		_w1304_,
		_w1321_,
		_w1322_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		_w1169_,
		_w1276_,
		_w1323_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		_w1322_,
		_w1323_,
		_w1324_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		_w1128_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1327_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w1326_,
		_w1327_,
		_w1328_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		_w1051_,
		_w1328_,
		_w1329_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		\u0_sp_tms_reg[10]/NET0131 ,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1331_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		\u5_state_reg[5]/NET0131 ,
		\u5_state_reg[6]/NET0131 ,
		_w1332_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		\u5_state_reg[1]/NET0131 ,
		_w1026_,
		_w1333_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w1196_,
		_w1333_,
		_w1334_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		_w996_,
		_w1030_,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		_w967_,
		_w1335_,
		_w1336_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		_w990_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		\u5_state_reg[33]/NET0131 ,
		_w991_,
		_w1338_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[36]/NET0131 ,
		_w1339_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		\u5_state_reg[37]/NET0131 ,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		\u5_state_reg[8]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w1341_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		_w978_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		_w969_,
		_w977_,
		_w1343_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		\u5_state_reg[7]/NET0131 ,
		_w970_,
		_w1345_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		_w1332_,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		_w964_,
		_w1008_,
		_w1347_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		_w1338_,
		_w1340_,
		_w1348_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		_w1347_,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		_w1005_,
		_w1346_,
		_w1350_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		_w1344_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		_w1334_,
		_w1349_,
		_w1352_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		_w1351_,
		_w1352_,
		_w1353_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		_w1337_,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w1331_,
		_w1354_,
		_w1355_
	);
	LUT2 #(
		.INIT('h2)
	) name397 (
		\u1_row_adr_reg[10]/P0001 ,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w1357_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		_w1293_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h2)
	) name400 (
		_w1124_,
		_w1358_,
		_w1359_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		_w1209_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		_w1361_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		_w1187_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		\u5_state_reg[7]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w1363_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		_w1251_,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w1362_,
		_w1364_,
		_w1365_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w1093_,
		_w1253_,
		_w1366_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w1108_,
		_w1263_,
		_w1367_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		_w1097_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w1365_,
		_w1366_,
		_w1369_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w1250_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w1360_,
		_w1371_,
		_w1372_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		\u0_sp_csc_reg[10]/NET0131 ,
		_w1051_,
		_w1373_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		\u0_csc_reg[10]/NET0131 ,
		_w1051_,
		_w1374_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w1373_,
		_w1374_,
		_w1375_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		_w1184_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w1377_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		wb_stb_i_pad,
		wb_we_i_pad,
		_w1378_
	);
	LUT2 #(
		.INIT('h2)
	) name420 (
		\u6_write_go_r1_reg/NET0131 ,
		_w1378_,
		_w1379_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w1380_
	);
	LUT2 #(
		.INIT('h4)
	) name422 (
		_w1049_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		_w1379_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		_w1377_,
		_w1382_,
		_w1383_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		_w1093_,
		_w1383_,
		_w1384_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		_w1376_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		_w1372_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		\u5_ap_en_reg/NET0131 ,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		_w1297_,
		_w1310_,
		_w1388_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		_w1078_,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w1259_,
		_w1266_,
		_w1391_
	);
	LUT2 #(
		.INIT('h4)
	) name433 (
		_w1230_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w1315_,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		_w1394_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		_w1212_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		_w1396_
	);
	LUT2 #(
		.INIT('h8)
	) name438 (
		_w1222_,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w1189_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		_w1399_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		_w1006_,
		_w1399_,
		_w1400_
	);
	LUT2 #(
		.INIT('h8)
	) name442 (
		_w1073_,
		_w1400_,
		_w1401_
	);
	LUT2 #(
		.INIT('h2)
	) name443 (
		_w1228_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w1169_,
		_w1402_,
		_w1403_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		_w1106_,
		_w1195_,
		_w1404_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w1272_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w1221_,
		_w1300_,
		_w1406_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		_w1395_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		_w1102_,
		_w1405_,
		_w1408_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		_w1288_,
		_w1390_,
		_w1409_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w1408_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		_w1088_,
		_w1407_,
		_w1411_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		_w1398_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		_w1388_,
		_w1410_,
		_w1413_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w1393_,
		_w1413_,
		_w1414_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		_w1412_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		_w1372_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h8)
	) name458 (
		_w1403_,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w1387_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h8)
	) name460 (
		\u5_tmr_done_reg/NET0131 ,
		_w1382_,
		_w1419_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		_w1253_,
		_w1419_,
		_w1420_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		_w1398_,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		_w1376_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w1217_,
		_w1423_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		\u5_tmr_done_reg/NET0131 ,
		_w1375_,
		_w1424_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		_w1302_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w1269_,
		_w1425_,
		_w1426_
	);
	LUT2 #(
		.INIT('h2)
	) name468 (
		\u5_cmd_a10_r_reg/P0001 ,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w1214_,
		_w1423_,
		_w1428_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		_w1077_,
		_w1428_,
		_w1429_
	);
	LUT2 #(
		.INIT('h4)
	) name471 (
		_w1427_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		_w1422_,
		_w1430_,
		_w1431_
	);
	LUT2 #(
		.INIT('h4)
	) name473 (
		_w1418_,
		_w1431_,
		_w1432_
	);
	LUT2 #(
		.INIT('h2)
	) name474 (
		_w1355_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w1329_,
		_w1356_,
		_w1434_
	);
	LUT2 #(
		.INIT('h4)
	) name476 (
		_w1433_,
		_w1434_,
		_w1435_
	);
	LUT2 #(
		.INIT('h2)
	) name477 (
		_w1062_,
		_w1330_,
		_w1436_
	);
	LUT2 #(
		.INIT('h4)
	) name478 (
		_w1435_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		_w1058_,
		_w1061_,
		_w1438_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		\u1_acs_addr_reg[10]/P0001 ,
		_w1438_,
		_w1439_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		_w1054_,
		_w1057_,
		_w1440_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		_w1061_,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		\u6_wr_hold_reg/NET0131 ,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		\wb_addr_i[12]_pad ,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		\u1_sram_addr_reg[10]/P0001 ,
		_w1442_,
		_w1444_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w1058_,
		_w1443_,
		_w1445_
	);
	LUT2 #(
		.INIT('h4)
	) name487 (
		_w1444_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w1439_,
		_w1447_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		_w1446_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h4)
	) name490 (
		_w1437_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		\u1_acs_addr_reg[0]/P0001 ,
		_w1438_,
		_w1450_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		\wb_addr_i[2]_pad ,
		_w1442_,
		_w1451_
	);
	LUT2 #(
		.INIT('h4)
	) name493 (
		\u1_sram_addr_reg[0]/P0001 ,
		_w1442_,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w1058_,
		_w1451_,
		_w1453_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		_w1452_,
		_w1453_,
		_w1454_
	);
	LUT2 #(
		.INIT('h4)
	) name496 (
		\u1_col_adr_reg[0]/P0001 ,
		_w1355_,
		_w1455_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		\u1_row_adr_reg[0]/P0001 ,
		_w1355_,
		_w1456_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		_w1455_,
		_w1456_,
		_w1457_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		_w1329_,
		_w1457_,
		_w1458_
	);
	LUT2 #(
		.INIT('h4)
	) name500 (
		\u0_sp_tms_reg[0]/NET0131 ,
		_w1329_,
		_w1459_
	);
	LUT2 #(
		.INIT('h2)
	) name501 (
		_w1062_,
		_w1458_,
		_w1460_
	);
	LUT2 #(
		.INIT('h4)
	) name502 (
		_w1459_,
		_w1460_,
		_w1461_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w1450_,
		_w1454_,
		_w1462_
	);
	LUT2 #(
		.INIT('h4)
	) name504 (
		_w1461_,
		_w1462_,
		_w1463_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		\u1_acs_addr_reg[11]/P0001 ,
		_w1438_,
		_w1464_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		\wb_addr_i[13]_pad ,
		_w1442_,
		_w1465_
	);
	LUT2 #(
		.INIT('h4)
	) name507 (
		\u1_sram_addr_reg[11]/P0001 ,
		_w1442_,
		_w1466_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w1058_,
		_w1465_,
		_w1467_
	);
	LUT2 #(
		.INIT('h4)
	) name509 (
		_w1466_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h4)
	) name510 (
		\u0_sp_tms_reg[11]/NET0131 ,
		_w1329_,
		_w1469_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\u1_row_adr_reg[11]/P0001 ,
		_w1355_,
		_w1470_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w1329_,
		_w1470_,
		_w1471_
	);
	LUT2 #(
		.INIT('h2)
	) name513 (
		_w1062_,
		_w1469_,
		_w1472_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		_w1471_,
		_w1472_,
		_w1473_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w1464_,
		_w1468_,
		_w1474_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w1473_,
		_w1474_,
		_w1475_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\u1_acs_addr_reg[12]/P0001 ,
		_w1438_,
		_w1476_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		\wb_addr_i[14]_pad ,
		_w1442_,
		_w1477_
	);
	LUT2 #(
		.INIT('h4)
	) name519 (
		\u1_sram_addr_reg[12]/P0001 ,
		_w1442_,
		_w1478_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		_w1058_,
		_w1477_,
		_w1479_
	);
	LUT2 #(
		.INIT('h4)
	) name521 (
		_w1478_,
		_w1479_,
		_w1480_
	);
	LUT2 #(
		.INIT('h4)
	) name522 (
		\u0_sp_tms_reg[12]/NET0131 ,
		_w1329_,
		_w1481_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		\u1_row_adr_reg[12]/P0001 ,
		_w1355_,
		_w1482_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w1329_,
		_w1482_,
		_w1483_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		_w1062_,
		_w1481_,
		_w1484_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w1483_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		_w1476_,
		_w1480_,
		_w1486_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		_w1485_,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		\u1_acs_addr_reg[1]/P0001 ,
		_w1438_,
		_w1488_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		\wb_addr_i[3]_pad ,
		_w1442_,
		_w1489_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		\u1_sram_addr_reg[1]/P0001 ,
		_w1442_,
		_w1490_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w1058_,
		_w1489_,
		_w1491_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		_w1490_,
		_w1491_,
		_w1492_
	);
	LUT2 #(
		.INIT('h4)
	) name534 (
		\u1_col_adr_reg[1]/P0001 ,
		_w1355_,
		_w1493_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		\u1_row_adr_reg[1]/P0001 ,
		_w1355_,
		_w1494_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w1493_,
		_w1494_,
		_w1495_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		_w1329_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		\u0_sp_tms_reg[1]/NET0131 ,
		_w1329_,
		_w1497_
	);
	LUT2 #(
		.INIT('h2)
	) name539 (
		_w1062_,
		_w1496_,
		_w1498_
	);
	LUT2 #(
		.INIT('h4)
	) name540 (
		_w1497_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w1488_,
		_w1492_,
		_w1500_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w1499_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		\u1_acs_addr_reg[2]/P0001 ,
		_w1438_,
		_w1502_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		\wb_addr_i[4]_pad ,
		_w1442_,
		_w1503_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		\u1_sram_addr_reg[2]/P0001 ,
		_w1442_,
		_w1504_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		_w1058_,
		_w1503_,
		_w1505_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		_w1504_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		\u1_col_adr_reg[2]/P0001 ,
		_w1355_,
		_w1507_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		\u1_row_adr_reg[2]/P0001 ,
		_w1355_,
		_w1508_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		_w1507_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		_w1329_,
		_w1509_,
		_w1510_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		\u0_sp_tms_reg[2]/NET0131 ,
		_w1329_,
		_w1511_
	);
	LUT2 #(
		.INIT('h2)
	) name553 (
		_w1062_,
		_w1510_,
		_w1512_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w1511_,
		_w1512_,
		_w1513_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w1502_,
		_w1506_,
		_w1514_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		_w1513_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		\u1_acs_addr_reg[3]/P0001 ,
		_w1438_,
		_w1516_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		\wb_addr_i[5]_pad ,
		_w1442_,
		_w1517_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		\u1_sram_addr_reg[3]/P0001 ,
		_w1442_,
		_w1518_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w1058_,
		_w1517_,
		_w1519_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		\u0_sp_tms_reg[3]/NET0131 ,
		_w1329_,
		_w1521_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		\u1_col_adr_reg[3]/P0001 ,
		_w1355_,
		_w1522_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		\u1_row_adr_reg[3]/P0001 ,
		_w1355_,
		_w1523_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		_w1522_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		_w1329_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		_w1062_,
		_w1521_,
		_w1526_
	);
	LUT2 #(
		.INIT('h4)
	) name568 (
		_w1525_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w1516_,
		_w1520_,
		_w1528_
	);
	LUT2 #(
		.INIT('h4)
	) name570 (
		_w1527_,
		_w1528_,
		_w1529_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		\u1_acs_addr_reg[4]/P0001 ,
		_w1438_,
		_w1530_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		\wb_addr_i[6]_pad ,
		_w1442_,
		_w1531_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		\u1_sram_addr_reg[4]/P0001 ,
		_w1442_,
		_w1532_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w1058_,
		_w1531_,
		_w1533_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		_w1532_,
		_w1533_,
		_w1534_
	);
	LUT2 #(
		.INIT('h4)
	) name576 (
		\u0_sp_tms_reg[4]/NET0131 ,
		_w1329_,
		_w1535_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		\u1_col_adr_reg[4]/P0001 ,
		_w1355_,
		_w1536_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		\u1_row_adr_reg[4]/P0001 ,
		_w1355_,
		_w1537_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w1329_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h2)
	) name581 (
		_w1062_,
		_w1535_,
		_w1540_
	);
	LUT2 #(
		.INIT('h4)
	) name582 (
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		_w1530_,
		_w1534_,
		_w1542_
	);
	LUT2 #(
		.INIT('h4)
	) name584 (
		_w1541_,
		_w1542_,
		_w1543_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		\u1_acs_addr_reg[5]/P0001 ,
		_w1438_,
		_w1544_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		\wb_addr_i[7]_pad ,
		_w1442_,
		_w1545_
	);
	LUT2 #(
		.INIT('h4)
	) name587 (
		\u1_sram_addr_reg[5]/P0001 ,
		_w1442_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w1058_,
		_w1545_,
		_w1547_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		_w1546_,
		_w1547_,
		_w1548_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		\u0_sp_tms_reg[5]/NET0131 ,
		_w1329_,
		_w1549_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		\u1_col_adr_reg[5]/P0001 ,
		_w1355_,
		_w1550_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		\u1_row_adr_reg[5]/P0001 ,
		_w1355_,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		_w1550_,
		_w1551_,
		_w1552_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		_w1329_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h2)
	) name595 (
		_w1062_,
		_w1549_,
		_w1554_
	);
	LUT2 #(
		.INIT('h4)
	) name596 (
		_w1553_,
		_w1554_,
		_w1555_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w1544_,
		_w1548_,
		_w1556_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		_w1555_,
		_w1556_,
		_w1557_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		\u1_acs_addr_reg[6]/P0001 ,
		_w1438_,
		_w1558_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		\wb_addr_i[8]_pad ,
		_w1442_,
		_w1559_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		\u1_sram_addr_reg[6]/P0001 ,
		_w1442_,
		_w1560_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		_w1058_,
		_w1559_,
		_w1561_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		_w1560_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h4)
	) name604 (
		\u0_sp_tms_reg[6]/NET0131 ,
		_w1329_,
		_w1563_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		\u1_col_adr_reg[6]/P0001 ,
		_w1355_,
		_w1564_
	);
	LUT2 #(
		.INIT('h1)
	) name606 (
		\u1_row_adr_reg[6]/P0001 ,
		_w1355_,
		_w1565_
	);
	LUT2 #(
		.INIT('h1)
	) name607 (
		_w1564_,
		_w1565_,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		_w1329_,
		_w1566_,
		_w1567_
	);
	LUT2 #(
		.INIT('h2)
	) name609 (
		_w1062_,
		_w1563_,
		_w1568_
	);
	LUT2 #(
		.INIT('h4)
	) name610 (
		_w1567_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w1558_,
		_w1562_,
		_w1570_
	);
	LUT2 #(
		.INIT('h4)
	) name612 (
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('h8)
	) name613 (
		\u1_acs_addr_reg[7]/P0001 ,
		_w1438_,
		_w1572_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		\wb_addr_i[9]_pad ,
		_w1442_,
		_w1573_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		\u1_sram_addr_reg[7]/P0001 ,
		_w1442_,
		_w1574_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		_w1058_,
		_w1573_,
		_w1575_
	);
	LUT2 #(
		.INIT('h4)
	) name617 (
		_w1574_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h4)
	) name618 (
		\u0_sp_tms_reg[7]/NET0131 ,
		_w1329_,
		_w1577_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		\u1_col_adr_reg[7]/P0001 ,
		_w1355_,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		\u1_row_adr_reg[7]/P0001 ,
		_w1355_,
		_w1579_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		_w1578_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		_w1329_,
		_w1580_,
		_w1581_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		_w1062_,
		_w1577_,
		_w1582_
	);
	LUT2 #(
		.INIT('h4)
	) name624 (
		_w1581_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		_w1572_,
		_w1576_,
		_w1584_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		_w1583_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h8)
	) name627 (
		\u1_acs_addr_reg[8]/P0001 ,
		_w1438_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		\wb_addr_i[10]_pad ,
		_w1442_,
		_w1587_
	);
	LUT2 #(
		.INIT('h4)
	) name629 (
		\u1_sram_addr_reg[8]/P0001 ,
		_w1442_,
		_w1588_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w1058_,
		_w1587_,
		_w1589_
	);
	LUT2 #(
		.INIT('h4)
	) name631 (
		_w1588_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h4)
	) name632 (
		\u0_sp_tms_reg[8]/NET0131 ,
		_w1329_,
		_w1591_
	);
	LUT2 #(
		.INIT('h4)
	) name633 (
		\u1_col_adr_reg[8]/P0001 ,
		_w1355_,
		_w1592_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		\u1_row_adr_reg[8]/P0001 ,
		_w1355_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w1592_,
		_w1593_,
		_w1594_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w1329_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h2)
	) name637 (
		_w1062_,
		_w1591_,
		_w1596_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		_w1595_,
		_w1596_,
		_w1597_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w1586_,
		_w1590_,
		_w1598_
	);
	LUT2 #(
		.INIT('h4)
	) name640 (
		_w1597_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		\u1_acs_addr_reg[9]/P0001 ,
		_w1438_,
		_w1600_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		\wb_addr_i[11]_pad ,
		_w1442_,
		_w1601_
	);
	LUT2 #(
		.INIT('h4)
	) name643 (
		\u1_sram_addr_reg[9]/P0001 ,
		_w1442_,
		_w1602_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w1058_,
		_w1601_,
		_w1603_
	);
	LUT2 #(
		.INIT('h4)
	) name645 (
		_w1602_,
		_w1603_,
		_w1604_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		\u1_col_adr_reg[9]/P0001 ,
		_w1355_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		\u1_row_adr_reg[9]/P0001 ,
		_w1355_,
		_w1606_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		_w1605_,
		_w1606_,
		_w1607_
	);
	LUT2 #(
		.INIT('h1)
	) name649 (
		_w1329_,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h4)
	) name650 (
		\u0_sp_tms_reg[9]/NET0131 ,
		_w1329_,
		_w1609_
	);
	LUT2 #(
		.INIT('h2)
	) name651 (
		_w1062_,
		_w1608_,
		_w1610_
	);
	LUT2 #(
		.INIT('h4)
	) name652 (
		_w1609_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w1600_,
		_w1604_,
		_w1612_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		_w1611_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h1)
	) name655 (
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		_w1614_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		_w1051_,
		_w1615_
	);
	LUT2 #(
		.INIT('h4)
	) name657 (
		\u0_cs_reg[0]/NET0131 ,
		_w1051_,
		_w1616_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		_w1615_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		_w1614_,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		\u0_u0_csc_reg[1]/NET0131 ,
		\u0_u0_csc_reg[2]/NET0131 ,
		_w1619_
	);
	LUT2 #(
		.INIT('h4)
	) name661 (
		\u0_u0_csc_reg[3]/NET0131 ,
		_w1619_,
		_w1620_
	);
	LUT2 #(
		.INIT('h8)
	) name662 (
		\u0_u0_csc_reg[0]/NET0131 ,
		_w1620_,
		_w1621_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		_w1614_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w1618_,
		_w1622_,
		_w1623_
	);
	LUT2 #(
		.INIT('h8)
	) name665 (
		\u5_cmd_del_reg[3]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1624_
	);
	LUT2 #(
		.INIT('h4)
	) name666 (
		\u5_cnt_reg/NET0131 ,
		_w1184_,
		_w1625_
	);
	LUT2 #(
		.INIT('h2)
	) name667 (
		\u5_cke_r_reg/NET0131 ,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		\u6_read_go_r1_reg/NET0131 ,
		_w1381_,
		_w1627_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		_w1382_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h2)
	) name670 (
		_w1377_,
		_w1628_,
		_w1629_
	);
	LUT2 #(
		.INIT('h2)
	) name671 (
		_w1625_,
		_w1629_,
		_w1630_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w1626_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		_w1358_,
		_w1362_,
		_w1632_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		_w1284_,
		_w1423_,
		_w1633_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w1217_,
		_w1279_,
		_w1634_
	);
	LUT2 #(
		.INIT('h1)
	) name676 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w1634_,
		_w1635_
	);
	LUT2 #(
		.INIT('h4)
	) name677 (
		\u4_rfr_req_reg/NET0131 ,
		_w1634_,
		_w1636_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		_w1284_,
		_w1635_,
		_w1637_
	);
	LUT2 #(
		.INIT('h4)
	) name679 (
		_w1636_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h2)
	) name680 (
		_w1632_,
		_w1633_,
		_w1639_
	);
	LUT2 #(
		.INIT('h4)
	) name681 (
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		\u5_mc_c_oe_reg/NET0131 ,
		_w1614_,
		_w1641_
	);
	LUT2 #(
		.INIT('h8)
	) name683 (
		_w1180_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		_w1640_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		\u5_burst_cnt_reg[0]/NET0131 ,
		\u5_burst_cnt_reg[1]/NET0131 ,
		_w1644_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		\u5_burst_cnt_reg[2]/NET0131 ,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		\u5_burst_cnt_reg[3]/NET0131 ,
		\u5_burst_cnt_reg[4]/NET0131 ,
		_w1646_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		\u5_burst_cnt_reg[5]/NET0131 ,
		\u5_burst_cnt_reg[6]/NET0131 ,
		_w1647_
	);
	LUT2 #(
		.INIT('h8)
	) name689 (
		_w1646_,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		_w1645_,
		_w1648_,
		_w1649_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		\u5_burst_cnt_reg[7]/NET0131 ,
		\u5_burst_cnt_reg[8]/NET0131 ,
		_w1650_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		_w1649_,
		_w1650_,
		_w1651_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		\u5_burst_cnt_reg[10]/NET0131 ,
		\u5_burst_cnt_reg[9]/NET0131 ,
		_w1652_
	);
	LUT2 #(
		.INIT('h8)
	) name694 (
		_w1651_,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w1643_,
		_w1653_,
		_w1654_
	);
	LUT2 #(
		.INIT('h8)
	) name696 (
		_w1184_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h4)
	) name697 (
		\u5_wb_write_go_r_reg/NET0131 ,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h4)
	) name698 (
		_w1631_,
		_w1656_,
		_w1657_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w1185_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h2)
	) name700 (
		_w1189_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h4)
	) name701 (
		_w1236_,
		_w1365_,
		_w1660_
	);
	LUT2 #(
		.INIT('h1)
	) name702 (
		_w1054_,
		_w1061_,
		_w1661_
	);
	LUT2 #(
		.INIT('h8)
	) name703 (
		_w1057_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h4)
	) name704 (
		_w1629_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		_w1382_,
		_w1629_,
		_w1664_
	);
	LUT2 #(
		.INIT('h8)
	) name706 (
		_w1440_,
		_w1664_,
		_w1665_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		_w1061_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		_w1663_,
		_w1666_,
		_w1667_
	);
	LUT2 #(
		.INIT('h2)
	) name709 (
		\u0_spec_req_cs_reg[1]/NET0131 ,
		_w1051_,
		_w1668_
	);
	LUT2 #(
		.INIT('h8)
	) name710 (
		\u0_cs_reg[1]/NET0131 ,
		_w1051_,
		_w1669_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w1668_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		_w1614_,
		_w1670_,
		_w1671_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		\u0_u1_csc_reg[1]/NET0131 ,
		\u0_u1_csc_reg[2]/NET0131 ,
		_w1672_
	);
	LUT2 #(
		.INIT('h4)
	) name714 (
		\u0_u1_csc_reg[3]/NET0131 ,
		_w1672_,
		_w1673_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		\u0_u1_csc_reg[0]/NET0131 ,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h4)
	) name716 (
		_w1614_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w1671_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h4)
	) name718 (
		_w1623_,
		_w1676_,
		_w1677_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		\u5_lookup_ready2_reg/NET0131 ,
		_w1677_,
		_w1678_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		_w1628_,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h2)
	) name721 (
		\u5_susp_req_r_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w1680_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		\u0_lmr_req_reg/NET0131 ,
		\u5_lookup_ready2_reg/NET0131 ,
		_w1681_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		\u0_init_req_reg/NET0131 ,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h4)
	) name724 (
		_w1680_,
		_w1682_,
		_w1683_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		\u4_rfr_req_reg/NET0131 ,
		_w1683_,
		_w1684_
	);
	LUT2 #(
		.INIT('h8)
	) name726 (
		_w1283_,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h8)
	) name727 (
		_w1679_,
		_w1685_,
		_w1686_
	);
	LUT2 #(
		.INIT('h4)
	) name728 (
		_w1667_,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name729 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1272_,
		_w1688_
	);
	LUT2 #(
		.INIT('h1)
	) name730 (
		_w1136_,
		_w1227_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		_w1244_,
		_w1292_,
		_w1690_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		\u0_tms_reg[19]/NET0131 ,
		_w1051_,
		_w1691_
	);
	LUT2 #(
		.INIT('h8)
	) name733 (
		_w1632_,
		_w1641_,
		_w1692_
	);
	LUT2 #(
		.INIT('h4)
	) name734 (
		_w1638_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h2)
	) name735 (
		\u0_sp_tms_reg[19]/NET0131 ,
		_w1051_,
		_w1694_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w1691_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		_w1693_,
		_w1695_,
		_w1696_
	);
	LUT2 #(
		.INIT('h8)
	) name738 (
		\u0_tms_reg[18]/NET0131 ,
		_w1051_,
		_w1697_
	);
	LUT2 #(
		.INIT('h2)
	) name739 (
		\u0_sp_tms_reg[18]/NET0131 ,
		_w1051_,
		_w1698_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		_w1697_,
		_w1698_,
		_w1699_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		_w1693_,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		\u0_tms_reg[17]/NET0131 ,
		_w1051_,
		_w1701_
	);
	LUT2 #(
		.INIT('h2)
	) name743 (
		\u0_sp_tms_reg[17]/NET0131 ,
		_w1051_,
		_w1702_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w1701_,
		_w1702_,
		_w1703_
	);
	LUT2 #(
		.INIT('h8)
	) name745 (
		_w1693_,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		\u0_tms_reg[16]/NET0131 ,
		_w1051_,
		_w1705_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		\u0_sp_tms_reg[16]/NET0131 ,
		_w1051_,
		_w1706_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h2)
	) name749 (
		_w1693_,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h8)
	) name750 (
		_w1696_,
		_w1700_,
		_w1709_
	);
	LUT2 #(
		.INIT('h8)
	) name751 (
		_w1704_,
		_w1708_,
		_w1710_
	);
	LUT2 #(
		.INIT('h8)
	) name752 (
		_w1709_,
		_w1710_,
		_w1711_
	);
	LUT2 #(
		.INIT('h2)
	) name753 (
		_w1087_,
		_w1711_,
		_w1712_
	);
	LUT2 #(
		.INIT('h2)
	) name754 (
		_w1103_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w1390_,
		_w1395_,
		_w1714_
	);
	LUT2 #(
		.INIT('h4)
	) name756 (
		\u5_wb_wait_r_reg/P0001 ,
		_w1300_,
		_w1715_
	);
	LUT2 #(
		.INIT('h8)
	) name757 (
		_w1302_,
		_w1424_,
		_w1716_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		_w1077_,
		_w1221_,
		_w1717_
	);
	LUT2 #(
		.INIT('h2)
	) name759 (
		_w1218_,
		_w1716_,
		_w1718_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		_w1717_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h4)
	) name761 (
		_w1715_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h4)
	) name762 (
		\u5_tmr_done_reg/NET0131 ,
		_w1238_,
		_w1721_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		_w1146_,
		_w1401_,
		_w1722_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w1358_,
		_w1688_,
		_w1723_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		_w1722_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h2)
	) name766 (
		_w1151_,
		_w1307_,
		_w1725_
	);
	LUT2 #(
		.INIT('h4)
	) name767 (
		_w1397_,
		_w1689_,
		_w1726_
	);
	LUT2 #(
		.INIT('h8)
	) name768 (
		_w1725_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h8)
	) name769 (
		_w1660_,
		_w1724_,
		_w1728_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		_w1690_,
		_w1714_,
		_w1729_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		_w1721_,
		_w1729_,
		_w1730_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		_w1727_,
		_w1728_,
		_w1731_
	);
	LUT2 #(
		.INIT('h2)
	) name773 (
		_w1393_,
		_w1687_,
		_w1732_
	);
	LUT2 #(
		.INIT('h8)
	) name774 (
		_w1731_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('h8)
	) name775 (
		_w1720_,
		_w1730_,
		_w1734_
	);
	LUT2 #(
		.INIT('h8)
	) name776 (
		_w1733_,
		_w1734_,
		_w1735_
	);
	LUT2 #(
		.INIT('h8)
	) name777 (
		_w1713_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h4)
	) name778 (
		_w1659_,
		_w1736_,
		_w1737_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1737_,
		_w1738_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w1624_,
		_w1738_,
		_w1739_
	);
	LUT2 #(
		.INIT('h2)
	) name781 (
		_w1623_,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		_w1676_,
		_w1739_,
		_w1741_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		_w1679_,
		_w1683_,
		_w1742_
	);
	LUT2 #(
		.INIT('h8)
	) name784 (
		_w1383_,
		_w1661_,
		_w1743_
	);
	LUT2 #(
		.INIT('h2)
	) name785 (
		_w1057_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		_w1742_,
		_w1744_,
		_w1745_
	);
	LUT2 #(
		.INIT('h2)
	) name787 (
		_w1283_,
		_w1745_,
		_w1746_
	);
	LUT2 #(
		.INIT('h8)
	) name788 (
		\u4_rfr_req_reg/NET0131 ,
		_w1283_,
		_w1747_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		\u5_tmr_done_reg/NET0131 ,
		_w1238_,
		_w1748_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		_w1279_,
		_w1287_,
		_w1749_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		_w1631_,
		_w1656_,
		_w1750_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		_w1190_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		_w1189_,
		_w1631_,
		_w1752_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		_w1185_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w1195_,
		_w1747_,
		_w1754_
	);
	LUT2 #(
		.INIT('h4)
	) name796 (
		_w1300_,
		_w1754_,
		_w1755_
	);
	LUT2 #(
		.INIT('h4)
	) name797 (
		_w1314_,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		_w1109_,
		_w1260_,
		_w1757_
	);
	LUT2 #(
		.INIT('h4)
	) name799 (
		_w1425_,
		_w1749_,
		_w1758_
	);
	LUT2 #(
		.INIT('h8)
	) name800 (
		_w1757_,
		_w1758_,
		_w1759_
	);
	LUT2 #(
		.INIT('h8)
	) name801 (
		_w1274_,
		_w1756_,
		_w1760_
	);
	LUT2 #(
		.INIT('h2)
	) name802 (
		_w1660_,
		_w1748_,
		_w1761_
	);
	LUT2 #(
		.INIT('h8)
	) name803 (
		_w1760_,
		_w1761_,
		_w1762_
	);
	LUT2 #(
		.INIT('h8)
	) name804 (
		_w1094_,
		_w1759_,
		_w1763_
	);
	LUT2 #(
		.INIT('h8)
	) name805 (
		_w1248_,
		_w1388_,
		_w1764_
	);
	LUT2 #(
		.INIT('h8)
	) name806 (
		_w1763_,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h4)
	) name807 (
		_w1746_,
		_w1762_,
		_w1766_
	);
	LUT2 #(
		.INIT('h4)
	) name808 (
		_w1753_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h8)
	) name809 (
		_w1360_,
		_w1765_,
		_w1768_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		_w1767_,
		_w1768_,
		_w1769_
	);
	LUT2 #(
		.INIT('h8)
	) name811 (
		_w1403_,
		_w1769_,
		_w1770_
	);
	LUT2 #(
		.INIT('h4)
	) name812 (
		_w1751_,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		\u5_mc_le_reg/NET0131 ,
		_w1737_,
		_w1772_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_mc_le_reg/NET0131 ,
		_w1773_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h8)
	) name816 (
		_w1383_,
		_w1662_,
		_w1775_
	);
	LUT2 #(
		.INIT('h8)
	) name817 (
		_w1686_,
		_w1775_,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		_w1102_,
		_w1776_,
		_w1777_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		_w1693_,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h2)
	) name820 (
		\u0_sp_tms_reg[14]/NET0131 ,
		_w1051_,
		_w1779_
	);
	LUT2 #(
		.INIT('h8)
	) name821 (
		\u0_tms_reg[14]/NET0131 ,
		_w1051_,
		_w1780_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w1779_,
		_w1780_,
		_w1781_
	);
	LUT2 #(
		.INIT('h4)
	) name823 (
		_w1777_,
		_w1781_,
		_w1782_
	);
	LUT2 #(
		.INIT('h2)
	) name824 (
		_w1141_,
		_w1266_,
		_w1783_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		\u5_tmr_done_reg/NET0131 ,
		_w1266_,
		_w1784_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w1783_,
		_w1784_,
		_w1785_
	);
	LUT2 #(
		.INIT('h2)
	) name827 (
		\u0_sp_tms_reg[10]/NET0131 ,
		_w1051_,
		_w1786_
	);
	LUT2 #(
		.INIT('h8)
	) name828 (
		\u0_tms_reg[10]/NET0131 ,
		_w1051_,
		_w1787_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w1786_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h4)
	) name830 (
		_w1785_,
		_w1788_,
		_w1789_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		\u5_state_reg[13]/NET0131 ,
		\u5_state_reg[14]/NET0131 ,
		_w1790_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		\u0_tms_reg[22]/NET0131 ,
		_w1051_,
		_w1791_
	);
	LUT2 #(
		.INIT('h2)
	) name833 (
		\u0_sp_tms_reg[22]/NET0131 ,
		_w1051_,
		_w1792_
	);
	LUT2 #(
		.INIT('h1)
	) name834 (
		_w1791_,
		_w1792_,
		_w1793_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		_w1693_,
		_w1793_,
		_w1794_
	);
	LUT2 #(
		.INIT('h4)
	) name836 (
		\u0_tms_reg[21]/NET0131 ,
		_w1051_,
		_w1795_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		\u0_sp_tms_reg[21]/NET0131 ,
		_w1051_,
		_w1796_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		_w1795_,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		_w1693_,
		_w1797_,
		_w1798_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		_w1708_,
		_w1798_,
		_w1799_
	);
	LUT2 #(
		.INIT('h8)
	) name841 (
		_w1708_,
		_w1798_,
		_w1800_
	);
	LUT2 #(
		.INIT('h2)
	) name842 (
		\u0_sp_tms_reg[15]/NET0131 ,
		_w1051_,
		_w1801_
	);
	LUT2 #(
		.INIT('h8)
	) name843 (
		\u0_tms_reg[15]/NET0131 ,
		_w1051_,
		_w1802_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		_w1801_,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('h2)
	) name845 (
		\u0_sp_tms_reg[20]/NET0131 ,
		_w1051_,
		_w1804_
	);
	LUT2 #(
		.INIT('h8)
	) name846 (
		\u0_tms_reg[20]/NET0131 ,
		_w1051_,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		_w1804_,
		_w1805_,
		_w1806_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w1803_,
		_w1806_,
		_w1807_
	);
	LUT2 #(
		.INIT('h2)
	) name849 (
		_w1693_,
		_w1807_,
		_w1808_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		_w1800_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w1799_,
		_w1809_,
		_w1810_
	);
	LUT2 #(
		.INIT('h8)
	) name852 (
		_w1794_,
		_w1810_,
		_w1811_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w1794_,
		_w1810_,
		_w1812_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w1811_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h1)
	) name855 (
		_w1790_,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h4)
	) name856 (
		_w1061_,
		_w1665_,
		_w1815_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		_w1686_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h1)
	) name858 (
		_w1236_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		\u5_state_reg[17]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w1818_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		\u5_state_reg[24]/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		_w1818_,
		_w1819_,
		_w1820_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		\u5_timer_reg[2]/NET0131 ,
		\u5_timer_reg[3]/NET0131 ,
		_w1821_
	);
	LUT2 #(
		.INIT('h1)
	) name863 (
		\u5_timer_reg[4]/NET0131 ,
		\u5_timer_reg[5]/NET0131 ,
		_w1822_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		_w1821_,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		\u5_timer_reg[0]/NET0131 ,
		\u5_timer_reg[1]/NET0131 ,
		_w1824_
	);
	LUT2 #(
		.INIT('h4)
	) name866 (
		\u5_timer_reg[6]/NET0131 ,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h8)
	) name867 (
		_w1823_,
		_w1825_,
		_w1826_
	);
	LUT2 #(
		.INIT('h4)
	) name868 (
		\u5_timer_reg[7]/NET0131 ,
		_w1826_,
		_w1827_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		\u5_mc_le_reg/NET0131 ,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h4)
	) name870 (
		\u5_timer_reg[0]/NET0131 ,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h4)
	) name871 (
		\u5_timer_reg[1]/NET0131 ,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		\u5_timer_reg[2]/NET0131 ,
		_w1830_,
		_w1831_
	);
	LUT2 #(
		.INIT('h2)
	) name873 (
		\u5_timer_reg[2]/NET0131 ,
		_w1830_,
		_w1832_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		_w1010_,
		_w1831_,
		_w1833_
	);
	LUT2 #(
		.INIT('h4)
	) name875 (
		_w1832_,
		_w1833_,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		\u5_state_reg[35]/NET0131 ,
		_w1834_,
		_w1835_
	);
	LUT2 #(
		.INIT('h2)
	) name877 (
		_w1820_,
		_w1835_,
		_w1836_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		\u5_state_reg[9]/NET0131 ,
		_w1720_,
		_w1837_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		\u0_sp_tms_reg[26]/NET0131 ,
		_w1051_,
		_w1838_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		\u0_tms_reg[26]/NET0131 ,
		_w1051_,
		_w1839_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w1820_,
		_w1838_,
		_w1840_
	);
	LUT2 #(
		.INIT('h4)
	) name882 (
		_w1839_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		_w1693_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w1836_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		_w1837_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('h8)
	) name886 (
		_w1715_,
		_w1719_,
		_w1845_
	);
	LUT2 #(
		.INIT('h4)
	) name887 (
		_w1696_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name888 (
		_w1719_,
		_w1794_,
		_w1847_
	);
	LUT2 #(
		.INIT('h2)
	) name889 (
		_w1790_,
		_w1846_,
		_w1848_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		_w1847_,
		_w1848_,
		_w1849_
	);
	LUT2 #(
		.INIT('h4)
	) name891 (
		_w1844_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h2)
	) name892 (
		_w1817_,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h4)
	) name893 (
		_w1814_,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w1175_,
		_w1693_,
		_w1853_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w1817_,
		_w1853_,
		_w1854_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		_w1785_,
		_w1854_,
		_w1855_
	);
	LUT2 #(
		.INIT('h4)
	) name897 (
		_w1852_,
		_w1855_,
		_w1856_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		_w1789_,
		_w1856_,
		_w1857_
	);
	LUT2 #(
		.INIT('h1)
	) name899 (
		_w1693_,
		_w1785_,
		_w1858_
	);
	LUT2 #(
		.INIT('h2)
	) name900 (
		_w1777_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h4)
	) name901 (
		_w1857_,
		_w1859_,
		_w1860_
	);
	LUT2 #(
		.INIT('h1)
	) name902 (
		_w1782_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w1778_,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h1)
	) name904 (
		_w1238_,
		_w1266_,
		_w1863_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		\u5_tmr_done_reg/NET0131 ,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h2)
	) name906 (
		_w1123_,
		_w1158_,
		_w1865_
	);
	LUT2 #(
		.INIT('h4)
	) name907 (
		\u5_mem_ack_r_reg/NET0131 ,
		_w1383_,
		_w1866_
	);
	LUT2 #(
		.INIT('h8)
	) name908 (
		_w1093_,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h1)
	) name909 (
		_w1864_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		_w1865_,
		_w1868_,
		_w1869_
	);
	LUT2 #(
		.INIT('h8)
	) name911 (
		wb_stb_i_pad,
		wb_we_i_pad,
		_w1870_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_ack_cnt_reg[1]/NET0131 ,
		_w1871_
	);
	LUT2 #(
		.INIT('h4)
	) name913 (
		\u5_ack_cnt_reg[2]/NET0131 ,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h4)
	) name914 (
		\u5_ack_cnt_reg[3]/NET0131 ,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('h2)
	) name915 (
		_w1627_,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		\u5_mem_ack_r_reg/NET0131 ,
		_w1629_,
		_w1875_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		_w1870_,
		_w1874_,
		_w1876_
	);
	LUT2 #(
		.INIT('h8)
	) name918 (
		_w1875_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h8)
	) name919 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1866_,
		_w1878_
	);
	LUT2 #(
		.INIT('h8)
	) name920 (
		_w1189_,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		_w1654_,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h8)
	) name922 (
		_w1383_,
		_w1441_,
		_w1881_
	);
	LUT2 #(
		.INIT('h8)
	) name923 (
		_w1686_,
		_w1881_,
		_w1882_
	);
	LUT2 #(
		.INIT('h8)
	) name924 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1312_,
		_w1883_
	);
	LUT2 #(
		.INIT('h8)
	) name925 (
		_w1866_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h4)
	) name926 (
		\u5_mem_ack_r_reg/NET0131 ,
		_w1420_,
		_w1885_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h4)
	) name928 (
		_w1882_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h8)
	) name929 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1397_,
		_w1888_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1866_,
		_w1889_
	);
	LUT2 #(
		.INIT('h8)
	) name931 (
		_w1888_,
		_w1889_,
		_w1890_
	);
	LUT2 #(
		.INIT('h8)
	) name932 (
		_w1654_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('h4)
	) name933 (
		_w1877_,
		_w1887_,
		_w1892_
	);
	LUT2 #(
		.INIT('h8)
	) name934 (
		_w1869_,
		_w1892_,
		_w1893_
	);
	LUT2 #(
		.INIT('h4)
	) name935 (
		_w1880_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('h4)
	) name936 (
		_w1891_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		_w1628_,
		_w1895_,
		_w1896_
	);
	LUT2 #(
		.INIT('h1)
	) name938 (
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		_w1897_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		_w1898_
	);
	LUT2 #(
		.INIT('h8)
	) name940 (
		_w1897_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		\u3_u0_r0_reg[13]/P0001 ,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h4)
	) name942 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		_w1901_
	);
	LUT2 #(
		.INIT('h8)
	) name943 (
		_w1897_,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		\u3_u0_r1_reg[13]/P0001 ,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		_w1904_
	);
	LUT2 #(
		.INIT('h4)
	) name946 (
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		_w1905_
	);
	LUT2 #(
		.INIT('h8)
	) name947 (
		_w1904_,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		\u3_u0_r3_reg[13]/P0001 ,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h2)
	) name949 (
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		_w1908_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		_w1904_,
		_w1908_,
		_w1909_
	);
	LUT2 #(
		.INIT('h8)
	) name951 (
		\u3_u0_r2_reg[13]/P0001 ,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h1)
	) name952 (
		_w1900_,
		_w1903_,
		_w1911_
	);
	LUT2 #(
		.INIT('h1)
	) name953 (
		_w1907_,
		_w1910_,
		_w1912_
	);
	LUT2 #(
		.INIT('h8)
	) name954 (
		_w1911_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h8)
	) name955 (
		\u3_u0_r0_reg[9]/P0001 ,
		_w1899_,
		_w1914_
	);
	LUT2 #(
		.INIT('h8)
	) name956 (
		\u3_u0_r1_reg[9]/P0001 ,
		_w1902_,
		_w1915_
	);
	LUT2 #(
		.INIT('h8)
	) name957 (
		\u3_u0_r3_reg[9]/P0001 ,
		_w1906_,
		_w1916_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		\u3_u0_r2_reg[9]/P0001 ,
		_w1909_,
		_w1917_
	);
	LUT2 #(
		.INIT('h1)
	) name959 (
		_w1914_,
		_w1915_,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		_w1916_,
		_w1917_,
		_w1919_
	);
	LUT2 #(
		.INIT('h8)
	) name961 (
		_w1918_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h2)
	) name962 (
		_w1913_,
		_w1920_,
		_w1921_
	);
	LUT2 #(
		.INIT('h4)
	) name963 (
		_w1913_,
		_w1920_,
		_w1922_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		_w1921_,
		_w1922_,
		_w1923_
	);
	LUT2 #(
		.INIT('h8)
	) name965 (
		\u3_u0_r0_reg[14]/P0001 ,
		_w1899_,
		_w1924_
	);
	LUT2 #(
		.INIT('h8)
	) name966 (
		\u3_u0_r1_reg[14]/P0001 ,
		_w1902_,
		_w1925_
	);
	LUT2 #(
		.INIT('h8)
	) name967 (
		\u3_u0_r3_reg[14]/P0001 ,
		_w1906_,
		_w1926_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		\u3_u0_r2_reg[14]/P0001 ,
		_w1909_,
		_w1927_
	);
	LUT2 #(
		.INIT('h1)
	) name969 (
		_w1924_,
		_w1925_,
		_w1928_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		_w1926_,
		_w1927_,
		_w1929_
	);
	LUT2 #(
		.INIT('h8)
	) name971 (
		_w1928_,
		_w1929_,
		_w1930_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		\u3_u0_r0_reg[11]/P0001 ,
		_w1899_,
		_w1931_
	);
	LUT2 #(
		.INIT('h8)
	) name973 (
		\u3_u0_r1_reg[11]/P0001 ,
		_w1902_,
		_w1932_
	);
	LUT2 #(
		.INIT('h8)
	) name974 (
		\u3_u0_r3_reg[11]/P0001 ,
		_w1906_,
		_w1933_
	);
	LUT2 #(
		.INIT('h8)
	) name975 (
		\u3_u0_r2_reg[11]/P0001 ,
		_w1909_,
		_w1934_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		_w1931_,
		_w1932_,
		_w1935_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		_w1933_,
		_w1934_,
		_w1936_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		_w1935_,
		_w1936_,
		_w1937_
	);
	LUT2 #(
		.INIT('h8)
	) name979 (
		\u3_u0_r0_reg[12]/P0001 ,
		_w1899_,
		_w1938_
	);
	LUT2 #(
		.INIT('h8)
	) name980 (
		\u3_u0_r1_reg[12]/P0001 ,
		_w1902_,
		_w1939_
	);
	LUT2 #(
		.INIT('h8)
	) name981 (
		\u3_u0_r3_reg[12]/P0001 ,
		_w1906_,
		_w1940_
	);
	LUT2 #(
		.INIT('h8)
	) name982 (
		\u3_u0_r2_reg[12]/P0001 ,
		_w1909_,
		_w1941_
	);
	LUT2 #(
		.INIT('h1)
	) name983 (
		_w1938_,
		_w1939_,
		_w1942_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		_w1940_,
		_w1941_,
		_w1943_
	);
	LUT2 #(
		.INIT('h8)
	) name985 (
		_w1942_,
		_w1943_,
		_w1944_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		_w1937_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		_w1937_,
		_w1944_,
		_w1946_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		_w1945_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h2)
	) name989 (
		_w1930_,
		_w1947_,
		_w1948_
	);
	LUT2 #(
		.INIT('h4)
	) name990 (
		_w1930_,
		_w1947_,
		_w1949_
	);
	LUT2 #(
		.INIT('h1)
	) name991 (
		_w1948_,
		_w1949_,
		_w1950_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		_w1923_,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('h1)
	) name993 (
		_w1923_,
		_w1950_,
		_w1952_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w1951_,
		_w1952_,
		_w1953_
	);
	LUT2 #(
		.INIT('h8)
	) name995 (
		\u3_u0_r0_reg[8]/P0001 ,
		_w1899_,
		_w1954_
	);
	LUT2 #(
		.INIT('h8)
	) name996 (
		\u3_u0_r1_reg[8]/P0001 ,
		_w1902_,
		_w1955_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		\u3_u0_r3_reg[8]/P0001 ,
		_w1906_,
		_w1956_
	);
	LUT2 #(
		.INIT('h8)
	) name998 (
		\u3_u0_r2_reg[8]/P0001 ,
		_w1909_,
		_w1957_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		_w1954_,
		_w1955_,
		_w1958_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w1956_,
		_w1957_,
		_w1959_
	);
	LUT2 #(
		.INIT('h8)
	) name1001 (
		_w1958_,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('h8)
	) name1002 (
		\u3_u0_r0_reg[15]/P0001 ,
		_w1899_,
		_w1961_
	);
	LUT2 #(
		.INIT('h8)
	) name1003 (
		\u3_u0_r1_reg[15]/P0001 ,
		_w1902_,
		_w1962_
	);
	LUT2 #(
		.INIT('h8)
	) name1004 (
		\u3_u0_r3_reg[15]/P0001 ,
		_w1906_,
		_w1963_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		\u3_u0_r2_reg[15]/P0001 ,
		_w1909_,
		_w1964_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		_w1961_,
		_w1962_,
		_w1965_
	);
	LUT2 #(
		.INIT('h1)
	) name1007 (
		_w1963_,
		_w1964_,
		_w1966_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		_w1965_,
		_w1966_,
		_w1967_
	);
	LUT2 #(
		.INIT('h2)
	) name1009 (
		_w1960_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		_w1960_,
		_w1967_,
		_w1969_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w1968_,
		_w1969_,
		_w1970_
	);
	LUT2 #(
		.INIT('h8)
	) name1012 (
		\u3_u0_r0_reg[33]/P0001 ,
		_w1899_,
		_w1971_
	);
	LUT2 #(
		.INIT('h8)
	) name1013 (
		\u3_u0_r1_reg[33]/P0001 ,
		_w1902_,
		_w1972_
	);
	LUT2 #(
		.INIT('h8)
	) name1014 (
		\u3_u0_r3_reg[33]/P0001 ,
		_w1906_,
		_w1973_
	);
	LUT2 #(
		.INIT('h8)
	) name1015 (
		\u3_u0_r2_reg[33]/P0001 ,
		_w1909_,
		_w1974_
	);
	LUT2 #(
		.INIT('h1)
	) name1016 (
		_w1971_,
		_w1972_,
		_w1975_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w1973_,
		_w1974_,
		_w1976_
	);
	LUT2 #(
		.INIT('h8)
	) name1018 (
		_w1975_,
		_w1976_,
		_w1977_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		\u3_u0_r0_reg[10]/P0001 ,
		_w1899_,
		_w1978_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		\u3_u0_r1_reg[10]/P0001 ,
		_w1902_,
		_w1979_
	);
	LUT2 #(
		.INIT('h8)
	) name1021 (
		\u3_u0_r3_reg[10]/P0001 ,
		_w1906_,
		_w1980_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		\u3_u0_r2_reg[10]/P0001 ,
		_w1909_,
		_w1981_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		_w1978_,
		_w1979_,
		_w1982_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w1980_,
		_w1981_,
		_w1983_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		_w1982_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h2)
	) name1026 (
		_w1977_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('h4)
	) name1027 (
		_w1977_,
		_w1984_,
		_w1986_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		_w1985_,
		_w1986_,
		_w1987_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		_w1970_,
		_w1987_,
		_w1988_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		_w1970_,
		_w1987_,
		_w1989_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w1988_,
		_w1989_,
		_w1990_
	);
	LUT2 #(
		.INIT('h4)
	) name1032 (
		_w1953_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('h2)
	) name1033 (
		_w1953_,
		_w1990_,
		_w1992_
	);
	LUT2 #(
		.INIT('h2)
	) name1034 (
		\wb_sel_i[1]_pad ,
		_w1991_,
		_w1993_
	);
	LUT2 #(
		.INIT('h4)
	) name1035 (
		_w1992_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		\u3_u0_r0_reg[30]/P0001 ,
		_w1899_,
		_w1995_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		\u3_u0_r1_reg[30]/P0001 ,
		_w1902_,
		_w1996_
	);
	LUT2 #(
		.INIT('h8)
	) name1038 (
		\u3_u0_r3_reg[30]/P0001 ,
		_w1906_,
		_w1997_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		\u3_u0_r2_reg[30]/P0001 ,
		_w1909_,
		_w1998_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		_w1995_,
		_w1996_,
		_w1999_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w1997_,
		_w1998_,
		_w2000_
	);
	LUT2 #(
		.INIT('h8)
	) name1042 (
		_w1999_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h8)
	) name1043 (
		\u3_u0_r3_reg[29]/P0001 ,
		_w1906_,
		_w2002_
	);
	LUT2 #(
		.INIT('h8)
	) name1044 (
		\u3_u0_r2_reg[29]/P0001 ,
		_w1909_,
		_w2003_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		\u3_u0_r1_reg[29]/P0001 ,
		_w1902_,
		_w2004_
	);
	LUT2 #(
		.INIT('h8)
	) name1046 (
		\u3_u0_r0_reg[29]/P0001 ,
		_w1899_,
		_w2005_
	);
	LUT2 #(
		.INIT('h1)
	) name1047 (
		_w2002_,
		_w2003_,
		_w2006_
	);
	LUT2 #(
		.INIT('h1)
	) name1048 (
		_w2004_,
		_w2005_,
		_w2007_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		_w2006_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		_w2001_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h4)
	) name1051 (
		_w2001_,
		_w2008_,
		_w2010_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w2009_,
		_w2010_,
		_w2011_
	);
	LUT2 #(
		.INIT('h8)
	) name1053 (
		\u3_u0_r0_reg[27]/P0001 ,
		_w1899_,
		_w2012_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		\u3_u0_r3_reg[27]/P0001 ,
		_w1906_,
		_w2013_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		\u3_u0_r1_reg[27]/P0001 ,
		_w1902_,
		_w2014_
	);
	LUT2 #(
		.INIT('h8)
	) name1056 (
		\u3_u0_r2_reg[27]/P0001 ,
		_w1909_,
		_w2015_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		_w2012_,
		_w2013_,
		_w2016_
	);
	LUT2 #(
		.INIT('h1)
	) name1058 (
		_w2014_,
		_w2015_,
		_w2017_
	);
	LUT2 #(
		.INIT('h8)
	) name1059 (
		_w2016_,
		_w2017_,
		_w2018_
	);
	LUT2 #(
		.INIT('h8)
	) name1060 (
		\u3_u0_r0_reg[25]/P0001 ,
		_w1899_,
		_w2019_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		\u3_u0_r1_reg[25]/P0001 ,
		_w1902_,
		_w2020_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		\u3_u0_r3_reg[25]/P0001 ,
		_w1906_,
		_w2021_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		\u3_u0_r2_reg[25]/P0001 ,
		_w1909_,
		_w2022_
	);
	LUT2 #(
		.INIT('h1)
	) name1064 (
		_w2019_,
		_w2020_,
		_w2023_
	);
	LUT2 #(
		.INIT('h1)
	) name1065 (
		_w2021_,
		_w2022_,
		_w2024_
	);
	LUT2 #(
		.INIT('h8)
	) name1066 (
		_w2023_,
		_w2024_,
		_w2025_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		\u3_u0_r0_reg[28]/P0001 ,
		_w1899_,
		_w2026_
	);
	LUT2 #(
		.INIT('h8)
	) name1068 (
		\u3_u0_r1_reg[28]/P0001 ,
		_w1902_,
		_w2027_
	);
	LUT2 #(
		.INIT('h8)
	) name1069 (
		\u3_u0_r3_reg[28]/P0001 ,
		_w1906_,
		_w2028_
	);
	LUT2 #(
		.INIT('h8)
	) name1070 (
		\u3_u0_r2_reg[28]/P0001 ,
		_w1909_,
		_w2029_
	);
	LUT2 #(
		.INIT('h1)
	) name1071 (
		_w2026_,
		_w2027_,
		_w2030_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w2028_,
		_w2029_,
		_w2031_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		_w2030_,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h1)
	) name1074 (
		_w2025_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h8)
	) name1075 (
		_w2025_,
		_w2032_,
		_w2034_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w2033_,
		_w2034_,
		_w2035_
	);
	LUT2 #(
		.INIT('h2)
	) name1077 (
		_w2018_,
		_w2035_,
		_w2036_
	);
	LUT2 #(
		.INIT('h4)
	) name1078 (
		_w2018_,
		_w2035_,
		_w2037_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w2036_,
		_w2037_,
		_w2038_
	);
	LUT2 #(
		.INIT('h8)
	) name1080 (
		_w2011_,
		_w2038_,
		_w2039_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w2011_,
		_w2038_,
		_w2040_
	);
	LUT2 #(
		.INIT('h1)
	) name1082 (
		_w2039_,
		_w2040_,
		_w2041_
	);
	LUT2 #(
		.INIT('h8)
	) name1083 (
		\u3_u0_r0_reg[24]/P0001 ,
		_w1899_,
		_w2042_
	);
	LUT2 #(
		.INIT('h8)
	) name1084 (
		\u3_u0_r2_reg[24]/P0001 ,
		_w1909_,
		_w2043_
	);
	LUT2 #(
		.INIT('h8)
	) name1085 (
		\u3_u0_r1_reg[24]/P0001 ,
		_w1902_,
		_w2044_
	);
	LUT2 #(
		.INIT('h8)
	) name1086 (
		\u3_u0_r3_reg[24]/P0001 ,
		_w1906_,
		_w2045_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		_w2042_,
		_w2043_,
		_w2046_
	);
	LUT2 #(
		.INIT('h1)
	) name1088 (
		_w2044_,
		_w2045_,
		_w2047_
	);
	LUT2 #(
		.INIT('h8)
	) name1089 (
		_w2046_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h8)
	) name1090 (
		\u3_u0_r0_reg[31]/P0001 ,
		_w1899_,
		_w2049_
	);
	LUT2 #(
		.INIT('h8)
	) name1091 (
		\u3_u0_r1_reg[31]/P0001 ,
		_w1902_,
		_w2050_
	);
	LUT2 #(
		.INIT('h8)
	) name1092 (
		\u3_u0_r3_reg[31]/P0001 ,
		_w1906_,
		_w2051_
	);
	LUT2 #(
		.INIT('h8)
	) name1093 (
		\u3_u0_r2_reg[31]/P0001 ,
		_w1909_,
		_w2052_
	);
	LUT2 #(
		.INIT('h1)
	) name1094 (
		_w2049_,
		_w2050_,
		_w2053_
	);
	LUT2 #(
		.INIT('h1)
	) name1095 (
		_w2051_,
		_w2052_,
		_w2054_
	);
	LUT2 #(
		.INIT('h8)
	) name1096 (
		_w2053_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h2)
	) name1097 (
		_w2048_,
		_w2055_,
		_w2056_
	);
	LUT2 #(
		.INIT('h4)
	) name1098 (
		_w2048_,
		_w2055_,
		_w2057_
	);
	LUT2 #(
		.INIT('h1)
	) name1099 (
		_w2056_,
		_w2057_,
		_w2058_
	);
	LUT2 #(
		.INIT('h8)
	) name1100 (
		\u3_u0_r1_reg[35]/P0001 ,
		_w1902_,
		_w2059_
	);
	LUT2 #(
		.INIT('h8)
	) name1101 (
		\u3_u0_r3_reg[35]/P0001 ,
		_w1906_,
		_w2060_
	);
	LUT2 #(
		.INIT('h8)
	) name1102 (
		\u3_u0_r0_reg[35]/P0001 ,
		_w1899_,
		_w2061_
	);
	LUT2 #(
		.INIT('h8)
	) name1103 (
		\u3_u0_r2_reg[35]/P0001 ,
		_w1909_,
		_w2062_
	);
	LUT2 #(
		.INIT('h1)
	) name1104 (
		_w2059_,
		_w2060_,
		_w2063_
	);
	LUT2 #(
		.INIT('h1)
	) name1105 (
		_w2061_,
		_w2062_,
		_w2064_
	);
	LUT2 #(
		.INIT('h8)
	) name1106 (
		_w2063_,
		_w2064_,
		_w2065_
	);
	LUT2 #(
		.INIT('h8)
	) name1107 (
		\u3_u0_r0_reg[26]/P0001 ,
		_w1899_,
		_w2066_
	);
	LUT2 #(
		.INIT('h8)
	) name1108 (
		\u3_u0_r1_reg[26]/P0001 ,
		_w1902_,
		_w2067_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		\u3_u0_r3_reg[26]/P0001 ,
		_w1906_,
		_w2068_
	);
	LUT2 #(
		.INIT('h8)
	) name1110 (
		\u3_u0_r2_reg[26]/P0001 ,
		_w1909_,
		_w2069_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w2066_,
		_w2067_,
		_w2070_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w2068_,
		_w2069_,
		_w2071_
	);
	LUT2 #(
		.INIT('h8)
	) name1113 (
		_w2070_,
		_w2071_,
		_w2072_
	);
	LUT2 #(
		.INIT('h2)
	) name1114 (
		_w2065_,
		_w2072_,
		_w2073_
	);
	LUT2 #(
		.INIT('h4)
	) name1115 (
		_w2065_,
		_w2072_,
		_w2074_
	);
	LUT2 #(
		.INIT('h1)
	) name1116 (
		_w2073_,
		_w2074_,
		_w2075_
	);
	LUT2 #(
		.INIT('h8)
	) name1117 (
		_w2058_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		_w2058_,
		_w2075_,
		_w2077_
	);
	LUT2 #(
		.INIT('h1)
	) name1119 (
		_w2076_,
		_w2077_,
		_w2078_
	);
	LUT2 #(
		.INIT('h4)
	) name1120 (
		_w2041_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h2)
	) name1121 (
		_w2041_,
		_w2078_,
		_w2080_
	);
	LUT2 #(
		.INIT('h2)
	) name1122 (
		\wb_sel_i[3]_pad ,
		_w2079_,
		_w2081_
	);
	LUT2 #(
		.INIT('h4)
	) name1123 (
		_w2080_,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h8)
	) name1124 (
		\u3_u0_r1_reg[21]/P0001 ,
		_w1902_,
		_w2083_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		\u3_u0_r0_reg[21]/P0001 ,
		_w1899_,
		_w2084_
	);
	LUT2 #(
		.INIT('h8)
	) name1126 (
		\u3_u0_r2_reg[21]/P0001 ,
		_w1909_,
		_w2085_
	);
	LUT2 #(
		.INIT('h8)
	) name1127 (
		\u3_u0_r3_reg[21]/P0001 ,
		_w1906_,
		_w2086_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w2083_,
		_w2084_,
		_w2087_
	);
	LUT2 #(
		.INIT('h1)
	) name1129 (
		_w2085_,
		_w2086_,
		_w2088_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		_w2087_,
		_w2088_,
		_w2089_
	);
	LUT2 #(
		.INIT('h8)
	) name1131 (
		\u3_u0_r0_reg[17]/P0001 ,
		_w1899_,
		_w2090_
	);
	LUT2 #(
		.INIT('h8)
	) name1132 (
		\u3_u0_r1_reg[17]/P0001 ,
		_w1902_,
		_w2091_
	);
	LUT2 #(
		.INIT('h8)
	) name1133 (
		\u3_u0_r3_reg[17]/P0001 ,
		_w1906_,
		_w2092_
	);
	LUT2 #(
		.INIT('h8)
	) name1134 (
		\u3_u0_r2_reg[17]/P0001 ,
		_w1909_,
		_w2093_
	);
	LUT2 #(
		.INIT('h1)
	) name1135 (
		_w2090_,
		_w2091_,
		_w2094_
	);
	LUT2 #(
		.INIT('h1)
	) name1136 (
		_w2092_,
		_w2093_,
		_w2095_
	);
	LUT2 #(
		.INIT('h8)
	) name1137 (
		_w2094_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('h2)
	) name1138 (
		_w2089_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h4)
	) name1139 (
		_w2089_,
		_w2096_,
		_w2098_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w2097_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h8)
	) name1141 (
		\u3_u0_r0_reg[22]/P0001 ,
		_w1899_,
		_w2100_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		\u3_u0_r1_reg[22]/P0001 ,
		_w1902_,
		_w2101_
	);
	LUT2 #(
		.INIT('h8)
	) name1143 (
		\u3_u0_r3_reg[22]/P0001 ,
		_w1906_,
		_w2102_
	);
	LUT2 #(
		.INIT('h8)
	) name1144 (
		\u3_u0_r2_reg[22]/P0001 ,
		_w1909_,
		_w2103_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		_w2100_,
		_w2101_,
		_w2104_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w2102_,
		_w2103_,
		_w2105_
	);
	LUT2 #(
		.INIT('h8)
	) name1147 (
		_w2104_,
		_w2105_,
		_w2106_
	);
	LUT2 #(
		.INIT('h8)
	) name1148 (
		\u3_u0_r0_reg[19]/P0001 ,
		_w1899_,
		_w2107_
	);
	LUT2 #(
		.INIT('h8)
	) name1149 (
		\u3_u0_r2_reg[19]/P0001 ,
		_w1909_,
		_w2108_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\u3_u0_r1_reg[19]/P0001 ,
		_w1902_,
		_w2109_
	);
	LUT2 #(
		.INIT('h8)
	) name1151 (
		\u3_u0_r3_reg[19]/P0001 ,
		_w1906_,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name1152 (
		_w2107_,
		_w2108_,
		_w2111_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		_w2109_,
		_w2110_,
		_w2112_
	);
	LUT2 #(
		.INIT('h8)
	) name1154 (
		_w2111_,
		_w2112_,
		_w2113_
	);
	LUT2 #(
		.INIT('h8)
	) name1155 (
		\u3_u0_r0_reg[20]/P0001 ,
		_w1899_,
		_w2114_
	);
	LUT2 #(
		.INIT('h8)
	) name1156 (
		\u3_u0_r3_reg[20]/P0001 ,
		_w1906_,
		_w2115_
	);
	LUT2 #(
		.INIT('h8)
	) name1157 (
		\u3_u0_r1_reg[20]/P0001 ,
		_w1902_,
		_w2116_
	);
	LUT2 #(
		.INIT('h8)
	) name1158 (
		\u3_u0_r2_reg[20]/P0001 ,
		_w1909_,
		_w2117_
	);
	LUT2 #(
		.INIT('h1)
	) name1159 (
		_w2114_,
		_w2115_,
		_w2118_
	);
	LUT2 #(
		.INIT('h1)
	) name1160 (
		_w2116_,
		_w2117_,
		_w2119_
	);
	LUT2 #(
		.INIT('h8)
	) name1161 (
		_w2118_,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		_w2113_,
		_w2120_,
		_w2121_
	);
	LUT2 #(
		.INIT('h8)
	) name1163 (
		_w2113_,
		_w2120_,
		_w2122_
	);
	LUT2 #(
		.INIT('h1)
	) name1164 (
		_w2121_,
		_w2122_,
		_w2123_
	);
	LUT2 #(
		.INIT('h2)
	) name1165 (
		_w2106_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		_w2106_,
		_w2123_,
		_w2125_
	);
	LUT2 #(
		.INIT('h1)
	) name1167 (
		_w2124_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h8)
	) name1168 (
		_w2099_,
		_w2126_,
		_w2127_
	);
	LUT2 #(
		.INIT('h1)
	) name1169 (
		_w2099_,
		_w2126_,
		_w2128_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		_w2127_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		\u3_u0_r0_reg[16]/P0001 ,
		_w1899_,
		_w2130_
	);
	LUT2 #(
		.INIT('h8)
	) name1172 (
		\u3_u0_r1_reg[16]/P0001 ,
		_w1902_,
		_w2131_
	);
	LUT2 #(
		.INIT('h8)
	) name1173 (
		\u3_u0_r3_reg[16]/P0001 ,
		_w1906_,
		_w2132_
	);
	LUT2 #(
		.INIT('h8)
	) name1174 (
		\u3_u0_r2_reg[16]/P0001 ,
		_w1909_,
		_w2133_
	);
	LUT2 #(
		.INIT('h1)
	) name1175 (
		_w2130_,
		_w2131_,
		_w2134_
	);
	LUT2 #(
		.INIT('h1)
	) name1176 (
		_w2132_,
		_w2133_,
		_w2135_
	);
	LUT2 #(
		.INIT('h8)
	) name1177 (
		_w2134_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		\u3_u0_r0_reg[23]/P0001 ,
		_w1899_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name1179 (
		\u3_u0_r1_reg[23]/P0001 ,
		_w1902_,
		_w2138_
	);
	LUT2 #(
		.INIT('h8)
	) name1180 (
		\u3_u0_r3_reg[23]/P0001 ,
		_w1906_,
		_w2139_
	);
	LUT2 #(
		.INIT('h8)
	) name1181 (
		\u3_u0_r2_reg[23]/P0001 ,
		_w1909_,
		_w2140_
	);
	LUT2 #(
		.INIT('h1)
	) name1182 (
		_w2137_,
		_w2138_,
		_w2141_
	);
	LUT2 #(
		.INIT('h1)
	) name1183 (
		_w2139_,
		_w2140_,
		_w2142_
	);
	LUT2 #(
		.INIT('h8)
	) name1184 (
		_w2141_,
		_w2142_,
		_w2143_
	);
	LUT2 #(
		.INIT('h2)
	) name1185 (
		_w2136_,
		_w2143_,
		_w2144_
	);
	LUT2 #(
		.INIT('h4)
	) name1186 (
		_w2136_,
		_w2143_,
		_w2145_
	);
	LUT2 #(
		.INIT('h1)
	) name1187 (
		_w2144_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h8)
	) name1188 (
		\u3_u0_r0_reg[34]/P0001 ,
		_w1899_,
		_w2147_
	);
	LUT2 #(
		.INIT('h8)
	) name1189 (
		\u3_u0_r1_reg[34]/P0001 ,
		_w1902_,
		_w2148_
	);
	LUT2 #(
		.INIT('h8)
	) name1190 (
		\u3_u0_r3_reg[34]/P0001 ,
		_w1906_,
		_w2149_
	);
	LUT2 #(
		.INIT('h8)
	) name1191 (
		\u3_u0_r2_reg[34]/P0001 ,
		_w1909_,
		_w2150_
	);
	LUT2 #(
		.INIT('h1)
	) name1192 (
		_w2147_,
		_w2148_,
		_w2151_
	);
	LUT2 #(
		.INIT('h1)
	) name1193 (
		_w2149_,
		_w2150_,
		_w2152_
	);
	LUT2 #(
		.INIT('h8)
	) name1194 (
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h8)
	) name1195 (
		\u3_u0_r0_reg[18]/P0001 ,
		_w1899_,
		_w2154_
	);
	LUT2 #(
		.INIT('h8)
	) name1196 (
		\u3_u0_r1_reg[18]/P0001 ,
		_w1902_,
		_w2155_
	);
	LUT2 #(
		.INIT('h8)
	) name1197 (
		\u3_u0_r3_reg[18]/P0001 ,
		_w1906_,
		_w2156_
	);
	LUT2 #(
		.INIT('h8)
	) name1198 (
		\u3_u0_r2_reg[18]/P0001 ,
		_w1909_,
		_w2157_
	);
	LUT2 #(
		.INIT('h1)
	) name1199 (
		_w2154_,
		_w2155_,
		_w2158_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w2156_,
		_w2157_,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1201 (
		_w2158_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h2)
	) name1202 (
		_w2153_,
		_w2160_,
		_w2161_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w2153_,
		_w2160_,
		_w2162_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		_w2161_,
		_w2162_,
		_w2163_
	);
	LUT2 #(
		.INIT('h8)
	) name1205 (
		_w2146_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w2146_,
		_w2163_,
		_w2165_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		_w2164_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		_w2129_,
		_w2166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h2)
	) name1209 (
		_w2129_,
		_w2166_,
		_w2168_
	);
	LUT2 #(
		.INIT('h2)
	) name1210 (
		\wb_sel_i[2]_pad ,
		_w2167_,
		_w2169_
	);
	LUT2 #(
		.INIT('h4)
	) name1211 (
		_w2168_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name1212 (
		\u3_u0_r0_reg[0]/P0001 ,
		_w1899_,
		_w2171_
	);
	LUT2 #(
		.INIT('h8)
	) name1213 (
		\u3_u0_r2_reg[0]/P0001 ,
		_w1909_,
		_w2172_
	);
	LUT2 #(
		.INIT('h8)
	) name1214 (
		\u3_u0_r1_reg[0]/P0001 ,
		_w1902_,
		_w2173_
	);
	LUT2 #(
		.INIT('h8)
	) name1215 (
		\u3_u0_r3_reg[0]/P0001 ,
		_w1906_,
		_w2174_
	);
	LUT2 #(
		.INIT('h1)
	) name1216 (
		_w2171_,
		_w2172_,
		_w2175_
	);
	LUT2 #(
		.INIT('h1)
	) name1217 (
		_w2173_,
		_w2174_,
		_w2176_
	);
	LUT2 #(
		.INIT('h8)
	) name1218 (
		_w2175_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		\u3_u0_r0_reg[2]/P0001 ,
		_w1899_,
		_w2178_
	);
	LUT2 #(
		.INIT('h8)
	) name1220 (
		\u3_u0_r1_reg[2]/P0001 ,
		_w1902_,
		_w2179_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		\u3_u0_r3_reg[2]/P0001 ,
		_w1906_,
		_w2180_
	);
	LUT2 #(
		.INIT('h8)
	) name1222 (
		\u3_u0_r2_reg[2]/P0001 ,
		_w1909_,
		_w2181_
	);
	LUT2 #(
		.INIT('h1)
	) name1223 (
		_w2178_,
		_w2179_,
		_w2182_
	);
	LUT2 #(
		.INIT('h1)
	) name1224 (
		_w2180_,
		_w2181_,
		_w2183_
	);
	LUT2 #(
		.INIT('h8)
	) name1225 (
		_w2182_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('h2)
	) name1226 (
		_w2177_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h4)
	) name1227 (
		_w2177_,
		_w2184_,
		_w2186_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		_w2185_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h8)
	) name1229 (
		\u3_u0_r0_reg[4]/P0001 ,
		_w1899_,
		_w2188_
	);
	LUT2 #(
		.INIT('h8)
	) name1230 (
		\u3_u0_r1_reg[4]/P0001 ,
		_w1902_,
		_w2189_
	);
	LUT2 #(
		.INIT('h8)
	) name1231 (
		\u3_u0_r3_reg[4]/P0001 ,
		_w1906_,
		_w2190_
	);
	LUT2 #(
		.INIT('h8)
	) name1232 (
		\u3_u0_r2_reg[4]/P0001 ,
		_w1909_,
		_w2191_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		_w2188_,
		_w2189_,
		_w2192_
	);
	LUT2 #(
		.INIT('h1)
	) name1234 (
		_w2190_,
		_w2191_,
		_w2193_
	);
	LUT2 #(
		.INIT('h8)
	) name1235 (
		_w2192_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h8)
	) name1236 (
		\u3_u0_r3_reg[7]/P0001 ,
		_w1906_,
		_w2195_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		\u3_u0_r2_reg[7]/P0001 ,
		_w1909_,
		_w2196_
	);
	LUT2 #(
		.INIT('h8)
	) name1238 (
		\u3_u0_r0_reg[7]/P0001 ,
		_w1899_,
		_w2197_
	);
	LUT2 #(
		.INIT('h8)
	) name1239 (
		\u3_u0_r1_reg[7]/P0001 ,
		_w1902_,
		_w2198_
	);
	LUT2 #(
		.INIT('h1)
	) name1240 (
		_w2195_,
		_w2196_,
		_w2199_
	);
	LUT2 #(
		.INIT('h1)
	) name1241 (
		_w2197_,
		_w2198_,
		_w2200_
	);
	LUT2 #(
		.INIT('h8)
	) name1242 (
		_w2199_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		\u3_u0_r1_reg[6]/P0001 ,
		_w1902_,
		_w2202_
	);
	LUT2 #(
		.INIT('h8)
	) name1244 (
		\u3_u0_r2_reg[6]/P0001 ,
		_w1909_,
		_w2203_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		\u3_u0_r0_reg[6]/P0001 ,
		_w1899_,
		_w2204_
	);
	LUT2 #(
		.INIT('h8)
	) name1246 (
		\u3_u0_r3_reg[6]/P0001 ,
		_w1906_,
		_w2205_
	);
	LUT2 #(
		.INIT('h1)
	) name1247 (
		_w2202_,
		_w2203_,
		_w2206_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w2204_,
		_w2205_,
		_w2207_
	);
	LUT2 #(
		.INIT('h8)
	) name1249 (
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h1)
	) name1250 (
		_w2201_,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h8)
	) name1251 (
		_w2201_,
		_w2208_,
		_w2210_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		_w2209_,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h2)
	) name1253 (
		_w2194_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h4)
	) name1254 (
		_w2194_,
		_w2211_,
		_w2213_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		_w2212_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h8)
	) name1256 (
		_w2187_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w2187_,
		_w2214_,
		_w2216_
	);
	LUT2 #(
		.INIT('h1)
	) name1258 (
		_w2215_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		\u3_u0_r3_reg[5]/P0001 ,
		_w1906_,
		_w2218_
	);
	LUT2 #(
		.INIT('h8)
	) name1260 (
		\u3_u0_r2_reg[5]/P0001 ,
		_w1909_,
		_w2219_
	);
	LUT2 #(
		.INIT('h8)
	) name1261 (
		\u3_u0_r0_reg[5]/P0001 ,
		_w1899_,
		_w2220_
	);
	LUT2 #(
		.INIT('h8)
	) name1262 (
		\u3_u0_r1_reg[5]/P0001 ,
		_w1902_,
		_w2221_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w2218_,
		_w2219_,
		_w2222_
	);
	LUT2 #(
		.INIT('h1)
	) name1264 (
		_w2220_,
		_w2221_,
		_w2223_
	);
	LUT2 #(
		.INIT('h8)
	) name1265 (
		_w2222_,
		_w2223_,
		_w2224_
	);
	LUT2 #(
		.INIT('h8)
	) name1266 (
		\u3_u0_r0_reg[3]/P0001 ,
		_w1899_,
		_w2225_
	);
	LUT2 #(
		.INIT('h8)
	) name1267 (
		\u3_u0_r2_reg[3]/P0001 ,
		_w1909_,
		_w2226_
	);
	LUT2 #(
		.INIT('h8)
	) name1268 (
		\u3_u0_r1_reg[3]/P0001 ,
		_w1902_,
		_w2227_
	);
	LUT2 #(
		.INIT('h8)
	) name1269 (
		\u3_u0_r3_reg[3]/P0001 ,
		_w1906_,
		_w2228_
	);
	LUT2 #(
		.INIT('h1)
	) name1270 (
		_w2225_,
		_w2226_,
		_w2229_
	);
	LUT2 #(
		.INIT('h1)
	) name1271 (
		_w2227_,
		_w2228_,
		_w2230_
	);
	LUT2 #(
		.INIT('h8)
	) name1272 (
		_w2229_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h2)
	) name1273 (
		_w2224_,
		_w2231_,
		_w2232_
	);
	LUT2 #(
		.INIT('h4)
	) name1274 (
		_w2224_,
		_w2231_,
		_w2233_
	);
	LUT2 #(
		.INIT('h1)
	) name1275 (
		_w2232_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name1276 (
		\u3_u0_r3_reg[32]/P0001 ,
		_w1906_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name1277 (
		\u3_u0_r2_reg[32]/P0001 ,
		_w1909_,
		_w2236_
	);
	LUT2 #(
		.INIT('h8)
	) name1278 (
		\u3_u0_r0_reg[32]/P0001 ,
		_w1899_,
		_w2237_
	);
	LUT2 #(
		.INIT('h8)
	) name1279 (
		\u3_u0_r1_reg[32]/P0001 ,
		_w1902_,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name1280 (
		_w2235_,
		_w2236_,
		_w2239_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w2237_,
		_w2238_,
		_w2240_
	);
	LUT2 #(
		.INIT('h8)
	) name1282 (
		_w2239_,
		_w2240_,
		_w2241_
	);
	LUT2 #(
		.INIT('h8)
	) name1283 (
		\u3_u0_r0_reg[1]/P0001 ,
		_w1899_,
		_w2242_
	);
	LUT2 #(
		.INIT('h8)
	) name1284 (
		\u3_u0_r1_reg[1]/P0001 ,
		_w1902_,
		_w2243_
	);
	LUT2 #(
		.INIT('h8)
	) name1285 (
		\u3_u0_r3_reg[1]/P0001 ,
		_w1906_,
		_w2244_
	);
	LUT2 #(
		.INIT('h8)
	) name1286 (
		\u3_u0_r2_reg[1]/P0001 ,
		_w1909_,
		_w2245_
	);
	LUT2 #(
		.INIT('h1)
	) name1287 (
		_w2242_,
		_w2243_,
		_w2246_
	);
	LUT2 #(
		.INIT('h1)
	) name1288 (
		_w2244_,
		_w2245_,
		_w2247_
	);
	LUT2 #(
		.INIT('h8)
	) name1289 (
		_w2246_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h2)
	) name1290 (
		_w2241_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h4)
	) name1291 (
		_w2241_,
		_w2248_,
		_w2250_
	);
	LUT2 #(
		.INIT('h1)
	) name1292 (
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		_w2234_,
		_w2251_,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		_w2234_,
		_w2251_,
		_w2253_
	);
	LUT2 #(
		.INIT('h1)
	) name1295 (
		_w2252_,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h4)
	) name1296 (
		_w2217_,
		_w2254_,
		_w2255_
	);
	LUT2 #(
		.INIT('h2)
	) name1297 (
		_w2217_,
		_w2254_,
		_w2256_
	);
	LUT2 #(
		.INIT('h2)
	) name1298 (
		\wb_sel_i[0]_pad ,
		_w2255_,
		_w2257_
	);
	LUT2 #(
		.INIT('h4)
	) name1299 (
		_w2256_,
		_w2257_,
		_w2258_
	);
	LUT2 #(
		.INIT('h1)
	) name1300 (
		_w1994_,
		_w2082_,
		_w2259_
	);
	LUT2 #(
		.INIT('h1)
	) name1301 (
		_w2170_,
		_w2258_,
		_w2260_
	);
	LUT2 #(
		.INIT('h8)
	) name1302 (
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h2)
	) name1303 (
		\u0_csc_reg[11]/NET0131 ,
		wb_we_i_pad,
		_w2262_
	);
	LUT2 #(
		.INIT('h4)
	) name1304 (
		_w2261_,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		_w1896_,
		_w2263_,
		_w2264_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		\u0_wp_err_reg/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w2265_
	);
	LUT2 #(
		.INIT('h4)
	) name1307 (
		_w2264_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h2)
	) name1308 (
		_w1046_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h1)
	) name1309 (
		\wb_addr_i[29]_pad ,
		\wb_addr_i[30]_pad ,
		_w2268_
	);
	LUT2 #(
		.INIT('h4)
	) name1310 (
		\wb_addr_i[31]_pad ,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h8)
	) name1311 (
		_w1896_,
		_w2269_,
		_w2270_
	);
	LUT2 #(
		.INIT('h4)
	) name1312 (
		_w2267_,
		_w2270_,
		_w2271_
	);
	LUT2 #(
		.INIT('h8)
	) name1313 (
		\wb_addr_i[29]_pad ,
		\wb_addr_i[30]_pad ,
		_w2272_
	);
	LUT2 #(
		.INIT('h4)
	) name1314 (
		\wb_addr_i[31]_pad ,
		_w2272_,
		_w2273_
	);
	LUT2 #(
		.INIT('h4)
	) name1315 (
		wb_ack_o_pad,
		_w1046_,
		_w2274_
	);
	LUT2 #(
		.INIT('h8)
	) name1316 (
		_w2273_,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h1)
	) name1317 (
		_w2271_,
		_w2275_,
		_w2276_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		_w1693_,
		_w1803_,
		_w2277_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		_w1777_,
		_w2277_,
		_w2278_
	);
	LUT2 #(
		.INIT('h8)
	) name1320 (
		\u0_tms_reg[23]/NET0131 ,
		_w1051_,
		_w2279_
	);
	LUT2 #(
		.INIT('h2)
	) name1321 (
		\u0_sp_tms_reg[23]/NET0131 ,
		_w1051_,
		_w2280_
	);
	LUT2 #(
		.INIT('h1)
	) name1322 (
		_w2279_,
		_w2280_,
		_w2281_
	);
	LUT2 #(
		.INIT('h8)
	) name1323 (
		_w1693_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h1)
	) name1324 (
		_w1719_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h2)
	) name1325 (
		\u5_timer_reg[3]/NET0131 ,
		_w1831_,
		_w2284_
	);
	LUT2 #(
		.INIT('h8)
	) name1326 (
		_w1821_,
		_w1830_,
		_w2285_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w2284_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h4)
	) name1328 (
		\u5_state_reg[35]/NET0131 ,
		_w1010_,
		_w2287_
	);
	LUT2 #(
		.INIT('h8)
	) name1329 (
		_w1820_,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('h4)
	) name1330 (
		_w2286_,
		_w2288_,
		_w2289_
	);
	LUT2 #(
		.INIT('h2)
	) name1331 (
		\u0_sp_tms_reg[27]/NET0131 ,
		_w1051_,
		_w2290_
	);
	LUT2 #(
		.INIT('h8)
	) name1332 (
		\u0_tms_reg[27]/NET0131 ,
		_w1051_,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name1333 (
		_w2290_,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h8)
	) name1334 (
		_w1693_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h1)
	) name1335 (
		_w1820_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('h1)
	) name1336 (
		_w2289_,
		_w2294_,
		_w2295_
	);
	LUT2 #(
		.INIT('h8)
	) name1337 (
		_w1790_,
		_w1837_,
		_w2296_
	);
	LUT2 #(
		.INIT('h4)
	) name1338 (
		_w2295_,
		_w2296_,
		_w2297_
	);
	LUT2 #(
		.INIT('h2)
	) name1339 (
		_w1812_,
		_w2282_,
		_w2298_
	);
	LUT2 #(
		.INIT('h4)
	) name1340 (
		_w1812_,
		_w2282_,
		_w2299_
	);
	LUT2 #(
		.INIT('h1)
	) name1341 (
		_w1790_,
		_w2298_,
		_w2300_
	);
	LUT2 #(
		.INIT('h4)
	) name1342 (
		_w2299_,
		_w2300_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name1343 (
		_w2283_,
		_w2297_,
		_w2302_
	);
	LUT2 #(
		.INIT('h4)
	) name1344 (
		_w2301_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h2)
	) name1345 (
		_w1817_,
		_w2303_,
		_w2304_
	);
	LUT2 #(
		.INIT('h8)
	) name1346 (
		\u0_tms_reg[3]/NET0131 ,
		_w1051_,
		_w2305_
	);
	LUT2 #(
		.INIT('h2)
	) name1347 (
		\u0_sp_tms_reg[3]/NET0131 ,
		_w1051_,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name1348 (
		_w2305_,
		_w2306_,
		_w2307_
	);
	LUT2 #(
		.INIT('h8)
	) name1349 (
		_w1693_,
		_w2307_,
		_w2308_
	);
	LUT2 #(
		.INIT('h1)
	) name1350 (
		_w1817_,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('h2)
	) name1351 (
		_w1785_,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h4)
	) name1352 (
		_w2304_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name1353 (
		\u0_tms_reg[11]/NET0131 ,
		_w1051_,
		_w2312_
	);
	LUT2 #(
		.INIT('h2)
	) name1354 (
		\u0_sp_tms_reg[11]/NET0131 ,
		_w1051_,
		_w2313_
	);
	LUT2 #(
		.INIT('h1)
	) name1355 (
		_w2312_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h8)
	) name1356 (
		_w1693_,
		_w2314_,
		_w2315_
	);
	LUT2 #(
		.INIT('h4)
	) name1357 (
		_w1785_,
		_w2315_,
		_w2316_
	);
	LUT2 #(
		.INIT('h2)
	) name1358 (
		_w1777_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('h4)
	) name1359 (
		_w2311_,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('h1)
	) name1360 (
		_w2278_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1221_,
		_w2320_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		\u5_state_reg[16]/NET0131 ,
		_w1631_,
		_w2321_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1184_,
		_w2322_
	);
	LUT2 #(
		.INIT('h1)
	) name1364 (
		\u5_ap_en_reg/NET0131 ,
		_w1654_,
		_w2323_
	);
	LUT2 #(
		.INIT('h4)
	) name1365 (
		\u5_wb_write_go_r_reg/NET0131 ,
		_w1627_,
		_w2324_
	);
	LUT2 #(
		.INIT('h2)
	) name1366 (
		\u5_state_reg[16]/NET0131 ,
		_w2324_,
		_w2325_
	);
	LUT2 #(
		.INIT('h8)
	) name1367 (
		_w1654_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h1)
	) name1368 (
		_w2323_,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h1)
	) name1369 (
		_w2322_,
		_w2327_,
		_w2328_
	);
	LUT2 #(
		.INIT('h8)
	) name1370 (
		_w1750_,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h1)
	) name1371 (
		_w2321_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h2)
	) name1372 (
		_w1189_,
		_w2330_,
		_w2331_
	);
	LUT2 #(
		.INIT('h1)
	) name1373 (
		_w1382_,
		_w1655_,
		_w2332_
	);
	LUT2 #(
		.INIT('h2)
	) name1374 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1654_,
		_w2333_
	);
	LUT2 #(
		.INIT('h4)
	) name1375 (
		\u5_ap_en_reg/NET0131 ,
		_w1888_,
		_w2334_
	);
	LUT2 #(
		.INIT('h4)
	) name1376 (
		_w2333_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h8)
	) name1377 (
		_w2332_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h2)
	) name1378 (
		\u5_state_reg[16]/NET0131 ,
		_w1875_,
		_w2337_
	);
	LUT2 #(
		.INIT('h4)
	) name1379 (
		\u5_ap_en_reg/NET0131 ,
		_w1375_,
		_w2338_
	);
	LUT2 #(
		.INIT('h1)
	) name1380 (
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT2 #(
		.INIT('h1)
	) name1381 (
		_w1382_,
		_w1873_,
		_w2340_
	);
	LUT2 #(
		.INIT('h2)
	) name1382 (
		_w1224_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('h4)
	) name1383 (
		_w2339_,
		_w2341_,
		_w2342_
	);
	LUT2 #(
		.INIT('h2)
	) name1384 (
		\u5_tmr_done_reg/NET0131 ,
		_w1375_,
		_w2343_
	);
	LUT2 #(
		.INIT('h2)
	) name1385 (
		_w1302_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1424_,
		_w2345_
	);
	LUT2 #(
		.INIT('h2)
	) name1387 (
		\u5_state_reg[16]/NET0131 ,
		_w2345_,
		_w2346_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		_w2344_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h1)
	) name1389 (
		_w2320_,
		_w2347_,
		_w2348_
	);
	LUT2 #(
		.INIT('h4)
	) name1390 (
		_w2342_,
		_w2348_,
		_w2349_
	);
	LUT2 #(
		.INIT('h4)
	) name1391 (
		_w2336_,
		_w2349_,
		_w2350_
	);
	LUT2 #(
		.INIT('h4)
	) name1392 (
		_w2331_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h2)
	) name1393 (
		\u0_sp_csc_reg[7]/NET0131 ,
		_w1051_,
		_w2352_
	);
	LUT2 #(
		.INIT('h8)
	) name1394 (
		\u0_csc_reg[7]/NET0131 ,
		_w1051_,
		_w2353_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		_w2352_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('h2)
	) name1396 (
		\u0_sp_csc_reg[6]/NET0131 ,
		_w1051_,
		_w2355_
	);
	LUT2 #(
		.INIT('h8)
	) name1397 (
		\u0_csc_reg[6]/NET0131 ,
		_w1051_,
		_w2356_
	);
	LUT2 #(
		.INIT('h1)
	) name1398 (
		_w2355_,
		_w2356_,
		_w2357_
	);
	LUT2 #(
		.INIT('h8)
	) name1399 (
		_w2354_,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('h2)
	) name1400 (
		\u0_sp_csc_reg[4]/NET0131 ,
		_w1051_,
		_w2359_
	);
	LUT2 #(
		.INIT('h8)
	) name1401 (
		\u0_csc_reg[4]/NET0131 ,
		_w1051_,
		_w2360_
	);
	LUT2 #(
		.INIT('h1)
	) name1402 (
		_w2359_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h2)
	) name1403 (
		_w2358_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h2)
	) name1404 (
		\u0_sp_csc_reg[5]/NET0131 ,
		_w1051_,
		_w2363_
	);
	LUT2 #(
		.INIT('h8)
	) name1405 (
		\u0_csc_reg[5]/NET0131 ,
		_w1051_,
		_w2364_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		_w2363_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h4)
	) name1407 (
		_w2362_,
		_w2365_,
		_w2366_
	);
	LUT2 #(
		.INIT('h2)
	) name1408 (
		\u5_state_reg[1]/NET0131 ,
		_w1853_,
		_w2367_
	);
	LUT2 #(
		.INIT('h4)
	) name1409 (
		_w2366_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h4)
	) name1410 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1044_,
		_w2369_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1887_,
		_w2370_
	);
	LUT2 #(
		.INIT('h8)
	) name1412 (
		_w1869_,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('h4)
	) name1413 (
		_w1880_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h4)
	) name1414 (
		_w1891_,
		_w2372_,
		_w2373_
	);
	LUT2 #(
		.INIT('h1)
	) name1415 (
		_w2369_,
		_w2373_,
		_w2374_
	);
	LUT2 #(
		.INIT('h8)
	) name1416 (
		_w1649_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h4)
	) name1417 (
		\u5_burst_cnt_reg[7]/NET0131 ,
		_w2375_,
		_w2376_
	);
	LUT2 #(
		.INIT('h2)
	) name1418 (
		\u5_burst_cnt_reg[8]/NET0131 ,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name1419 (
		_w1651_,
		_w2374_,
		_w2378_
	);
	LUT2 #(
		.INIT('h1)
	) name1420 (
		_w2377_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h1)
	) name1421 (
		\u5_state_reg[1]/NET0131 ,
		_w2379_,
		_w2380_
	);
	LUT2 #(
		.INIT('h1)
	) name1422 (
		_w2368_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('h1)
	) name1423 (
		\u5_state_reg[52]/NET0131 ,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h4)
	) name1424 (
		\u5_burst_cnt_reg[9]/NET0131 ,
		_w2378_,
		_w2383_
	);
	LUT2 #(
		.INIT('h2)
	) name1425 (
		\u5_burst_cnt_reg[10]/NET0131 ,
		_w2383_,
		_w2384_
	);
	LUT2 #(
		.INIT('h8)
	) name1426 (
		_w1653_,
		_w2374_,
		_w2385_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h1)
	) name1428 (
		\u5_state_reg[1]/NET0131 ,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('h8)
	) name1429 (
		_w2361_,
		_w2365_,
		_w2388_
	);
	LUT2 #(
		.INIT('h4)
	) name1430 (
		_w2358_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		_w2367_,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h1)
	) name1432 (
		_w2387_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name1433 (
		\u5_state_reg[52]/NET0131 ,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h4)
	) name1434 (
		\u5_burst_cnt_reg[0]/NET0131 ,
		_w2374_,
		_w2393_
	);
	LUT2 #(
		.INIT('h2)
	) name1435 (
		\u5_burst_cnt_reg[0]/NET0131 ,
		_w2374_,
		_w2394_
	);
	LUT2 #(
		.INIT('h1)
	) name1436 (
		_w2393_,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		\u5_state_reg[1]/NET0131 ,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h8)
	) name1438 (
		_w1179_,
		_w1693_,
		_w2397_
	);
	LUT2 #(
		.INIT('h8)
	) name1439 (
		\u5_state_reg[1]/NET0131 ,
		_w2397_,
		_w2398_
	);
	LUT2 #(
		.INIT('h8)
	) name1440 (
		_w1176_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h1)
	) name1441 (
		_w2396_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		\u5_state_reg[52]/NET0131 ,
		_w2400_,
		_w2401_
	);
	LUT2 #(
		.INIT('h1)
	) name1443 (
		\u5_state_reg[17]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2402_
	);
	LUT2 #(
		.INIT('h4)
	) name1444 (
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2403_
	);
	LUT2 #(
		.INIT('h2)
	) name1445 (
		_w1279_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h1)
	) name1446 (
		_w1195_,
		_w2404_,
		_w2405_
	);
	LUT2 #(
		.INIT('h1)
	) name1447 (
		_w2402_,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('h4)
	) name1448 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1362_,
		_w2407_
	);
	LUT2 #(
		.INIT('h1)
	) name1449 (
		_w2406_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h4)
	) name1450 (
		wb_err_o_pad,
		_w2269_,
		_w2409_
	);
	LUT2 #(
		.INIT('h8)
	) name1451 (
		_w2267_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h4)
	) name1452 (
		\u5_cs_le_r_reg/P0001 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w2411_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		\u5_state_reg[1]/NET0131 ,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('h8)
	) name1454 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1629_,
		_w2413_
	);
	LUT2 #(
		.INIT('h2)
	) name1455 (
		\u5_tmr2_done_reg/NET0131 ,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h8)
	) name1456 (
		_w1106_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h4)
	) name1457 (
		_w2412_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h1)
	) name1458 (
		\u5_state_reg[1]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2417_
	);
	LUT2 #(
		.INIT('h1)
	) name1459 (
		_w1269_,
		_w1309_,
		_w2418_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w2417_,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h4)
	) name1461 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2420_
	);
	LUT2 #(
		.INIT('h4)
	) name1462 (
		_w1679_,
		_w2420_,
		_w2421_
	);
	LUT2 #(
		.INIT('h2)
	) name1463 (
		\u5_lookup_ready2_reg/NET0131 ,
		_w1629_,
		_w2422_
	);
	LUT2 #(
		.INIT('h2)
	) name1464 (
		_w1062_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h1)
	) name1465 (
		_w1438_,
		_w1440_,
		_w2424_
	);
	LUT2 #(
		.INIT('h2)
	) name1466 (
		_w1629_,
		_w2424_,
		_w2425_
	);
	LUT2 #(
		.INIT('h1)
	) name1467 (
		_w2423_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h8)
	) name1468 (
		_w1679_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h2)
	) name1469 (
		_w1685_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h4)
	) name1470 (
		_w2421_,
		_w2428_,
		_w2429_
	);
	LUT2 #(
		.INIT('h8)
	) name1471 (
		_w1302_,
		_w2343_,
		_w2430_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		_w1108_,
		_w2419_,
		_w2431_
	);
	LUT2 #(
		.INIT('h4)
	) name1473 (
		_w2416_,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h4)
	) name1474 (
		_w2430_,
		_w2432_,
		_w2433_
	);
	LUT2 #(
		.INIT('h4)
	) name1475 (
		_w2429_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h4)
	) name1476 (
		_w1172_,
		_w1853_,
		_w2435_
	);
	LUT2 #(
		.INIT('h8)
	) name1477 (
		_w2398_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('h4)
	) name1478 (
		\u5_burst_cnt_reg[1]/NET0131 ,
		_w2393_,
		_w2437_
	);
	LUT2 #(
		.INIT('h2)
	) name1479 (
		\u5_burst_cnt_reg[2]/NET0131 ,
		_w2437_,
		_w2438_
	);
	LUT2 #(
		.INIT('h8)
	) name1480 (
		_w1645_,
		_w2374_,
		_w2439_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		_w2438_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h1)
	) name1482 (
		\u5_state_reg[1]/NET0131 ,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('h1)
	) name1483 (
		\u5_state_reg[52]/NET0131 ,
		_w2436_,
		_w2442_
	);
	LUT2 #(
		.INIT('h4)
	) name1484 (
		_w2441_,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('h2)
	) name1485 (
		\u5_burst_cnt_reg[9]/NET0131 ,
		_w2378_,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		_w2383_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h1)
	) name1487 (
		\u5_state_reg[1]/NET0131 ,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h2)
	) name1488 (
		_w2358_,
		_w2388_,
		_w2447_
	);
	LUT2 #(
		.INIT('h4)
	) name1489 (
		_w2358_,
		_w2361_,
		_w2448_
	);
	LUT2 #(
		.INIT('h1)
	) name1490 (
		_w2447_,
		_w2448_,
		_w2449_
	);
	LUT2 #(
		.INIT('h8)
	) name1491 (
		_w2367_,
		_w2449_,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name1492 (
		_w2446_,
		_w2450_,
		_w2451_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		\u5_state_reg[52]/NET0131 ,
		_w2451_,
		_w2452_
	);
	LUT2 #(
		.INIT('h2)
	) name1494 (
		\u5_data_oe_reg/NET0131 ,
		\u7_mc_dqm_r2_reg[0]/P0001 ,
		_w2453_
	);
	LUT2 #(
		.INIT('h2)
	) name1495 (
		\u5_wb_cycle_reg/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w2454_
	);
	LUT2 #(
		.INIT('h1)
	) name1496 (
		\u5_data_oe_reg/NET0131 ,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h1)
	) name1497 (
		\u5_susp_sel_r_reg/NET0131 ,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h4)
	) name1498 (
		_w2453_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h2)
	) name1499 (
		\u5_data_oe_reg/NET0131 ,
		\u7_mc_dqm_r2_reg[1]/P0001 ,
		_w2458_
	);
	LUT2 #(
		.INIT('h2)
	) name1500 (
		_w2456_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('h2)
	) name1501 (
		\u5_data_oe_reg/NET0131 ,
		\u7_mc_dqm_r2_reg[2]/P0001 ,
		_w2460_
	);
	LUT2 #(
		.INIT('h2)
	) name1502 (
		_w2456_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('h2)
	) name1503 (
		\u5_data_oe_reg/NET0131 ,
		\u7_mc_dqm_r2_reg[3]/P0001 ,
		_w2462_
	);
	LUT2 #(
		.INIT('h2)
	) name1504 (
		_w2456_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		\u5_state_reg[2]/NET0131 ,
		_w1631_,
		_w2464_
	);
	LUT2 #(
		.INIT('h1)
	) name1506 (
		\u5_state_reg[2]/NET0131 ,
		_w2324_,
		_w2465_
	);
	LUT2 #(
		.INIT('h8)
	) name1507 (
		_w1654_,
		_w2465_,
		_w2466_
	);
	LUT2 #(
		.INIT('h1)
	) name1508 (
		_w2323_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h8)
	) name1509 (
		_w1750_,
		_w2467_,
		_w2468_
	);
	LUT2 #(
		.INIT('h4)
	) name1510 (
		_w1631_,
		_w2322_,
		_w2469_
	);
	LUT2 #(
		.INIT('h1)
	) name1511 (
		_w2464_,
		_w2469_,
		_w2470_
	);
	LUT2 #(
		.INIT('h4)
	) name1512 (
		_w2468_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h2)
	) name1513 (
		_w1189_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h8)
	) name1514 (
		\u5_ap_en_reg/NET0131 ,
		_w2332_,
		_w2473_
	);
	LUT2 #(
		.INIT('h1)
	) name1515 (
		_w2333_,
		_w2473_,
		_w2474_
	);
	LUT2 #(
		.INIT('h2)
	) name1516 (
		_w1888_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h1)
	) name1517 (
		\u5_tmr_done_reg/NET0131 ,
		_w1270_,
		_w2476_
	);
	LUT2 #(
		.INIT('h2)
	) name1518 (
		_w1714_,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h2)
	) name1519 (
		\u5_state_reg[2]/NET0131 ,
		_w2477_,
		_w2478_
	);
	LUT2 #(
		.INIT('h4)
	) name1520 (
		_w1362_,
		_w1714_,
		_w2479_
	);
	LUT2 #(
		.INIT('h2)
	) name1521 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h4)
	) name1522 (
		\u5_state_reg[2]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2481_
	);
	LUT2 #(
		.INIT('h2)
	) name1523 (
		_w1168_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('h1)
	) name1524 (
		\u5_state_reg[2]/NET0131 ,
		_w2345_,
		_w2483_
	);
	LUT2 #(
		.INIT('h2)
	) name1525 (
		_w2344_,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('h1)
	) name1526 (
		\u5_state_reg[2]/NET0131 ,
		_w1875_,
		_w2485_
	);
	LUT2 #(
		.INIT('h1)
	) name1527 (
		_w2338_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('h8)
	) name1528 (
		_w2341_,
		_w2486_,
		_w2487_
	);
	LUT2 #(
		.INIT('h1)
	) name1529 (
		_w1141_,
		_w1748_,
		_w2488_
	);
	LUT2 #(
		.INIT('h1)
	) name1530 (
		_w2482_,
		_w2484_,
		_w2489_
	);
	LUT2 #(
		.INIT('h8)
	) name1531 (
		_w2488_,
		_w2489_,
		_w2490_
	);
	LUT2 #(
		.INIT('h4)
	) name1532 (
		_w2487_,
		_w2490_,
		_w2491_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		_w2478_,
		_w2480_,
		_w2492_
	);
	LUT2 #(
		.INIT('h8)
	) name1534 (
		_w2491_,
		_w2492_,
		_w2493_
	);
	LUT2 #(
		.INIT('h4)
	) name1535 (
		_w2475_,
		_w2493_,
		_w2494_
	);
	LUT2 #(
		.INIT('h4)
	) name1536 (
		_w2472_,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h8)
	) name1537 (
		_w1287_,
		_w1664_,
		_w2496_
	);
	LUT2 #(
		.INIT('h4)
	) name1538 (
		\u5_state_reg[57]/NET0131 ,
		_w1382_,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		_w1629_,
		_w2497_,
		_w2498_
	);
	LUT2 #(
		.INIT('h8)
	) name1540 (
		_w1883_,
		_w2498_,
		_w2499_
	);
	LUT2 #(
		.INIT('h2)
	) name1541 (
		\u5_state_reg[57]/NET0131 ,
		_w1873_,
		_w2500_
	);
	LUT2 #(
		.INIT('h2)
	) name1542 (
		_w1627_,
		_w2500_,
		_w2501_
	);
	LUT2 #(
		.INIT('h2)
	) name1543 (
		_w1139_,
		_w2501_,
		_w2502_
	);
	LUT2 #(
		.INIT('h8)
	) name1544 (
		\u5_state_reg[57]/NET0131 ,
		_w1377_,
		_w2503_
	);
	LUT2 #(
		.INIT('h2)
	) name1545 (
		_w1627_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('h2)
	) name1546 (
		_w1241_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h1)
	) name1547 (
		_w2496_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h4)
	) name1548 (
		_w2499_,
		_w2506_,
		_w2507_
	);
	LUT2 #(
		.INIT('h4)
	) name1549 (
		_w2502_,
		_w2507_,
		_w2508_
	);
	LUT2 #(
		.INIT('h1)
	) name1550 (
		_w1287_,
		_w1883_,
		_w2509_
	);
	LUT2 #(
		.INIT('h2)
	) name1551 (
		_w1629_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h8)
	) name1552 (
		\u5_state_reg[59]/NET0131 ,
		_w1382_,
		_w2511_
	);
	LUT2 #(
		.INIT('h8)
	) name1553 (
		_w1883_,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		_w2510_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('h1)
	) name1555 (
		_w1817_,
		_w2397_,
		_w2514_
	);
	LUT2 #(
		.INIT('h4)
	) name1556 (
		_w1704_,
		_w1845_,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name1557 (
		\u0_tms_reg[24]/NET0131 ,
		_w1051_,
		_w2516_
	);
	LUT2 #(
		.INIT('h1)
	) name1558 (
		\u0_sp_tms_reg[24]/NET0131 ,
		_w1051_,
		_w2517_
	);
	LUT2 #(
		.INIT('h1)
	) name1559 (
		_w2516_,
		_w2517_,
		_w2518_
	);
	LUT2 #(
		.INIT('h2)
	) name1560 (
		_w1693_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h4)
	) name1561 (
		_w1820_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h2)
	) name1562 (
		\u5_timer_reg[0]/NET0131 ,
		_w1828_,
		_w2521_
	);
	LUT2 #(
		.INIT('h4)
	) name1563 (
		_w1829_,
		_w2288_,
		_w2522_
	);
	LUT2 #(
		.INIT('h4)
	) name1564 (
		_w2521_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h1)
	) name1565 (
		_w2520_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h1)
	) name1566 (
		\u5_state_reg[9]/NET0131 ,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h8)
	) name1567 (
		\u0_tms_reg[4]/NET0131 ,
		_w1051_,
		_w2526_
	);
	LUT2 #(
		.INIT('h2)
	) name1568 (
		\u0_sp_tms_reg[4]/NET0131 ,
		_w1051_,
		_w2527_
	);
	LUT2 #(
		.INIT('h1)
	) name1569 (
		_w2526_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h8)
	) name1570 (
		_w1693_,
		_w2528_,
		_w2529_
	);
	LUT2 #(
		.INIT('h8)
	) name1571 (
		\u5_state_reg[9]/NET0131 ,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h2)
	) name1572 (
		_w1720_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h4)
	) name1573 (
		_w2525_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('h8)
	) name1574 (
		_w1693_,
		_w1806_,
		_w2533_
	);
	LUT2 #(
		.INIT('h1)
	) name1575 (
		_w1719_,
		_w2533_,
		_w2534_
	);
	LUT2 #(
		.INIT('h2)
	) name1576 (
		_w1790_,
		_w2515_,
		_w2535_
	);
	LUT2 #(
		.INIT('h4)
	) name1577 (
		_w2534_,
		_w2535_,
		_w2536_
	);
	LUT2 #(
		.INIT('h4)
	) name1578 (
		_w2532_,
		_w2536_,
		_w2537_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		_w1806_,
		_w2277_,
		_w2538_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		_w1808_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h1)
	) name1581 (
		_w1790_,
		_w2539_,
		_w2540_
	);
	LUT2 #(
		.INIT('h2)
	) name1582 (
		_w1817_,
		_w2540_,
		_w2541_
	);
	LUT2 #(
		.INIT('h4)
	) name1583 (
		_w2537_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h1)
	) name1584 (
		_w2514_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h2)
	) name1585 (
		_w1785_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('h8)
	) name1586 (
		\u0_tms_reg[8]/NET0131 ,
		_w1051_,
		_w2545_
	);
	LUT2 #(
		.INIT('h2)
	) name1587 (
		\u0_sp_tms_reg[8]/NET0131 ,
		_w1051_,
		_w2546_
	);
	LUT2 #(
		.INIT('h1)
	) name1588 (
		_w2545_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h8)
	) name1589 (
		_w1693_,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w1785_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h1)
	) name1591 (
		_w2544_,
		_w2549_,
		_w2550_
	);
	LUT2 #(
		.INIT('h2)
	) name1592 (
		_w1777_,
		_w2550_,
		_w2551_
	);
	LUT2 #(
		.INIT('h8)
	) name1593 (
		\u0_tms_reg[12]/NET0131 ,
		_w1051_,
		_w2552_
	);
	LUT2 #(
		.INIT('h2)
	) name1594 (
		\u0_sp_tms_reg[12]/NET0131 ,
		_w1051_,
		_w2553_
	);
	LUT2 #(
		.INIT('h1)
	) name1595 (
		_w2552_,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h8)
	) name1596 (
		_w1693_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h1)
	) name1597 (
		_w1777_,
		_w2555_,
		_w2556_
	);
	LUT2 #(
		.INIT('h1)
	) name1598 (
		_w2551_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name1599 (
		\u0_sp_tms_reg[13]/NET0131 ,
		_w1051_,
		_w2558_
	);
	LUT2 #(
		.INIT('h8)
	) name1600 (
		\u0_tms_reg[13]/NET0131 ,
		_w1051_,
		_w2559_
	);
	LUT2 #(
		.INIT('h1)
	) name1601 (
		_w2558_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h4)
	) name1602 (
		_w1777_,
		_w2560_,
		_w2561_
	);
	LUT2 #(
		.INIT('h8)
	) name1603 (
		_w1183_,
		_w1693_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name1604 (
		_w1785_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h8)
	) name1605 (
		_w1172_,
		_w1693_,
		_w2564_
	);
	LUT2 #(
		.INIT('h4)
	) name1606 (
		_w1817_,
		_w2564_,
		_w2565_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w1799_,
		_w1800_,
		_w2566_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w1808_,
		_w2566_,
		_w2567_
	);
	LUT2 #(
		.INIT('h8)
	) name1609 (
		_w1808_,
		_w2566_,
		_w2568_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		_w1790_,
		_w2567_,
		_w2569_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		_w2568_,
		_w2569_,
		_w2570_
	);
	LUT2 #(
		.INIT('h4)
	) name1612 (
		\u0_tms_reg[25]/NET0131 ,
		_w1051_,
		_w2571_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		\u0_sp_tms_reg[25]/NET0131 ,
		_w1051_,
		_w2572_
	);
	LUT2 #(
		.INIT('h1)
	) name1614 (
		_w2571_,
		_w2572_,
		_w2573_
	);
	LUT2 #(
		.INIT('h2)
	) name1615 (
		_w1693_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h4)
	) name1616 (
		_w1820_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h2)
	) name1617 (
		\u5_timer_reg[1]/NET0131 ,
		_w1829_,
		_w2576_
	);
	LUT2 #(
		.INIT('h4)
	) name1618 (
		_w1830_,
		_w2288_,
		_w2577_
	);
	LUT2 #(
		.INIT('h4)
	) name1619 (
		_w2576_,
		_w2577_,
		_w2578_
	);
	LUT2 #(
		.INIT('h1)
	) name1620 (
		_w2575_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h1)
	) name1621 (
		\u5_state_reg[9]/NET0131 ,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name1622 (
		\u0_tms_reg[5]/NET0131 ,
		_w1051_,
		_w2581_
	);
	LUT2 #(
		.INIT('h2)
	) name1623 (
		\u0_sp_tms_reg[5]/NET0131 ,
		_w1051_,
		_w2582_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		_w2581_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h8)
	) name1625 (
		_w1693_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h8)
	) name1626 (
		\u5_state_reg[9]/NET0131 ,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h2)
	) name1627 (
		_w1720_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h4)
	) name1628 (
		_w2580_,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('h1)
	) name1629 (
		_w1719_,
		_w1798_,
		_w2588_
	);
	LUT2 #(
		.INIT('h4)
	) name1630 (
		_w1700_,
		_w1845_,
		_w2589_
	);
	LUT2 #(
		.INIT('h2)
	) name1631 (
		_w1790_,
		_w2588_,
		_w2590_
	);
	LUT2 #(
		.INIT('h4)
	) name1632 (
		_w2589_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('h4)
	) name1633 (
		_w2587_,
		_w2591_,
		_w2592_
	);
	LUT2 #(
		.INIT('h1)
	) name1634 (
		_w2570_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h2)
	) name1635 (
		_w1817_,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h2)
	) name1636 (
		_w1785_,
		_w2565_,
		_w2595_
	);
	LUT2 #(
		.INIT('h4)
	) name1637 (
		_w2594_,
		_w2595_,
		_w2596_
	);
	LUT2 #(
		.INIT('h2)
	) name1638 (
		_w1777_,
		_w2563_,
		_w2597_
	);
	LUT2 #(
		.INIT('h4)
	) name1639 (
		_w2596_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name1640 (
		_w2561_,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h1)
	) name1641 (
		_w1778_,
		_w2599_,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		\u5_state_reg[41]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2601_
	);
	LUT2 #(
		.INIT('h2)
	) name1643 (
		\u5_tmr2_done_reg/NET0131 ,
		_w2388_,
		_w2602_
	);
	LUT2 #(
		.INIT('h1)
	) name1644 (
		_w2601_,
		_w2602_,
		_w2603_
	);
	LUT2 #(
		.INIT('h8)
	) name1645 (
		_w1292_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h1)
	) name1646 (
		\u5_state_reg[45]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2605_
	);
	LUT2 #(
		.INIT('h4)
	) name1647 (
		_w2361_,
		_w2365_,
		_w2606_
	);
	LUT2 #(
		.INIT('h2)
	) name1648 (
		\u5_tmr2_done_reg/NET0131 ,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h2)
	) name1649 (
		_w1292_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h1)
	) name1650 (
		_w1136_,
		_w2608_,
		_w2609_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		_w2605_,
		_w2609_,
		_w2610_
	);
	LUT2 #(
		.INIT('h1)
	) name1652 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1689_,
		_w2611_
	);
	LUT2 #(
		.INIT('h8)
	) name1653 (
		\u5_state_reg[46]/NET0131 ,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h1)
	) name1654 (
		_w1148_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h2)
	) name1655 (
		\u5_state_reg[47]/NET0131 ,
		_w2426_,
		_w2614_
	);
	LUT2 #(
		.INIT('h8)
	) name1656 (
		_w1383_,
		_w1438_,
		_w2615_
	);
	LUT2 #(
		.INIT('h1)
	) name1657 (
		_w2614_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h2)
	) name1658 (
		_w1679_,
		_w2616_,
		_w2617_
	);
	LUT2 #(
		.INIT('h1)
	) name1659 (
		_w1679_,
		_w2420_,
		_w2618_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		\u5_state_reg[47]/NET0131 ,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		_w2617_,
		_w2619_,
		_w2620_
	);
	LUT2 #(
		.INIT('h2)
	) name1662 (
		_w1685_,
		_w2620_,
		_w2621_
	);
	LUT2 #(
		.INIT('h4)
	) name1663 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1314_,
		_w2622_
	);
	LUT2 #(
		.INIT('h8)
	) name1664 (
		_w1666_,
		_w1679_,
		_w2623_
	);
	LUT2 #(
		.INIT('h2)
	) name1665 (
		\u5_state_reg[52]/NET0131 ,
		_w2421_,
		_w2624_
	);
	LUT2 #(
		.INIT('h4)
	) name1666 (
		_w2427_,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h1)
	) name1667 (
		_w2623_,
		_w2625_,
		_w2626_
	);
	LUT2 #(
		.INIT('h2)
	) name1668 (
		_w1685_,
		_w2626_,
		_w2627_
	);
	LUT2 #(
		.INIT('h4)
	) name1669 (
		_w1377_,
		_w1627_,
		_w2628_
	);
	LUT2 #(
		.INIT('h8)
	) name1670 (
		_w1241_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h1)
	) name1671 (
		_w2622_,
		_w2629_,
		_w2630_
	);
	LUT2 #(
		.INIT('h4)
	) name1672 (
		_w2627_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h4)
	) name1673 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1312_,
		_w2632_
	);
	LUT2 #(
		.INIT('h2)
	) name1674 (
		\u5_state_reg[58]/NET0131 ,
		_w2426_,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name1675 (
		_w1881_,
		_w2633_,
		_w2634_
	);
	LUT2 #(
		.INIT('h2)
	) name1676 (
		_w1679_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h8)
	) name1677 (
		\u5_state_reg[58]/NET0131 ,
		_w2618_,
		_w2636_
	);
	LUT2 #(
		.INIT('h1)
	) name1678 (
		_w2635_,
		_w2636_,
		_w2637_
	);
	LUT2 #(
		.INIT('h2)
	) name1679 (
		_w1685_,
		_w2637_,
		_w2638_
	);
	LUT2 #(
		.INIT('h1)
	) name1680 (
		_w1287_,
		_w1312_,
		_w2639_
	);
	LUT2 #(
		.INIT('h2)
	) name1681 (
		_w1383_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		_w2632_,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('h4)
	) name1683 (
		_w2638_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		_w2643_
	);
	LUT2 #(
		.INIT('h2)
	) name1685 (
		_w1217_,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h1)
	) name1686 (
		_w1279_,
		_w1295_,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name1687 (
		\u5_tmr_done_reg/NET0131 ,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name1688 (
		\u5_state_reg[5]/NET0131 ,
		_w2646_,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		_w2644_,
		_w2647_,
		_w2648_
	);
	LUT2 #(
		.INIT('h2)
	) name1690 (
		\u5_state_reg[60]/NET0131 ,
		_w2426_,
		_w2649_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w1815_,
		_w2649_,
		_w2650_
	);
	LUT2 #(
		.INIT('h2)
	) name1692 (
		_w1679_,
		_w2650_,
		_w2651_
	);
	LUT2 #(
		.INIT('h8)
	) name1693 (
		\u5_state_reg[60]/NET0131 ,
		_w2618_,
		_w2652_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w2651_,
		_w2652_,
		_w2653_
	);
	LUT2 #(
		.INIT('h2)
	) name1695 (
		_w1685_,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h2)
	) name1696 (
		\u5_state_reg[60]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2655_
	);
	LUT2 #(
		.INIT('h4)
	) name1697 (
		\u7_mc_ack_r_reg/NET0131 ,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h8)
	) name1698 (
		_w1236_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h1)
	) name1699 (
		_w2654_,
		_w2657_,
		_w2658_
	);
	LUT2 #(
		.INIT('h2)
	) name1700 (
		\u5_state_reg[63]/NET0131 ,
		_w2426_,
		_w2659_
	);
	LUT2 #(
		.INIT('h1)
	) name1701 (
		_w1775_,
		_w2659_,
		_w2660_
	);
	LUT2 #(
		.INIT('h2)
	) name1702 (
		_w1679_,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h8)
	) name1703 (
		\u5_state_reg[63]/NET0131 ,
		_w2618_,
		_w2662_
	);
	LUT2 #(
		.INIT('h1)
	) name1704 (
		_w2661_,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('h2)
	) name1705 (
		_w1685_,
		_w2663_,
		_w2664_
	);
	LUT2 #(
		.INIT('h2)
	) name1706 (
		\u5_state_reg[63]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2665_
	);
	LUT2 #(
		.INIT('h4)
	) name1707 (
		\u7_mc_ack_r_reg/NET0131 ,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h8)
	) name1708 (
		_w1102_,
		_w2666_,
		_w2667_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w2664_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h1)
	) name1710 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		_w2669_
	);
	LUT2 #(
		.INIT('h2)
	) name1711 (
		_w1300_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h2)
	) name1712 (
		\u5_tmr_done_reg/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w2671_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		\u5_state_reg[7]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2672_
	);
	LUT2 #(
		.INIT('h1)
	) name1714 (
		_w2671_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h4)
	) name1715 (
		_w1419_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h8)
	) name1716 (
		_w1253_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h1)
	) name1717 (
		_w2670_,
		_w2675_,
		_w2676_
	);
	LUT2 #(
		.INIT('h2)
	) name1718 (
		\u5_state_reg[8]/NET0131 ,
		_w2426_,
		_w2677_
	);
	LUT2 #(
		.INIT('h8)
	) name1719 (
		_w1062_,
		_w2422_,
		_w2678_
	);
	LUT2 #(
		.INIT('h2)
	) name1720 (
		\u2_bank_open_reg/P0001 ,
		_w1375_,
		_w2679_
	);
	LUT2 #(
		.INIT('h8)
	) name1721 (
		\u2_row_same_reg/P0001 ,
		_w2679_,
		_w2680_
	);
	LUT2 #(
		.INIT('h8)
	) name1722 (
		_w2678_,
		_w2680_,
		_w2681_
	);
	LUT2 #(
		.INIT('h1)
	) name1723 (
		_w2677_,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('h2)
	) name1724 (
		_w1679_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h8)
	) name1725 (
		\u5_state_reg[8]/NET0131 ,
		_w2618_,
		_w2684_
	);
	LUT2 #(
		.INIT('h1)
	) name1726 (
		_w2683_,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('h2)
	) name1727 (
		_w1685_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h2)
	) name1728 (
		\u5_wb_wait_r_reg/P0001 ,
		_w1375_,
		_w2687_
	);
	LUT2 #(
		.INIT('h1)
	) name1729 (
		_w1629_,
		_w2687_,
		_w2688_
	);
	LUT2 #(
		.INIT('h2)
	) name1730 (
		_w1093_,
		_w1383_,
		_w2689_
	);
	LUT2 #(
		.INIT('h4)
	) name1731 (
		_w2688_,
		_w2689_,
		_w2690_
	);
	LUT2 #(
		.INIT('h1)
	) name1732 (
		_w2686_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h1)
	) name1733 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1365_,
		_w2692_
	);
	LUT2 #(
		.INIT('h1)
	) name1734 (
		_w2689_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h2)
	) name1735 (
		\u5_state_reg[9]/NET0131 ,
		_w2693_,
		_w2694_
	);
	LUT2 #(
		.INIT('h8)
	) name1736 (
		_w1253_,
		_w2671_,
		_w2695_
	);
	LUT2 #(
		.INIT('h8)
	) name1737 (
		_w1093_,
		_w2688_,
		_w2696_
	);
	LUT2 #(
		.INIT('h1)
	) name1738 (
		_w2695_,
		_w2696_,
		_w2697_
	);
	LUT2 #(
		.INIT('h1)
	) name1739 (
		_w1382_,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w2694_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h8)
	) name1741 (
		_w1119_,
		_w1257_,
		_w2700_
	);
	LUT2 #(
		.INIT('h4)
	) name1742 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1146_,
		_w2701_
	);
	LUT2 #(
		.INIT('h1)
	) name1743 (
		_w2700_,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h8)
	) name1744 (
		\u7_mc_ack_r_reg/NET0131 ,
		_w1102_,
		_w2703_
	);
	LUT2 #(
		.INIT('h1)
	) name1745 (
		_w1721_,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h1)
	) name1746 (
		_w1102_,
		_w1236_,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name1747 (
		\u5_state_reg[65]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2706_
	);
	LUT2 #(
		.INIT('h1)
	) name1748 (
		\u7_mc_ack_r_reg/NET0131 ,
		_w2706_,
		_w2707_
	);
	LUT2 #(
		.INIT('h4)
	) name1749 (
		_w2705_,
		_w2707_,
		_w2708_
	);
	LUT2 #(
		.INIT('h4)
	) name1750 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1300_,
		_w2709_
	);
	LUT2 #(
		.INIT('h2)
	) name1751 (
		\u5_state_reg[6]/NET0131 ,
		_w2426_,
		_w2710_
	);
	LUT2 #(
		.INIT('h2)
	) name1752 (
		_w2678_,
		_w2679_,
		_w2711_
	);
	LUT2 #(
		.INIT('h1)
	) name1753 (
		_w2710_,
		_w2711_,
		_w2712_
	);
	LUT2 #(
		.INIT('h2)
	) name1754 (
		_w1679_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h8)
	) name1755 (
		\u5_state_reg[6]/NET0131 ,
		_w2618_,
		_w2714_
	);
	LUT2 #(
		.INIT('h1)
	) name1756 (
		_w2713_,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h2)
	) name1757 (
		_w1685_,
		_w2715_,
		_w2716_
	);
	LUT2 #(
		.INIT('h2)
	) name1758 (
		\u5_state_reg[6]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2717_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w2403_,
		_w2717_,
		_w2718_
	);
	LUT2 #(
		.INIT('h2)
	) name1760 (
		_w1279_,
		_w2718_,
		_w2719_
	);
	LUT2 #(
		.INIT('h1)
	) name1761 (
		_w2709_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h4)
	) name1762 (
		_w2716_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h1)
	) name1763 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1654_,
		_w2722_
	);
	LUT2 #(
		.INIT('h2)
	) name1764 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1382_,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name1765 (
		_w2722_,
		_w2723_,
		_w2724_
	);
	LUT2 #(
		.INIT('h2)
	) name1766 (
		_w1039_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h8)
	) name1767 (
		_w1654_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h8)
	) name1768 (
		\u5_tmr_done_reg/NET0131 ,
		_w1246_,
		_w2727_
	);
	LUT2 #(
		.INIT('h1)
	) name1769 (
		_w2726_,
		_w2727_,
		_w2728_
	);
	LUT2 #(
		.INIT('h1)
	) name1770 (
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[52]/NET0131 ,
		_w2729_
	);
	LUT2 #(
		.INIT('h2)
	) name1771 (
		\u5_burst_cnt_reg[1]/NET0131 ,
		_w2393_,
		_w2730_
	);
	LUT2 #(
		.INIT('h1)
	) name1772 (
		_w2437_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h2)
	) name1773 (
		_w2729_,
		_w2731_,
		_w2732_
	);
	LUT2 #(
		.INIT('h2)
	) name1774 (
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[52]/NET0131 ,
		_w2733_
	);
	LUT2 #(
		.INIT('h4)
	) name1775 (
		_w2397_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('h8)
	) name1776 (
		_w1175_,
		_w2564_,
		_w2735_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		_w2734_,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('h1)
	) name1778 (
		_w2732_,
		_w2736_,
		_w2737_
	);
	LUT2 #(
		.INIT('h8)
	) name1779 (
		_w2435_,
		_w2734_,
		_w2738_
	);
	LUT2 #(
		.INIT('h4)
	) name1780 (
		\u5_burst_cnt_reg[3]/NET0131 ,
		_w2439_,
		_w2739_
	);
	LUT2 #(
		.INIT('h2)
	) name1781 (
		\u5_burst_cnt_reg[3]/NET0131 ,
		_w2439_,
		_w2740_
	);
	LUT2 #(
		.INIT('h1)
	) name1782 (
		_w2739_,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('h2)
	) name1783 (
		_w2729_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h1)
	) name1784 (
		_w2738_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h8)
	) name1785 (
		\u5_resume_req_r_reg/NET0131 ,
		_w1206_,
		_w2744_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1314_,
		_w2745_
	);
	LUT2 #(
		.INIT('h4)
	) name1787 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1113_,
		_w2746_
	);
	LUT2 #(
		.INIT('h1)
	) name1788 (
		_w2745_,
		_w2746_,
		_w2747_
	);
	LUT2 #(
		.INIT('h4)
	) name1789 (
		\u5_burst_cnt_reg[4]/NET0131 ,
		_w2739_,
		_w2748_
	);
	LUT2 #(
		.INIT('h2)
	) name1790 (
		\u5_burst_cnt_reg[5]/NET0131 ,
		_w2748_,
		_w2749_
	);
	LUT2 #(
		.INIT('h4)
	) name1791 (
		\u5_burst_cnt_reg[5]/NET0131 ,
		_w2748_,
		_w2750_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		_w2749_,
		_w2750_,
		_w2751_
	);
	LUT2 #(
		.INIT('h2)
	) name1793 (
		_w2729_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h2)
	) name1794 (
		\u5_burst_cnt_reg[6]/NET0131 ,
		_w2750_,
		_w2753_
	);
	LUT2 #(
		.INIT('h1)
	) name1795 (
		_w2375_,
		_w2753_,
		_w2754_
	);
	LUT2 #(
		.INIT('h2)
	) name1796 (
		_w2729_,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('h1)
	) name1797 (
		\u5_oe__reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		_w2756_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		\u5_burst_cnt_reg[7]/NET0131 ,
		_w2375_,
		_w2757_
	);
	LUT2 #(
		.INIT('h1)
	) name1799 (
		_w2376_,
		_w2757_,
		_w2758_
	);
	LUT2 #(
		.INIT('h2)
	) name1800 (
		_w2729_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h2)
	) name1801 (
		\u5_burst_cnt_reg[4]/NET0131 ,
		_w2739_,
		_w2760_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		_w2748_,
		_w2760_,
		_w2761_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		_w2729_,
		_w2761_,
		_w2762_
	);
	LUT2 #(
		.INIT('h1)
	) name1804 (
		_w1097_,
		_w1113_,
		_w2763_
	);
	LUT2 #(
		.INIT('h2)
	) name1805 (
		\u5_state_reg[48]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2764_
	);
	LUT2 #(
		.INIT('h4)
	) name1806 (
		_w2763_,
		_w2764_,
		_w2765_
	);
	LUT2 #(
		.INIT('h1)
	) name1807 (
		_w1230_,
		_w2765_,
		_w2766_
	);
	LUT2 #(
		.INIT('h4)
	) name1808 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1221_,
		_w2767_
	);
	LUT2 #(
		.INIT('h8)
	) name1809 (
		_w1189_,
		_w1657_,
		_w2768_
	);
	LUT2 #(
		.INIT('h8)
	) name1810 (
		\u5_state_reg[15]/NET0131 ,
		_w1654_,
		_w2769_
	);
	LUT2 #(
		.INIT('h1)
	) name1811 (
		_w2724_,
		_w2769_,
		_w2770_
	);
	LUT2 #(
		.INIT('h2)
	) name1812 (
		_w1039_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h4)
	) name1813 (
		_w1382_,
		_w1888_,
		_w2772_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		_w1655_,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h1)
	) name1815 (
		_w2767_,
		_w2773_,
		_w2774_
	);
	LUT2 #(
		.INIT('h4)
	) name1816 (
		_w2768_,
		_w2774_,
		_w2775_
	);
	LUT2 #(
		.INIT('h4)
	) name1817 (
		_w2771_,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('h8)
	) name1818 (
		_w1139_,
		_w1874_,
		_w2777_
	);
	LUT2 #(
		.INIT('h8)
	) name1819 (
		_w1627_,
		_w1654_,
		_w2778_
	);
	LUT2 #(
		.INIT('h2)
	) name1820 (
		_w1023_,
		_w2778_,
		_w2779_
	);
	LUT2 #(
		.INIT('h1)
	) name1821 (
		_w2777_,
		_w2779_,
		_w2780_
	);
	LUT2 #(
		.INIT('h4)
	) name1822 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[14]/NET0131 ,
		_w2781_
	);
	LUT2 #(
		.INIT('h8)
	) name1823 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1382_,
		_w2782_
	);
	LUT2 #(
		.INIT('h4)
	) name1824 (
		_w2333_,
		_w2782_,
		_w2783_
	);
	LUT2 #(
		.INIT('h1)
	) name1825 (
		_w2781_,
		_w2783_,
		_w2784_
	);
	LUT2 #(
		.INIT('h2)
	) name1826 (
		_w1397_,
		_w2784_,
		_w2785_
	);
	LUT2 #(
		.INIT('h2)
	) name1827 (
		_w1189_,
		_w2324_,
		_w2786_
	);
	LUT2 #(
		.INIT('h4)
	) name1828 (
		_w2322_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h8)
	) name1829 (
		_w1654_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h8)
	) name1830 (
		_w1750_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h1)
	) name1831 (
		_w1752_,
		_w2785_,
		_w2790_
	);
	LUT2 #(
		.INIT('h4)
	) name1832 (
		_w2789_,
		_w2790_,
		_w2791_
	);
	LUT2 #(
		.INIT('h8)
	) name1833 (
		\u5_data_oe_reg/NET0131 ,
		\u5_mc_c_oe_reg/NET0131 ,
		_w2792_
	);
	LUT2 #(
		.INIT('h4)
	) name1834 (
		\u5_susp_sel_r_reg/NET0131 ,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h1)
	) name1835 (
		\u5_state_reg[24]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name1836 (
		\u5_ir_cnt_done_reg/P0001 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2795_
	);
	LUT2 #(
		.INIT('h2)
	) name1837 (
		_w1131_,
		_w2795_,
		_w2796_
	);
	LUT2 #(
		.INIT('h1)
	) name1838 (
		_w1203_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w2794_,
		_w2797_,
		_w2798_
	);
	LUT2 #(
		.INIT('h4)
	) name1840 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1401_,
		_w2799_
	);
	LUT2 #(
		.INIT('h1)
	) name1841 (
		_w2798_,
		_w2799_,
		_w2800_
	);
	LUT2 #(
		.INIT('h2)
	) name1842 (
		\u6_wb_first_r_reg/NET0131 ,
		wb_ack_o_pad,
		_w2801_
	);
	LUT2 #(
		.INIT('h4)
	) name1843 (
		wb_err_o_pad,
		_w2801_,
		_w2802_
	);
	LUT2 #(
		.INIT('h1)
	) name1844 (
		\u6_read_go_r_reg/NET0131 ,
		\u6_write_go_r_reg/NET0131 ,
		_w2803_
	);
	LUT2 #(
		.INIT('h8)
	) name1845 (
		_w1046_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h8)
	) name1846 (
		_w2269_,
		_w2804_,
		_w2805_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		_w2802_,
		_w2805_,
		_w2806_
	);
	LUT2 #(
		.INIT('h2)
	) name1848 (
		wb_stb_i_pad,
		_w2806_,
		_w2807_
	);
	LUT2 #(
		.INIT('h1)
	) name1849 (
		\u5_wb_stb_first_reg/NET0131 ,
		_w2807_,
		_w2808_
	);
	LUT2 #(
		.INIT('h1)
	) name1850 (
		_w1896_,
		_w2808_,
		_w2809_
	);
	LUT2 #(
		.INIT('h1)
	) name1851 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		_w2810_
	);
	LUT2 #(
		.INIT('h2)
	) name1852 (
		_w1070_,
		_w2810_,
		_w2811_
	);
	LUT2 #(
		.INIT('h4)
	) name1853 (
		\u5_tmr_done_reg/NET0131 ,
		_w1080_,
		_w2812_
	);
	LUT2 #(
		.INIT('h1)
	) name1854 (
		_w2811_,
		_w2812_,
		_w2813_
	);
	LUT2 #(
		.INIT('h8)
	) name1855 (
		_w1023_,
		_w2778_,
		_w2814_
	);
	LUT2 #(
		.INIT('h1)
	) name1856 (
		\u5_state_reg[54]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2815_
	);
	LUT2 #(
		.INIT('h2)
	) name1857 (
		_w1113_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('h1)
	) name1858 (
		_w2814_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h8)
	) name1859 (
		_w1283_,
		_w1662_,
		_w2818_
	);
	LUT2 #(
		.INIT('h8)
	) name1860 (
		_w1700_,
		_w2818_,
		_w2819_
	);
	LUT2 #(
		.INIT('h4)
	) name1861 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1097_,
		_w2820_
	);
	LUT2 #(
		.INIT('h1)
	) name1862 (
		_w1230_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('h8)
	) name1863 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1097_,
		_w2822_
	);
	LUT2 #(
		.INIT('h8)
	) name1864 (
		_w2821_,
		_w2822_,
		_w2823_
	);
	LUT2 #(
		.INIT('h4)
	) name1865 (
		_w1704_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h8)
	) name1866 (
		_w1283_,
		_w1440_,
		_w2825_
	);
	LUT2 #(
		.INIT('h1)
	) name1867 (
		_w1314_,
		_w2825_,
		_w2826_
	);
	LUT2 #(
		.INIT('h2)
	) name1868 (
		_w1693_,
		_w2821_,
		_w2827_
	);
	LUT2 #(
		.INIT('h8)
	) name1869 (
		_w1781_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h2)
	) name1870 (
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w2829_
	);
	LUT2 #(
		.INIT('h4)
	) name1871 (
		_w2562_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h1)
	) name1872 (
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w2831_
	);
	LUT2 #(
		.INIT('h4)
	) name1873 (
		\u5_state_reg[36]/NET0131 ,
		_w987_,
		_w2832_
	);
	LUT2 #(
		.INIT('h4)
	) name1874 (
		\u5_state_reg[41]/NET0131 ,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h1)
	) name1875 (
		_w2564_,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h1)
	) name1876 (
		\u5_timer2_reg[0]/P0001 ,
		\u5_timer2_reg[1]/P0001 ,
		_w2835_
	);
	LUT2 #(
		.INIT('h4)
	) name1877 (
		\u5_timer2_reg[2]/P0001 ,
		_w2835_,
		_w2836_
	);
	LUT2 #(
		.INIT('h4)
	) name1878 (
		\u5_timer2_reg[3]/P0001 ,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h4)
	) name1879 (
		\u5_timer2_reg[4]/P0001 ,
		_w2837_,
		_w2838_
	);
	LUT2 #(
		.INIT('h4)
	) name1880 (
		\u5_timer2_reg[5]/P0001 ,
		_w2838_,
		_w2839_
	);
	LUT2 #(
		.INIT('h4)
	) name1881 (
		\u5_timer2_reg[6]/P0001 ,
		_w2839_,
		_w2840_
	);
	LUT2 #(
		.INIT('h4)
	) name1882 (
		\u5_timer2_reg[7]/P0001 ,
		_w2840_,
		_w2841_
	);
	LUT2 #(
		.INIT('h4)
	) name1883 (
		\u5_timer2_reg[8]/P0001 ,
		_w2841_,
		_w2842_
	);
	LUT2 #(
		.INIT('h2)
	) name1884 (
		_w2833_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h2)
	) name1885 (
		\u5_timer2_reg[2]/P0001 ,
		_w2835_,
		_w2844_
	);
	LUT2 #(
		.INIT('h1)
	) name1886 (
		_w2836_,
		_w2844_,
		_w2845_
	);
	LUT2 #(
		.INIT('h2)
	) name1887 (
		_w2843_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h1)
	) name1888 (
		_w2834_,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('h2)
	) name1889 (
		_w2831_,
		_w2847_,
		_w2848_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		_w2830_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h1)
	) name1891 (
		_w2822_,
		_w2849_,
		_w2850_
	);
	LUT2 #(
		.INIT('h2)
	) name1892 (
		\u5_state_reg[51]/NET0131 ,
		_w1794_,
		_w2851_
	);
	LUT2 #(
		.INIT('h2)
	) name1893 (
		_w2821_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h4)
	) name1894 (
		_w2850_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('h1)
	) name1895 (
		_w2828_,
		_w2853_,
		_w2854_
	);
	LUT2 #(
		.INIT('h4)
	) name1896 (
		_w2824_,
		_w2826_,
		_w2855_
	);
	LUT2 #(
		.INIT('h4)
	) name1897 (
		_w2854_,
		_w2855_,
		_w2856_
	);
	LUT2 #(
		.INIT('h1)
	) name1898 (
		_w2819_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('h1)
	) name1899 (
		\u5_cs_le_reg/P0001 ,
		wb_we_i_pad,
		_w2858_
	);
	LUT2 #(
		.INIT('h8)
	) name1900 (
		\u5_state_reg[37]/NET0131 ,
		_w2365_,
		_w2859_
	);
	LUT2 #(
		.INIT('h2)
	) name1901 (
		_w988_,
		_w2859_,
		_w2860_
	);
	LUT2 #(
		.INIT('h2)
	) name1902 (
		\u5_tmr2_done_reg/NET0131 ,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h8)
	) name1903 (
		\u1_u0_out_r_reg[12]/P0001 ,
		_w2861_,
		_w2862_
	);
	LUT2 #(
		.INIT('h8)
	) name1904 (
		\u1_acs_addr_reg[12]/P0001 ,
		_w2862_,
		_w2863_
	);
	LUT2 #(
		.INIT('h8)
	) name1905 (
		\u1_acs_addr_reg[13]/P0001 ,
		_w2863_,
		_w2864_
	);
	LUT2 #(
		.INIT('h8)
	) name1906 (
		\u1_acs_addr_reg[14]/P0001 ,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h8)
	) name1907 (
		\u1_acs_addr_reg[15]/P0001 ,
		_w2865_,
		_w2866_
	);
	LUT2 #(
		.INIT('h8)
	) name1908 (
		\u1_acs_addr_reg[16]/P0001 ,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h8)
	) name1909 (
		\u1_acs_addr_reg[17]/P0001 ,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('h8)
	) name1910 (
		\u1_acs_addr_reg[18]/P0001 ,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		\u1_acs_addr_reg[19]/P0001 ,
		_w2869_,
		_w2870_
	);
	LUT2 #(
		.INIT('h8)
	) name1912 (
		\u1_acs_addr_reg[20]/P0001 ,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h8)
	) name1913 (
		\u1_acs_addr_reg[21]/P0001 ,
		_w2871_,
		_w2872_
	);
	LUT2 #(
		.INIT('h8)
	) name1914 (
		\u1_acs_addr_reg[22]/P0001 ,
		_w2872_,
		_w2873_
	);
	LUT2 #(
		.INIT('h2)
	) name1915 (
		\u1_acs_addr_reg[23]/P0001 ,
		_w2873_,
		_w2874_
	);
	LUT2 #(
		.INIT('h4)
	) name1916 (
		\u1_acs_addr_reg[23]/P0001 ,
		_w2873_,
		_w2875_
	);
	LUT2 #(
		.INIT('h2)
	) name1917 (
		_w2858_,
		_w2874_,
		_w2876_
	);
	LUT2 #(
		.INIT('h4)
	) name1918 (
		_w2875_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('h2)
	) name1919 (
		_w2361_,
		_w2365_,
		_w2878_
	);
	LUT2 #(
		.INIT('h8)
	) name1920 (
		\wb_addr_i[25]_pad ,
		_w2878_,
		_w2879_
	);
	LUT2 #(
		.INIT('h8)
	) name1921 (
		\wb_addr_i[24]_pad ,
		_w2606_,
		_w2880_
	);
	LUT2 #(
		.INIT('h8)
	) name1922 (
		\wb_addr_i[23]_pad ,
		_w2388_,
		_w2881_
	);
	LUT2 #(
		.INIT('h1)
	) name1923 (
		_w2858_,
		_w2879_,
		_w2882_
	);
	LUT2 #(
		.INIT('h1)
	) name1924 (
		_w2880_,
		_w2881_,
		_w2883_
	);
	LUT2 #(
		.INIT('h8)
	) name1925 (
		_w2882_,
		_w2883_,
		_w2884_
	);
	LUT2 #(
		.INIT('h1)
	) name1926 (
		_w2877_,
		_w2884_,
		_w2885_
	);
	LUT2 #(
		.INIT('h4)
	) name1927 (
		_w1704_,
		_w2818_,
		_w2886_
	);
	LUT2 #(
		.INIT('h4)
	) name1928 (
		_w1708_,
		_w2823_,
		_w2887_
	);
	LUT2 #(
		.INIT('h8)
	) name1929 (
		_w2560_,
		_w2827_,
		_w2888_
	);
	LUT2 #(
		.INIT('h1)
	) name1930 (
		_w2397_,
		_w2833_,
		_w2889_
	);
	LUT2 #(
		.INIT('h8)
	) name1931 (
		\u5_timer2_reg[0]/P0001 ,
		\u5_timer2_reg[1]/P0001 ,
		_w2890_
	);
	LUT2 #(
		.INIT('h1)
	) name1932 (
		_w2835_,
		_w2890_,
		_w2891_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		_w2843_,
		_w2891_,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name1934 (
		_w2889_,
		_w2892_,
		_w2893_
	);
	LUT2 #(
		.INIT('h2)
	) name1935 (
		_w2831_,
		_w2893_,
		_w2894_
	);
	LUT2 #(
		.INIT('h4)
	) name1936 (
		_w2548_,
		_w2829_,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name1937 (
		_w2894_,
		_w2895_,
		_w2896_
	);
	LUT2 #(
		.INIT('h1)
	) name1938 (
		_w2822_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h2)
	) name1939 (
		\u5_state_reg[51]/NET0131 ,
		_w1798_,
		_w2898_
	);
	LUT2 #(
		.INIT('h2)
	) name1940 (
		_w2821_,
		_w2898_,
		_w2899_
	);
	LUT2 #(
		.INIT('h4)
	) name1941 (
		_w2897_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('h1)
	) name1942 (
		_w2888_,
		_w2900_,
		_w2901_
	);
	LUT2 #(
		.INIT('h1)
	) name1943 (
		_w2887_,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('h2)
	) name1944 (
		_w2826_,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h1)
	) name1945 (
		_w2886_,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h4)
	) name1946 (
		_w1696_,
		_w2818_,
		_w2905_
	);
	LUT2 #(
		.INIT('h2)
	) name1947 (
		_w2277_,
		_w2821_,
		_w2906_
	);
	LUT2 #(
		.INIT('h4)
	) name1948 (
		_w1700_,
		_w2822_,
		_w2907_
	);
	LUT2 #(
		.INIT('h2)
	) name1949 (
		\u5_state_reg[51]/NET0131 ,
		_w2282_,
		_w2908_
	);
	LUT2 #(
		.INIT('h8)
	) name1950 (
		_w1693_,
		_w1788_,
		_w2909_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		_w2829_,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h2)
	) name1952 (
		_w2836_,
		_w2842_,
		_w2911_
	);
	LUT2 #(
		.INIT('h2)
	) name1953 (
		\u5_timer2_reg[3]/P0001 ,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h2)
	) name1954 (
		_w2837_,
		_w2842_,
		_w2913_
	);
	LUT2 #(
		.INIT('h2)
	) name1955 (
		_w2833_,
		_w2913_,
		_w2914_
	);
	LUT2 #(
		.INIT('h4)
	) name1956 (
		_w2912_,
		_w2914_,
		_w2915_
	);
	LUT2 #(
		.INIT('h2)
	) name1957 (
		_w1853_,
		_w2833_,
		_w2916_
	);
	LUT2 #(
		.INIT('h2)
	) name1958 (
		_w2831_,
		_w2915_,
		_w2917_
	);
	LUT2 #(
		.INIT('h4)
	) name1959 (
		_w2916_,
		_w2917_,
		_w2918_
	);
	LUT2 #(
		.INIT('h1)
	) name1960 (
		_w2910_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name1961 (
		_w2822_,
		_w2919_,
		_w2920_
	);
	LUT2 #(
		.INIT('h2)
	) name1962 (
		_w2821_,
		_w2907_,
		_w2921_
	);
	LUT2 #(
		.INIT('h4)
	) name1963 (
		_w2908_,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h4)
	) name1964 (
		_w2920_,
		_w2922_,
		_w2923_
	);
	LUT2 #(
		.INIT('h2)
	) name1965 (
		_w2826_,
		_w2906_,
		_w2924_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		_w2923_,
		_w2924_,
		_w2925_
	);
	LUT2 #(
		.INIT('h1)
	) name1967 (
		_w2905_,
		_w2925_,
		_w2926_
	);
	LUT2 #(
		.INIT('h2)
	) name1968 (
		_w1686_,
		_w2424_,
		_w2927_
	);
	LUT2 #(
		.INIT('h1)
	) name1969 (
		_w1093_,
		_w1287_,
		_w2928_
	);
	LUT2 #(
		.INIT('h4)
	) name1970 (
		_w2927_,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('h2)
	) name1971 (
		_w1383_,
		_w2929_,
		_w2930_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		_w1230_,
		_w1312_,
		_w2931_
	);
	LUT2 #(
		.INIT('h4)
	) name1973 (
		_w1238_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h8)
	) name1974 (
		_w1398_,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h4)
	) name1975 (
		_w2930_,
		_w2933_,
		_w2934_
	);
	LUT2 #(
		.INIT('h8)
	) name1976 (
		_w1713_,
		_w2934_,
		_w2935_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		\u5_wr_cycle_reg/NET0131 ,
		_w2935_,
		_w2936_
	);
	LUT2 #(
		.INIT('h8)
	) name1978 (
		\u5_data_oe_r2_reg/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w2937_
	);
	LUT2 #(
		.INIT('h1)
	) name1979 (
		_w2936_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h2)
	) name1980 (
		_w1303_,
		_w1358_,
		_w2939_
	);
	LUT2 #(
		.INIT('h1)
	) name1981 (
		_w1214_,
		_w1401_,
		_w2940_
	);
	LUT2 #(
		.INIT('h2)
	) name1982 (
		_w1276_,
		_w1364_,
		_w2941_
	);
	LUT2 #(
		.INIT('h4)
	) name1983 (
		_w1217_,
		_w2479_,
		_w2942_
	);
	LUT2 #(
		.INIT('h8)
	) name1984 (
		_w1128_,
		_w2942_,
		_w2943_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		_w2941_,
		_w2943_,
		_w2944_
	);
	LUT2 #(
		.INIT('h8)
	) name1986 (
		_w2940_,
		_w2944_,
		_w2945_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		_w1232_,
		_w1397_,
		_w2946_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		_w1164_,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('h1)
	) name1989 (
		_w1195_,
		_w1203_,
		_w2948_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		_w1039_,
		_w1189_,
		_w2949_
	);
	LUT2 #(
		.INIT('h8)
	) name1991 (
		_w2948_,
		_w2949_,
		_w2950_
	);
	LUT2 #(
		.INIT('h8)
	) name1992 (
		_w1316_,
		_w2950_,
		_w2951_
	);
	LUT2 #(
		.INIT('h4)
	) name1993 (
		_w1168_,
		_w1201_,
		_w2952_
	);
	LUT2 #(
		.INIT('h8)
	) name1994 (
		_w2951_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h8)
	) name1995 (
		_w2947_,
		_w2953_,
		_w2954_
	);
	LUT2 #(
		.INIT('h8)
	) name1996 (
		_w1298_,
		_w2939_,
		_w2955_
	);
	LUT2 #(
		.INIT('h8)
	) name1997 (
		_w2954_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h8)
	) name1998 (
		_w2945_,
		_w2956_,
		_w2957_
	);
	LUT2 #(
		.INIT('h1)
	) name1999 (
		_w1039_,
		_w2957_,
		_w2958_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		\u5_cnt_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w2959_
	);
	LUT2 #(
		.INIT('h8)
	) name2001 (
		_w1654_,
		_w2959_,
		_w2960_
	);
	LUT2 #(
		.INIT('h8)
	) name2002 (
		_w1629_,
		_w2960_,
		_w2961_
	);
	LUT2 #(
		.INIT('h1)
	) name2003 (
		mc_cke_pad_o__pad,
		_w2960_,
		_w2962_
	);
	LUT2 #(
		.INIT('h2)
	) name2004 (
		_w1039_,
		_w2961_,
		_w2963_
	);
	LUT2 #(
		.INIT('h4)
	) name2005 (
		_w2962_,
		_w2963_,
		_w2964_
	);
	LUT2 #(
		.INIT('h1)
	) name2006 (
		_w2958_,
		_w2964_,
		_w2965_
	);
	LUT2 #(
		.INIT('h2)
	) name2007 (
		\u5_cke_r_reg/NET0131 ,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h4)
	) name2008 (
		_w1309_,
		_w2948_,
		_w2967_
	);
	LUT2 #(
		.INIT('h1)
	) name2009 (
		\u5_tmr_done_reg/NET0131 ,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('h8)
	) name2010 (
		\u5_state_reg[0]/NET0131 ,
		_w2968_,
		_w2969_
	);
	LUT2 #(
		.INIT('h8)
	) name2011 (
		\wb_addr_i[20]_pad ,
		_w2606_,
		_w2970_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		\wb_addr_i[19]_pad ,
		_w2388_,
		_w2971_
	);
	LUT2 #(
		.INIT('h8)
	) name2013 (
		\wb_addr_i[21]_pad ,
		_w2878_,
		_w2972_
	);
	LUT2 #(
		.INIT('h1)
	) name2014 (
		_w2970_,
		_w2971_,
		_w2973_
	);
	LUT2 #(
		.INIT('h4)
	) name2015 (
		_w2972_,
		_w2973_,
		_w2974_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		_w2858_,
		_w2974_,
		_w2975_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		\u1_acs_addr_reg[19]/P0001 ,
		_w2869_,
		_w2976_
	);
	LUT2 #(
		.INIT('h2)
	) name2018 (
		_w2858_,
		_w2870_,
		_w2977_
	);
	LUT2 #(
		.INIT('h4)
	) name2019 (
		_w2976_,
		_w2977_,
		_w2978_
	);
	LUT2 #(
		.INIT('h1)
	) name2020 (
		_w2975_,
		_w2978_,
		_w2979_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		\wb_addr_i[22]_pad ,
		_w2388_,
		_w2980_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		\wb_addr_i[24]_pad ,
		_w2878_,
		_w2981_
	);
	LUT2 #(
		.INIT('h8)
	) name2023 (
		\wb_addr_i[23]_pad ,
		_w2606_,
		_w2982_
	);
	LUT2 #(
		.INIT('h1)
	) name2024 (
		_w2980_,
		_w2981_,
		_w2983_
	);
	LUT2 #(
		.INIT('h4)
	) name2025 (
		_w2982_,
		_w2983_,
		_w2984_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		_w2858_,
		_w2984_,
		_w2985_
	);
	LUT2 #(
		.INIT('h1)
	) name2027 (
		\u1_acs_addr_reg[22]/P0001 ,
		_w2872_,
		_w2986_
	);
	LUT2 #(
		.INIT('h2)
	) name2028 (
		_w2858_,
		_w2873_,
		_w2987_
	);
	LUT2 #(
		.INIT('h4)
	) name2029 (
		_w2986_,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h1)
	) name2030 (
		_w2985_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h8)
	) name2031 (
		_w1040_,
		_w1654_,
		_w2990_
	);
	LUT2 #(
		.INIT('h8)
	) name2032 (
		_w1629_,
		_w2990_,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name2033 (
		\u5_cke_r_reg/NET0131 ,
		_w2990_,
		_w2992_
	);
	LUT2 #(
		.INIT('h1)
	) name2034 (
		_w1189_,
		_w2991_,
		_w2993_
	);
	LUT2 #(
		.INIT('h4)
	) name2035 (
		_w2992_,
		_w2993_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name2036 (
		\u5_cnt_reg/NET0131 ,
		_w1629_,
		_w2995_
	);
	LUT2 #(
		.INIT('h8)
	) name2037 (
		\u5_cke_r_reg/NET0131 ,
		\u5_cnt_reg/NET0131 ,
		_w2996_
	);
	LUT2 #(
		.INIT('h1)
	) name2038 (
		_w2995_,
		_w2996_,
		_w2997_
	);
	LUT2 #(
		.INIT('h8)
	) name2039 (
		_w1189_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h1)
	) name2040 (
		_w1397_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h1)
	) name2041 (
		_w2994_,
		_w2999_,
		_w3000_
	);
	LUT2 #(
		.INIT('h4)
	) name2042 (
		_w1206_,
		_w2954_,
		_w3001_
	);
	LUT2 #(
		.INIT('h8)
	) name2043 (
		_w1304_,
		_w1398_,
		_w3002_
	);
	LUT2 #(
		.INIT('h8)
	) name2044 (
		_w3001_,
		_w3002_,
		_w3003_
	);
	LUT2 #(
		.INIT('h8)
	) name2045 (
		_w2945_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h1)
	) name2046 (
		_w3000_,
		_w3004_,
		_w3005_
	);
	LUT2 #(
		.INIT('h4)
	) name2047 (
		_w1798_,
		_w2818_,
		_w3006_
	);
	LUT2 #(
		.INIT('h8)
	) name2048 (
		_w2821_,
		_w2826_,
		_w3007_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		_w2822_,
		_w3007_,
		_w3008_
	);
	LUT2 #(
		.INIT('h8)
	) name2050 (
		\u5_state_reg[51]/NET0131 ,
		_w2574_,
		_w3009_
	);
	LUT2 #(
		.INIT('h2)
	) name2051 (
		\u5_timer2_reg[5]/P0001 ,
		_w2838_,
		_w3010_
	);
	LUT2 #(
		.INIT('h1)
	) name2052 (
		_w2839_,
		_w3010_,
		_w3011_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		\u5_state_reg[40]/NET0131 ,
		_w3011_,
		_w3012_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		_w2843_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h1)
	) name2055 (
		\u5_state_reg[40]/NET0131 ,
		_w2833_,
		_w3014_
	);
	LUT2 #(
		.INIT('h4)
	) name2056 (
		_w2529_,
		_w3014_,
		_w3015_
	);
	LUT2 #(
		.INIT('h1)
	) name2057 (
		\u5_state_reg[51]/NET0131 ,
		_w3013_,
		_w3016_
	);
	LUT2 #(
		.INIT('h4)
	) name2058 (
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT2 #(
		.INIT('h2)
	) name2059 (
		_w3008_,
		_w3009_,
		_w3018_
	);
	LUT2 #(
		.INIT('h4)
	) name2060 (
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h1)
	) name2061 (
		_w3006_,
		_w3019_,
		_w3020_
	);
	LUT2 #(
		.INIT('h1)
	) name2062 (
		\u1_acs_addr_reg[20]/P0001 ,
		_w2870_,
		_w3021_
	);
	LUT2 #(
		.INIT('h1)
	) name2063 (
		_w2871_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h2)
	) name2064 (
		_w2858_,
		_w3022_,
		_w3023_
	);
	LUT2 #(
		.INIT('h8)
	) name2065 (
		\wb_addr_i[22]_pad ,
		_w2878_,
		_w3024_
	);
	LUT2 #(
		.INIT('h8)
	) name2066 (
		\wb_addr_i[21]_pad ,
		_w2606_,
		_w3025_
	);
	LUT2 #(
		.INIT('h8)
	) name2067 (
		\wb_addr_i[20]_pad ,
		_w2388_,
		_w3026_
	);
	LUT2 #(
		.INIT('h1)
	) name2068 (
		_w2858_,
		_w3024_,
		_w3027_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		_w3025_,
		_w3026_,
		_w3028_
	);
	LUT2 #(
		.INIT('h8)
	) name2070 (
		_w3027_,
		_w3028_,
		_w3029_
	);
	LUT2 #(
		.INIT('h1)
	) name2071 (
		_w3023_,
		_w3029_,
		_w3030_
	);
	LUT2 #(
		.INIT('h4)
	) name2072 (
		_w1696_,
		_w2822_,
		_w3031_
	);
	LUT2 #(
		.INIT('h1)
	) name2073 (
		\u5_state_reg[51]/NET0131 ,
		_w2822_,
		_w3032_
	);
	LUT2 #(
		.INIT('h4)
	) name2074 (
		_w2308_,
		_w3014_,
		_w3033_
	);
	LUT2 #(
		.INIT('h2)
	) name2075 (
		\u5_state_reg[40]/NET0131 ,
		_w2315_,
		_w3034_
	);
	LUT2 #(
		.INIT('h8)
	) name2076 (
		_w985_,
		_w2832_,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name2077 (
		\u5_timer2_reg[4]/P0001 ,
		_w2913_,
		_w3036_
	);
	LUT2 #(
		.INIT('h8)
	) name2078 (
		\u5_timer2_reg[4]/P0001 ,
		_w2913_,
		_w3037_
	);
	LUT2 #(
		.INIT('h2)
	) name2079 (
		_w3035_,
		_w3036_,
		_w3038_
	);
	LUT2 #(
		.INIT('h4)
	) name2080 (
		_w3037_,
		_w3038_,
		_w3039_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w3033_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h4)
	) name2082 (
		_w3034_,
		_w3040_,
		_w3041_
	);
	LUT2 #(
		.INIT('h2)
	) name2083 (
		_w3032_,
		_w3041_,
		_w3042_
	);
	LUT2 #(
		.INIT('h2)
	) name2084 (
		\u5_state_reg[51]/NET0131 ,
		_w2519_,
		_w3043_
	);
	LUT2 #(
		.INIT('h1)
	) name2085 (
		_w3031_,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h4)
	) name2086 (
		_w3042_,
		_w3044_,
		_w3045_
	);
	LUT2 #(
		.INIT('h2)
	) name2087 (
		_w3007_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('h4)
	) name2088 (
		_w2533_,
		_w2818_,
		_w3047_
	);
	LUT2 #(
		.INIT('h1)
	) name2089 (
		_w3046_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h2)
	) name2090 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		_w3049_
	);
	LUT2 #(
		.INIT('h2)
	) name2091 (
		\u5_state_reg[7]/NET0131 ,
		_w1375_,
		_w3050_
	);
	LUT2 #(
		.INIT('h8)
	) name2092 (
		_w1623_,
		_w3050_,
		_w3051_
	);
	LUT2 #(
		.INIT('h8)
	) name2093 (
		_w3049_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		_w960_,
		_w996_,
		_w3053_
	);
	LUT2 #(
		.INIT('h8)
	) name2095 (
		_w992_,
		_w1143_,
		_w3054_
	);
	LUT2 #(
		.INIT('h8)
	) name2096 (
		_w3053_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h1)
	) name2097 (
		\u5_state_reg[22]/NET0131 ,
		_w1213_,
		_w3056_
	);
	LUT2 #(
		.INIT('h4)
	) name2098 (
		_w1394_,
		_w3056_,
		_w3057_
	);
	LUT2 #(
		.INIT('h8)
	) name2099 (
		_w1133_,
		_w1155_,
		_w3058_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		\u5_state_reg[22]/NET0131 ,
		_w1000_,
		_w3059_
	);
	LUT2 #(
		.INIT('h4)
	) name2101 (
		\u5_state_reg[21]/NET0131 ,
		_w991_,
		_w3060_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		_w999_,
		_w3060_,
		_w3061_
	);
	LUT2 #(
		.INIT('h8)
	) name2103 (
		_w1011_,
		_w1074_,
		_w3062_
	);
	LUT2 #(
		.INIT('h4)
	) name2104 (
		_w3059_,
		_w3062_,
		_w3063_
	);
	LUT2 #(
		.INIT('h4)
	) name2105 (
		_w3057_,
		_w3061_,
		_w3064_
	);
	LUT2 #(
		.INIT('h8)
	) name2106 (
		_w3063_,
		_w3064_,
		_w3065_
	);
	LUT2 #(
		.INIT('h8)
	) name2107 (
		_w3055_,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('h8)
	) name2108 (
		_w3058_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h1)
	) name2109 (
		\u5_state_reg[20]/NET0131 ,
		_w3067_,
		_w3068_
	);
	LUT2 #(
		.INIT('h2)
	) name2110 (
		_w1002_,
		_w3068_,
		_w3069_
	);
	LUT2 #(
		.INIT('h1)
	) name2111 (
		_w1069_,
		_w3069_,
		_w3070_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		\u5_state_reg[21]/NET0131 ,
		\u5_state_reg[23]/NET0131 ,
		_w3071_
	);
	LUT2 #(
		.INIT('h8)
	) name2113 (
		_w1007_,
		_w3071_,
		_w3072_
	);
	LUT2 #(
		.INIT('h8)
	) name2114 (
		_w1338_,
		_w3072_,
		_w3073_
	);
	LUT2 #(
		.INIT('h1)
	) name2115 (
		\u5_state_reg[25]/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w3074_
	);
	LUT2 #(
		.INIT('h4)
	) name2116 (
		\u5_state_reg[27]/NET0131 ,
		_w999_,
		_w3075_
	);
	LUT2 #(
		.INIT('h8)
	) name2117 (
		_w3058_,
		_w3075_,
		_w3076_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		_w1196_,
		_w3074_,
		_w3077_
	);
	LUT2 #(
		.INIT('h8)
	) name2119 (
		_w3073_,
		_w3077_,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name2120 (
		_w3055_,
		_w3078_,
		_w3079_
	);
	LUT2 #(
		.INIT('h8)
	) name2121 (
		_w3076_,
		_w3079_,
		_w3080_
	);
	LUT2 #(
		.INIT('h4)
	) name2122 (
		_w3070_,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h4)
	) name2123 (
		\u5_state_reg[20]/NET0131 ,
		_w3069_,
		_w3082_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		_w3081_,
		_w3082_,
		_w3083_
	);
	LUT2 #(
		.INIT('h4)
	) name2125 (
		\u5_state_reg[7]/NET0131 ,
		_w977_,
		_w3084_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		_w1016_,
		_w1332_,
		_w3085_
	);
	LUT2 #(
		.INIT('h8)
	) name2127 (
		_w3084_,
		_w3085_,
		_w3086_
	);
	LUT2 #(
		.INIT('h8)
	) name2128 (
		_w971_,
		_w1026_,
		_w3087_
	);
	LUT2 #(
		.INIT('h8)
	) name2129 (
		_w1342_,
		_w3087_,
		_w3088_
	);
	LUT2 #(
		.INIT('h8)
	) name2130 (
		_w3086_,
		_w3088_,
		_w3089_
	);
	LUT2 #(
		.INIT('h4)
	) name2131 (
		_w3083_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h8)
	) name2132 (
		_w1623_,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h1)
	) name2133 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3091_,
		_w3092_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		_w3093_
	);
	LUT2 #(
		.INIT('h8)
	) name2135 (
		\u5_state_reg[4]/NET0131 ,
		_w3093_,
		_w3094_
	);
	LUT2 #(
		.INIT('h2)
	) name2136 (
		\u5_state_reg[16]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		_w3095_
	);
	LUT2 #(
		.INIT('h8)
	) name2137 (
		_w1424_,
		_w3095_,
		_w3096_
	);
	LUT2 #(
		.INIT('h1)
	) name2138 (
		_w3094_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h2)
	) name2139 (
		_w1623_,
		_w3097_,
		_w3098_
	);
	LUT2 #(
		.INIT('h8)
	) name2140 (
		_w3049_,
		_w3098_,
		_w3099_
	);
	LUT2 #(
		.INIT('h2)
	) name2141 (
		\u2_u0_bank1_open_reg/NET0131 ,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h8)
	) name2142 (
		_w3092_,
		_w3100_,
		_w3101_
	);
	LUT2 #(
		.INIT('h1)
	) name2143 (
		_w3052_,
		_w3101_,
		_w3102_
	);
	LUT2 #(
		.INIT('h4)
	) name2144 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name2145 (
		_w3051_,
		_w3103_,
		_w3104_
	);
	LUT2 #(
		.INIT('h8)
	) name2146 (
		_w3098_,
		_w3103_,
		_w3105_
	);
	LUT2 #(
		.INIT('h2)
	) name2147 (
		\u2_u0_bank2_open_reg/NET0131 ,
		_w3105_,
		_w3106_
	);
	LUT2 #(
		.INIT('h8)
	) name2148 (
		_w3092_,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h1)
	) name2149 (
		_w3104_,
		_w3107_,
		_w3108_
	);
	LUT2 #(
		.INIT('h4)
	) name2150 (
		_w1676_,
		_w3050_,
		_w3109_
	);
	LUT2 #(
		.INIT('h8)
	) name2151 (
		_w3103_,
		_w3109_,
		_w3110_
	);
	LUT2 #(
		.INIT('h4)
	) name2152 (
		_w1676_,
		_w3090_,
		_w3111_
	);
	LUT2 #(
		.INIT('h1)
	) name2153 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3111_,
		_w3112_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		_w1676_,
		_w3097_,
		_w3113_
	);
	LUT2 #(
		.INIT('h8)
	) name2155 (
		_w3103_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h2)
	) name2156 (
		\u2_u1_bank2_open_reg/NET0131 ,
		_w3114_,
		_w3115_
	);
	LUT2 #(
		.INIT('h8)
	) name2157 (
		_w3112_,
		_w3115_,
		_w3116_
	);
	LUT2 #(
		.INIT('h1)
	) name2158 (
		_w3110_,
		_w3116_,
		_w3117_
	);
	LUT2 #(
		.INIT('h8)
	) name2159 (
		_w3049_,
		_w3109_,
		_w3118_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		_w3049_,
		_w3113_,
		_w3119_
	);
	LUT2 #(
		.INIT('h2)
	) name2161 (
		\u2_u1_bank1_open_reg/NET0131 ,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h8)
	) name2162 (
		_w3112_,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h1)
	) name2163 (
		_w3118_,
		_w3121_,
		_w3122_
	);
	LUT2 #(
		.INIT('h1)
	) name2164 (
		\u1_acs_addr_reg[16]/P0001 ,
		_w2866_,
		_w3123_
	);
	LUT2 #(
		.INIT('h1)
	) name2165 (
		_w2867_,
		_w3123_,
		_w3124_
	);
	LUT2 #(
		.INIT('h2)
	) name2166 (
		_w2858_,
		_w3124_,
		_w3125_
	);
	LUT2 #(
		.INIT('h8)
	) name2167 (
		\wb_addr_i[16]_pad ,
		_w2388_,
		_w3126_
	);
	LUT2 #(
		.INIT('h8)
	) name2168 (
		\wb_addr_i[18]_pad ,
		_w2878_,
		_w3127_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		\wb_addr_i[17]_pad ,
		_w2606_,
		_w3128_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w2858_,
		_w3126_,
		_w3129_
	);
	LUT2 #(
		.INIT('h1)
	) name2171 (
		_w3127_,
		_w3128_,
		_w3130_
	);
	LUT2 #(
		.INIT('h8)
	) name2172 (
		_w3129_,
		_w3130_,
		_w3131_
	);
	LUT2 #(
		.INIT('h1)
	) name2173 (
		_w3125_,
		_w3131_,
		_w3132_
	);
	LUT2 #(
		.INIT('h8)
	) name2174 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name2175 (
		_w3051_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h8)
	) name2176 (
		_w3098_,
		_w3133_,
		_w3135_
	);
	LUT2 #(
		.INIT('h2)
	) name2177 (
		\u2_u0_bank3_open_reg/NET0131 ,
		_w3135_,
		_w3136_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		_w3092_,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w3134_,
		_w3137_,
		_w3138_
	);
	LUT2 #(
		.INIT('h8)
	) name2180 (
		_w3109_,
		_w3133_,
		_w3139_
	);
	LUT2 #(
		.INIT('h8)
	) name2181 (
		_w3113_,
		_w3133_,
		_w3140_
	);
	LUT2 #(
		.INIT('h2)
	) name2182 (
		\u2_u1_bank3_open_reg/NET0131 ,
		_w3140_,
		_w3141_
	);
	LUT2 #(
		.INIT('h8)
	) name2183 (
		_w3112_,
		_w3141_,
		_w3142_
	);
	LUT2 #(
		.INIT('h1)
	) name2184 (
		_w3139_,
		_w3142_,
		_w3143_
	);
	LUT2 #(
		.INIT('h8)
	) name2185 (
		\wb_addr_i[18]_pad ,
		_w2388_,
		_w3144_
	);
	LUT2 #(
		.INIT('h8)
	) name2186 (
		\wb_addr_i[20]_pad ,
		_w2878_,
		_w3145_
	);
	LUT2 #(
		.INIT('h8)
	) name2187 (
		\wb_addr_i[19]_pad ,
		_w2606_,
		_w3146_
	);
	LUT2 #(
		.INIT('h1)
	) name2188 (
		_w3144_,
		_w3145_,
		_w3147_
	);
	LUT2 #(
		.INIT('h4)
	) name2189 (
		_w3146_,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h1)
	) name2190 (
		_w2858_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h1)
	) name2191 (
		\u1_acs_addr_reg[18]/P0001 ,
		_w2868_,
		_w3150_
	);
	LUT2 #(
		.INIT('h2)
	) name2192 (
		_w2858_,
		_w2869_,
		_w3151_
	);
	LUT2 #(
		.INIT('h4)
	) name2193 (
		_w3150_,
		_w3151_,
		_w3152_
	);
	LUT2 #(
		.INIT('h1)
	) name2194 (
		_w3149_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h4)
	) name2195 (
		_w1708_,
		_w2818_,
		_w3154_
	);
	LUT2 #(
		.INIT('h2)
	) name2196 (
		_w2555_,
		_w2821_,
		_w3155_
	);
	LUT2 #(
		.INIT('h8)
	) name2197 (
		\u5_state_reg[51]/NET0131 ,
		_w2533_,
		_w3156_
	);
	LUT2 #(
		.INIT('h1)
	) name2198 (
		\u5_timer2_reg[0]/P0001 ,
		_w2842_,
		_w3157_
	);
	LUT2 #(
		.INIT('h8)
	) name2199 (
		\u5_timer2_reg[0]/P0001 ,
		_w2842_,
		_w3158_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		_w2831_,
		_w2833_,
		_w3159_
	);
	LUT2 #(
		.INIT('h4)
	) name2201 (
		_w3157_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h4)
	) name2202 (
		_w3158_,
		_w3160_,
		_w3161_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		_w2822_,
		_w3161_,
		_w3162_
	);
	LUT2 #(
		.INIT('h4)
	) name2204 (
		_w3156_,
		_w3162_,
		_w3163_
	);
	LUT2 #(
		.INIT('h2)
	) name2205 (
		_w2821_,
		_w3163_,
		_w3164_
	);
	LUT2 #(
		.INIT('h2)
	) name2206 (
		_w2826_,
		_w3155_,
		_w3165_
	);
	LUT2 #(
		.INIT('h4)
	) name2207 (
		_w3164_,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('h1)
	) name2208 (
		_w3154_,
		_w3166_,
		_w3167_
	);
	LUT2 #(
		.INIT('h4)
	) name2209 (
		_w1794_,
		_w2818_,
		_w3168_
	);
	LUT2 #(
		.INIT('h2)
	) name2210 (
		_w2840_,
		_w2842_,
		_w3169_
	);
	LUT2 #(
		.INIT('h2)
	) name2211 (
		\u5_timer2_reg[6]/P0001 ,
		_w2839_,
		_w3170_
	);
	LUT2 #(
		.INIT('h2)
	) name2212 (
		_w2833_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h4)
	) name2213 (
		_w3169_,
		_w3171_,
		_w3172_
	);
	LUT2 #(
		.INIT('h8)
	) name2214 (
		_w2831_,
		_w3008_,
		_w3173_
	);
	LUT2 #(
		.INIT('h2)
	) name2215 (
		_w2584_,
		_w2833_,
		_w3174_
	);
	LUT2 #(
		.INIT('h1)
	) name2216 (
		_w3172_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h8)
	) name2217 (
		_w3173_,
		_w3175_,
		_w3176_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		_w3168_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('h4)
	) name2219 (
		\u4_rfr_req_reg/NET0131 ,
		_w1283_,
		_w3178_
	);
	LUT2 #(
		.INIT('h4)
	) name2220 (
		_w1057_,
		_w1679_,
		_w3179_
	);
	LUT2 #(
		.INIT('h2)
	) name2221 (
		\u5_wb_stb_first_reg/NET0131 ,
		_w3179_,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name2222 (
		_w1377_,
		_w1628_,
		_w3181_
	);
	LUT2 #(
		.INIT('h4)
	) name2223 (
		_w2424_,
		_w3181_,
		_w3182_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		_w1678_,
		_w3182_,
		_w3183_
	);
	LUT2 #(
		.INIT('h2)
	) name2225 (
		_w1683_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h4)
	) name2226 (
		_w3180_,
		_w3184_,
		_w3185_
	);
	LUT2 #(
		.INIT('h2)
	) name2227 (
		_w3178_,
		_w3185_,
		_w3186_
	);
	LUT2 #(
		.INIT('h8)
	) name2228 (
		\u5_wb_stb_first_reg/NET0131 ,
		_w1747_,
		_w3187_
	);
	LUT2 #(
		.INIT('h2)
	) name2229 (
		\u5_tmr_done_reg/NET0131 ,
		_w1629_,
		_w3188_
	);
	LUT2 #(
		.INIT('h8)
	) name2230 (
		_w1269_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h1)
	) name2231 (
		_w1108_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h4)
	) name2232 (
		_w2415_,
		_w3190_,
		_w3191_
	);
	LUT2 #(
		.INIT('h2)
	) name2233 (
		\u5_wb_cycle_reg/NET0131 ,
		_w3191_,
		_w3192_
	);
	LUT2 #(
		.INIT('h8)
	) name2234 (
		_w2430_,
		_w3181_,
		_w3193_
	);
	LUT2 #(
		.INIT('h1)
	) name2235 (
		_w1263_,
		_w1362_,
		_w3194_
	);
	LUT2 #(
		.INIT('h4)
	) name2236 (
		_w3187_,
		_w3194_,
		_w3195_
	);
	LUT2 #(
		.INIT('h1)
	) name2237 (
		_w1168_,
		_w1200_,
		_w3196_
	);
	LUT2 #(
		.INIT('h4)
	) name2238 (
		_w2629_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h4)
	) name2239 (
		_w3193_,
		_w3195_,
		_w3198_
	);
	LUT2 #(
		.INIT('h8)
	) name2240 (
		_w3197_,
		_w3198_,
		_w3199_
	);
	LUT2 #(
		.INIT('h4)
	) name2241 (
		_w3192_,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h4)
	) name2242 (
		_w3186_,
		_w3200_,
		_w3201_
	);
	LUT2 #(
		.INIT('h4)
	) name2243 (
		\u0_rf_we_reg/NET0131 ,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('h2)
	) name2244 (
		_w1046_,
		_w3202_,
		_w3203_
	);
	LUT2 #(
		.INIT('h2)
	) name2245 (
		\u0_sp_tms_reg[0]/NET0131 ,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h8)
	) name2246 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[0]/P0001 ,
		_w3205_
	);
	LUT2 #(
		.INIT('h4)
	) name2247 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		_w3206_
	);
	LUT2 #(
		.INIT('h8)
	) name2248 (
		\u0_u1_tms_reg[0]/P0001 ,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name2249 (
		_w3205_,
		_w3207_,
		_w3208_
	);
	LUT2 #(
		.INIT('h2)
	) name2250 (
		_w3203_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h1)
	) name2251 (
		_w3204_,
		_w3209_,
		_w3210_
	);
	LUT2 #(
		.INIT('h2)
	) name2252 (
		\u0_sp_tms_reg[10]/NET0131 ,
		_w3203_,
		_w3211_
	);
	LUT2 #(
		.INIT('h8)
	) name2253 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[10]/P0001 ,
		_w3212_
	);
	LUT2 #(
		.INIT('h8)
	) name2254 (
		\u0_u1_tms_reg[10]/P0001 ,
		_w3206_,
		_w3213_
	);
	LUT2 #(
		.INIT('h1)
	) name2255 (
		_w3212_,
		_w3213_,
		_w3214_
	);
	LUT2 #(
		.INIT('h2)
	) name2256 (
		_w3203_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('h1)
	) name2257 (
		_w3211_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h2)
	) name2258 (
		\u0_sp_tms_reg[11]/NET0131 ,
		_w3203_,
		_w3217_
	);
	LUT2 #(
		.INIT('h8)
	) name2259 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[11]/P0001 ,
		_w3218_
	);
	LUT2 #(
		.INIT('h8)
	) name2260 (
		\u0_u1_tms_reg[11]/P0001 ,
		_w3206_,
		_w3219_
	);
	LUT2 #(
		.INIT('h1)
	) name2261 (
		_w3218_,
		_w3219_,
		_w3220_
	);
	LUT2 #(
		.INIT('h2)
	) name2262 (
		_w3203_,
		_w3220_,
		_w3221_
	);
	LUT2 #(
		.INIT('h1)
	) name2263 (
		_w3217_,
		_w3221_,
		_w3222_
	);
	LUT2 #(
		.INIT('h2)
	) name2264 (
		\u0_sp_tms_reg[12]/NET0131 ,
		_w3203_,
		_w3223_
	);
	LUT2 #(
		.INIT('h8)
	) name2265 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[12]/P0001 ,
		_w3224_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		\u0_u1_tms_reg[12]/P0001 ,
		_w3206_,
		_w3225_
	);
	LUT2 #(
		.INIT('h1)
	) name2267 (
		_w3224_,
		_w3225_,
		_w3226_
	);
	LUT2 #(
		.INIT('h2)
	) name2268 (
		_w3203_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h1)
	) name2269 (
		_w3223_,
		_w3227_,
		_w3228_
	);
	LUT2 #(
		.INIT('h2)
	) name2270 (
		\u0_sp_tms_reg[14]/NET0131 ,
		_w3203_,
		_w3229_
	);
	LUT2 #(
		.INIT('h8)
	) name2271 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[14]/P0001 ,
		_w3230_
	);
	LUT2 #(
		.INIT('h8)
	) name2272 (
		\u0_u1_tms_reg[14]/P0001 ,
		_w3206_,
		_w3231_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w3230_,
		_w3231_,
		_w3232_
	);
	LUT2 #(
		.INIT('h2)
	) name2274 (
		_w3203_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h1)
	) name2275 (
		_w3229_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h2)
	) name2276 (
		\u0_sp_tms_reg[13]/NET0131 ,
		_w3203_,
		_w3235_
	);
	LUT2 #(
		.INIT('h8)
	) name2277 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[13]/P0001 ,
		_w3236_
	);
	LUT2 #(
		.INIT('h8)
	) name2278 (
		\u0_u1_tms_reg[13]/P0001 ,
		_w3206_,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name2279 (
		_w3236_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h2)
	) name2280 (
		_w3203_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('h1)
	) name2281 (
		_w3235_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h2)
	) name2282 (
		\u0_sp_tms_reg[16]/NET0131 ,
		_w3203_,
		_w3241_
	);
	LUT2 #(
		.INIT('h8)
	) name2283 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[16]/P0001 ,
		_w3242_
	);
	LUT2 #(
		.INIT('h8)
	) name2284 (
		\u0_u1_tms_reg[16]/P0001 ,
		_w3206_,
		_w3243_
	);
	LUT2 #(
		.INIT('h1)
	) name2285 (
		_w3242_,
		_w3243_,
		_w3244_
	);
	LUT2 #(
		.INIT('h2)
	) name2286 (
		_w3203_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('h1)
	) name2287 (
		_w3241_,
		_w3245_,
		_w3246_
	);
	LUT2 #(
		.INIT('h2)
	) name2288 (
		\u0_sp_tms_reg[17]/NET0131 ,
		_w3203_,
		_w3247_
	);
	LUT2 #(
		.INIT('h8)
	) name2289 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[17]/P0001 ,
		_w3248_
	);
	LUT2 #(
		.INIT('h8)
	) name2290 (
		\u0_u1_tms_reg[17]/P0001 ,
		_w3206_,
		_w3249_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w3248_,
		_w3249_,
		_w3250_
	);
	LUT2 #(
		.INIT('h2)
	) name2292 (
		_w3203_,
		_w3250_,
		_w3251_
	);
	LUT2 #(
		.INIT('h1)
	) name2293 (
		_w3247_,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('h2)
	) name2294 (
		\u0_sp_tms_reg[18]/NET0131 ,
		_w3203_,
		_w3253_
	);
	LUT2 #(
		.INIT('h8)
	) name2295 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[18]/P0001 ,
		_w3254_
	);
	LUT2 #(
		.INIT('h8)
	) name2296 (
		\u0_u1_tms_reg[18]/P0001 ,
		_w3206_,
		_w3255_
	);
	LUT2 #(
		.INIT('h1)
	) name2297 (
		_w3254_,
		_w3255_,
		_w3256_
	);
	LUT2 #(
		.INIT('h2)
	) name2298 (
		_w3203_,
		_w3256_,
		_w3257_
	);
	LUT2 #(
		.INIT('h1)
	) name2299 (
		_w3253_,
		_w3257_,
		_w3258_
	);
	LUT2 #(
		.INIT('h2)
	) name2300 (
		\u0_sp_tms_reg[19]/NET0131 ,
		_w3203_,
		_w3259_
	);
	LUT2 #(
		.INIT('h8)
	) name2301 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[19]/P0001 ,
		_w3260_
	);
	LUT2 #(
		.INIT('h8)
	) name2302 (
		\u0_u1_tms_reg[19]/P0001 ,
		_w3206_,
		_w3261_
	);
	LUT2 #(
		.INIT('h1)
	) name2303 (
		_w3260_,
		_w3261_,
		_w3262_
	);
	LUT2 #(
		.INIT('h2)
	) name2304 (
		_w3203_,
		_w3262_,
		_w3263_
	);
	LUT2 #(
		.INIT('h1)
	) name2305 (
		_w3259_,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h2)
	) name2306 (
		\u0_sp_tms_reg[15]/NET0131 ,
		_w3203_,
		_w3265_
	);
	LUT2 #(
		.INIT('h8)
	) name2307 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[15]/P0001 ,
		_w3266_
	);
	LUT2 #(
		.INIT('h8)
	) name2308 (
		\u0_u1_tms_reg[15]/P0001 ,
		_w3206_,
		_w3267_
	);
	LUT2 #(
		.INIT('h1)
	) name2309 (
		_w3266_,
		_w3267_,
		_w3268_
	);
	LUT2 #(
		.INIT('h2)
	) name2310 (
		_w3203_,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h1)
	) name2311 (
		_w3265_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h2)
	) name2312 (
		\u0_sp_tms_reg[1]/NET0131 ,
		_w3203_,
		_w3271_
	);
	LUT2 #(
		.INIT('h8)
	) name2313 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[1]/P0001 ,
		_w3272_
	);
	LUT2 #(
		.INIT('h8)
	) name2314 (
		\u0_u1_tms_reg[1]/P0001 ,
		_w3206_,
		_w3273_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w3272_,
		_w3273_,
		_w3274_
	);
	LUT2 #(
		.INIT('h2)
	) name2316 (
		_w3203_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		_w3271_,
		_w3275_,
		_w3276_
	);
	LUT2 #(
		.INIT('h2)
	) name2318 (
		\u0_sp_tms_reg[21]/NET0131 ,
		_w3203_,
		_w3277_
	);
	LUT2 #(
		.INIT('h8)
	) name2319 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[21]/P0001 ,
		_w3278_
	);
	LUT2 #(
		.INIT('h8)
	) name2320 (
		\u0_u1_tms_reg[21]/P0001 ,
		_w3206_,
		_w3279_
	);
	LUT2 #(
		.INIT('h1)
	) name2321 (
		_w3278_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h2)
	) name2322 (
		_w3203_,
		_w3280_,
		_w3281_
	);
	LUT2 #(
		.INIT('h1)
	) name2323 (
		_w3277_,
		_w3281_,
		_w3282_
	);
	LUT2 #(
		.INIT('h2)
	) name2324 (
		\u0_sp_tms_reg[20]/NET0131 ,
		_w3203_,
		_w3283_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[20]/P0001 ,
		_w3284_
	);
	LUT2 #(
		.INIT('h8)
	) name2326 (
		\u0_u1_tms_reg[20]/P0001 ,
		_w3206_,
		_w3285_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		_w3284_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h2)
	) name2328 (
		_w3203_,
		_w3286_,
		_w3287_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		_w3283_,
		_w3287_,
		_w3288_
	);
	LUT2 #(
		.INIT('h2)
	) name2330 (
		\u0_sp_tms_reg[22]/NET0131 ,
		_w3203_,
		_w3289_
	);
	LUT2 #(
		.INIT('h8)
	) name2331 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[22]/P0001 ,
		_w3290_
	);
	LUT2 #(
		.INIT('h8)
	) name2332 (
		\u0_u1_tms_reg[22]/P0001 ,
		_w3206_,
		_w3291_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		_w3290_,
		_w3291_,
		_w3292_
	);
	LUT2 #(
		.INIT('h2)
	) name2334 (
		_w3203_,
		_w3292_,
		_w3293_
	);
	LUT2 #(
		.INIT('h1)
	) name2335 (
		_w3289_,
		_w3293_,
		_w3294_
	);
	LUT2 #(
		.INIT('h2)
	) name2336 (
		\u0_sp_tms_reg[23]/NET0131 ,
		_w3203_,
		_w3295_
	);
	LUT2 #(
		.INIT('h8)
	) name2337 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[23]/P0001 ,
		_w3296_
	);
	LUT2 #(
		.INIT('h8)
	) name2338 (
		\u0_u1_tms_reg[23]/P0001 ,
		_w3206_,
		_w3297_
	);
	LUT2 #(
		.INIT('h1)
	) name2339 (
		_w3296_,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h2)
	) name2340 (
		_w3203_,
		_w3298_,
		_w3299_
	);
	LUT2 #(
		.INIT('h1)
	) name2341 (
		_w3295_,
		_w3299_,
		_w3300_
	);
	LUT2 #(
		.INIT('h2)
	) name2342 (
		\u0_sp_tms_reg[24]/NET0131 ,
		_w3203_,
		_w3301_
	);
	LUT2 #(
		.INIT('h8)
	) name2343 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[24]/P0001 ,
		_w3302_
	);
	LUT2 #(
		.INIT('h8)
	) name2344 (
		\u0_u1_tms_reg[24]/P0001 ,
		_w3206_,
		_w3303_
	);
	LUT2 #(
		.INIT('h1)
	) name2345 (
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h2)
	) name2346 (
		_w3203_,
		_w3304_,
		_w3305_
	);
	LUT2 #(
		.INIT('h1)
	) name2347 (
		_w3301_,
		_w3305_,
		_w3306_
	);
	LUT2 #(
		.INIT('h2)
	) name2348 (
		\u0_sp_tms_reg[25]/NET0131 ,
		_w3203_,
		_w3307_
	);
	LUT2 #(
		.INIT('h8)
	) name2349 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[25]/P0001 ,
		_w3308_
	);
	LUT2 #(
		.INIT('h8)
	) name2350 (
		\u0_u1_tms_reg[25]/P0001 ,
		_w3206_,
		_w3309_
	);
	LUT2 #(
		.INIT('h1)
	) name2351 (
		_w3308_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h2)
	) name2352 (
		_w3203_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h1)
	) name2353 (
		_w3307_,
		_w3311_,
		_w3312_
	);
	LUT2 #(
		.INIT('h2)
	) name2354 (
		\u0_sp_tms_reg[26]/NET0131 ,
		_w3203_,
		_w3313_
	);
	LUT2 #(
		.INIT('h8)
	) name2355 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[26]/P0001 ,
		_w3314_
	);
	LUT2 #(
		.INIT('h8)
	) name2356 (
		\u0_u1_tms_reg[26]/P0001 ,
		_w3206_,
		_w3315_
	);
	LUT2 #(
		.INIT('h1)
	) name2357 (
		_w3314_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h2)
	) name2358 (
		_w3203_,
		_w3316_,
		_w3317_
	);
	LUT2 #(
		.INIT('h1)
	) name2359 (
		_w3313_,
		_w3317_,
		_w3318_
	);
	LUT2 #(
		.INIT('h2)
	) name2360 (
		\u0_sp_tms_reg[27]/NET0131 ,
		_w3203_,
		_w3319_
	);
	LUT2 #(
		.INIT('h8)
	) name2361 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[27]/P0001 ,
		_w3320_
	);
	LUT2 #(
		.INIT('h8)
	) name2362 (
		\u0_u1_tms_reg[27]/P0001 ,
		_w3206_,
		_w3321_
	);
	LUT2 #(
		.INIT('h1)
	) name2363 (
		_w3320_,
		_w3321_,
		_w3322_
	);
	LUT2 #(
		.INIT('h2)
	) name2364 (
		_w3203_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		_w3319_,
		_w3323_,
		_w3324_
	);
	LUT2 #(
		.INIT('h2)
	) name2366 (
		\u0_sp_tms_reg[2]/NET0131 ,
		_w3203_,
		_w3325_
	);
	LUT2 #(
		.INIT('h8)
	) name2367 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[2]/P0001 ,
		_w3326_
	);
	LUT2 #(
		.INIT('h8)
	) name2368 (
		\u0_u1_tms_reg[2]/P0001 ,
		_w3206_,
		_w3327_
	);
	LUT2 #(
		.INIT('h1)
	) name2369 (
		_w3326_,
		_w3327_,
		_w3328_
	);
	LUT2 #(
		.INIT('h2)
	) name2370 (
		_w3203_,
		_w3328_,
		_w3329_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w3325_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h2)
	) name2372 (
		\u0_sp_tms_reg[3]/NET0131 ,
		_w3203_,
		_w3331_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[3]/P0001 ,
		_w3332_
	);
	LUT2 #(
		.INIT('h8)
	) name2374 (
		\u0_u1_tms_reg[3]/P0001 ,
		_w3206_,
		_w3333_
	);
	LUT2 #(
		.INIT('h1)
	) name2375 (
		_w3332_,
		_w3333_,
		_w3334_
	);
	LUT2 #(
		.INIT('h2)
	) name2376 (
		_w3203_,
		_w3334_,
		_w3335_
	);
	LUT2 #(
		.INIT('h1)
	) name2377 (
		_w3331_,
		_w3335_,
		_w3336_
	);
	LUT2 #(
		.INIT('h2)
	) name2378 (
		\u0_sp_tms_reg[4]/NET0131 ,
		_w3203_,
		_w3337_
	);
	LUT2 #(
		.INIT('h8)
	) name2379 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[4]/P0001 ,
		_w3338_
	);
	LUT2 #(
		.INIT('h8)
	) name2380 (
		\u0_u1_tms_reg[4]/P0001 ,
		_w3206_,
		_w3339_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		_w3338_,
		_w3339_,
		_w3340_
	);
	LUT2 #(
		.INIT('h2)
	) name2382 (
		_w3203_,
		_w3340_,
		_w3341_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w3337_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h2)
	) name2384 (
		\u0_sp_tms_reg[5]/NET0131 ,
		_w3203_,
		_w3343_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[5]/P0001 ,
		_w3344_
	);
	LUT2 #(
		.INIT('h8)
	) name2386 (
		\u0_u1_tms_reg[5]/P0001 ,
		_w3206_,
		_w3345_
	);
	LUT2 #(
		.INIT('h1)
	) name2387 (
		_w3344_,
		_w3345_,
		_w3346_
	);
	LUT2 #(
		.INIT('h2)
	) name2388 (
		_w3203_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h1)
	) name2389 (
		_w3343_,
		_w3347_,
		_w3348_
	);
	LUT2 #(
		.INIT('h2)
	) name2390 (
		\u0_sp_tms_reg[7]/NET0131 ,
		_w3203_,
		_w3349_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[7]/P0001 ,
		_w3350_
	);
	LUT2 #(
		.INIT('h8)
	) name2392 (
		\u0_u1_tms_reg[7]/P0001 ,
		_w3206_,
		_w3351_
	);
	LUT2 #(
		.INIT('h1)
	) name2393 (
		_w3350_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h2)
	) name2394 (
		_w3203_,
		_w3352_,
		_w3353_
	);
	LUT2 #(
		.INIT('h1)
	) name2395 (
		_w3349_,
		_w3353_,
		_w3354_
	);
	LUT2 #(
		.INIT('h2)
	) name2396 (
		\u0_sp_tms_reg[6]/NET0131 ,
		_w3203_,
		_w3355_
	);
	LUT2 #(
		.INIT('h8)
	) name2397 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[6]/P0001 ,
		_w3356_
	);
	LUT2 #(
		.INIT('h8)
	) name2398 (
		\u0_u1_tms_reg[6]/P0001 ,
		_w3206_,
		_w3357_
	);
	LUT2 #(
		.INIT('h1)
	) name2399 (
		_w3356_,
		_w3357_,
		_w3358_
	);
	LUT2 #(
		.INIT('h2)
	) name2400 (
		_w3203_,
		_w3358_,
		_w3359_
	);
	LUT2 #(
		.INIT('h1)
	) name2401 (
		_w3355_,
		_w3359_,
		_w3360_
	);
	LUT2 #(
		.INIT('h2)
	) name2402 (
		\u0_sp_tms_reg[8]/NET0131 ,
		_w3203_,
		_w3361_
	);
	LUT2 #(
		.INIT('h8)
	) name2403 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[8]/P0001 ,
		_w3362_
	);
	LUT2 #(
		.INIT('h8)
	) name2404 (
		\u0_u1_tms_reg[8]/P0001 ,
		_w3206_,
		_w3363_
	);
	LUT2 #(
		.INIT('h1)
	) name2405 (
		_w3362_,
		_w3363_,
		_w3364_
	);
	LUT2 #(
		.INIT('h2)
	) name2406 (
		_w3203_,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h1)
	) name2407 (
		_w3361_,
		_w3365_,
		_w3366_
	);
	LUT2 #(
		.INIT('h2)
	) name2408 (
		\u0_sp_tms_reg[9]/NET0131 ,
		_w3203_,
		_w3367_
	);
	LUT2 #(
		.INIT('h8)
	) name2409 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_tms_reg[9]/P0001 ,
		_w3368_
	);
	LUT2 #(
		.INIT('h8)
	) name2410 (
		\u0_u1_tms_reg[9]/P0001 ,
		_w3206_,
		_w3369_
	);
	LUT2 #(
		.INIT('h1)
	) name2411 (
		_w3368_,
		_w3369_,
		_w3370_
	);
	LUT2 #(
		.INIT('h2)
	) name2412 (
		_w3203_,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h1)
	) name2413 (
		_w3367_,
		_w3371_,
		_w3372_
	);
	LUT2 #(
		.INIT('h2)
	) name2414 (
		\u0_tms_reg[10]/NET0131 ,
		_w3203_,
		_w3373_
	);
	LUT2 #(
		.INIT('h8)
	) name2415 (
		\u0_u0_csc_reg[8]/P0001 ,
		wb_we_i_pad,
		_w3374_
	);
	LUT2 #(
		.INIT('h1)
	) name2416 (
		\u0_u0_csc_reg[18]/P0001 ,
		\wb_addr_i[23]_pad ,
		_w3375_
	);
	LUT2 #(
		.INIT('h8)
	) name2417 (
		\u0_u0_csc_reg[18]/P0001 ,
		\wb_addr_i[23]_pad ,
		_w3376_
	);
	LUT2 #(
		.INIT('h2)
	) name2418 (
		\u0_csc_mask_r_reg[2]/NET0131 ,
		_w3375_,
		_w3377_
	);
	LUT2 #(
		.INIT('h4)
	) name2419 (
		_w3376_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h2)
	) name2420 (
		\u0_u0_csc_reg[20]/P0001 ,
		\wb_addr_i[25]_pad ,
		_w3379_
	);
	LUT2 #(
		.INIT('h4)
	) name2421 (
		\u0_u0_csc_reg[20]/P0001 ,
		\wb_addr_i[25]_pad ,
		_w3380_
	);
	LUT2 #(
		.INIT('h1)
	) name2422 (
		_w3379_,
		_w3380_,
		_w3381_
	);
	LUT2 #(
		.INIT('h2)
	) name2423 (
		\u0_csc_mask_r_reg[4]/NET0131 ,
		_w3381_,
		_w3382_
	);
	LUT2 #(
		.INIT('h1)
	) name2424 (
		\u0_u0_csc_reg[22]/P0001 ,
		\wb_addr_i[27]_pad ,
		_w3383_
	);
	LUT2 #(
		.INIT('h8)
	) name2425 (
		\u0_u0_csc_reg[22]/P0001 ,
		\wb_addr_i[27]_pad ,
		_w3384_
	);
	LUT2 #(
		.INIT('h2)
	) name2426 (
		\u0_csc_mask_r_reg[6]/NET0131 ,
		_w3383_,
		_w3385_
	);
	LUT2 #(
		.INIT('h4)
	) name2427 (
		_w3384_,
		_w3385_,
		_w3386_
	);
	LUT2 #(
		.INIT('h1)
	) name2428 (
		\u0_u0_csc_reg[23]/P0001 ,
		\wb_addr_i[28]_pad ,
		_w3387_
	);
	LUT2 #(
		.INIT('h8)
	) name2429 (
		\u0_u0_csc_reg[23]/P0001 ,
		\wb_addr_i[28]_pad ,
		_w3388_
	);
	LUT2 #(
		.INIT('h2)
	) name2430 (
		\u0_csc_mask_r_reg[7]/NET0131 ,
		_w3387_,
		_w3389_
	);
	LUT2 #(
		.INIT('h4)
	) name2431 (
		_w3388_,
		_w3389_,
		_w3390_
	);
	LUT2 #(
		.INIT('h1)
	) name2432 (
		\u0_u0_csc_reg[17]/P0001 ,
		\wb_addr_i[22]_pad ,
		_w3391_
	);
	LUT2 #(
		.INIT('h8)
	) name2433 (
		\u0_u0_csc_reg[17]/P0001 ,
		\wb_addr_i[22]_pad ,
		_w3392_
	);
	LUT2 #(
		.INIT('h2)
	) name2434 (
		\u0_csc_mask_r_reg[1]/NET0131 ,
		_w3391_,
		_w3393_
	);
	LUT2 #(
		.INIT('h4)
	) name2435 (
		_w3392_,
		_w3393_,
		_w3394_
	);
	LUT2 #(
		.INIT('h1)
	) name2436 (
		\u0_u0_csc_reg[16]/P0001 ,
		\wb_addr_i[21]_pad ,
		_w3395_
	);
	LUT2 #(
		.INIT('h8)
	) name2437 (
		\u0_u0_csc_reg[16]/P0001 ,
		\wb_addr_i[21]_pad ,
		_w3396_
	);
	LUT2 #(
		.INIT('h2)
	) name2438 (
		\u0_csc_mask_r_reg[0]/NET0131 ,
		_w3395_,
		_w3397_
	);
	LUT2 #(
		.INIT('h4)
	) name2439 (
		_w3396_,
		_w3397_,
		_w3398_
	);
	LUT2 #(
		.INIT('h1)
	) name2440 (
		\u0_u0_csc_reg[19]/P0001 ,
		\wb_addr_i[24]_pad ,
		_w3399_
	);
	LUT2 #(
		.INIT('h8)
	) name2441 (
		\u0_u0_csc_reg[19]/P0001 ,
		\wb_addr_i[24]_pad ,
		_w3400_
	);
	LUT2 #(
		.INIT('h2)
	) name2442 (
		\u0_csc_mask_r_reg[3]/NET0131 ,
		_w3399_,
		_w3401_
	);
	LUT2 #(
		.INIT('h4)
	) name2443 (
		_w3400_,
		_w3401_,
		_w3402_
	);
	LUT2 #(
		.INIT('h1)
	) name2444 (
		\u0_u0_csc_reg[21]/P0001 ,
		\wb_addr_i[26]_pad ,
		_w3403_
	);
	LUT2 #(
		.INIT('h8)
	) name2445 (
		\u0_u0_csc_reg[21]/P0001 ,
		\wb_addr_i[26]_pad ,
		_w3404_
	);
	LUT2 #(
		.INIT('h2)
	) name2446 (
		\u0_csc_mask_r_reg[5]/NET0131 ,
		_w3403_,
		_w3405_
	);
	LUT2 #(
		.INIT('h4)
	) name2447 (
		_w3404_,
		_w3405_,
		_w3406_
	);
	LUT2 #(
		.INIT('h2)
	) name2448 (
		\u0_u0_csc_reg[0]/NET0131 ,
		_w3378_,
		_w3407_
	);
	LUT2 #(
		.INIT('h1)
	) name2449 (
		_w3382_,
		_w3386_,
		_w3408_
	);
	LUT2 #(
		.INIT('h1)
	) name2450 (
		_w3390_,
		_w3394_,
		_w3409_
	);
	LUT2 #(
		.INIT('h1)
	) name2451 (
		_w3398_,
		_w3402_,
		_w3410_
	);
	LUT2 #(
		.INIT('h4)
	) name2452 (
		_w3406_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h8)
	) name2453 (
		_w3408_,
		_w3409_,
		_w3412_
	);
	LUT2 #(
		.INIT('h8)
	) name2454 (
		_w3407_,
		_w3412_,
		_w3413_
	);
	LUT2 #(
		.INIT('h8)
	) name2455 (
		_w3411_,
		_w3413_,
		_w3414_
	);
	LUT2 #(
		.INIT('h4)
	) name2456 (
		_w3374_,
		_w3414_,
		_w3415_
	);
	LUT2 #(
		.INIT('h8)
	) name2457 (
		\u0_u1_csc_reg[8]/P0001 ,
		wb_we_i_pad,
		_w3416_
	);
	LUT2 #(
		.INIT('h1)
	) name2458 (
		\u0_u1_csc_reg[17]/P0001 ,
		\wb_addr_i[22]_pad ,
		_w3417_
	);
	LUT2 #(
		.INIT('h8)
	) name2459 (
		\u0_u1_csc_reg[17]/P0001 ,
		\wb_addr_i[22]_pad ,
		_w3418_
	);
	LUT2 #(
		.INIT('h2)
	) name2460 (
		\u0_csc_mask_r_reg[1]/NET0131 ,
		_w3417_,
		_w3419_
	);
	LUT2 #(
		.INIT('h4)
	) name2461 (
		_w3418_,
		_w3419_,
		_w3420_
	);
	LUT2 #(
		.INIT('h2)
	) name2462 (
		\u0_u1_csc_reg[21]/P0001 ,
		\wb_addr_i[26]_pad ,
		_w3421_
	);
	LUT2 #(
		.INIT('h4)
	) name2463 (
		\u0_u1_csc_reg[21]/P0001 ,
		\wb_addr_i[26]_pad ,
		_w3422_
	);
	LUT2 #(
		.INIT('h1)
	) name2464 (
		_w3421_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h2)
	) name2465 (
		\u0_csc_mask_r_reg[5]/NET0131 ,
		_w3423_,
		_w3424_
	);
	LUT2 #(
		.INIT('h1)
	) name2466 (
		\u0_u1_csc_reg[22]/P0001 ,
		\wb_addr_i[27]_pad ,
		_w3425_
	);
	LUT2 #(
		.INIT('h8)
	) name2467 (
		\u0_u1_csc_reg[22]/P0001 ,
		\wb_addr_i[27]_pad ,
		_w3426_
	);
	LUT2 #(
		.INIT('h2)
	) name2468 (
		\u0_csc_mask_r_reg[6]/NET0131 ,
		_w3425_,
		_w3427_
	);
	LUT2 #(
		.INIT('h4)
	) name2469 (
		_w3426_,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h1)
	) name2470 (
		\u0_u1_csc_reg[19]/P0001 ,
		\wb_addr_i[24]_pad ,
		_w3429_
	);
	LUT2 #(
		.INIT('h8)
	) name2471 (
		\u0_u1_csc_reg[19]/P0001 ,
		\wb_addr_i[24]_pad ,
		_w3430_
	);
	LUT2 #(
		.INIT('h2)
	) name2472 (
		\u0_csc_mask_r_reg[3]/NET0131 ,
		_w3429_,
		_w3431_
	);
	LUT2 #(
		.INIT('h4)
	) name2473 (
		_w3430_,
		_w3431_,
		_w3432_
	);
	LUT2 #(
		.INIT('h1)
	) name2474 (
		\u0_u1_csc_reg[16]/P0001 ,
		\wb_addr_i[21]_pad ,
		_w3433_
	);
	LUT2 #(
		.INIT('h8)
	) name2475 (
		\u0_u1_csc_reg[16]/P0001 ,
		\wb_addr_i[21]_pad ,
		_w3434_
	);
	LUT2 #(
		.INIT('h2)
	) name2476 (
		\u0_csc_mask_r_reg[0]/NET0131 ,
		_w3433_,
		_w3435_
	);
	LUT2 #(
		.INIT('h4)
	) name2477 (
		_w3434_,
		_w3435_,
		_w3436_
	);
	LUT2 #(
		.INIT('h1)
	) name2478 (
		\u0_u1_csc_reg[18]/P0001 ,
		\wb_addr_i[23]_pad ,
		_w3437_
	);
	LUT2 #(
		.INIT('h8)
	) name2479 (
		\u0_u1_csc_reg[18]/P0001 ,
		\wb_addr_i[23]_pad ,
		_w3438_
	);
	LUT2 #(
		.INIT('h2)
	) name2480 (
		\u0_csc_mask_r_reg[2]/NET0131 ,
		_w3437_,
		_w3439_
	);
	LUT2 #(
		.INIT('h4)
	) name2481 (
		_w3438_,
		_w3439_,
		_w3440_
	);
	LUT2 #(
		.INIT('h1)
	) name2482 (
		\u0_u1_csc_reg[23]/P0001 ,
		\wb_addr_i[28]_pad ,
		_w3441_
	);
	LUT2 #(
		.INIT('h8)
	) name2483 (
		\u0_u1_csc_reg[23]/P0001 ,
		\wb_addr_i[28]_pad ,
		_w3442_
	);
	LUT2 #(
		.INIT('h2)
	) name2484 (
		\u0_csc_mask_r_reg[7]/NET0131 ,
		_w3441_,
		_w3443_
	);
	LUT2 #(
		.INIT('h4)
	) name2485 (
		_w3442_,
		_w3443_,
		_w3444_
	);
	LUT2 #(
		.INIT('h1)
	) name2486 (
		\u0_u1_csc_reg[20]/P0001 ,
		\wb_addr_i[25]_pad ,
		_w3445_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		\u0_u1_csc_reg[20]/P0001 ,
		\wb_addr_i[25]_pad ,
		_w3446_
	);
	LUT2 #(
		.INIT('h2)
	) name2488 (
		\u0_csc_mask_r_reg[4]/NET0131 ,
		_w3445_,
		_w3447_
	);
	LUT2 #(
		.INIT('h4)
	) name2489 (
		_w3446_,
		_w3447_,
		_w3448_
	);
	LUT2 #(
		.INIT('h2)
	) name2490 (
		\u0_u1_csc_reg[0]/NET0131 ,
		_w3420_,
		_w3449_
	);
	LUT2 #(
		.INIT('h1)
	) name2491 (
		_w3424_,
		_w3428_,
		_w3450_
	);
	LUT2 #(
		.INIT('h1)
	) name2492 (
		_w3432_,
		_w3436_,
		_w3451_
	);
	LUT2 #(
		.INIT('h1)
	) name2493 (
		_w3440_,
		_w3444_,
		_w3452_
	);
	LUT2 #(
		.INIT('h4)
	) name2494 (
		_w3448_,
		_w3452_,
		_w3453_
	);
	LUT2 #(
		.INIT('h8)
	) name2495 (
		_w3450_,
		_w3451_,
		_w3454_
	);
	LUT2 #(
		.INIT('h8)
	) name2496 (
		_w3449_,
		_w3454_,
		_w3455_
	);
	LUT2 #(
		.INIT('h8)
	) name2497 (
		_w3453_,
		_w3455_,
		_w3456_
	);
	LUT2 #(
		.INIT('h4)
	) name2498 (
		_w3416_,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('h4)
	) name2499 (
		_w3415_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h8)
	) name2500 (
		\u0_u1_tms_reg[10]/P0001 ,
		_w3458_,
		_w3459_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		\u0_u0_tms_reg[10]/P0001 ,
		_w3415_,
		_w3460_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		_w3459_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h2)
	) name2503 (
		_w3203_,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h1)
	) name2504 (
		_w3373_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h2)
	) name2505 (
		\u0_tms_reg[11]/NET0131 ,
		_w3203_,
		_w3464_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		\u0_u1_tms_reg[11]/P0001 ,
		_w3458_,
		_w3465_
	);
	LUT2 #(
		.INIT('h8)
	) name2507 (
		\u0_u0_tms_reg[11]/P0001 ,
		_w3415_,
		_w3466_
	);
	LUT2 #(
		.INIT('h1)
	) name2508 (
		_w3465_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h2)
	) name2509 (
		_w3203_,
		_w3467_,
		_w3468_
	);
	LUT2 #(
		.INIT('h1)
	) name2510 (
		_w3464_,
		_w3468_,
		_w3469_
	);
	LUT2 #(
		.INIT('h2)
	) name2511 (
		\u0_tms_reg[12]/NET0131 ,
		_w3203_,
		_w3470_
	);
	LUT2 #(
		.INIT('h8)
	) name2512 (
		\u0_u1_tms_reg[12]/P0001 ,
		_w3458_,
		_w3471_
	);
	LUT2 #(
		.INIT('h8)
	) name2513 (
		\u0_u0_tms_reg[12]/P0001 ,
		_w3415_,
		_w3472_
	);
	LUT2 #(
		.INIT('h1)
	) name2514 (
		_w3471_,
		_w3472_,
		_w3473_
	);
	LUT2 #(
		.INIT('h2)
	) name2515 (
		_w3203_,
		_w3473_,
		_w3474_
	);
	LUT2 #(
		.INIT('h1)
	) name2516 (
		_w3470_,
		_w3474_,
		_w3475_
	);
	LUT2 #(
		.INIT('h2)
	) name2517 (
		\u0_tms_reg[13]/NET0131 ,
		_w3203_,
		_w3476_
	);
	LUT2 #(
		.INIT('h8)
	) name2518 (
		\u0_u1_tms_reg[13]/P0001 ,
		_w3458_,
		_w3477_
	);
	LUT2 #(
		.INIT('h8)
	) name2519 (
		\u0_u0_tms_reg[13]/P0001 ,
		_w3415_,
		_w3478_
	);
	LUT2 #(
		.INIT('h1)
	) name2520 (
		_w3477_,
		_w3478_,
		_w3479_
	);
	LUT2 #(
		.INIT('h2)
	) name2521 (
		_w3203_,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h1)
	) name2522 (
		_w3476_,
		_w3480_,
		_w3481_
	);
	LUT2 #(
		.INIT('h2)
	) name2523 (
		\u0_tms_reg[0]/NET0131 ,
		_w3203_,
		_w3482_
	);
	LUT2 #(
		.INIT('h8)
	) name2524 (
		\u0_u1_tms_reg[0]/P0001 ,
		_w3458_,
		_w3483_
	);
	LUT2 #(
		.INIT('h8)
	) name2525 (
		\u0_u0_tms_reg[0]/P0001 ,
		_w3415_,
		_w3484_
	);
	LUT2 #(
		.INIT('h1)
	) name2526 (
		_w3483_,
		_w3484_,
		_w3485_
	);
	LUT2 #(
		.INIT('h2)
	) name2527 (
		_w3203_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h1)
	) name2528 (
		_w3482_,
		_w3486_,
		_w3487_
	);
	LUT2 #(
		.INIT('h2)
	) name2529 (
		\u0_tms_reg[14]/NET0131 ,
		_w3203_,
		_w3488_
	);
	LUT2 #(
		.INIT('h8)
	) name2530 (
		\u0_u1_tms_reg[14]/P0001 ,
		_w3458_,
		_w3489_
	);
	LUT2 #(
		.INIT('h8)
	) name2531 (
		\u0_u0_tms_reg[14]/P0001 ,
		_w3415_,
		_w3490_
	);
	LUT2 #(
		.INIT('h1)
	) name2532 (
		_w3489_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h2)
	) name2533 (
		_w3203_,
		_w3491_,
		_w3492_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w3488_,
		_w3492_,
		_w3493_
	);
	LUT2 #(
		.INIT('h2)
	) name2535 (
		\u0_tms_reg[15]/NET0131 ,
		_w3203_,
		_w3494_
	);
	LUT2 #(
		.INIT('h8)
	) name2536 (
		\u0_u1_tms_reg[15]/P0001 ,
		_w3458_,
		_w3495_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		\u0_u0_tms_reg[15]/P0001 ,
		_w3415_,
		_w3496_
	);
	LUT2 #(
		.INIT('h1)
	) name2538 (
		_w3495_,
		_w3496_,
		_w3497_
	);
	LUT2 #(
		.INIT('h2)
	) name2539 (
		_w3203_,
		_w3497_,
		_w3498_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		_w3494_,
		_w3498_,
		_w3499_
	);
	LUT2 #(
		.INIT('h2)
	) name2541 (
		\u0_tms_reg[16]/NET0131 ,
		_w3203_,
		_w3500_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		\u0_u1_tms_reg[16]/P0001 ,
		_w3458_,
		_w3501_
	);
	LUT2 #(
		.INIT('h8)
	) name2543 (
		\u0_u0_tms_reg[16]/P0001 ,
		_w3415_,
		_w3502_
	);
	LUT2 #(
		.INIT('h1)
	) name2544 (
		_w3501_,
		_w3502_,
		_w3503_
	);
	LUT2 #(
		.INIT('h2)
	) name2545 (
		_w3203_,
		_w3503_,
		_w3504_
	);
	LUT2 #(
		.INIT('h1)
	) name2546 (
		_w3500_,
		_w3504_,
		_w3505_
	);
	LUT2 #(
		.INIT('h2)
	) name2547 (
		\u0_tms_reg[17]/NET0131 ,
		_w3203_,
		_w3506_
	);
	LUT2 #(
		.INIT('h8)
	) name2548 (
		\u0_u1_tms_reg[17]/P0001 ,
		_w3458_,
		_w3507_
	);
	LUT2 #(
		.INIT('h8)
	) name2549 (
		\u0_u0_tms_reg[17]/P0001 ,
		_w3415_,
		_w3508_
	);
	LUT2 #(
		.INIT('h1)
	) name2550 (
		_w3507_,
		_w3508_,
		_w3509_
	);
	LUT2 #(
		.INIT('h2)
	) name2551 (
		_w3203_,
		_w3509_,
		_w3510_
	);
	LUT2 #(
		.INIT('h1)
	) name2552 (
		_w3506_,
		_w3510_,
		_w3511_
	);
	LUT2 #(
		.INIT('h2)
	) name2553 (
		\u0_tms_reg[18]/NET0131 ,
		_w3203_,
		_w3512_
	);
	LUT2 #(
		.INIT('h8)
	) name2554 (
		\u0_u1_tms_reg[18]/P0001 ,
		_w3458_,
		_w3513_
	);
	LUT2 #(
		.INIT('h8)
	) name2555 (
		\u0_u0_tms_reg[18]/P0001 ,
		_w3415_,
		_w3514_
	);
	LUT2 #(
		.INIT('h1)
	) name2556 (
		_w3513_,
		_w3514_,
		_w3515_
	);
	LUT2 #(
		.INIT('h2)
	) name2557 (
		_w3203_,
		_w3515_,
		_w3516_
	);
	LUT2 #(
		.INIT('h1)
	) name2558 (
		_w3512_,
		_w3516_,
		_w3517_
	);
	LUT2 #(
		.INIT('h2)
	) name2559 (
		\u0_tms_reg[19]/NET0131 ,
		_w3203_,
		_w3518_
	);
	LUT2 #(
		.INIT('h8)
	) name2560 (
		\u0_u1_tms_reg[19]/P0001 ,
		_w3458_,
		_w3519_
	);
	LUT2 #(
		.INIT('h8)
	) name2561 (
		\u0_u0_tms_reg[19]/P0001 ,
		_w3415_,
		_w3520_
	);
	LUT2 #(
		.INIT('h1)
	) name2562 (
		_w3519_,
		_w3520_,
		_w3521_
	);
	LUT2 #(
		.INIT('h2)
	) name2563 (
		_w3203_,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h1)
	) name2564 (
		_w3518_,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h2)
	) name2565 (
		\u0_tms_reg[1]/NET0131 ,
		_w3203_,
		_w3524_
	);
	LUT2 #(
		.INIT('h8)
	) name2566 (
		\u0_u1_tms_reg[1]/P0001 ,
		_w3458_,
		_w3525_
	);
	LUT2 #(
		.INIT('h8)
	) name2567 (
		\u0_u0_tms_reg[1]/P0001 ,
		_w3415_,
		_w3526_
	);
	LUT2 #(
		.INIT('h1)
	) name2568 (
		_w3525_,
		_w3526_,
		_w3527_
	);
	LUT2 #(
		.INIT('h2)
	) name2569 (
		_w3203_,
		_w3527_,
		_w3528_
	);
	LUT2 #(
		.INIT('h1)
	) name2570 (
		_w3524_,
		_w3528_,
		_w3529_
	);
	LUT2 #(
		.INIT('h2)
	) name2571 (
		\u0_tms_reg[20]/NET0131 ,
		_w3203_,
		_w3530_
	);
	LUT2 #(
		.INIT('h8)
	) name2572 (
		\u0_u1_tms_reg[20]/P0001 ,
		_w3458_,
		_w3531_
	);
	LUT2 #(
		.INIT('h8)
	) name2573 (
		\u0_u0_tms_reg[20]/P0001 ,
		_w3415_,
		_w3532_
	);
	LUT2 #(
		.INIT('h1)
	) name2574 (
		_w3531_,
		_w3532_,
		_w3533_
	);
	LUT2 #(
		.INIT('h2)
	) name2575 (
		_w3203_,
		_w3533_,
		_w3534_
	);
	LUT2 #(
		.INIT('h1)
	) name2576 (
		_w3530_,
		_w3534_,
		_w3535_
	);
	LUT2 #(
		.INIT('h2)
	) name2577 (
		\u0_tms_reg[21]/NET0131 ,
		_w3203_,
		_w3536_
	);
	LUT2 #(
		.INIT('h8)
	) name2578 (
		\u0_u1_tms_reg[21]/P0001 ,
		_w3458_,
		_w3537_
	);
	LUT2 #(
		.INIT('h8)
	) name2579 (
		\u0_u0_tms_reg[21]/P0001 ,
		_w3415_,
		_w3538_
	);
	LUT2 #(
		.INIT('h1)
	) name2580 (
		_w3537_,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h2)
	) name2581 (
		_w3203_,
		_w3539_,
		_w3540_
	);
	LUT2 #(
		.INIT('h1)
	) name2582 (
		_w3536_,
		_w3540_,
		_w3541_
	);
	LUT2 #(
		.INIT('h2)
	) name2583 (
		\u0_tms_reg[23]/NET0131 ,
		_w3203_,
		_w3542_
	);
	LUT2 #(
		.INIT('h8)
	) name2584 (
		\u0_u1_tms_reg[23]/P0001 ,
		_w3458_,
		_w3543_
	);
	LUT2 #(
		.INIT('h8)
	) name2585 (
		\u0_u0_tms_reg[23]/P0001 ,
		_w3415_,
		_w3544_
	);
	LUT2 #(
		.INIT('h1)
	) name2586 (
		_w3543_,
		_w3544_,
		_w3545_
	);
	LUT2 #(
		.INIT('h2)
	) name2587 (
		_w3203_,
		_w3545_,
		_w3546_
	);
	LUT2 #(
		.INIT('h1)
	) name2588 (
		_w3542_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h2)
	) name2589 (
		\u0_tms_reg[24]/NET0131 ,
		_w3203_,
		_w3548_
	);
	LUT2 #(
		.INIT('h8)
	) name2590 (
		\u0_u1_tms_reg[24]/P0001 ,
		_w3458_,
		_w3549_
	);
	LUT2 #(
		.INIT('h8)
	) name2591 (
		\u0_u0_tms_reg[24]/P0001 ,
		_w3415_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name2592 (
		_w3549_,
		_w3550_,
		_w3551_
	);
	LUT2 #(
		.INIT('h2)
	) name2593 (
		_w3203_,
		_w3551_,
		_w3552_
	);
	LUT2 #(
		.INIT('h1)
	) name2594 (
		_w3548_,
		_w3552_,
		_w3553_
	);
	LUT2 #(
		.INIT('h2)
	) name2595 (
		\u0_tms_reg[22]/NET0131 ,
		_w3203_,
		_w3554_
	);
	LUT2 #(
		.INIT('h8)
	) name2596 (
		\u0_u1_tms_reg[22]/P0001 ,
		_w3458_,
		_w3555_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		\u0_u0_tms_reg[22]/P0001 ,
		_w3415_,
		_w3556_
	);
	LUT2 #(
		.INIT('h1)
	) name2598 (
		_w3555_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h2)
	) name2599 (
		_w3203_,
		_w3557_,
		_w3558_
	);
	LUT2 #(
		.INIT('h1)
	) name2600 (
		_w3554_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h2)
	) name2601 (
		\u0_tms_reg[25]/NET0131 ,
		_w3203_,
		_w3560_
	);
	LUT2 #(
		.INIT('h8)
	) name2602 (
		\u0_u1_tms_reg[25]/P0001 ,
		_w3458_,
		_w3561_
	);
	LUT2 #(
		.INIT('h8)
	) name2603 (
		\u0_u0_tms_reg[25]/P0001 ,
		_w3415_,
		_w3562_
	);
	LUT2 #(
		.INIT('h1)
	) name2604 (
		_w3561_,
		_w3562_,
		_w3563_
	);
	LUT2 #(
		.INIT('h2)
	) name2605 (
		_w3203_,
		_w3563_,
		_w3564_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		_w3560_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h2)
	) name2607 (
		\u0_tms_reg[26]/NET0131 ,
		_w3203_,
		_w3566_
	);
	LUT2 #(
		.INIT('h8)
	) name2608 (
		\u0_u1_tms_reg[26]/P0001 ,
		_w3458_,
		_w3567_
	);
	LUT2 #(
		.INIT('h8)
	) name2609 (
		\u0_u0_tms_reg[26]/P0001 ,
		_w3415_,
		_w3568_
	);
	LUT2 #(
		.INIT('h1)
	) name2610 (
		_w3567_,
		_w3568_,
		_w3569_
	);
	LUT2 #(
		.INIT('h2)
	) name2611 (
		_w3203_,
		_w3569_,
		_w3570_
	);
	LUT2 #(
		.INIT('h1)
	) name2612 (
		_w3566_,
		_w3570_,
		_w3571_
	);
	LUT2 #(
		.INIT('h2)
	) name2613 (
		\u0_tms_reg[27]/NET0131 ,
		_w3203_,
		_w3572_
	);
	LUT2 #(
		.INIT('h8)
	) name2614 (
		\u0_u1_tms_reg[27]/P0001 ,
		_w3458_,
		_w3573_
	);
	LUT2 #(
		.INIT('h8)
	) name2615 (
		\u0_u0_tms_reg[27]/P0001 ,
		_w3415_,
		_w3574_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		_w3573_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h2)
	) name2617 (
		_w3203_,
		_w3575_,
		_w3576_
	);
	LUT2 #(
		.INIT('h1)
	) name2618 (
		_w3572_,
		_w3576_,
		_w3577_
	);
	LUT2 #(
		.INIT('h2)
	) name2619 (
		\u0_tms_reg[2]/NET0131 ,
		_w3203_,
		_w3578_
	);
	LUT2 #(
		.INIT('h8)
	) name2620 (
		\u0_u1_tms_reg[2]/P0001 ,
		_w3458_,
		_w3579_
	);
	LUT2 #(
		.INIT('h8)
	) name2621 (
		\u0_u0_tms_reg[2]/P0001 ,
		_w3415_,
		_w3580_
	);
	LUT2 #(
		.INIT('h1)
	) name2622 (
		_w3579_,
		_w3580_,
		_w3581_
	);
	LUT2 #(
		.INIT('h2)
	) name2623 (
		_w3203_,
		_w3581_,
		_w3582_
	);
	LUT2 #(
		.INIT('h1)
	) name2624 (
		_w3578_,
		_w3582_,
		_w3583_
	);
	LUT2 #(
		.INIT('h2)
	) name2625 (
		\u0_tms_reg[3]/NET0131 ,
		_w3203_,
		_w3584_
	);
	LUT2 #(
		.INIT('h8)
	) name2626 (
		\u0_u1_tms_reg[3]/P0001 ,
		_w3458_,
		_w3585_
	);
	LUT2 #(
		.INIT('h8)
	) name2627 (
		\u0_u0_tms_reg[3]/P0001 ,
		_w3415_,
		_w3586_
	);
	LUT2 #(
		.INIT('h1)
	) name2628 (
		_w3585_,
		_w3586_,
		_w3587_
	);
	LUT2 #(
		.INIT('h2)
	) name2629 (
		_w3203_,
		_w3587_,
		_w3588_
	);
	LUT2 #(
		.INIT('h1)
	) name2630 (
		_w3584_,
		_w3588_,
		_w3589_
	);
	LUT2 #(
		.INIT('h2)
	) name2631 (
		\u0_tms_reg[4]/NET0131 ,
		_w3203_,
		_w3590_
	);
	LUT2 #(
		.INIT('h8)
	) name2632 (
		\u0_u1_tms_reg[4]/P0001 ,
		_w3458_,
		_w3591_
	);
	LUT2 #(
		.INIT('h8)
	) name2633 (
		\u0_u0_tms_reg[4]/P0001 ,
		_w3415_,
		_w3592_
	);
	LUT2 #(
		.INIT('h1)
	) name2634 (
		_w3591_,
		_w3592_,
		_w3593_
	);
	LUT2 #(
		.INIT('h2)
	) name2635 (
		_w3203_,
		_w3593_,
		_w3594_
	);
	LUT2 #(
		.INIT('h1)
	) name2636 (
		_w3590_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h2)
	) name2637 (
		\u0_tms_reg[5]/NET0131 ,
		_w3203_,
		_w3596_
	);
	LUT2 #(
		.INIT('h8)
	) name2638 (
		\u0_u1_tms_reg[5]/P0001 ,
		_w3458_,
		_w3597_
	);
	LUT2 #(
		.INIT('h8)
	) name2639 (
		\u0_u0_tms_reg[5]/P0001 ,
		_w3415_,
		_w3598_
	);
	LUT2 #(
		.INIT('h1)
	) name2640 (
		_w3597_,
		_w3598_,
		_w3599_
	);
	LUT2 #(
		.INIT('h2)
	) name2641 (
		_w3203_,
		_w3599_,
		_w3600_
	);
	LUT2 #(
		.INIT('h1)
	) name2642 (
		_w3596_,
		_w3600_,
		_w3601_
	);
	LUT2 #(
		.INIT('h2)
	) name2643 (
		\u0_tms_reg[6]/NET0131 ,
		_w3203_,
		_w3602_
	);
	LUT2 #(
		.INIT('h8)
	) name2644 (
		\u0_u1_tms_reg[6]/P0001 ,
		_w3458_,
		_w3603_
	);
	LUT2 #(
		.INIT('h8)
	) name2645 (
		\u0_u0_tms_reg[6]/P0001 ,
		_w3415_,
		_w3604_
	);
	LUT2 #(
		.INIT('h1)
	) name2646 (
		_w3603_,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('h2)
	) name2647 (
		_w3203_,
		_w3605_,
		_w3606_
	);
	LUT2 #(
		.INIT('h1)
	) name2648 (
		_w3602_,
		_w3606_,
		_w3607_
	);
	LUT2 #(
		.INIT('h2)
	) name2649 (
		\u0_tms_reg[7]/NET0131 ,
		_w3203_,
		_w3608_
	);
	LUT2 #(
		.INIT('h8)
	) name2650 (
		\u0_u1_tms_reg[7]/P0001 ,
		_w3458_,
		_w3609_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		\u0_u0_tms_reg[7]/P0001 ,
		_w3415_,
		_w3610_
	);
	LUT2 #(
		.INIT('h1)
	) name2652 (
		_w3609_,
		_w3610_,
		_w3611_
	);
	LUT2 #(
		.INIT('h2)
	) name2653 (
		_w3203_,
		_w3611_,
		_w3612_
	);
	LUT2 #(
		.INIT('h1)
	) name2654 (
		_w3608_,
		_w3612_,
		_w3613_
	);
	LUT2 #(
		.INIT('h2)
	) name2655 (
		\u0_tms_reg[8]/NET0131 ,
		_w3203_,
		_w3614_
	);
	LUT2 #(
		.INIT('h8)
	) name2656 (
		\u0_u1_tms_reg[8]/P0001 ,
		_w3458_,
		_w3615_
	);
	LUT2 #(
		.INIT('h8)
	) name2657 (
		\u0_u0_tms_reg[8]/P0001 ,
		_w3415_,
		_w3616_
	);
	LUT2 #(
		.INIT('h1)
	) name2658 (
		_w3615_,
		_w3616_,
		_w3617_
	);
	LUT2 #(
		.INIT('h2)
	) name2659 (
		_w3203_,
		_w3617_,
		_w3618_
	);
	LUT2 #(
		.INIT('h1)
	) name2660 (
		_w3614_,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('h2)
	) name2661 (
		\u0_tms_reg[9]/NET0131 ,
		_w3203_,
		_w3620_
	);
	LUT2 #(
		.INIT('h8)
	) name2662 (
		\u0_u1_tms_reg[9]/P0001 ,
		_w3458_,
		_w3621_
	);
	LUT2 #(
		.INIT('h8)
	) name2663 (
		\u0_u0_tms_reg[9]/P0001 ,
		_w3415_,
		_w3622_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		_w3621_,
		_w3622_,
		_w3623_
	);
	LUT2 #(
		.INIT('h2)
	) name2665 (
		_w3203_,
		_w3623_,
		_w3624_
	);
	LUT2 #(
		.INIT('h1)
	) name2666 (
		_w3620_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('h4)
	) name2667 (
		_w2282_,
		_w2818_,
		_w3626_
	);
	LUT2 #(
		.INIT('h8)
	) name2668 (
		\u0_tms_reg[6]/NET0131 ,
		_w1051_,
		_w3627_
	);
	LUT2 #(
		.INIT('h2)
	) name2669 (
		\u0_sp_tms_reg[6]/NET0131 ,
		_w1051_,
		_w3628_
	);
	LUT2 #(
		.INIT('h1)
	) name2670 (
		_w3627_,
		_w3628_,
		_w3629_
	);
	LUT2 #(
		.INIT('h8)
	) name2671 (
		_w1693_,
		_w3629_,
		_w3630_
	);
	LUT2 #(
		.INIT('h4)
	) name2672 (
		_w2833_,
		_w3630_,
		_w3631_
	);
	LUT2 #(
		.INIT('h1)
	) name2673 (
		\u5_timer2_reg[7]/P0001 ,
		_w3169_,
		_w3632_
	);
	LUT2 #(
		.INIT('h8)
	) name2674 (
		\u5_timer2_reg[7]/P0001 ,
		_w2840_,
		_w3633_
	);
	LUT2 #(
		.INIT('h1)
	) name2675 (
		_w3632_,
		_w3633_,
		_w3634_
	);
	LUT2 #(
		.INIT('h2)
	) name2676 (
		_w2833_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('h1)
	) name2677 (
		_w3631_,
		_w3635_,
		_w3636_
	);
	LUT2 #(
		.INIT('h8)
	) name2678 (
		_w3173_,
		_w3636_,
		_w3637_
	);
	LUT2 #(
		.INIT('h1)
	) name2679 (
		_w3626_,
		_w3637_,
		_w3638_
	);
	LUT2 #(
		.INIT('h4)
	) name2680 (
		_w2519_,
		_w2818_,
		_w3639_
	);
	LUT2 #(
		.INIT('h2)
	) name2681 (
		\u5_timer2_reg[8]/P0001 ,
		_w2841_,
		_w3640_
	);
	LUT2 #(
		.INIT('h2)
	) name2682 (
		_w2833_,
		_w3640_,
		_w3641_
	);
	LUT2 #(
		.INIT('h8)
	) name2683 (
		\u0_tms_reg[7]/NET0131 ,
		_w1051_,
		_w3642_
	);
	LUT2 #(
		.INIT('h2)
	) name2684 (
		\u0_sp_tms_reg[7]/NET0131 ,
		_w1051_,
		_w3643_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		_w3642_,
		_w3643_,
		_w3644_
	);
	LUT2 #(
		.INIT('h8)
	) name2686 (
		_w1693_,
		_w3644_,
		_w3645_
	);
	LUT2 #(
		.INIT('h4)
	) name2687 (
		_w2833_,
		_w3645_,
		_w3646_
	);
	LUT2 #(
		.INIT('h1)
	) name2688 (
		_w3641_,
		_w3646_,
		_w3647_
	);
	LUT2 #(
		.INIT('h8)
	) name2689 (
		_w3173_,
		_w3647_,
		_w3648_
	);
	LUT2 #(
		.INIT('h1)
	) name2690 (
		_w3639_,
		_w3648_,
		_w3649_
	);
	LUT2 #(
		.INIT('h8)
	) name2691 (
		\wb_addr_i[15]_pad ,
		_w2388_,
		_w3650_
	);
	LUT2 #(
		.INIT('h8)
	) name2692 (
		\wb_addr_i[17]_pad ,
		_w2878_,
		_w3651_
	);
	LUT2 #(
		.INIT('h8)
	) name2693 (
		\wb_addr_i[16]_pad ,
		_w2606_,
		_w3652_
	);
	LUT2 #(
		.INIT('h1)
	) name2694 (
		_w3650_,
		_w3651_,
		_w3653_
	);
	LUT2 #(
		.INIT('h4)
	) name2695 (
		_w3652_,
		_w3653_,
		_w3654_
	);
	LUT2 #(
		.INIT('h1)
	) name2696 (
		_w2858_,
		_w3654_,
		_w3655_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		\u1_acs_addr_reg[15]/P0001 ,
		_w2865_,
		_w3656_
	);
	LUT2 #(
		.INIT('h2)
	) name2698 (
		_w2858_,
		_w2866_,
		_w3657_
	);
	LUT2 #(
		.INIT('h4)
	) name2699 (
		_w3656_,
		_w3657_,
		_w3658_
	);
	LUT2 #(
		.INIT('h1)
	) name2700 (
		_w3655_,
		_w3658_,
		_w3659_
	);
	LUT2 #(
		.INIT('h2)
	) name2701 (
		_w1046_,
		_w3201_,
		_w3660_
	);
	LUT2 #(
		.INIT('h8)
	) name2702 (
		\u0_u1_csc_reg[4]/P0001 ,
		_w3660_,
		_w3661_
	);
	LUT2 #(
		.INIT('h8)
	) name2703 (
		_w3458_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h8)
	) name2704 (
		_w3415_,
		_w3660_,
		_w3663_
	);
	LUT2 #(
		.INIT('h8)
	) name2705 (
		\u0_u0_csc_reg[4]/P0001 ,
		_w3663_,
		_w3664_
	);
	LUT2 #(
		.INIT('h2)
	) name2706 (
		\u0_csc_reg[4]/NET0131 ,
		_w3660_,
		_w3665_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		_w3662_,
		_w3665_,
		_w3666_
	);
	LUT2 #(
		.INIT('h4)
	) name2708 (
		_w3664_,
		_w3666_,
		_w3667_
	);
	LUT2 #(
		.INIT('h8)
	) name2709 (
		\u0_u1_csc_reg[5]/P0001 ,
		_w3660_,
		_w3668_
	);
	LUT2 #(
		.INIT('h8)
	) name2710 (
		_w3458_,
		_w3668_,
		_w3669_
	);
	LUT2 #(
		.INIT('h8)
	) name2711 (
		\u0_u0_csc_reg[5]/P0001 ,
		_w3663_,
		_w3670_
	);
	LUT2 #(
		.INIT('h2)
	) name2712 (
		\u0_csc_reg[5]/NET0131 ,
		_w3660_,
		_w3671_
	);
	LUT2 #(
		.INIT('h1)
	) name2713 (
		_w3669_,
		_w3671_,
		_w3672_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		_w3670_,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('h8)
	) name2715 (
		\u0_u0_csc_reg[6]/P0001 ,
		_w3663_,
		_w3674_
	);
	LUT2 #(
		.INIT('h8)
	) name2716 (
		\u0_u1_csc_reg[6]/P0001 ,
		_w3660_,
		_w3675_
	);
	LUT2 #(
		.INIT('h8)
	) name2717 (
		_w3458_,
		_w3675_,
		_w3676_
	);
	LUT2 #(
		.INIT('h2)
	) name2718 (
		\u0_csc_reg[6]/NET0131 ,
		_w3660_,
		_w3677_
	);
	LUT2 #(
		.INIT('h1)
	) name2719 (
		_w3674_,
		_w3677_,
		_w3678_
	);
	LUT2 #(
		.INIT('h4)
	) name2720 (
		_w3676_,
		_w3678_,
		_w3679_
	);
	LUT2 #(
		.INIT('h8)
	) name2721 (
		\u0_u0_csc_reg[9]/P0001 ,
		_w3663_,
		_w3680_
	);
	LUT2 #(
		.INIT('h8)
	) name2722 (
		\u0_u1_csc_reg[9]/P0001 ,
		_w3660_,
		_w3681_
	);
	LUT2 #(
		.INIT('h8)
	) name2723 (
		_w3458_,
		_w3681_,
		_w3682_
	);
	LUT2 #(
		.INIT('h2)
	) name2724 (
		\u0_csc_reg[9]/NET0131 ,
		_w3660_,
		_w3683_
	);
	LUT2 #(
		.INIT('h1)
	) name2725 (
		_w3680_,
		_w3683_,
		_w3684_
	);
	LUT2 #(
		.INIT('h4)
	) name2726 (
		_w3682_,
		_w3684_,
		_w3685_
	);
	LUT2 #(
		.INIT('h8)
	) name2727 (
		\u0_u0_csc_reg[7]/P0001 ,
		_w3663_,
		_w3686_
	);
	LUT2 #(
		.INIT('h8)
	) name2728 (
		\u0_u1_csc_reg[7]/P0001 ,
		_w3660_,
		_w3687_
	);
	LUT2 #(
		.INIT('h8)
	) name2729 (
		_w3458_,
		_w3687_,
		_w3688_
	);
	LUT2 #(
		.INIT('h2)
	) name2730 (
		\u0_csc_reg[7]/NET0131 ,
		_w3660_,
		_w3689_
	);
	LUT2 #(
		.INIT('h1)
	) name2731 (
		_w3686_,
		_w3689_,
		_w3690_
	);
	LUT2 #(
		.INIT('h4)
	) name2732 (
		_w3688_,
		_w3690_,
		_w3691_
	);
	LUT2 #(
		.INIT('h8)
	) name2733 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		_w3660_,
		_w3692_
	);
	LUT2 #(
		.INIT('h8)
	) name2734 (
		\u0_u0_csc_reg[10]/P0001 ,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h8)
	) name2735 (
		\u0_u1_csc_reg[10]/P0001 ,
		_w3660_,
		_w3694_
	);
	LUT2 #(
		.INIT('h8)
	) name2736 (
		_w3206_,
		_w3694_,
		_w3695_
	);
	LUT2 #(
		.INIT('h2)
	) name2737 (
		\u0_sp_csc_reg[10]/NET0131 ,
		_w3660_,
		_w3696_
	);
	LUT2 #(
		.INIT('h1)
	) name2738 (
		_w3693_,
		_w3696_,
		_w3697_
	);
	LUT2 #(
		.INIT('h4)
	) name2739 (
		_w3695_,
		_w3697_,
		_w3698_
	);
	LUT2 #(
		.INIT('h8)
	) name2740 (
		\u0_u0_csc_reg[4]/P0001 ,
		_w3692_,
		_w3699_
	);
	LUT2 #(
		.INIT('h8)
	) name2741 (
		_w3206_,
		_w3661_,
		_w3700_
	);
	LUT2 #(
		.INIT('h2)
	) name2742 (
		\u0_sp_csc_reg[4]/NET0131 ,
		_w3660_,
		_w3701_
	);
	LUT2 #(
		.INIT('h1)
	) name2743 (
		_w3699_,
		_w3701_,
		_w3702_
	);
	LUT2 #(
		.INIT('h4)
	) name2744 (
		_w3700_,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h8)
	) name2745 (
		\u0_u0_csc_reg[5]/P0001 ,
		_w3692_,
		_w3704_
	);
	LUT2 #(
		.INIT('h8)
	) name2746 (
		_w3206_,
		_w3668_,
		_w3705_
	);
	LUT2 #(
		.INIT('h2)
	) name2747 (
		\u0_sp_csc_reg[5]/NET0131 ,
		_w3660_,
		_w3706_
	);
	LUT2 #(
		.INIT('h1)
	) name2748 (
		_w3704_,
		_w3706_,
		_w3707_
	);
	LUT2 #(
		.INIT('h4)
	) name2749 (
		_w3705_,
		_w3707_,
		_w3708_
	);
	LUT2 #(
		.INIT('h8)
	) name2750 (
		\u0_u0_csc_reg[6]/P0001 ,
		_w3692_,
		_w3709_
	);
	LUT2 #(
		.INIT('h8)
	) name2751 (
		_w3206_,
		_w3675_,
		_w3710_
	);
	LUT2 #(
		.INIT('h2)
	) name2752 (
		\u0_sp_csc_reg[6]/NET0131 ,
		_w3660_,
		_w3711_
	);
	LUT2 #(
		.INIT('h1)
	) name2753 (
		_w3709_,
		_w3711_,
		_w3712_
	);
	LUT2 #(
		.INIT('h4)
	) name2754 (
		_w3710_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('h8)
	) name2755 (
		\u0_u0_csc_reg[7]/P0001 ,
		_w3692_,
		_w3714_
	);
	LUT2 #(
		.INIT('h8)
	) name2756 (
		_w3206_,
		_w3687_,
		_w3715_
	);
	LUT2 #(
		.INIT('h2)
	) name2757 (
		\u0_sp_csc_reg[7]/NET0131 ,
		_w3660_,
		_w3716_
	);
	LUT2 #(
		.INIT('h1)
	) name2758 (
		_w3714_,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h4)
	) name2759 (
		_w3715_,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h8)
	) name2760 (
		\u0_u0_csc_reg[9]/P0001 ,
		_w3692_,
		_w3719_
	);
	LUT2 #(
		.INIT('h8)
	) name2761 (
		_w3206_,
		_w3681_,
		_w3720_
	);
	LUT2 #(
		.INIT('h2)
	) name2762 (
		\u0_sp_csc_reg[9]/NET0131 ,
		_w3660_,
		_w3721_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		_w3719_,
		_w3721_,
		_w3722_
	);
	LUT2 #(
		.INIT('h4)
	) name2764 (
		_w3720_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h8)
	) name2765 (
		_w3458_,
		_w3694_,
		_w3724_
	);
	LUT2 #(
		.INIT('h8)
	) name2766 (
		\u0_u0_csc_reg[10]/P0001 ,
		_w3663_,
		_w3725_
	);
	LUT2 #(
		.INIT('h2)
	) name2767 (
		\u0_csc_reg[10]/NET0131 ,
		_w3660_,
		_w3726_
	);
	LUT2 #(
		.INIT('h1)
	) name2768 (
		_w3724_,
		_w3726_,
		_w3727_
	);
	LUT2 #(
		.INIT('h4)
	) name2769 (
		_w3725_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h2)
	) name2770 (
		\u5_ap_en_reg/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w3729_
	);
	LUT2 #(
		.INIT('h8)
	) name2771 (
		_w1375_,
		_w2399_,
		_w3730_
	);
	LUT2 #(
		.INIT('h1)
	) name2772 (
		_w3729_,
		_w3730_,
		_w3731_
	);
	LUT2 #(
		.INIT('h2)
	) name2773 (
		\u0_sp_csc_reg[2]/NET0131 ,
		_w3660_,
		_w3732_
	);
	LUT2 #(
		.INIT('h8)
	) name2774 (
		\u0_u0_csc_reg[2]/NET0131 ,
		_w3692_,
		_w3733_
	);
	LUT2 #(
		.INIT('h8)
	) name2775 (
		\u0_u1_csc_reg[2]/NET0131 ,
		_w3206_,
		_w3734_
	);
	LUT2 #(
		.INIT('h8)
	) name2776 (
		_w3660_,
		_w3734_,
		_w3735_
	);
	LUT2 #(
		.INIT('h1)
	) name2777 (
		_w3732_,
		_w3735_,
		_w3736_
	);
	LUT2 #(
		.INIT('h4)
	) name2778 (
		_w3733_,
		_w3736_,
		_w3737_
	);
	LUT2 #(
		.INIT('h2)
	) name2779 (
		\u0_sp_csc_reg[1]/NET0131 ,
		_w3660_,
		_w3738_
	);
	LUT2 #(
		.INIT('h8)
	) name2780 (
		\u0_u0_csc_reg[1]/NET0131 ,
		_w3692_,
		_w3739_
	);
	LUT2 #(
		.INIT('h8)
	) name2781 (
		\u0_u1_csc_reg[1]/NET0131 ,
		_w3206_,
		_w3740_
	);
	LUT2 #(
		.INIT('h8)
	) name2782 (
		_w3660_,
		_w3740_,
		_w3741_
	);
	LUT2 #(
		.INIT('h1)
	) name2783 (
		_w3738_,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('h4)
	) name2784 (
		_w3739_,
		_w3742_,
		_w3743_
	);
	LUT2 #(
		.INIT('h2)
	) name2785 (
		\u0_sp_csc_reg[3]/NET0131 ,
		_w3660_,
		_w3744_
	);
	LUT2 #(
		.INIT('h8)
	) name2786 (
		\u0_u0_csc_reg[3]/NET0131 ,
		_w3692_,
		_w3745_
	);
	LUT2 #(
		.INIT('h8)
	) name2787 (
		\u0_u1_csc_reg[3]/NET0131 ,
		_w3206_,
		_w3746_
	);
	LUT2 #(
		.INIT('h8)
	) name2788 (
		_w3660_,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h1)
	) name2789 (
		_w3744_,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h4)
	) name2790 (
		_w3745_,
		_w3748_,
		_w3749_
	);
	LUT2 #(
		.INIT('h8)
	) name2791 (
		_w1777_,
		_w1785_,
		_w3750_
	);
	LUT2 #(
		.INIT('h1)
	) name2792 (
		_w1817_,
		_w2529_,
		_w3751_
	);
	LUT2 #(
		.INIT('h2)
	) name2793 (
		\u5_timer_reg[4]/NET0131 ,
		_w2285_,
		_w3752_
	);
	LUT2 #(
		.INIT('h4)
	) name2794 (
		\u5_timer_reg[4]/NET0131 ,
		_w2285_,
		_w3753_
	);
	LUT2 #(
		.INIT('h1)
	) name2795 (
		_w3752_,
		_w3753_,
		_w3754_
	);
	LUT2 #(
		.INIT('h8)
	) name2796 (
		_w1817_,
		_w2288_,
		_w3755_
	);
	LUT2 #(
		.INIT('h8)
	) name2797 (
		_w2296_,
		_w3755_,
		_w3756_
	);
	LUT2 #(
		.INIT('h4)
	) name2798 (
		_w3754_,
		_w3756_,
		_w3757_
	);
	LUT2 #(
		.INIT('h1)
	) name2799 (
		_w3751_,
		_w3757_,
		_w3758_
	);
	LUT2 #(
		.INIT('h2)
	) name2800 (
		_w3750_,
		_w3758_,
		_w3759_
	);
	LUT2 #(
		.INIT('h1)
	) name2801 (
		_w1817_,
		_w2584_,
		_w3760_
	);
	LUT2 #(
		.INIT('h2)
	) name2802 (
		\u5_timer_reg[5]/NET0131 ,
		_w3753_,
		_w3761_
	);
	LUT2 #(
		.INIT('h8)
	) name2803 (
		_w1823_,
		_w1830_,
		_w3762_
	);
	LUT2 #(
		.INIT('h1)
	) name2804 (
		_w3761_,
		_w3762_,
		_w3763_
	);
	LUT2 #(
		.INIT('h2)
	) name2805 (
		_w3756_,
		_w3763_,
		_w3764_
	);
	LUT2 #(
		.INIT('h1)
	) name2806 (
		_w3760_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h2)
	) name2807 (
		_w3750_,
		_w3765_,
		_w3766_
	);
	LUT2 #(
		.INIT('h2)
	) name2808 (
		\u5_timer_reg[6]/NET0131 ,
		_w3762_,
		_w3767_
	);
	LUT2 #(
		.INIT('h4)
	) name2809 (
		\u5_mc_le_reg/NET0131 ,
		_w1826_,
		_w3768_
	);
	LUT2 #(
		.INIT('h4)
	) name2810 (
		_w1827_,
		_w3768_,
		_w3769_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w3767_,
		_w3769_,
		_w3770_
	);
	LUT2 #(
		.INIT('h2)
	) name2812 (
		_w3756_,
		_w3770_,
		_w3771_
	);
	LUT2 #(
		.INIT('h1)
	) name2813 (
		_w1817_,
		_w3630_,
		_w3772_
	);
	LUT2 #(
		.INIT('h1)
	) name2814 (
		_w3771_,
		_w3772_,
		_w3773_
	);
	LUT2 #(
		.INIT('h2)
	) name2815 (
		_w3750_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('h1)
	) name2816 (
		_w1817_,
		_w3645_,
		_w3775_
	);
	LUT2 #(
		.INIT('h2)
	) name2817 (
		\u5_timer_reg[7]/NET0131 ,
		_w3768_,
		_w3776_
	);
	LUT2 #(
		.INIT('h8)
	) name2818 (
		_w3756_,
		_w3776_,
		_w3777_
	);
	LUT2 #(
		.INIT('h1)
	) name2819 (
		_w3775_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h2)
	) name2820 (
		_w3750_,
		_w3778_,
		_w3779_
	);
	LUT2 #(
		.INIT('h2)
	) name2821 (
		\u0_csc_reg[11]/NET0131 ,
		_w3660_,
		_w3780_
	);
	LUT2 #(
		.INIT('h8)
	) name2822 (
		\u0_u1_csc_reg[11]/P0001 ,
		_w3458_,
		_w3781_
	);
	LUT2 #(
		.INIT('h8)
	) name2823 (
		\u0_u0_csc_reg[11]/P0001 ,
		_w3415_,
		_w3782_
	);
	LUT2 #(
		.INIT('h1)
	) name2824 (
		_w3781_,
		_w3782_,
		_w3783_
	);
	LUT2 #(
		.INIT('h2)
	) name2825 (
		_w3660_,
		_w3783_,
		_w3784_
	);
	LUT2 #(
		.INIT('h1)
	) name2826 (
		_w3780_,
		_w3784_,
		_w3785_
	);
	LUT2 #(
		.INIT('h8)
	) name2827 (
		\wb_addr_i[14]_pad ,
		_w2388_,
		_w3786_
	);
	LUT2 #(
		.INIT('h8)
	) name2828 (
		\wb_addr_i[16]_pad ,
		_w2878_,
		_w3787_
	);
	LUT2 #(
		.INIT('h8)
	) name2829 (
		\wb_addr_i[15]_pad ,
		_w2606_,
		_w3788_
	);
	LUT2 #(
		.INIT('h1)
	) name2830 (
		_w3786_,
		_w3787_,
		_w3789_
	);
	LUT2 #(
		.INIT('h4)
	) name2831 (
		_w3788_,
		_w3789_,
		_w3790_
	);
	LUT2 #(
		.INIT('h1)
	) name2832 (
		_w2858_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('h1)
	) name2833 (
		\u1_acs_addr_reg[14]/P0001 ,
		_w2864_,
		_w3792_
	);
	LUT2 #(
		.INIT('h2)
	) name2834 (
		_w2858_,
		_w2865_,
		_w3793_
	);
	LUT2 #(
		.INIT('h4)
	) name2835 (
		_w3792_,
		_w3793_,
		_w3794_
	);
	LUT2 #(
		.INIT('h1)
	) name2836 (
		_w3791_,
		_w3794_,
		_w3795_
	);
	LUT2 #(
		.INIT('h8)
	) name2837 (
		_w1666_,
		_w1686_,
		_w3796_
	);
	LUT2 #(
		.INIT('h1)
	) name2838 (
		_w1139_,
		_w1241_,
		_w3797_
	);
	LUT2 #(
		.INIT('h1)
	) name2839 (
		_w1627_,
		_w3797_,
		_w3798_
	);
	LUT2 #(
		.INIT('h1)
	) name2840 (
		_w1139_,
		_w1664_,
		_w3799_
	);
	LUT2 #(
		.INIT('h2)
	) name2841 (
		_w1287_,
		_w3799_,
		_w3800_
	);
	LUT2 #(
		.INIT('h4)
	) name2842 (
		_w1108_,
		_w1315_,
		_w3801_
	);
	LUT2 #(
		.INIT('h4)
	) name2843 (
		_w3796_,
		_w3801_,
		_w3802_
	);
	LUT2 #(
		.INIT('h1)
	) name2844 (
		_w3798_,
		_w3800_,
		_w3803_
	);
	LUT2 #(
		.INIT('h8)
	) name2845 (
		_w3802_,
		_w3803_,
		_w3804_
	);
	LUT2 #(
		.INIT('h8)
	) name2846 (
		\u5_cmd_del_reg[2]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w3805_
	);
	LUT2 #(
		.INIT('h8)
	) name2847 (
		\u5_wb_wait_r_reg/P0001 ,
		_w1300_,
		_w3806_
	);
	LUT2 #(
		.INIT('h1)
	) name2848 (
		_w1425_,
		_w3806_,
		_w3807_
	);
	LUT2 #(
		.INIT('h8)
	) name2849 (
		_w1298_,
		_w3807_,
		_w3808_
	);
	LUT2 #(
		.INIT('h8)
	) name2850 (
		_w1127_,
		_w3808_,
		_w3809_
	);
	LUT2 #(
		.INIT('h8)
	) name2851 (
		_w2941_,
		_w3809_,
		_w3810_
	);
	LUT2 #(
		.INIT('h8)
	) name2852 (
		_w3001_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h1)
	) name2853 (
		\u5_wr_cycle_reg/NET0131 ,
		_w3811_,
		_w3812_
	);
	LUT2 #(
		.INIT('h1)
	) name2854 (
		_w3805_,
		_w3812_,
		_w3813_
	);
	LUT2 #(
		.INIT('h8)
	) name2855 (
		\wb_addr_i[21]_pad ,
		_w2388_,
		_w3814_
	);
	LUT2 #(
		.INIT('h8)
	) name2856 (
		\wb_addr_i[23]_pad ,
		_w2878_,
		_w3815_
	);
	LUT2 #(
		.INIT('h8)
	) name2857 (
		\wb_addr_i[22]_pad ,
		_w2606_,
		_w3816_
	);
	LUT2 #(
		.INIT('h1)
	) name2858 (
		_w3814_,
		_w3815_,
		_w3817_
	);
	LUT2 #(
		.INIT('h4)
	) name2859 (
		_w3816_,
		_w3817_,
		_w3818_
	);
	LUT2 #(
		.INIT('h1)
	) name2860 (
		_w2858_,
		_w3818_,
		_w3819_
	);
	LUT2 #(
		.INIT('h1)
	) name2861 (
		\u1_acs_addr_reg[21]/P0001 ,
		_w2871_,
		_w3820_
	);
	LUT2 #(
		.INIT('h2)
	) name2862 (
		_w2858_,
		_w2872_,
		_w3821_
	);
	LUT2 #(
		.INIT('h4)
	) name2863 (
		_w3820_,
		_w3821_,
		_w3822_
	);
	LUT2 #(
		.INIT('h1)
	) name2864 (
		_w3819_,
		_w3822_,
		_w3823_
	);
	LUT2 #(
		.INIT('h1)
	) name2865 (
		\u4_rfr_clr_reg/P0001 ,
		\u4_rfr_req_reg/NET0131 ,
		_w3824_
	);
	LUT2 #(
		.INIT('h1)
	) name2866 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('h8)
	) name2867 (
		\wb_addr_i[13]_pad ,
		_w2388_,
		_w3826_
	);
	LUT2 #(
		.INIT('h8)
	) name2868 (
		\wb_addr_i[15]_pad ,
		_w2878_,
		_w3827_
	);
	LUT2 #(
		.INIT('h8)
	) name2869 (
		\wb_addr_i[14]_pad ,
		_w2606_,
		_w3828_
	);
	LUT2 #(
		.INIT('h1)
	) name2870 (
		_w3826_,
		_w3827_,
		_w3829_
	);
	LUT2 #(
		.INIT('h4)
	) name2871 (
		_w3828_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h1)
	) name2872 (
		_w2858_,
		_w3830_,
		_w3831_
	);
	LUT2 #(
		.INIT('h1)
	) name2873 (
		\u1_acs_addr_reg[13]/P0001 ,
		_w2863_,
		_w3832_
	);
	LUT2 #(
		.INIT('h2)
	) name2874 (
		_w2858_,
		_w2864_,
		_w3833_
	);
	LUT2 #(
		.INIT('h4)
	) name2875 (
		_w3832_,
		_w3833_,
		_w3834_
	);
	LUT2 #(
		.INIT('h1)
	) name2876 (
		_w3831_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h1)
	) name2877 (
		\u1_acs_addr_reg[11]/P0001 ,
		_w2861_,
		_w3836_
	);
	LUT2 #(
		.INIT('h4)
	) name2878 (
		\u1_u0_out_r_reg[11]/P0001 ,
		_w2861_,
		_w3837_
	);
	LUT2 #(
		.INIT('h2)
	) name2879 (
		_w2858_,
		_w3836_,
		_w3838_
	);
	LUT2 #(
		.INIT('h4)
	) name2880 (
		_w3837_,
		_w3838_,
		_w3839_
	);
	LUT2 #(
		.INIT('h8)
	) name2881 (
		\wb_addr_i[11]_pad ,
		_w2388_,
		_w3840_
	);
	LUT2 #(
		.INIT('h8)
	) name2882 (
		\wb_addr_i[12]_pad ,
		_w2606_,
		_w3841_
	);
	LUT2 #(
		.INIT('h8)
	) name2883 (
		\wb_addr_i[13]_pad ,
		_w2878_,
		_w3842_
	);
	LUT2 #(
		.INIT('h1)
	) name2884 (
		_w3840_,
		_w3841_,
		_w3843_
	);
	LUT2 #(
		.INIT('h4)
	) name2885 (
		_w3842_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h1)
	) name2886 (
		_w2858_,
		_w3844_,
		_w3845_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		_w3839_,
		_w3845_,
		_w3846_
	);
	LUT2 #(
		.INIT('h8)
	) name2888 (
		\wb_addr_i[17]_pad ,
		_w2388_,
		_w3847_
	);
	LUT2 #(
		.INIT('h8)
	) name2889 (
		\wb_addr_i[19]_pad ,
		_w2878_,
		_w3848_
	);
	LUT2 #(
		.INIT('h8)
	) name2890 (
		\wb_addr_i[18]_pad ,
		_w2606_,
		_w3849_
	);
	LUT2 #(
		.INIT('h1)
	) name2891 (
		_w3847_,
		_w3848_,
		_w3850_
	);
	LUT2 #(
		.INIT('h4)
	) name2892 (
		_w3849_,
		_w3850_,
		_w3851_
	);
	LUT2 #(
		.INIT('h1)
	) name2893 (
		_w2858_,
		_w3851_,
		_w3852_
	);
	LUT2 #(
		.INIT('h1)
	) name2894 (
		\u1_acs_addr_reg[17]/P0001 ,
		_w2867_,
		_w3853_
	);
	LUT2 #(
		.INIT('h2)
	) name2895 (
		_w2858_,
		_w2868_,
		_w3854_
	);
	LUT2 #(
		.INIT('h4)
	) name2896 (
		_w3853_,
		_w3854_,
		_w3855_
	);
	LUT2 #(
		.INIT('h1)
	) name2897 (
		_w3852_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h8)
	) name2898 (
		_w1684_,
		_w2421_,
		_w3857_
	);
	LUT2 #(
		.INIT('h2)
	) name2899 (
		_w1283_,
		_w3857_,
		_w3858_
	);
	LUT2 #(
		.INIT('h8)
	) name2900 (
		\u7_mc_br_r_reg/P0001 ,
		_w1168_,
		_w3859_
	);
	LUT2 #(
		.INIT('h4)
	) name2901 (
		_w1206_,
		_w1749_,
		_w3860_
	);
	LUT2 #(
		.INIT('h8)
	) name2902 (
		_w2940_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h8)
	) name2903 (
		_w1297_,
		_w2939_,
		_w3862_
	);
	LUT2 #(
		.INIT('h4)
	) name2904 (
		_w3859_,
		_w3862_,
		_w3863_
	);
	LUT2 #(
		.INIT('h8)
	) name2905 (
		_w3861_,
		_w3863_,
		_w3864_
	);
	LUT2 #(
		.INIT('h2)
	) name2906 (
		_w2951_,
		_w3858_,
		_w3865_
	);
	LUT2 #(
		.INIT('h8)
	) name2907 (
		_w3864_,
		_w3865_,
		_w3866_
	);
	LUT2 #(
		.INIT('h8)
	) name2908 (
		_w2947_,
		_w3866_,
		_w3867_
	);
	LUT2 #(
		.INIT('h8)
	) name2909 (
		_w2944_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		\wb_addr_i[8]_pad ,
		_w2606_,
		_w3869_
	);
	LUT2 #(
		.INIT('h8)
	) name2911 (
		\wb_addr_i[9]_pad ,
		_w2878_,
		_w3870_
	);
	LUT2 #(
		.INIT('h8)
	) name2912 (
		\wb_addr_i[7]_pad ,
		_w2388_,
		_w3871_
	);
	LUT2 #(
		.INIT('h1)
	) name2913 (
		_w3869_,
		_w3870_,
		_w3872_
	);
	LUT2 #(
		.INIT('h4)
	) name2914 (
		_w3871_,
		_w3872_,
		_w3873_
	);
	LUT2 #(
		.INIT('h1)
	) name2915 (
		_w2858_,
		_w3873_,
		_w3874_
	);
	LUT2 #(
		.INIT('h1)
	) name2916 (
		\u1_acs_addr_reg[7]/P0001 ,
		_w2861_,
		_w3875_
	);
	LUT2 #(
		.INIT('h4)
	) name2917 (
		\u1_u0_out_r_reg[7]/P0001 ,
		_w2861_,
		_w3876_
	);
	LUT2 #(
		.INIT('h2)
	) name2918 (
		_w2858_,
		_w3875_,
		_w3877_
	);
	LUT2 #(
		.INIT('h4)
	) name2919 (
		_w3876_,
		_w3877_,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name2920 (
		_w3874_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h4)
	) name2921 (
		\u5_state_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w3880_
	);
	LUT2 #(
		.INIT('h1)
	) name2922 (
		_w1382_,
		_w1870_,
		_w3881_
	);
	LUT2 #(
		.INIT('h8)
	) name2923 (
		_w1686_,
		_w2678_,
		_w3882_
	);
	LUT2 #(
		.INIT('h2)
	) name2924 (
		_w1366_,
		_w3882_,
		_w3883_
	);
	LUT2 #(
		.INIT('h1)
	) name2925 (
		_w3881_,
		_w3883_,
		_w3884_
	);
	LUT2 #(
		.INIT('h1)
	) name2926 (
		_w3880_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h2)
	) name2927 (
		\u0_csr_r_reg[8]/NET0131 ,
		\u4_rfr_cnt_reg[1]/NET0131 ,
		_w3886_
	);
	LUT2 #(
		.INIT('h1)
	) name2928 (
		\u0_csr_r_reg[10]/NET0131 ,
		\u0_csr_r_reg[9]/NET0131 ,
		_w3887_
	);
	LUT2 #(
		.INIT('h4)
	) name2929 (
		_w3886_,
		_w3887_,
		_w3888_
	);
	LUT2 #(
		.INIT('h2)
	) name2930 (
		\u0_csr_r_reg[8]/NET0131 ,
		\u4_rfr_cnt_reg[3]/NET0131 ,
		_w3889_
	);
	LUT2 #(
		.INIT('h1)
	) name2931 (
		\u0_csr_r_reg[10]/NET0131 ,
		_w3889_,
		_w3890_
	);
	LUT2 #(
		.INIT('h2)
	) name2932 (
		\u0_csr_r_reg[8]/NET0131 ,
		\u4_rfr_cnt_reg[5]/NET0131 ,
		_w3891_
	);
	LUT2 #(
		.INIT('h1)
	) name2933 (
		\u0_csr_r_reg[9]/NET0131 ,
		_w3891_,
		_w3892_
	);
	LUT2 #(
		.INIT('h2)
	) name2934 (
		\u0_csr_r_reg[8]/NET0131 ,
		\u4_rfr_cnt_reg[7]/NET0131 ,
		_w3893_
	);
	LUT2 #(
		.INIT('h8)
	) name2935 (
		\u4_rfr_cnt_reg[5]/NET0131 ,
		\u4_rfr_cnt_reg[6]/NET0131 ,
		_w3894_
	);
	LUT2 #(
		.INIT('h4)
	) name2936 (
		_w3893_,
		_w3894_,
		_w3895_
	);
	LUT2 #(
		.INIT('h1)
	) name2937 (
		_w3892_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h8)
	) name2938 (
		\u4_rfr_cnt_reg[3]/NET0131 ,
		\u4_rfr_cnt_reg[4]/NET0131 ,
		_w3897_
	);
	LUT2 #(
		.INIT('h4)
	) name2939 (
		_w3896_,
		_w3897_,
		_w3898_
	);
	LUT2 #(
		.INIT('h1)
	) name2940 (
		_w3890_,
		_w3898_,
		_w3899_
	);
	LUT2 #(
		.INIT('h8)
	) name2941 (
		\u4_rfr_cnt_reg[1]/NET0131 ,
		\u4_rfr_cnt_reg[2]/NET0131 ,
		_w3900_
	);
	LUT2 #(
		.INIT('h4)
	) name2942 (
		_w3899_,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h1)
	) name2943 (
		_w3888_,
		_w3901_,
		_w3902_
	);
	LUT2 #(
		.INIT('h8)
	) name2944 (
		\u4_rfr_cnt_reg[0]/NET0131 ,
		\u4_rfr_early_reg/NET0131 ,
		_w3903_
	);
	LUT2 #(
		.INIT('h4)
	) name2945 (
		_w3902_,
		_w3903_,
		_w3904_
	);
	LUT2 #(
		.INIT('h8)
	) name2946 (
		\wb_addr_i[12]_pad ,
		_w2388_,
		_w3905_
	);
	LUT2 #(
		.INIT('h8)
	) name2947 (
		\wb_addr_i[14]_pad ,
		_w2878_,
		_w3906_
	);
	LUT2 #(
		.INIT('h8)
	) name2948 (
		\wb_addr_i[13]_pad ,
		_w2606_,
		_w3907_
	);
	LUT2 #(
		.INIT('h1)
	) name2949 (
		_w3905_,
		_w3906_,
		_w3908_
	);
	LUT2 #(
		.INIT('h4)
	) name2950 (
		_w3907_,
		_w3908_,
		_w3909_
	);
	LUT2 #(
		.INIT('h1)
	) name2951 (
		_w2858_,
		_w3909_,
		_w3910_
	);
	LUT2 #(
		.INIT('h1)
	) name2952 (
		\u1_acs_addr_reg[12]/P0001 ,
		_w2862_,
		_w3911_
	);
	LUT2 #(
		.INIT('h2)
	) name2953 (
		_w2858_,
		_w2863_,
		_w3912_
	);
	LUT2 #(
		.INIT('h4)
	) name2954 (
		_w3911_,
		_w3912_,
		_w3913_
	);
	LUT2 #(
		.INIT('h1)
	) name2955 (
		_w3910_,
		_w3913_,
		_w3914_
	);
	LUT2 #(
		.INIT('h1)
	) name2956 (
		_w1044_,
		_w1877_,
		_w3915_
	);
	LUT2 #(
		.INIT('h8)
	) name2957 (
		_w1044_,
		_w1877_,
		_w3916_
	);
	LUT2 #(
		.INIT('h1)
	) name2958 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		_w3916_,
		_w3917_
	);
	LUT2 #(
		.INIT('h4)
	) name2959 (
		_w3915_,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w3915_,
		_w3916_,
		_w3919_
	);
	LUT2 #(
		.INIT('h2)
	) name2961 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('h1)
	) name2962 (
		\u5_no_wb_cycle_reg/NET0131 ,
		_w3918_,
		_w3921_
	);
	LUT2 #(
		.INIT('h4)
	) name2963 (
		_w3920_,
		_w3921_,
		_w3922_
	);
	LUT2 #(
		.INIT('h1)
	) name2964 (
		_w3915_,
		_w3917_,
		_w3923_
	);
	LUT2 #(
		.INIT('h8)
	) name2965 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_ack_cnt_reg[1]/NET0131 ,
		_w3924_
	);
	LUT2 #(
		.INIT('h1)
	) name2966 (
		_w1871_,
		_w3924_,
		_w3925_
	);
	LUT2 #(
		.INIT('h1)
	) name2967 (
		_w3923_,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('h8)
	) name2968 (
		_w3923_,
		_w3925_,
		_w3927_
	);
	LUT2 #(
		.INIT('h1)
	) name2969 (
		\u5_no_wb_cycle_reg/NET0131 ,
		_w3926_,
		_w3928_
	);
	LUT2 #(
		.INIT('h4)
	) name2970 (
		_w3927_,
		_w3928_,
		_w3929_
	);
	LUT2 #(
		.INIT('h1)
	) name2971 (
		\u5_ack_cnt_reg[2]/NET0131 ,
		_w3924_,
		_w3930_
	);
	LUT2 #(
		.INIT('h8)
	) name2972 (
		\u5_ack_cnt_reg[2]/NET0131 ,
		_w3924_,
		_w3931_
	);
	LUT2 #(
		.INIT('h1)
	) name2973 (
		_w3930_,
		_w3931_,
		_w3932_
	);
	LUT2 #(
		.INIT('h2)
	) name2974 (
		_w3915_,
		_w3932_,
		_w3933_
	);
	LUT2 #(
		.INIT('h8)
	) name2975 (
		_w1871_,
		_w3916_,
		_w3934_
	);
	LUT2 #(
		.INIT('h2)
	) name2976 (
		\u5_ack_cnt_reg[2]/NET0131 ,
		_w3934_,
		_w3935_
	);
	LUT2 #(
		.INIT('h8)
	) name2977 (
		_w1872_,
		_w3916_,
		_w3936_
	);
	LUT2 #(
		.INIT('h1)
	) name2978 (
		_w3915_,
		_w3936_,
		_w3937_
	);
	LUT2 #(
		.INIT('h4)
	) name2979 (
		_w3935_,
		_w3937_,
		_w3938_
	);
	LUT2 #(
		.INIT('h1)
	) name2980 (
		\u5_no_wb_cycle_reg/NET0131 ,
		_w3933_,
		_w3939_
	);
	LUT2 #(
		.INIT('h4)
	) name2981 (
		_w3938_,
		_w3939_,
		_w3940_
	);
	LUT2 #(
		.INIT('h8)
	) name2982 (
		_w1873_,
		_w3916_,
		_w3941_
	);
	LUT2 #(
		.INIT('h2)
	) name2983 (
		\u5_ack_cnt_reg[3]/NET0131 ,
		_w3936_,
		_w3942_
	);
	LUT2 #(
		.INIT('h1)
	) name2984 (
		_w3915_,
		_w3941_,
		_w3943_
	);
	LUT2 #(
		.INIT('h4)
	) name2985 (
		_w3942_,
		_w3943_,
		_w3944_
	);
	LUT2 #(
		.INIT('h2)
	) name2986 (
		\u5_ack_cnt_reg[3]/NET0131 ,
		_w3931_,
		_w3945_
	);
	LUT2 #(
		.INIT('h4)
	) name2987 (
		\u5_ack_cnt_reg[3]/NET0131 ,
		_w3931_,
		_w3946_
	);
	LUT2 #(
		.INIT('h1)
	) name2988 (
		_w3945_,
		_w3946_,
		_w3947_
	);
	LUT2 #(
		.INIT('h8)
	) name2989 (
		_w3915_,
		_w3947_,
		_w3948_
	);
	LUT2 #(
		.INIT('h1)
	) name2990 (
		\u5_no_wb_cycle_reg/NET0131 ,
		_w3948_,
		_w3949_
	);
	LUT2 #(
		.INIT('h4)
	) name2991 (
		_w3944_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('h8)
	) name2992 (
		\wb_addr_i[5]_pad ,
		_w2606_,
		_w3951_
	);
	LUT2 #(
		.INIT('h8)
	) name2993 (
		\wb_addr_i[6]_pad ,
		_w2878_,
		_w3952_
	);
	LUT2 #(
		.INIT('h8)
	) name2994 (
		\wb_addr_i[4]_pad ,
		_w2388_,
		_w3953_
	);
	LUT2 #(
		.INIT('h1)
	) name2995 (
		_w3951_,
		_w3952_,
		_w3954_
	);
	LUT2 #(
		.INIT('h4)
	) name2996 (
		_w3953_,
		_w3954_,
		_w3955_
	);
	LUT2 #(
		.INIT('h1)
	) name2997 (
		_w2858_,
		_w3955_,
		_w3956_
	);
	LUT2 #(
		.INIT('h1)
	) name2998 (
		\u1_acs_addr_reg[4]/P0001 ,
		_w2861_,
		_w3957_
	);
	LUT2 #(
		.INIT('h4)
	) name2999 (
		\u1_u0_out_r_reg[4]/P0001 ,
		_w2861_,
		_w3958_
	);
	LUT2 #(
		.INIT('h2)
	) name3000 (
		_w2858_,
		_w3957_,
		_w3959_
	);
	LUT2 #(
		.INIT('h4)
	) name3001 (
		_w3958_,
		_w3959_,
		_w3960_
	);
	LUT2 #(
		.INIT('h1)
	) name3002 (
		_w3956_,
		_w3960_,
		_w3961_
	);
	LUT2 #(
		.INIT('h1)
	) name3003 (
		\u1_acs_addr_reg[8]/P0001 ,
		_w2861_,
		_w3962_
	);
	LUT2 #(
		.INIT('h4)
	) name3004 (
		\u1_u0_out_r_reg[8]/P0001 ,
		_w2861_,
		_w3963_
	);
	LUT2 #(
		.INIT('h2)
	) name3005 (
		_w2858_,
		_w3962_,
		_w3964_
	);
	LUT2 #(
		.INIT('h4)
	) name3006 (
		_w3963_,
		_w3964_,
		_w3965_
	);
	LUT2 #(
		.INIT('h8)
	) name3007 (
		\wb_addr_i[9]_pad ,
		_w2606_,
		_w3966_
	);
	LUT2 #(
		.INIT('h8)
	) name3008 (
		\wb_addr_i[10]_pad ,
		_w2878_,
		_w3967_
	);
	LUT2 #(
		.INIT('h8)
	) name3009 (
		\wb_addr_i[8]_pad ,
		_w2388_,
		_w3968_
	);
	LUT2 #(
		.INIT('h1)
	) name3010 (
		_w3966_,
		_w3967_,
		_w3969_
	);
	LUT2 #(
		.INIT('h4)
	) name3011 (
		_w3968_,
		_w3969_,
		_w3970_
	);
	LUT2 #(
		.INIT('h1)
	) name3012 (
		_w2858_,
		_w3970_,
		_w3971_
	);
	LUT2 #(
		.INIT('h1)
	) name3013 (
		_w3965_,
		_w3971_,
		_w3972_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		_w3026_,
		_w3146_,
		_w3973_
	);
	LUT2 #(
		.INIT('h2)
	) name3015 (
		_w2358_,
		_w3973_,
		_w3974_
	);
	LUT2 #(
		.INIT('h2)
	) name3016 (
		_w2354_,
		_w2357_,
		_w3975_
	);
	LUT2 #(
		.INIT('h4)
	) name3017 (
		_w2354_,
		_w2357_,
		_w3976_
	);
	LUT2 #(
		.INIT('h1)
	) name3018 (
		_w3975_,
		_w3976_,
		_w3977_
	);
	LUT2 #(
		.INIT('h1)
	) name3019 (
		_w2970_,
		_w3814_,
		_w3978_
	);
	LUT2 #(
		.INIT('h1)
	) name3020 (
		_w3977_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('h1)
	) name3021 (
		_w2354_,
		_w2357_,
		_w3980_
	);
	LUT2 #(
		.INIT('h2)
	) name3022 (
		_w3848_,
		_w3980_,
		_w3981_
	);
	LUT2 #(
		.INIT('h1)
	) name3023 (
		_w3974_,
		_w3981_,
		_w3982_
	);
	LUT2 #(
		.INIT('h4)
	) name3024 (
		_w3979_,
		_w3982_,
		_w3983_
	);
	LUT2 #(
		.INIT('h2)
	) name3025 (
		\u0_sp_csc_reg[9]/NET0131 ,
		_w1051_,
		_w3984_
	);
	LUT2 #(
		.INIT('h8)
	) name3026 (
		\u0_csc_reg[9]/NET0131 ,
		_w1051_,
		_w3985_
	);
	LUT2 #(
		.INIT('h1)
	) name3027 (
		_w3984_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h2)
	) name3028 (
		_w3983_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h8)
	) name3029 (
		_w2358_,
		_w2972_,
		_w3988_
	);
	LUT2 #(
		.INIT('h8)
	) name3030 (
		_w2358_,
		_w3025_,
		_w3989_
	);
	LUT2 #(
		.INIT('h2)
	) name3031 (
		\wb_addr_i[23]_pad ,
		_w3977_,
		_w3990_
	);
	LUT2 #(
		.INIT('h8)
	) name3032 (
		\wb_addr_i[22]_pad ,
		_w2358_,
		_w3991_
	);
	LUT2 #(
		.INIT('h1)
	) name3033 (
		_w3990_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h2)
	) name3034 (
		_w2388_,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h1)
	) name3035 (
		_w2972_,
		_w3816_,
		_w3994_
	);
	LUT2 #(
		.INIT('h1)
	) name3036 (
		_w3977_,
		_w3994_,
		_w3995_
	);
	LUT2 #(
		.INIT('h1)
	) name3037 (
		_w3989_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h4)
	) name3038 (
		_w3993_,
		_w3996_,
		_w3997_
	);
	LUT2 #(
		.INIT('h2)
	) name3039 (
		_w3986_,
		_w3988_,
		_w3998_
	);
	LUT2 #(
		.INIT('h8)
	) name3040 (
		_w3997_,
		_w3998_,
		_w3999_
	);
	LUT2 #(
		.INIT('h1)
	) name3041 (
		_w3987_,
		_w3999_,
		_w4000_
	);
	LUT2 #(
		.INIT('h8)
	) name3042 (
		\u1_acs_addr_reg[0]/P0001 ,
		\u1_acs_addr_reg[1]/P0001 ,
		_w4001_
	);
	LUT2 #(
		.INIT('h8)
	) name3043 (
		\u1_acs_addr_reg[2]/P0001 ,
		_w4001_,
		_w4002_
	);
	LUT2 #(
		.INIT('h8)
	) name3044 (
		\u1_acs_addr_reg[3]/P0001 ,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('h8)
	) name3045 (
		\u1_acs_addr_reg[4]/P0001 ,
		_w4003_,
		_w4004_
	);
	LUT2 #(
		.INIT('h8)
	) name3046 (
		\u1_acs_addr_reg[5]/P0001 ,
		_w4004_,
		_w4005_
	);
	LUT2 #(
		.INIT('h8)
	) name3047 (
		\u1_acs_addr_reg[6]/P0001 ,
		_w4005_,
		_w4006_
	);
	LUT2 #(
		.INIT('h8)
	) name3048 (
		\u1_acs_addr_reg[7]/P0001 ,
		_w4006_,
		_w4007_
	);
	LUT2 #(
		.INIT('h8)
	) name3049 (
		\u1_acs_addr_reg[8]/P0001 ,
		_w4007_,
		_w4008_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		\u1_acs_addr_reg[9]/P0001 ,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h8)
	) name3051 (
		\u1_acs_addr_reg[10]/P0001 ,
		_w4009_,
		_w4010_
	);
	LUT2 #(
		.INIT('h8)
	) name3052 (
		\u1_acs_addr_reg[11]/P0001 ,
		_w4010_,
		_w4011_
	);
	LUT2 #(
		.INIT('h1)
	) name3053 (
		\u1_acs_addr_reg[11]/P0001 ,
		_w4010_,
		_w4012_
	);
	LUT2 #(
		.INIT('h1)
	) name3054 (
		_w4011_,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('h2)
	) name3055 (
		_w3967_,
		_w3980_,
		_w4014_
	);
	LUT2 #(
		.INIT('h8)
	) name3056 (
		\wb_addr_i[11]_pad ,
		_w2606_,
		_w4015_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		_w3905_,
		_w4015_,
		_w4016_
	);
	LUT2 #(
		.INIT('h1)
	) name3058 (
		_w3977_,
		_w4016_,
		_w4017_
	);
	LUT2 #(
		.INIT('h8)
	) name3059 (
		\wb_addr_i[10]_pad ,
		_w2606_,
		_w4018_
	);
	LUT2 #(
		.INIT('h1)
	) name3060 (
		_w3840_,
		_w4018_,
		_w4019_
	);
	LUT2 #(
		.INIT('h2)
	) name3061 (
		_w2358_,
		_w4019_,
		_w4020_
	);
	LUT2 #(
		.INIT('h1)
	) name3062 (
		_w4014_,
		_w4017_,
		_w4021_
	);
	LUT2 #(
		.INIT('h4)
	) name3063 (
		_w4020_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h2)
	) name3064 (
		_w3986_,
		_w4022_,
		_w4023_
	);
	LUT2 #(
		.INIT('h1)
	) name3065 (
		_w2881_,
		_w3816_,
		_w4024_
	);
	LUT2 #(
		.INIT('h2)
	) name3066 (
		_w2358_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h8)
	) name3067 (
		\wb_addr_i[24]_pad ,
		_w2388_,
		_w4026_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		_w2982_,
		_w4026_,
		_w4027_
	);
	LUT2 #(
		.INIT('h2)
	) name3069 (
		_w3975_,
		_w4027_,
		_w4028_
	);
	LUT2 #(
		.INIT('h1)
	) name3070 (
		_w4025_,
		_w4028_,
		_w4029_
	);
	LUT2 #(
		.INIT('h8)
	) name3071 (
		_w3024_,
		_w3975_,
		_w4030_
	);
	LUT2 #(
		.INIT('h8)
	) name3072 (
		\wb_addr_i[25]_pad ,
		_w2388_,
		_w4031_
	);
	LUT2 #(
		.INIT('h1)
	) name3073 (
		_w2880_,
		_w3815_,
		_w4032_
	);
	LUT2 #(
		.INIT('h4)
	) name3074 (
		_w4031_,
		_w4032_,
		_w4033_
	);
	LUT2 #(
		.INIT('h2)
	) name3075 (
		_w3976_,
		_w4033_,
		_w4034_
	);
	LUT2 #(
		.INIT('h1)
	) name3076 (
		_w3988_,
		_w4030_,
		_w4035_
	);
	LUT2 #(
		.INIT('h8)
	) name3077 (
		_w4029_,
		_w4035_,
		_w4036_
	);
	LUT2 #(
		.INIT('h4)
	) name3078 (
		_w4034_,
		_w4036_,
		_w4037_
	);
	LUT2 #(
		.INIT('h1)
	) name3079 (
		_w3986_,
		_w4037_,
		_w4038_
	);
	LUT2 #(
		.INIT('h1)
	) name3080 (
		_w4023_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h2)
	) name3081 (
		_w2358_,
		_w4016_,
		_w4040_
	);
	LUT2 #(
		.INIT('h1)
	) name3082 (
		_w3826_,
		_w3841_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name3083 (
		_w3977_,
		_w4041_,
		_w4042_
	);
	LUT2 #(
		.INIT('h8)
	) name3084 (
		\wb_addr_i[11]_pad ,
		_w2878_,
		_w4043_
	);
	LUT2 #(
		.INIT('h4)
	) name3085 (
		_w3980_,
		_w4043_,
		_w4044_
	);
	LUT2 #(
		.INIT('h1)
	) name3086 (
		_w4040_,
		_w4044_,
		_w4045_
	);
	LUT2 #(
		.INIT('h4)
	) name3087 (
		_w4042_,
		_w4045_,
		_w4046_
	);
	LUT2 #(
		.INIT('h2)
	) name3088 (
		_w3986_,
		_w4046_,
		_w4047_
	);
	LUT2 #(
		.INIT('h8)
	) name3089 (
		_w2358_,
		_w2982_,
		_w4048_
	);
	LUT2 #(
		.INIT('h2)
	) name3090 (
		_w3975_,
		_w4033_,
		_w4049_
	);
	LUT2 #(
		.INIT('h1)
	) name3091 (
		_w4048_,
		_w4049_,
		_w4050_
	);
	LUT2 #(
		.INIT('h1)
	) name3092 (
		_w3024_,
		_w4026_,
		_w4051_
	);
	LUT2 #(
		.INIT('h2)
	) name3093 (
		_w2358_,
		_w4051_,
		_w4052_
	);
	LUT2 #(
		.INIT('h8)
	) name3094 (
		\wb_addr_i[26]_pad ,
		_w2388_,
		_w4053_
	);
	LUT2 #(
		.INIT('h8)
	) name3095 (
		\wb_addr_i[25]_pad ,
		_w2606_,
		_w4054_
	);
	LUT2 #(
		.INIT('h1)
	) name3096 (
		_w2981_,
		_w4053_,
		_w4055_
	);
	LUT2 #(
		.INIT('h4)
	) name3097 (
		_w4054_,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h2)
	) name3098 (
		_w3976_,
		_w4056_,
		_w4057_
	);
	LUT2 #(
		.INIT('h1)
	) name3099 (
		_w4052_,
		_w4057_,
		_w4058_
	);
	LUT2 #(
		.INIT('h8)
	) name3100 (
		_w4050_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h1)
	) name3101 (
		_w3986_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h1)
	) name3102 (
		_w4047_,
		_w4060_,
		_w4061_
	);
	LUT2 #(
		.INIT('h2)
	) name3103 (
		_w2358_,
		_w4041_,
		_w4062_
	);
	LUT2 #(
		.INIT('h1)
	) name3104 (
		_w3786_,
		_w3907_,
		_w4063_
	);
	LUT2 #(
		.INIT('h1)
	) name3105 (
		_w3977_,
		_w4063_,
		_w4064_
	);
	LUT2 #(
		.INIT('h8)
	) name3106 (
		\wb_addr_i[12]_pad ,
		_w2878_,
		_w4065_
	);
	LUT2 #(
		.INIT('h4)
	) name3107 (
		_w3980_,
		_w4065_,
		_w4066_
	);
	LUT2 #(
		.INIT('h1)
	) name3108 (
		_w4062_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h4)
	) name3109 (
		_w4064_,
		_w4067_,
		_w4068_
	);
	LUT2 #(
		.INIT('h2)
	) name3110 (
		_w3986_,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('h1)
	) name3111 (
		_w3986_,
		_w4022_,
		_w4070_
	);
	LUT2 #(
		.INIT('h1)
	) name3112 (
		_w4069_,
		_w4070_,
		_w4071_
	);
	LUT2 #(
		.INIT('h2)
	) name3113 (
		_w3145_,
		_w3980_,
		_w4072_
	);
	LUT2 #(
		.INIT('h2)
	) name3114 (
		_w2358_,
		_w3978_,
		_w4073_
	);
	LUT2 #(
		.INIT('h1)
	) name3115 (
		_w2980_,
		_w3025_,
		_w4074_
	);
	LUT2 #(
		.INIT('h1)
	) name3116 (
		_w3977_,
		_w4074_,
		_w4075_
	);
	LUT2 #(
		.INIT('h1)
	) name3117 (
		_w4072_,
		_w4073_,
		_w4076_
	);
	LUT2 #(
		.INIT('h4)
	) name3118 (
		_w4075_,
		_w4076_,
		_w4077_
	);
	LUT2 #(
		.INIT('h1)
	) name3119 (
		_w3986_,
		_w4077_,
		_w4078_
	);
	LUT2 #(
		.INIT('h8)
	) name3120 (
		_w2354_,
		_w3024_,
		_w4079_
	);
	LUT2 #(
		.INIT('h4)
	) name3121 (
		_w3024_,
		_w4027_,
		_w4080_
	);
	LUT2 #(
		.INIT('h2)
	) name3122 (
		_w3976_,
		_w4080_,
		_w4081_
	);
	LUT2 #(
		.INIT('h2)
	) name3123 (
		_w4029_,
		_w4079_,
		_w4082_
	);
	LUT2 #(
		.INIT('h4)
	) name3124 (
		_w4081_,
		_w4082_,
		_w4083_
	);
	LUT2 #(
		.INIT('h2)
	) name3125 (
		_w3986_,
		_w4083_,
		_w4084_
	);
	LUT2 #(
		.INIT('h1)
	) name3126 (
		_w4078_,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h2)
	) name3127 (
		_w2358_,
		_w4063_,
		_w4086_
	);
	LUT2 #(
		.INIT('h1)
	) name3128 (
		_w3650_,
		_w3828_,
		_w4087_
	);
	LUT2 #(
		.INIT('h1)
	) name3129 (
		_w3977_,
		_w4087_,
		_w4088_
	);
	LUT2 #(
		.INIT('h2)
	) name3130 (
		_w3842_,
		_w3980_,
		_w4089_
	);
	LUT2 #(
		.INIT('h1)
	) name3131 (
		_w4086_,
		_w4089_,
		_w4090_
	);
	LUT2 #(
		.INIT('h4)
	) name3132 (
		_w4088_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h2)
	) name3133 (
		_w3986_,
		_w4091_,
		_w4092_
	);
	LUT2 #(
		.INIT('h1)
	) name3134 (
		_w3986_,
		_w4046_,
		_w4093_
	);
	LUT2 #(
		.INIT('h1)
	) name3135 (
		_w4092_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h2)
	) name3136 (
		_w2358_,
		_w4087_,
		_w4095_
	);
	LUT2 #(
		.INIT('h1)
	) name3137 (
		_w3126_,
		_w3788_,
		_w4096_
	);
	LUT2 #(
		.INIT('h1)
	) name3138 (
		_w3977_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h2)
	) name3139 (
		_w3906_,
		_w3980_,
		_w4098_
	);
	LUT2 #(
		.INIT('h1)
	) name3140 (
		_w4095_,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h4)
	) name3141 (
		_w4097_,
		_w4099_,
		_w4100_
	);
	LUT2 #(
		.INIT('h2)
	) name3142 (
		_w3986_,
		_w4100_,
		_w4101_
	);
	LUT2 #(
		.INIT('h1)
	) name3143 (
		_w3986_,
		_w4068_,
		_w4102_
	);
	LUT2 #(
		.INIT('h1)
	) name3144 (
		_w4101_,
		_w4102_,
		_w4103_
	);
	LUT2 #(
		.INIT('h2)
	) name3145 (
		_w2358_,
		_w4096_,
		_w4104_
	);
	LUT2 #(
		.INIT('h1)
	) name3146 (
		_w3652_,
		_w3847_,
		_w4105_
	);
	LUT2 #(
		.INIT('h1)
	) name3147 (
		_w3977_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h2)
	) name3148 (
		_w3827_,
		_w3980_,
		_w4107_
	);
	LUT2 #(
		.INIT('h1)
	) name3149 (
		_w4104_,
		_w4107_,
		_w4108_
	);
	LUT2 #(
		.INIT('h4)
	) name3150 (
		_w4106_,
		_w4108_,
		_w4109_
	);
	LUT2 #(
		.INIT('h2)
	) name3151 (
		_w3986_,
		_w4109_,
		_w4110_
	);
	LUT2 #(
		.INIT('h1)
	) name3152 (
		_w3986_,
		_w4091_,
		_w4111_
	);
	LUT2 #(
		.INIT('h1)
	) name3153 (
		_w4110_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h2)
	) name3154 (
		_w2358_,
		_w4105_,
		_w4113_
	);
	LUT2 #(
		.INIT('h1)
	) name3155 (
		_w3128_,
		_w3144_,
		_w4114_
	);
	LUT2 #(
		.INIT('h1)
	) name3156 (
		_w3977_,
		_w4114_,
		_w4115_
	);
	LUT2 #(
		.INIT('h2)
	) name3157 (
		_w3787_,
		_w3980_,
		_w4116_
	);
	LUT2 #(
		.INIT('h1)
	) name3158 (
		_w4113_,
		_w4116_,
		_w4117_
	);
	LUT2 #(
		.INIT('h4)
	) name3159 (
		_w4115_,
		_w4117_,
		_w4118_
	);
	LUT2 #(
		.INIT('h2)
	) name3160 (
		_w3986_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h1)
	) name3161 (
		_w3986_,
		_w4100_,
		_w4120_
	);
	LUT2 #(
		.INIT('h1)
	) name3162 (
		_w4119_,
		_w4120_,
		_w4121_
	);
	LUT2 #(
		.INIT('h2)
	) name3163 (
		_w2358_,
		_w4114_,
		_w4122_
	);
	LUT2 #(
		.INIT('h1)
	) name3164 (
		_w2971_,
		_w3849_,
		_w4123_
	);
	LUT2 #(
		.INIT('h1)
	) name3165 (
		_w3977_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h2)
	) name3166 (
		_w3651_,
		_w3980_,
		_w4125_
	);
	LUT2 #(
		.INIT('h1)
	) name3167 (
		_w4122_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h4)
	) name3168 (
		_w4124_,
		_w4126_,
		_w4127_
	);
	LUT2 #(
		.INIT('h2)
	) name3169 (
		_w3986_,
		_w4127_,
		_w4128_
	);
	LUT2 #(
		.INIT('h1)
	) name3170 (
		_w3986_,
		_w4109_,
		_w4129_
	);
	LUT2 #(
		.INIT('h1)
	) name3171 (
		_w4128_,
		_w4129_,
		_w4130_
	);
	LUT2 #(
		.INIT('h2)
	) name3172 (
		_w2358_,
		_w4123_,
		_w4131_
	);
	LUT2 #(
		.INIT('h1)
	) name3173 (
		_w3973_,
		_w3977_,
		_w4132_
	);
	LUT2 #(
		.INIT('h2)
	) name3174 (
		_w3127_,
		_w3980_,
		_w4133_
	);
	LUT2 #(
		.INIT('h1)
	) name3175 (
		_w4131_,
		_w4133_,
		_w4134_
	);
	LUT2 #(
		.INIT('h4)
	) name3176 (
		_w4132_,
		_w4134_,
		_w4135_
	);
	LUT2 #(
		.INIT('h2)
	) name3177 (
		_w3986_,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h1)
	) name3178 (
		_w3986_,
		_w4118_,
		_w4137_
	);
	LUT2 #(
		.INIT('h1)
	) name3179 (
		_w4136_,
		_w4137_,
		_w4138_
	);
	LUT2 #(
		.INIT('h4)
	) name3180 (
		_w3986_,
		_w4127_,
		_w4139_
	);
	LUT2 #(
		.INIT('h8)
	) name3181 (
		_w3983_,
		_w3986_,
		_w4140_
	);
	LUT2 #(
		.INIT('h1)
	) name3182 (
		_w4139_,
		_w4140_,
		_w4141_
	);
	LUT2 #(
		.INIT('h1)
	) name3183 (
		_w3986_,
		_w4135_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name3184 (
		_w3986_,
		_w4077_,
		_w4143_
	);
	LUT2 #(
		.INIT('h1)
	) name3185 (
		_w4142_,
		_w4143_,
		_w4144_
	);
	LUT2 #(
		.INIT('h1)
	) name3186 (
		_w3986_,
		_w3997_,
		_w4145_
	);
	LUT2 #(
		.INIT('h8)
	) name3187 (
		_w2358_,
		_w4026_,
		_w4146_
	);
	LUT2 #(
		.INIT('h1)
	) name3188 (
		_w4034_,
		_w4146_,
		_w4147_
	);
	LUT2 #(
		.INIT('h8)
	) name3189 (
		_w4050_,
		_w4147_,
		_w4148_
	);
	LUT2 #(
		.INIT('h2)
	) name3190 (
		_w3986_,
		_w4148_,
		_w4149_
	);
	LUT2 #(
		.INIT('h1)
	) name3191 (
		_w4145_,
		_w4149_,
		_w4150_
	);
	LUT2 #(
		.INIT('h1)
	) name3192 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		_w4151_
	);
	LUT2 #(
		.INIT('h8)
	) name3193 (
		\u5_pack_le1_reg/P0001 ,
		_w4151_,
		_w4152_
	);
	LUT2 #(
		.INIT('h2)
	) name3194 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		_w4153_
	);
	LUT2 #(
		.INIT('h8)
	) name3195 (
		\u5_pack_le0_reg/P0001 ,
		_w4153_,
		_w4154_
	);
	LUT2 #(
		.INIT('h2)
	) name3196 (
		\u3_byte1_reg[0]/P0001 ,
		_w4154_,
		_w4155_
	);
	LUT2 #(
		.INIT('h8)
	) name3197 (
		\u7_mc_data_ir_reg[8]/P0001 ,
		_w4154_,
		_w4156_
	);
	LUT2 #(
		.INIT('h1)
	) name3198 (
		_w4155_,
		_w4156_,
		_w4157_
	);
	LUT2 #(
		.INIT('h1)
	) name3199 (
		_w4152_,
		_w4157_,
		_w4158_
	);
	LUT2 #(
		.INIT('h8)
	) name3200 (
		\u7_mc_data_ir_reg[0]/P0001 ,
		_w4152_,
		_w4159_
	);
	LUT2 #(
		.INIT('h1)
	) name3201 (
		_w4158_,
		_w4159_,
		_w4160_
	);
	LUT2 #(
		.INIT('h2)
	) name3202 (
		\u3_byte1_reg[2]/P0001 ,
		_w4154_,
		_w4161_
	);
	LUT2 #(
		.INIT('h8)
	) name3203 (
		\u7_mc_data_ir_reg[10]/P0001 ,
		_w4154_,
		_w4162_
	);
	LUT2 #(
		.INIT('h1)
	) name3204 (
		_w4161_,
		_w4162_,
		_w4163_
	);
	LUT2 #(
		.INIT('h1)
	) name3205 (
		_w4152_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h8)
	) name3206 (
		\u7_mc_data_ir_reg[2]/P0001 ,
		_w4152_,
		_w4165_
	);
	LUT2 #(
		.INIT('h1)
	) name3207 (
		_w4164_,
		_w4165_,
		_w4166_
	);
	LUT2 #(
		.INIT('h2)
	) name3208 (
		\u3_byte1_reg[1]/P0001 ,
		_w4154_,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name3209 (
		\u7_mc_data_ir_reg[9]/P0001 ,
		_w4154_,
		_w4168_
	);
	LUT2 #(
		.INIT('h1)
	) name3210 (
		_w4167_,
		_w4168_,
		_w4169_
	);
	LUT2 #(
		.INIT('h1)
	) name3211 (
		_w4152_,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h8)
	) name3212 (
		\u7_mc_data_ir_reg[1]/P0001 ,
		_w4152_,
		_w4171_
	);
	LUT2 #(
		.INIT('h1)
	) name3213 (
		_w4170_,
		_w4171_,
		_w4172_
	);
	LUT2 #(
		.INIT('h2)
	) name3214 (
		\u3_byte1_reg[3]/P0001 ,
		_w4154_,
		_w4173_
	);
	LUT2 #(
		.INIT('h8)
	) name3215 (
		\u7_mc_data_ir_reg[11]/P0001 ,
		_w4154_,
		_w4174_
	);
	LUT2 #(
		.INIT('h1)
	) name3216 (
		_w4173_,
		_w4174_,
		_w4175_
	);
	LUT2 #(
		.INIT('h1)
	) name3217 (
		_w4152_,
		_w4175_,
		_w4176_
	);
	LUT2 #(
		.INIT('h8)
	) name3218 (
		\u7_mc_data_ir_reg[3]/P0001 ,
		_w4152_,
		_w4177_
	);
	LUT2 #(
		.INIT('h1)
	) name3219 (
		_w4176_,
		_w4177_,
		_w4178_
	);
	LUT2 #(
		.INIT('h2)
	) name3220 (
		\u3_byte1_reg[4]/P0001 ,
		_w4154_,
		_w4179_
	);
	LUT2 #(
		.INIT('h8)
	) name3221 (
		\u7_mc_data_ir_reg[12]/P0001 ,
		_w4154_,
		_w4180_
	);
	LUT2 #(
		.INIT('h1)
	) name3222 (
		_w4179_,
		_w4180_,
		_w4181_
	);
	LUT2 #(
		.INIT('h1)
	) name3223 (
		_w4152_,
		_w4181_,
		_w4182_
	);
	LUT2 #(
		.INIT('h8)
	) name3224 (
		\u7_mc_data_ir_reg[4]/P0001 ,
		_w4152_,
		_w4183_
	);
	LUT2 #(
		.INIT('h1)
	) name3225 (
		_w4182_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h2)
	) name3226 (
		\u3_byte1_reg[5]/P0001 ,
		_w4154_,
		_w4185_
	);
	LUT2 #(
		.INIT('h8)
	) name3227 (
		\u7_mc_data_ir_reg[13]/P0001 ,
		_w4154_,
		_w4186_
	);
	LUT2 #(
		.INIT('h1)
	) name3228 (
		_w4185_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h1)
	) name3229 (
		_w4152_,
		_w4187_,
		_w4188_
	);
	LUT2 #(
		.INIT('h8)
	) name3230 (
		\u7_mc_data_ir_reg[5]/P0001 ,
		_w4152_,
		_w4189_
	);
	LUT2 #(
		.INIT('h1)
	) name3231 (
		_w4188_,
		_w4189_,
		_w4190_
	);
	LUT2 #(
		.INIT('h2)
	) name3232 (
		\u3_byte1_reg[6]/P0001 ,
		_w4154_,
		_w4191_
	);
	LUT2 #(
		.INIT('h8)
	) name3233 (
		\u7_mc_data_ir_reg[14]/P0001 ,
		_w4154_,
		_w4192_
	);
	LUT2 #(
		.INIT('h1)
	) name3234 (
		_w4191_,
		_w4192_,
		_w4193_
	);
	LUT2 #(
		.INIT('h1)
	) name3235 (
		_w4152_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h8)
	) name3236 (
		\u7_mc_data_ir_reg[6]/P0001 ,
		_w4152_,
		_w4195_
	);
	LUT2 #(
		.INIT('h1)
	) name3237 (
		_w4194_,
		_w4195_,
		_w4196_
	);
	LUT2 #(
		.INIT('h2)
	) name3238 (
		\u3_byte1_reg[7]/P0001 ,
		_w4154_,
		_w4197_
	);
	LUT2 #(
		.INIT('h8)
	) name3239 (
		\u7_mc_data_ir_reg[15]/P0001 ,
		_w4154_,
		_w4198_
	);
	LUT2 #(
		.INIT('h1)
	) name3240 (
		_w4197_,
		_w4198_,
		_w4199_
	);
	LUT2 #(
		.INIT('h1)
	) name3241 (
		_w4152_,
		_w4199_,
		_w4200_
	);
	LUT2 #(
		.INIT('h8)
	) name3242 (
		\u7_mc_data_ir_reg[7]/P0001 ,
		_w4152_,
		_w4201_
	);
	LUT2 #(
		.INIT('h1)
	) name3243 (
		_w4200_,
		_w4201_,
		_w4202_
	);
	LUT2 #(
		.INIT('h2)
	) name3244 (
		wb_cyc_i_pad,
		_w1870_,
		_w4203_
	);
	LUT2 #(
		.INIT('h8)
	) name3245 (
		\u3_u0_wr_adr_reg[0]/NET0131 ,
		_w1044_,
		_w4204_
	);
	LUT2 #(
		.INIT('h4)
	) name3246 (
		_w1045_,
		_w4203_,
		_w4205_
	);
	LUT2 #(
		.INIT('h4)
	) name3247 (
		_w4204_,
		_w4205_,
		_w4206_
	);
	LUT2 #(
		.INIT('h8)
	) name3248 (
		\u3_u0_wr_adr_reg[2]/NET0131 ,
		_w1044_,
		_w4207_
	);
	LUT2 #(
		.INIT('h2)
	) name3249 (
		\u3_u0_wr_adr_reg[1]/NET0131 ,
		_w1044_,
		_w4208_
	);
	LUT2 #(
		.INIT('h1)
	) name3250 (
		_w4207_,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h2)
	) name3251 (
		_w4203_,
		_w4209_,
		_w4210_
	);
	LUT2 #(
		.INIT('h8)
	) name3252 (
		\u3_u0_wr_adr_reg[3]/NET0131 ,
		_w1044_,
		_w4211_
	);
	LUT2 #(
		.INIT('h2)
	) name3253 (
		\u3_u0_wr_adr_reg[2]/NET0131 ,
		_w1044_,
		_w4212_
	);
	LUT2 #(
		.INIT('h1)
	) name3254 (
		_w4211_,
		_w4212_,
		_w4213_
	);
	LUT2 #(
		.INIT('h2)
	) name3255 (
		_w4203_,
		_w4213_,
		_w4214_
	);
	LUT2 #(
		.INIT('h4)
	) name3256 (
		\u0_init_req_reg/NET0131 ,
		_w1681_,
		_w4215_
	);
	LUT2 #(
		.INIT('h4)
	) name3257 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w4216_
	);
	LUT2 #(
		.INIT('h8)
	) name3258 (
		_w4215_,
		_w4216_,
		_w4217_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		_w1079_,
		_w1389_,
		_w4218_
	);
	LUT2 #(
		.INIT('h1)
	) name3260 (
		\u5_state_reg[18]/NET0131 ,
		_w4218_,
		_w4219_
	);
	LUT2 #(
		.INIT('h1)
	) name3261 (
		_w1069_,
		_w4219_,
		_w4220_
	);
	LUT2 #(
		.INIT('h2)
	) name3262 (
		_w3089_,
		_w4220_,
		_w4221_
	);
	LUT2 #(
		.INIT('h8)
	) name3263 (
		_w3080_,
		_w4221_,
		_w4222_
	);
	LUT2 #(
		.INIT('h1)
	) name3264 (
		_w4217_,
		_w4222_,
		_w4223_
	);
	LUT2 #(
		.INIT('h8)
	) name3265 (
		\wb_addr_i[2]_pad ,
		_w2878_,
		_w4224_
	);
	LUT2 #(
		.INIT('h8)
	) name3266 (
		\wb_addr_i[1]_pad ,
		_w2606_,
		_w4225_
	);
	LUT2 #(
		.INIT('h8)
	) name3267 (
		\wb_addr_i[0]_pad ,
		_w2388_,
		_w4226_
	);
	LUT2 #(
		.INIT('h1)
	) name3268 (
		_w4224_,
		_w4225_,
		_w4227_
	);
	LUT2 #(
		.INIT('h4)
	) name3269 (
		_w4226_,
		_w4227_,
		_w4228_
	);
	LUT2 #(
		.INIT('h1)
	) name3270 (
		_w2858_,
		_w4228_,
		_w4229_
	);
	LUT2 #(
		.INIT('h1)
	) name3271 (
		\u1_acs_addr_reg[0]/P0001 ,
		_w2861_,
		_w4230_
	);
	LUT2 #(
		.INIT('h4)
	) name3272 (
		\u1_u0_out_r_reg[0]/P0001 ,
		_w2861_,
		_w4231_
	);
	LUT2 #(
		.INIT('h2)
	) name3273 (
		_w2858_,
		_w4230_,
		_w4232_
	);
	LUT2 #(
		.INIT('h4)
	) name3274 (
		_w4231_,
		_w4232_,
		_w4233_
	);
	LUT2 #(
		.INIT('h1)
	) name3275 (
		_w4229_,
		_w4233_,
		_w4234_
	);
	LUT2 #(
		.INIT('h1)
	) name3276 (
		\u1_acs_addr_reg[10]/P0001 ,
		_w2861_,
		_w4235_
	);
	LUT2 #(
		.INIT('h4)
	) name3277 (
		\u1_u0_out_r_reg[10]/P0001 ,
		_w2861_,
		_w4236_
	);
	LUT2 #(
		.INIT('h2)
	) name3278 (
		_w2858_,
		_w4235_,
		_w4237_
	);
	LUT2 #(
		.INIT('h4)
	) name3279 (
		_w4236_,
		_w4237_,
		_w4238_
	);
	LUT2 #(
		.INIT('h8)
	) name3280 (
		\wb_addr_i[10]_pad ,
		_w2388_,
		_w4239_
	);
	LUT2 #(
		.INIT('h1)
	) name3281 (
		_w4015_,
		_w4065_,
		_w4240_
	);
	LUT2 #(
		.INIT('h4)
	) name3282 (
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h1)
	) name3283 (
		_w2858_,
		_w4241_,
		_w4242_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		_w4238_,
		_w4242_,
		_w4243_
	);
	LUT2 #(
		.INIT('h8)
	) name3285 (
		\wb_addr_i[3]_pad ,
		_w2878_,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name3286 (
		\wb_addr_i[1]_pad ,
		_w2388_,
		_w4245_
	);
	LUT2 #(
		.INIT('h8)
	) name3287 (
		\wb_addr_i[2]_pad ,
		_w2606_,
		_w4246_
	);
	LUT2 #(
		.INIT('h1)
	) name3288 (
		_w4244_,
		_w4245_,
		_w4247_
	);
	LUT2 #(
		.INIT('h4)
	) name3289 (
		_w4246_,
		_w4247_,
		_w4248_
	);
	LUT2 #(
		.INIT('h1)
	) name3290 (
		_w2858_,
		_w4248_,
		_w4249_
	);
	LUT2 #(
		.INIT('h1)
	) name3291 (
		\u1_acs_addr_reg[1]/P0001 ,
		_w2861_,
		_w4250_
	);
	LUT2 #(
		.INIT('h4)
	) name3292 (
		\u1_u0_out_r_reg[1]/P0001 ,
		_w2861_,
		_w4251_
	);
	LUT2 #(
		.INIT('h2)
	) name3293 (
		_w2858_,
		_w4250_,
		_w4252_
	);
	LUT2 #(
		.INIT('h4)
	) name3294 (
		_w4251_,
		_w4252_,
		_w4253_
	);
	LUT2 #(
		.INIT('h1)
	) name3295 (
		_w4249_,
		_w4253_,
		_w4254_
	);
	LUT2 #(
		.INIT('h8)
	) name3296 (
		\wb_addr_i[3]_pad ,
		_w2606_,
		_w4255_
	);
	LUT2 #(
		.INIT('h8)
	) name3297 (
		\wb_addr_i[4]_pad ,
		_w2878_,
		_w4256_
	);
	LUT2 #(
		.INIT('h8)
	) name3298 (
		\wb_addr_i[2]_pad ,
		_w2388_,
		_w4257_
	);
	LUT2 #(
		.INIT('h1)
	) name3299 (
		_w4255_,
		_w4256_,
		_w4258_
	);
	LUT2 #(
		.INIT('h4)
	) name3300 (
		_w4257_,
		_w4258_,
		_w4259_
	);
	LUT2 #(
		.INIT('h1)
	) name3301 (
		_w2858_,
		_w4259_,
		_w4260_
	);
	LUT2 #(
		.INIT('h1)
	) name3302 (
		\u1_acs_addr_reg[2]/P0001 ,
		_w2861_,
		_w4261_
	);
	LUT2 #(
		.INIT('h4)
	) name3303 (
		\u1_u0_out_r_reg[2]/P0001 ,
		_w2861_,
		_w4262_
	);
	LUT2 #(
		.INIT('h2)
	) name3304 (
		_w2858_,
		_w4261_,
		_w4263_
	);
	LUT2 #(
		.INIT('h4)
	) name3305 (
		_w4262_,
		_w4263_,
		_w4264_
	);
	LUT2 #(
		.INIT('h1)
	) name3306 (
		_w4260_,
		_w4264_,
		_w4265_
	);
	LUT2 #(
		.INIT('h8)
	) name3307 (
		\wb_addr_i[4]_pad ,
		_w2606_,
		_w4266_
	);
	LUT2 #(
		.INIT('h8)
	) name3308 (
		\wb_addr_i[5]_pad ,
		_w2878_,
		_w4267_
	);
	LUT2 #(
		.INIT('h8)
	) name3309 (
		\wb_addr_i[3]_pad ,
		_w2388_,
		_w4268_
	);
	LUT2 #(
		.INIT('h1)
	) name3310 (
		_w4266_,
		_w4267_,
		_w4269_
	);
	LUT2 #(
		.INIT('h4)
	) name3311 (
		_w4268_,
		_w4269_,
		_w4270_
	);
	LUT2 #(
		.INIT('h1)
	) name3312 (
		_w2858_,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('h1)
	) name3313 (
		\u1_acs_addr_reg[3]/P0001 ,
		_w2861_,
		_w4272_
	);
	LUT2 #(
		.INIT('h4)
	) name3314 (
		\u1_u0_out_r_reg[3]/P0001 ,
		_w2861_,
		_w4273_
	);
	LUT2 #(
		.INIT('h2)
	) name3315 (
		_w2858_,
		_w4272_,
		_w4274_
	);
	LUT2 #(
		.INIT('h4)
	) name3316 (
		_w4273_,
		_w4274_,
		_w4275_
	);
	LUT2 #(
		.INIT('h1)
	) name3317 (
		_w4271_,
		_w4275_,
		_w4276_
	);
	LUT2 #(
		.INIT('h8)
	) name3318 (
		\wb_addr_i[6]_pad ,
		_w2606_,
		_w4277_
	);
	LUT2 #(
		.INIT('h8)
	) name3319 (
		\wb_addr_i[7]_pad ,
		_w2878_,
		_w4278_
	);
	LUT2 #(
		.INIT('h8)
	) name3320 (
		\wb_addr_i[5]_pad ,
		_w2388_,
		_w4279_
	);
	LUT2 #(
		.INIT('h1)
	) name3321 (
		_w4277_,
		_w4278_,
		_w4280_
	);
	LUT2 #(
		.INIT('h4)
	) name3322 (
		_w4279_,
		_w4280_,
		_w4281_
	);
	LUT2 #(
		.INIT('h1)
	) name3323 (
		_w2858_,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h1)
	) name3324 (
		\u1_acs_addr_reg[5]/P0001 ,
		_w2861_,
		_w4283_
	);
	LUT2 #(
		.INIT('h4)
	) name3325 (
		\u1_u0_out_r_reg[5]/P0001 ,
		_w2861_,
		_w4284_
	);
	LUT2 #(
		.INIT('h2)
	) name3326 (
		_w2858_,
		_w4283_,
		_w4285_
	);
	LUT2 #(
		.INIT('h4)
	) name3327 (
		_w4284_,
		_w4285_,
		_w4286_
	);
	LUT2 #(
		.INIT('h1)
	) name3328 (
		_w4282_,
		_w4286_,
		_w4287_
	);
	LUT2 #(
		.INIT('h8)
	) name3329 (
		\wb_addr_i[7]_pad ,
		_w2606_,
		_w4288_
	);
	LUT2 #(
		.INIT('h8)
	) name3330 (
		\wb_addr_i[8]_pad ,
		_w2878_,
		_w4289_
	);
	LUT2 #(
		.INIT('h8)
	) name3331 (
		\wb_addr_i[6]_pad ,
		_w2388_,
		_w4290_
	);
	LUT2 #(
		.INIT('h1)
	) name3332 (
		_w4288_,
		_w4289_,
		_w4291_
	);
	LUT2 #(
		.INIT('h4)
	) name3333 (
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT2 #(
		.INIT('h1)
	) name3334 (
		_w2858_,
		_w4292_,
		_w4293_
	);
	LUT2 #(
		.INIT('h1)
	) name3335 (
		\u1_acs_addr_reg[6]/P0001 ,
		_w2861_,
		_w4294_
	);
	LUT2 #(
		.INIT('h4)
	) name3336 (
		\u1_u0_out_r_reg[6]/P0001 ,
		_w2861_,
		_w4295_
	);
	LUT2 #(
		.INIT('h2)
	) name3337 (
		_w2858_,
		_w4294_,
		_w4296_
	);
	LUT2 #(
		.INIT('h4)
	) name3338 (
		_w4295_,
		_w4296_,
		_w4297_
	);
	LUT2 #(
		.INIT('h1)
	) name3339 (
		_w4293_,
		_w4297_,
		_w4298_
	);
	LUT2 #(
		.INIT('h1)
	) name3340 (
		\u1_acs_addr_reg[9]/P0001 ,
		_w2861_,
		_w4299_
	);
	LUT2 #(
		.INIT('h4)
	) name3341 (
		\u1_u0_out_r_reg[9]/P0001 ,
		_w2861_,
		_w4300_
	);
	LUT2 #(
		.INIT('h2)
	) name3342 (
		_w2858_,
		_w4299_,
		_w4301_
	);
	LUT2 #(
		.INIT('h4)
	) name3343 (
		_w4300_,
		_w4301_,
		_w4302_
	);
	LUT2 #(
		.INIT('h8)
	) name3344 (
		\wb_addr_i[9]_pad ,
		_w2388_,
		_w4303_
	);
	LUT2 #(
		.INIT('h1)
	) name3345 (
		_w4018_,
		_w4043_,
		_w4304_
	);
	LUT2 #(
		.INIT('h4)
	) name3346 (
		_w4303_,
		_w4304_,
		_w4305_
	);
	LUT2 #(
		.INIT('h1)
	) name3347 (
		_w2858_,
		_w4305_,
		_w4306_
	);
	LUT2 #(
		.INIT('h1)
	) name3348 (
		_w4302_,
		_w4306_,
		_w4307_
	);
	LUT2 #(
		.INIT('h4)
	) name3349 (
		_w1039_,
		_w1398_,
		_w4308_
	);
	LUT2 #(
		.INIT('h1)
	) name3350 (
		\u5_cnt_reg/NET0131 ,
		_w4308_,
		_w4309_
	);
	LUT2 #(
		.INIT('h2)
	) name3351 (
		wb_stb_i_pad,
		_w2269_,
		_w4310_
	);
	LUT2 #(
		.INIT('h8)
	) name3352 (
		\u5_wb_cycle_reg/NET0131 ,
		wb_cyc_i_pad,
		_w4311_
	);
	LUT2 #(
		.INIT('h4)
	) name3353 (
		_w4310_,
		_w4311_,
		_w4312_
	);
	LUT2 #(
		.INIT('h1)
	) name3354 (
		_w1686_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('h8)
	) name3355 (
		\mem_ack_r_reg/P0001 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w4314_
	);
	LUT2 #(
		.INIT('h4)
	) name3356 (
		\u5_wr_cycle_reg/NET0131 ,
		wb_stb_i_pad,
		_w4315_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w4314_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h8)
	) name3358 (
		\u1_col_adr_reg[8]/P0001 ,
		_w4316_,
		_w4317_
	);
	LUT2 #(
		.INIT('h2)
	) name3359 (
		\wb_addr_i[10]_pad ,
		_w4316_,
		_w4318_
	);
	LUT2 #(
		.INIT('h4)
	) name3360 (
		_w3980_,
		_w4318_,
		_w4319_
	);
	LUT2 #(
		.INIT('h8)
	) name3361 (
		_w2366_,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h1)
	) name3362 (
		_w4317_,
		_w4320_,
		_w4321_
	);
	LUT2 #(
		.INIT('h1)
	) name3363 (
		\u1_acs_addr_reg[7]/P0001 ,
		_w4006_,
		_w4322_
	);
	LUT2 #(
		.INIT('h1)
	) name3364 (
		_w4007_,
		_w4322_,
		_w4323_
	);
	LUT2 #(
		.INIT('h2)
	) name3365 (
		\u5_state_reg[61]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w4324_
	);
	LUT2 #(
		.INIT('h1)
	) name3366 (
		\u7_mc_ack_r_reg/NET0131 ,
		_w4324_,
		_w4325_
	);
	LUT2 #(
		.INIT('h2)
	) name3367 (
		_w1236_,
		_w4325_,
		_w4326_
	);
	LUT2 #(
		.INIT('h4)
	) name3368 (
		_w1238_,
		_w1270_,
		_w4327_
	);
	LUT2 #(
		.INIT('h2)
	) name3369 (
		\u5_state_reg[61]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w4328_
	);
	LUT2 #(
		.INIT('h4)
	) name3370 (
		_w4327_,
		_w4328_,
		_w4329_
	);
	LUT2 #(
		.INIT('h1)
	) name3371 (
		_w4326_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h8)
	) name3372 (
		\u4_ps_cnt_reg[0]/NET0131 ,
		\u4_rfr_en_reg/NET0131 ,
		_w4331_
	);
	LUT2 #(
		.INIT('h8)
	) name3373 (
		\u4_ps_cnt_reg[1]/NET0131 ,
		_w4331_,
		_w4332_
	);
	LUT2 #(
		.INIT('h8)
	) name3374 (
		\u4_ps_cnt_reg[2]/NET0131 ,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h8)
	) name3375 (
		\u4_ps_cnt_reg[3]/NET0131 ,
		_w4333_,
		_w4334_
	);
	LUT2 #(
		.INIT('h8)
	) name3376 (
		\u4_ps_cnt_reg[4]/NET0131 ,
		_w4334_,
		_w4335_
	);
	LUT2 #(
		.INIT('h1)
	) name3377 (
		\u4_ps_cnt_reg[4]/NET0131 ,
		_w4334_,
		_w4336_
	);
	LUT2 #(
		.INIT('h4)
	) name3378 (
		\u0_csr_r2_reg[1]/NET0131 ,
		\u4_ps_cnt_reg[1]/NET0131 ,
		_w4337_
	);
	LUT2 #(
		.INIT('h1)
	) name3379 (
		\u0_csr_r2_reg[5]/NET0131 ,
		\u4_ps_cnt_reg[5]/NET0131 ,
		_w4338_
	);
	LUT2 #(
		.INIT('h8)
	) name3380 (
		\u0_csr_r2_reg[5]/NET0131 ,
		\u4_ps_cnt_reg[5]/NET0131 ,
		_w4339_
	);
	LUT2 #(
		.INIT('h1)
	) name3381 (
		_w4338_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h2)
	) name3382 (
		\u0_csr_r2_reg[4]/NET0131 ,
		\u4_ps_cnt_reg[4]/NET0131 ,
		_w4341_
	);
	LUT2 #(
		.INIT('h4)
	) name3383 (
		\u0_csr_r2_reg[4]/NET0131 ,
		\u4_ps_cnt_reg[4]/NET0131 ,
		_w4342_
	);
	LUT2 #(
		.INIT('h1)
	) name3384 (
		\u0_csr_r2_reg[7]/NET0131 ,
		\u4_ps_cnt_reg[7]/NET0131 ,
		_w4343_
	);
	LUT2 #(
		.INIT('h8)
	) name3385 (
		\u0_csr_r2_reg[7]/NET0131 ,
		\u4_ps_cnt_reg[7]/NET0131 ,
		_w4344_
	);
	LUT2 #(
		.INIT('h1)
	) name3386 (
		_w4343_,
		_w4344_,
		_w4345_
	);
	LUT2 #(
		.INIT('h4)
	) name3387 (
		\u0_csr_r2_reg[2]/NET0131 ,
		\u4_ps_cnt_reg[2]/NET0131 ,
		_w4346_
	);
	LUT2 #(
		.INIT('h2)
	) name3388 (
		\u0_csr_r2_reg[2]/NET0131 ,
		\u4_ps_cnt_reg[2]/NET0131 ,
		_w4347_
	);
	LUT2 #(
		.INIT('h2)
	) name3389 (
		\u0_csr_r2_reg[6]/NET0131 ,
		\u4_ps_cnt_reg[6]/NET0131 ,
		_w4348_
	);
	LUT2 #(
		.INIT('h4)
	) name3390 (
		\u0_csr_r2_reg[6]/NET0131 ,
		\u4_ps_cnt_reg[6]/NET0131 ,
		_w4349_
	);
	LUT2 #(
		.INIT('h4)
	) name3391 (
		\u0_csr_r2_reg[3]/NET0131 ,
		\u4_ps_cnt_reg[3]/NET0131 ,
		_w4350_
	);
	LUT2 #(
		.INIT('h2)
	) name3392 (
		\u0_csr_r2_reg[0]/NET0131 ,
		\u4_ps_cnt_reg[0]/NET0131 ,
		_w4351_
	);
	LUT2 #(
		.INIT('h2)
	) name3393 (
		\u0_csr_r2_reg[3]/NET0131 ,
		\u4_ps_cnt_reg[3]/NET0131 ,
		_w4352_
	);
	LUT2 #(
		.INIT('h4)
	) name3394 (
		\u0_csr_r2_reg[0]/NET0131 ,
		\u4_ps_cnt_reg[0]/NET0131 ,
		_w4353_
	);
	LUT2 #(
		.INIT('h2)
	) name3395 (
		\u0_csr_r2_reg[1]/NET0131 ,
		\u4_ps_cnt_reg[1]/NET0131 ,
		_w4354_
	);
	LUT2 #(
		.INIT('h1)
	) name3396 (
		_w4337_,
		_w4341_,
		_w4355_
	);
	LUT2 #(
		.INIT('h1)
	) name3397 (
		_w4342_,
		_w4346_,
		_w4356_
	);
	LUT2 #(
		.INIT('h1)
	) name3398 (
		_w4347_,
		_w4348_,
		_w4357_
	);
	LUT2 #(
		.INIT('h1)
	) name3399 (
		_w4349_,
		_w4350_,
		_w4358_
	);
	LUT2 #(
		.INIT('h1)
	) name3400 (
		_w4351_,
		_w4352_,
		_w4359_
	);
	LUT2 #(
		.INIT('h1)
	) name3401 (
		_w4353_,
		_w4354_,
		_w4360_
	);
	LUT2 #(
		.INIT('h8)
	) name3402 (
		_w4359_,
		_w4360_,
		_w4361_
	);
	LUT2 #(
		.INIT('h8)
	) name3403 (
		_w4357_,
		_w4358_,
		_w4362_
	);
	LUT2 #(
		.INIT('h8)
	) name3404 (
		_w4355_,
		_w4356_,
		_w4363_
	);
	LUT2 #(
		.INIT('h1)
	) name3405 (
		_w4340_,
		_w4345_,
		_w4364_
	);
	LUT2 #(
		.INIT('h8)
	) name3406 (
		_w4363_,
		_w4364_,
		_w4365_
	);
	LUT2 #(
		.INIT('h8)
	) name3407 (
		_w4361_,
		_w4362_,
		_w4366_
	);
	LUT2 #(
		.INIT('h8)
	) name3408 (
		_w4365_,
		_w4366_,
		_w4367_
	);
	LUT2 #(
		.INIT('h1)
	) name3409 (
		\u0_csr_r2_reg[0]/NET0131 ,
		\u0_csr_r2_reg[1]/NET0131 ,
		_w4368_
	);
	LUT2 #(
		.INIT('h1)
	) name3410 (
		\u0_csr_r2_reg[2]/NET0131 ,
		\u0_csr_r2_reg[3]/NET0131 ,
		_w4369_
	);
	LUT2 #(
		.INIT('h1)
	) name3411 (
		\u0_csr_r2_reg[4]/NET0131 ,
		\u0_csr_r2_reg[5]/NET0131 ,
		_w4370_
	);
	LUT2 #(
		.INIT('h1)
	) name3412 (
		\u0_csr_r2_reg[6]/NET0131 ,
		\u0_csr_r2_reg[7]/NET0131 ,
		_w4371_
	);
	LUT2 #(
		.INIT('h8)
	) name3413 (
		_w4370_,
		_w4371_,
		_w4372_
	);
	LUT2 #(
		.INIT('h8)
	) name3414 (
		_w4368_,
		_w4369_,
		_w4373_
	);
	LUT2 #(
		.INIT('h8)
	) name3415 (
		_w4372_,
		_w4373_,
		_w4374_
	);
	LUT2 #(
		.INIT('h2)
	) name3416 (
		_w4367_,
		_w4374_,
		_w4375_
	);
	LUT2 #(
		.INIT('h1)
	) name3417 (
		_w4335_,
		_w4336_,
		_w4376_
	);
	LUT2 #(
		.INIT('h4)
	) name3418 (
		_w4375_,
		_w4376_,
		_w4377_
	);
	LUT2 #(
		.INIT('h8)
	) name3419 (
		\u4_rfr_ce_reg/NET0131 ,
		\u4_rfr_cnt_reg[0]/NET0131 ,
		_w4378_
	);
	LUT2 #(
		.INIT('h1)
	) name3420 (
		\u4_rfr_cnt_reg[1]/NET0131 ,
		_w4378_,
		_w4379_
	);
	LUT2 #(
		.INIT('h8)
	) name3421 (
		\u4_rfr_cnt_reg[1]/NET0131 ,
		_w4378_,
		_w4380_
	);
	LUT2 #(
		.INIT('h1)
	) name3422 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w4379_,
		_w4381_
	);
	LUT2 #(
		.INIT('h4)
	) name3423 (
		_w4380_,
		_w4381_,
		_w4382_
	);
	LUT2 #(
		.INIT('h4)
	) name3424 (
		\u5_state_reg[7]/NET0131 ,
		_w970_,
		_w4383_
	);
	LUT2 #(
		.INIT('h8)
	) name3425 (
		_w1261_,
		_w4383_,
		_w4384_
	);
	LUT2 #(
		.INIT('h8)
	) name3426 (
		_w1344_,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h8)
	) name3427 (
		_w1334_,
		_w4385_,
		_w4386_
	);
	LUT2 #(
		.INIT('h8)
	) name3428 (
		\u5_state_reg[33]/NET0131 ,
		\u5_state_reg[34]/NET0131 ,
		_w4387_
	);
	LUT2 #(
		.INIT('h8)
	) name3429 (
		_w1332_,
		_w3074_,
		_w4388_
	);
	LUT2 #(
		.INIT('h1)
	) name3430 (
		\u5_state_reg[33]/NET0131 ,
		\u5_state_reg[34]/NET0131 ,
		_w4389_
	);
	LUT2 #(
		.INIT('h1)
	) name3431 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		_w4390_
	);
	LUT2 #(
		.INIT('h4)
	) name3432 (
		_w4387_,
		_w4390_,
		_w4391_
	);
	LUT2 #(
		.INIT('h4)
	) name3433 (
		_w4389_,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h8)
	) name3434 (
		_w3072_,
		_w4388_,
		_w4393_
	);
	LUT2 #(
		.INIT('h8)
	) name3435 (
		_w4392_,
		_w4393_,
		_w4394_
	);
	LUT2 #(
		.INIT('h8)
	) name3436 (
		_w3055_,
		_w4394_,
		_w4395_
	);
	LUT2 #(
		.INIT('h8)
	) name3437 (
		_w4386_,
		_w4395_,
		_w4396_
	);
	LUT2 #(
		.INIT('h8)
	) name3438 (
		_w3076_,
		_w4396_,
		_w4397_
	);
	LUT2 #(
		.INIT('h1)
	) name3439 (
		\u0_init_req_reg/NET0131 ,
		\u0_lmr_req_reg/NET0131 ,
		_w4398_
	);
	LUT2 #(
		.INIT('h4)
	) name3440 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		_w4399_
	);
	LUT2 #(
		.INIT('h4)
	) name3441 (
		\u5_susp_req_r_reg/NET0131 ,
		_w4399_,
		_w4400_
	);
	LUT2 #(
		.INIT('h8)
	) name3442 (
		_w4398_,
		_w4400_,
		_w4401_
	);
	LUT2 #(
		.INIT('h8)
	) name3443 (
		_w1628_,
		_w4401_,
		_w4402_
	);
	LUT2 #(
		.INIT('h1)
	) name3444 (
		_w4397_,
		_w4402_,
		_w4403_
	);
	LUT2 #(
		.INIT('h1)
	) name3445 (
		\u4_rfr_ce_reg/NET0131 ,
		\u4_rfr_cnt_reg[0]/NET0131 ,
		_w4404_
	);
	LUT2 #(
		.INIT('h1)
	) name3446 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w4378_,
		_w4405_
	);
	LUT2 #(
		.INIT('h4)
	) name3447 (
		_w4404_,
		_w4405_,
		_w4406_
	);
	LUT2 #(
		.INIT('h1)
	) name3448 (
		\u4_rfr_cnt_reg[2]/NET0131 ,
		_w4380_,
		_w4407_
	);
	LUT2 #(
		.INIT('h8)
	) name3449 (
		\u4_rfr_cnt_reg[2]/NET0131 ,
		_w4380_,
		_w4408_
	);
	LUT2 #(
		.INIT('h1)
	) name3450 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w4407_,
		_w4409_
	);
	LUT2 #(
		.INIT('h4)
	) name3451 (
		_w4408_,
		_w4409_,
		_w4410_
	);
	LUT2 #(
		.INIT('h8)
	) name3452 (
		\u4_rfr_cnt_reg[3]/NET0131 ,
		_w4408_,
		_w4411_
	);
	LUT2 #(
		.INIT('h1)
	) name3453 (
		\u4_rfr_cnt_reg[3]/NET0131 ,
		_w4408_,
		_w4412_
	);
	LUT2 #(
		.INIT('h1)
	) name3454 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w4411_,
		_w4413_
	);
	LUT2 #(
		.INIT('h4)
	) name3455 (
		_w4412_,
		_w4413_,
		_w4414_
	);
	LUT2 #(
		.INIT('h1)
	) name3456 (
		\u4_rfr_cnt_reg[4]/NET0131 ,
		_w4411_,
		_w4415_
	);
	LUT2 #(
		.INIT('h8)
	) name3457 (
		\u4_rfr_cnt_reg[4]/NET0131 ,
		_w4411_,
		_w4416_
	);
	LUT2 #(
		.INIT('h1)
	) name3458 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w4415_,
		_w4417_
	);
	LUT2 #(
		.INIT('h4)
	) name3459 (
		_w4416_,
		_w4417_,
		_w4418_
	);
	LUT2 #(
		.INIT('h1)
	) name3460 (
		\u4_rfr_cnt_reg[5]/NET0131 ,
		_w4416_,
		_w4419_
	);
	LUT2 #(
		.INIT('h8)
	) name3461 (
		\u4_rfr_cnt_reg[5]/NET0131 ,
		_w4416_,
		_w4420_
	);
	LUT2 #(
		.INIT('h1)
	) name3462 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w4419_,
		_w4421_
	);
	LUT2 #(
		.INIT('h4)
	) name3463 (
		_w4420_,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h1)
	) name3464 (
		\u4_rfr_cnt_reg[6]/NET0131 ,
		_w4420_,
		_w4423_
	);
	LUT2 #(
		.INIT('h8)
	) name3465 (
		\u4_rfr_cnt_reg[6]/NET0131 ,
		_w4420_,
		_w4424_
	);
	LUT2 #(
		.INIT('h1)
	) name3466 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w4423_,
		_w4425_
	);
	LUT2 #(
		.INIT('h4)
	) name3467 (
		_w4424_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h1)
	) name3468 (
		\u4_rfr_cnt_reg[7]/NET0131 ,
		_w4424_,
		_w4427_
	);
	LUT2 #(
		.INIT('h8)
	) name3469 (
		\u4_rfr_cnt_reg[7]/NET0131 ,
		_w4424_,
		_w4428_
	);
	LUT2 #(
		.INIT('h1)
	) name3470 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w4427_,
		_w4429_
	);
	LUT2 #(
		.INIT('h4)
	) name3471 (
		_w4428_,
		_w4429_,
		_w4430_
	);
	LUT2 #(
		.INIT('h8)
	) name3472 (
		\u5_cs_le_reg/P0001 ,
		_w1046_,
		_w4431_
	);
	LUT2 #(
		.INIT('h8)
	) name3473 (
		\u0_wp_err_reg/NET0131 ,
		wb_cyc_i_pad,
		_w4432_
	);
	LUT2 #(
		.INIT('h4)
	) name3474 (
		_w4431_,
		_w4432_,
		_w4433_
	);
	LUT2 #(
		.INIT('h8)
	) name3475 (
		\u0_u0_csc_reg[8]/P0001 ,
		_w3414_,
		_w4434_
	);
	LUT2 #(
		.INIT('h8)
	) name3476 (
		\u0_u1_csc_reg[8]/P0001 ,
		_w3456_,
		_w4435_
	);
	LUT2 #(
		.INIT('h1)
	) name3477 (
		_w4434_,
		_w4435_,
		_w4436_
	);
	LUT2 #(
		.INIT('h8)
	) name3478 (
		\u5_cs_le_reg/P0001 ,
		_w1047_,
		_w4437_
	);
	LUT2 #(
		.INIT('h4)
	) name3479 (
		_w4436_,
		_w4437_,
		_w4438_
	);
	LUT2 #(
		.INIT('h1)
	) name3480 (
		_w4433_,
		_w4438_,
		_w4439_
	);
	LUT2 #(
		.INIT('h8)
	) name3481 (
		\u5_mc_adv_r1_reg/NET0131 ,
		\u5_mc_le_reg/NET0131 ,
		_w4440_
	);
	LUT2 #(
		.INIT('h2)
	) name3482 (
		_w1629_,
		_w2746_,
		_w4441_
	);
	LUT2 #(
		.INIT('h8)
	) name3483 (
		_w1023_,
		_w1113_,
		_w4442_
	);
	LUT2 #(
		.INIT('h1)
	) name3484 (
		_w1114_,
		_w4441_,
		_w4443_
	);
	LUT2 #(
		.INIT('h4)
	) name3485 (
		_w4442_,
		_w4443_,
		_w4444_
	);
	LUT2 #(
		.INIT('h4)
	) name3486 (
		\u5_mc_le_reg/NET0131 ,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('h1)
	) name3487 (
		_w4440_,
		_w4445_,
		_w4446_
	);
	LUT2 #(
		.INIT('h2)
	) name3488 (
		_w3986_,
		_w4057_,
		_w4447_
	);
	LUT2 #(
		.INIT('h1)
	) name3489 (
		_w3986_,
		_w4081_,
		_w4448_
	);
	LUT2 #(
		.INIT('h1)
	) name3490 (
		_w4447_,
		_w4448_,
		_w4449_
	);
	LUT2 #(
		.INIT('h8)
	) name3491 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1401_,
		_w4450_
	);
	LUT2 #(
		.INIT('h4)
	) name3492 (
		\u5_ir_cnt_reg[0]/P0001 ,
		_w4450_,
		_w4451_
	);
	LUT2 #(
		.INIT('h2)
	) name3493 (
		\u5_ir_cnt_reg[1]/P0001 ,
		_w4451_,
		_w4452_
	);
	LUT2 #(
		.INIT('h1)
	) name3494 (
		\u5_ir_cnt_reg[0]/P0001 ,
		\u5_ir_cnt_reg[1]/P0001 ,
		_w4453_
	);
	LUT2 #(
		.INIT('h8)
	) name3495 (
		_w4450_,
		_w4453_,
		_w4454_
	);
	LUT2 #(
		.INIT('h1)
	) name3496 (
		\u5_state_reg[22]/NET0131 ,
		_w4454_,
		_w4455_
	);
	LUT2 #(
		.INIT('h4)
	) name3497 (
		_w4452_,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h8)
	) name3498 (
		\u4_ps_cnt_reg[5]/NET0131 ,
		_w4335_,
		_w4457_
	);
	LUT2 #(
		.INIT('h8)
	) name3499 (
		\u4_ps_cnt_reg[6]/NET0131 ,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h1)
	) name3500 (
		\u4_ps_cnt_reg[7]/NET0131 ,
		_w4458_,
		_w4459_
	);
	LUT2 #(
		.INIT('h8)
	) name3501 (
		\u4_ps_cnt_reg[7]/NET0131 ,
		_w4458_,
		_w4460_
	);
	LUT2 #(
		.INIT('h1)
	) name3502 (
		_w4375_,
		_w4459_,
		_w4461_
	);
	LUT2 #(
		.INIT('h4)
	) name3503 (
		_w4460_,
		_w4461_,
		_w4462_
	);
	LUT2 #(
		.INIT('h4)
	) name3504 (
		\u5_ir_cnt_reg[2]/P0001 ,
		_w4454_,
		_w4463_
	);
	LUT2 #(
		.INIT('h2)
	) name3505 (
		\u5_ir_cnt_reg[3]/P0001 ,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h1)
	) name3506 (
		\u5_ir_cnt_reg[2]/P0001 ,
		\u5_ir_cnt_reg[3]/P0001 ,
		_w4465_
	);
	LUT2 #(
		.INIT('h8)
	) name3507 (
		_w4453_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h8)
	) name3508 (
		_w4450_,
		_w4466_,
		_w4467_
	);
	LUT2 #(
		.INIT('h1)
	) name3509 (
		_w4464_,
		_w4467_,
		_w4468_
	);
	LUT2 #(
		.INIT('h1)
	) name3510 (
		\u5_state_reg[22]/NET0131 ,
		_w4468_,
		_w4469_
	);
	LUT2 #(
		.INIT('h2)
	) name3511 (
		\u5_ir_cnt_reg[0]/P0001 ,
		_w4450_,
		_w4470_
	);
	LUT2 #(
		.INIT('h1)
	) name3512 (
		_w4451_,
		_w4470_,
		_w4471_
	);
	LUT2 #(
		.INIT('h1)
	) name3513 (
		\u5_state_reg[22]/NET0131 ,
		_w4471_,
		_w4472_
	);
	LUT2 #(
		.INIT('h2)
	) name3514 (
		\u5_ir_cnt_reg[2]/P0001 ,
		_w4454_,
		_w4473_
	);
	LUT2 #(
		.INIT('h1)
	) name3515 (
		_w4463_,
		_w4473_,
		_w4474_
	);
	LUT2 #(
		.INIT('h1)
	) name3516 (
		\u5_state_reg[22]/NET0131 ,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h2)
	) name3517 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b3_last_row_reg[3]/P0001 ,
		_w4476_
	);
	LUT2 #(
		.INIT('h2)
	) name3518 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b3_last_row_reg[11]/P0001 ,
		_w4477_
	);
	LUT2 #(
		.INIT('h4)
	) name3519 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u1_b3_last_row_reg[0]/P0001 ,
		_w4478_
	);
	LUT2 #(
		.INIT('h2)
	) name3520 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b3_last_row_reg[2]/P0001 ,
		_w4479_
	);
	LUT2 #(
		.INIT('h2)
	) name3521 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b3_last_row_reg[12]/P0001 ,
		_w4480_
	);
	LUT2 #(
		.INIT('h2)
	) name3522 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b3_last_row_reg[9]/P0001 ,
		_w4481_
	);
	LUT2 #(
		.INIT('h1)
	) name3523 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u1_b3_last_row_reg[10]/P0001 ,
		_w4482_
	);
	LUT2 #(
		.INIT('h8)
	) name3524 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u1_b3_last_row_reg[10]/P0001 ,
		_w4483_
	);
	LUT2 #(
		.INIT('h1)
	) name3525 (
		_w4482_,
		_w4483_,
		_w4484_
	);
	LUT2 #(
		.INIT('h2)
	) name3526 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b3_last_row_reg[5]/P0001 ,
		_w4485_
	);
	LUT2 #(
		.INIT('h4)
	) name3527 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b3_last_row_reg[3]/P0001 ,
		_w4486_
	);
	LUT2 #(
		.INIT('h2)
	) name3528 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b3_last_row_reg[6]/P0001 ,
		_w4487_
	);
	LUT2 #(
		.INIT('h4)
	) name3529 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b3_last_row_reg[5]/P0001 ,
		_w4488_
	);
	LUT2 #(
		.INIT('h4)
	) name3530 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b3_last_row_reg[9]/P0001 ,
		_w4489_
	);
	LUT2 #(
		.INIT('h4)
	) name3531 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b3_last_row_reg[2]/P0001 ,
		_w4490_
	);
	LUT2 #(
		.INIT('h2)
	) name3532 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b3_last_row_reg[4]/P0001 ,
		_w4491_
	);
	LUT2 #(
		.INIT('h4)
	) name3533 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b3_last_row_reg[1]/P0001 ,
		_w4492_
	);
	LUT2 #(
		.INIT('h4)
	) name3534 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b3_last_row_reg[12]/P0001 ,
		_w4493_
	);
	LUT2 #(
		.INIT('h2)
	) name3535 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b3_last_row_reg[1]/P0001 ,
		_w4494_
	);
	LUT2 #(
		.INIT('h4)
	) name3536 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b3_last_row_reg[4]/P0001 ,
		_w4495_
	);
	LUT2 #(
		.INIT('h2)
	) name3537 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u1_b3_last_row_reg[0]/P0001 ,
		_w4496_
	);
	LUT2 #(
		.INIT('h2)
	) name3538 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b3_last_row_reg[8]/P0001 ,
		_w4497_
	);
	LUT2 #(
		.INIT('h4)
	) name3539 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b3_last_row_reg[11]/P0001 ,
		_w4498_
	);
	LUT2 #(
		.INIT('h4)
	) name3540 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b3_last_row_reg[8]/P0001 ,
		_w4499_
	);
	LUT2 #(
		.INIT('h2)
	) name3541 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b3_last_row_reg[7]/P0001 ,
		_w4500_
	);
	LUT2 #(
		.INIT('h4)
	) name3542 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b3_last_row_reg[7]/P0001 ,
		_w4501_
	);
	LUT2 #(
		.INIT('h4)
	) name3543 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b3_last_row_reg[6]/P0001 ,
		_w4502_
	);
	LUT2 #(
		.INIT('h2)
	) name3544 (
		_w3133_,
		_w4476_,
		_w4503_
	);
	LUT2 #(
		.INIT('h1)
	) name3545 (
		_w4477_,
		_w4478_,
		_w4504_
	);
	LUT2 #(
		.INIT('h1)
	) name3546 (
		_w4479_,
		_w4480_,
		_w4505_
	);
	LUT2 #(
		.INIT('h1)
	) name3547 (
		_w4481_,
		_w4485_,
		_w4506_
	);
	LUT2 #(
		.INIT('h1)
	) name3548 (
		_w4486_,
		_w4487_,
		_w4507_
	);
	LUT2 #(
		.INIT('h1)
	) name3549 (
		_w4488_,
		_w4489_,
		_w4508_
	);
	LUT2 #(
		.INIT('h1)
	) name3550 (
		_w4490_,
		_w4491_,
		_w4509_
	);
	LUT2 #(
		.INIT('h1)
	) name3551 (
		_w4492_,
		_w4493_,
		_w4510_
	);
	LUT2 #(
		.INIT('h1)
	) name3552 (
		_w4494_,
		_w4495_,
		_w4511_
	);
	LUT2 #(
		.INIT('h1)
	) name3553 (
		_w4496_,
		_w4497_,
		_w4512_
	);
	LUT2 #(
		.INIT('h1)
	) name3554 (
		_w4498_,
		_w4499_,
		_w4513_
	);
	LUT2 #(
		.INIT('h1)
	) name3555 (
		_w4500_,
		_w4501_,
		_w4514_
	);
	LUT2 #(
		.INIT('h4)
	) name3556 (
		_w4502_,
		_w4514_,
		_w4515_
	);
	LUT2 #(
		.INIT('h8)
	) name3557 (
		_w4512_,
		_w4513_,
		_w4516_
	);
	LUT2 #(
		.INIT('h8)
	) name3558 (
		_w4510_,
		_w4511_,
		_w4517_
	);
	LUT2 #(
		.INIT('h8)
	) name3559 (
		_w4508_,
		_w4509_,
		_w4518_
	);
	LUT2 #(
		.INIT('h8)
	) name3560 (
		_w4506_,
		_w4507_,
		_w4519_
	);
	LUT2 #(
		.INIT('h8)
	) name3561 (
		_w4504_,
		_w4505_,
		_w4520_
	);
	LUT2 #(
		.INIT('h4)
	) name3562 (
		_w4484_,
		_w4503_,
		_w4521_
	);
	LUT2 #(
		.INIT('h8)
	) name3563 (
		_w4520_,
		_w4521_,
		_w4522_
	);
	LUT2 #(
		.INIT('h8)
	) name3564 (
		_w4518_,
		_w4519_,
		_w4523_
	);
	LUT2 #(
		.INIT('h8)
	) name3565 (
		_w4516_,
		_w4517_,
		_w4524_
	);
	LUT2 #(
		.INIT('h8)
	) name3566 (
		_w4515_,
		_w4524_,
		_w4525_
	);
	LUT2 #(
		.INIT('h8)
	) name3567 (
		_w4522_,
		_w4523_,
		_w4526_
	);
	LUT2 #(
		.INIT('h8)
	) name3568 (
		_w4525_,
		_w4526_,
		_w4527_
	);
	LUT2 #(
		.INIT('h2)
	) name3569 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b2_last_row_reg[12]/P0001 ,
		_w4528_
	);
	LUT2 #(
		.INIT('h2)
	) name3570 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b2_last_row_reg[6]/P0001 ,
		_w4529_
	);
	LUT2 #(
		.INIT('h2)
	) name3571 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b2_last_row_reg[5]/P0001 ,
		_w4530_
	);
	LUT2 #(
		.INIT('h2)
	) name3572 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b2_last_row_reg[1]/P0001 ,
		_w4531_
	);
	LUT2 #(
		.INIT('h4)
	) name3573 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b2_last_row_reg[11]/P0001 ,
		_w4532_
	);
	LUT2 #(
		.INIT('h2)
	) name3574 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b2_last_row_reg[11]/P0001 ,
		_w4533_
	);
	LUT2 #(
		.INIT('h2)
	) name3575 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b2_last_row_reg[9]/P0001 ,
		_w4534_
	);
	LUT2 #(
		.INIT('h4)
	) name3576 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u1_b2_last_row_reg[10]/P0001 ,
		_w4535_
	);
	LUT2 #(
		.INIT('h4)
	) name3577 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b2_last_row_reg[1]/P0001 ,
		_w4536_
	);
	LUT2 #(
		.INIT('h4)
	) name3578 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b2_last_row_reg[6]/P0001 ,
		_w4537_
	);
	LUT2 #(
		.INIT('h4)
	) name3579 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b2_last_row_reg[12]/P0001 ,
		_w4538_
	);
	LUT2 #(
		.INIT('h4)
	) name3580 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b2_last_row_reg[5]/P0001 ,
		_w4539_
	);
	LUT2 #(
		.INIT('h4)
	) name3581 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b2_last_row_reg[9]/P0001 ,
		_w4540_
	);
	LUT2 #(
		.INIT('h2)
	) name3582 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u1_b2_last_row_reg[10]/P0001 ,
		_w4541_
	);
	LUT2 #(
		.INIT('h2)
	) name3583 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b2_last_row_reg[4]/P0001 ,
		_w4542_
	);
	LUT2 #(
		.INIT('h4)
	) name3584 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b2_last_row_reg[7]/P0001 ,
		_w4543_
	);
	LUT2 #(
		.INIT('h2)
	) name3585 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b2_last_row_reg[2]/P0001 ,
		_w4544_
	);
	LUT2 #(
		.INIT('h2)
	) name3586 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b2_last_row_reg[7]/P0001 ,
		_w4545_
	);
	LUT2 #(
		.INIT('h2)
	) name3587 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u1_b2_last_row_reg[0]/P0001 ,
		_w4546_
	);
	LUT2 #(
		.INIT('h4)
	) name3588 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b2_last_row_reg[4]/P0001 ,
		_w4547_
	);
	LUT2 #(
		.INIT('h4)
	) name3589 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b2_last_row_reg[2]/P0001 ,
		_w4548_
	);
	LUT2 #(
		.INIT('h2)
	) name3590 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b2_last_row_reg[8]/P0001 ,
		_w4549_
	);
	LUT2 #(
		.INIT('h4)
	) name3591 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u1_b2_last_row_reg[0]/P0001 ,
		_w4550_
	);
	LUT2 #(
		.INIT('h2)
	) name3592 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b2_last_row_reg[3]/P0001 ,
		_w4551_
	);
	LUT2 #(
		.INIT('h4)
	) name3593 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b2_last_row_reg[8]/P0001 ,
		_w4552_
	);
	LUT2 #(
		.INIT('h4)
	) name3594 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b2_last_row_reg[3]/P0001 ,
		_w4553_
	);
	LUT2 #(
		.INIT('h2)
	) name3595 (
		_w3103_,
		_w4528_,
		_w4554_
	);
	LUT2 #(
		.INIT('h1)
	) name3596 (
		_w4529_,
		_w4530_,
		_w4555_
	);
	LUT2 #(
		.INIT('h1)
	) name3597 (
		_w4531_,
		_w4532_,
		_w4556_
	);
	LUT2 #(
		.INIT('h1)
	) name3598 (
		_w4533_,
		_w4534_,
		_w4557_
	);
	LUT2 #(
		.INIT('h1)
	) name3599 (
		_w4535_,
		_w4536_,
		_w4558_
	);
	LUT2 #(
		.INIT('h1)
	) name3600 (
		_w4537_,
		_w4538_,
		_w4559_
	);
	LUT2 #(
		.INIT('h1)
	) name3601 (
		_w4539_,
		_w4540_,
		_w4560_
	);
	LUT2 #(
		.INIT('h1)
	) name3602 (
		_w4541_,
		_w4542_,
		_w4561_
	);
	LUT2 #(
		.INIT('h1)
	) name3603 (
		_w4543_,
		_w4544_,
		_w4562_
	);
	LUT2 #(
		.INIT('h1)
	) name3604 (
		_w4545_,
		_w4546_,
		_w4563_
	);
	LUT2 #(
		.INIT('h1)
	) name3605 (
		_w4547_,
		_w4548_,
		_w4564_
	);
	LUT2 #(
		.INIT('h1)
	) name3606 (
		_w4549_,
		_w4550_,
		_w4565_
	);
	LUT2 #(
		.INIT('h1)
	) name3607 (
		_w4551_,
		_w4552_,
		_w4566_
	);
	LUT2 #(
		.INIT('h4)
	) name3608 (
		_w4553_,
		_w4566_,
		_w4567_
	);
	LUT2 #(
		.INIT('h8)
	) name3609 (
		_w4564_,
		_w4565_,
		_w4568_
	);
	LUT2 #(
		.INIT('h8)
	) name3610 (
		_w4562_,
		_w4563_,
		_w4569_
	);
	LUT2 #(
		.INIT('h8)
	) name3611 (
		_w4560_,
		_w4561_,
		_w4570_
	);
	LUT2 #(
		.INIT('h8)
	) name3612 (
		_w4558_,
		_w4559_,
		_w4571_
	);
	LUT2 #(
		.INIT('h8)
	) name3613 (
		_w4556_,
		_w4557_,
		_w4572_
	);
	LUT2 #(
		.INIT('h8)
	) name3614 (
		_w4554_,
		_w4555_,
		_w4573_
	);
	LUT2 #(
		.INIT('h8)
	) name3615 (
		_w4572_,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h8)
	) name3616 (
		_w4570_,
		_w4571_,
		_w4575_
	);
	LUT2 #(
		.INIT('h8)
	) name3617 (
		_w4568_,
		_w4569_,
		_w4576_
	);
	LUT2 #(
		.INIT('h8)
	) name3618 (
		_w4567_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h8)
	) name3619 (
		_w4574_,
		_w4575_,
		_w4578_
	);
	LUT2 #(
		.INIT('h8)
	) name3620 (
		_w4577_,
		_w4578_,
		_w4579_
	);
	LUT2 #(
		.INIT('h4)
	) name3621 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u1_b0_last_row_reg[10]/P0001 ,
		_w4580_
	);
	LUT2 #(
		.INIT('h1)
	) name3622 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b0_last_row_reg[7]/P0001 ,
		_w4581_
	);
	LUT2 #(
		.INIT('h8)
	) name3623 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b0_last_row_reg[7]/P0001 ,
		_w4582_
	);
	LUT2 #(
		.INIT('h1)
	) name3624 (
		_w4581_,
		_w4582_,
		_w4583_
	);
	LUT2 #(
		.INIT('h2)
	) name3625 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b0_last_row_reg[12]/P0001 ,
		_w4584_
	);
	LUT2 #(
		.INIT('h2)
	) name3626 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b0_last_row_reg[4]/P0001 ,
		_w4585_
	);
	LUT2 #(
		.INIT('h1)
	) name3627 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u1_b0_last_row_reg[0]/P0001 ,
		_w4586_
	);
	LUT2 #(
		.INIT('h8)
	) name3628 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u1_b0_last_row_reg[0]/P0001 ,
		_w4587_
	);
	LUT2 #(
		.INIT('h1)
	) name3629 (
		_w4586_,
		_w4587_,
		_w4588_
	);
	LUT2 #(
		.INIT('h4)
	) name3630 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b0_last_row_reg[8]/P0001 ,
		_w4589_
	);
	LUT2 #(
		.INIT('h4)
	) name3631 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b0_last_row_reg[3]/P0001 ,
		_w4590_
	);
	LUT2 #(
		.INIT('h4)
	) name3632 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b0_last_row_reg[12]/P0001 ,
		_w4591_
	);
	LUT2 #(
		.INIT('h2)
	) name3633 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b0_last_row_reg[8]/P0001 ,
		_w4592_
	);
	LUT2 #(
		.INIT('h4)
	) name3634 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b0_last_row_reg[6]/P0001 ,
		_w4593_
	);
	LUT2 #(
		.INIT('h4)
	) name3635 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b0_last_row_reg[5]/P0001 ,
		_w4594_
	);
	LUT2 #(
		.INIT('h4)
	) name3636 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b0_last_row_reg[11]/P0001 ,
		_w4595_
	);
	LUT2 #(
		.INIT('h4)
	) name3637 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b0_last_row_reg[1]/P0001 ,
		_w4596_
	);
	LUT2 #(
		.INIT('h4)
	) name3638 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b0_last_row_reg[2]/P0001 ,
		_w4597_
	);
	LUT2 #(
		.INIT('h2)
	) name3639 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b0_last_row_reg[6]/P0001 ,
		_w4598_
	);
	LUT2 #(
		.INIT('h2)
	) name3640 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b0_last_row_reg[11]/P0001 ,
		_w4599_
	);
	LUT2 #(
		.INIT('h2)
	) name3641 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b0_last_row_reg[3]/P0001 ,
		_w4600_
	);
	LUT2 #(
		.INIT('h4)
	) name3642 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b0_last_row_reg[9]/P0001 ,
		_w4601_
	);
	LUT2 #(
		.INIT('h2)
	) name3643 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b0_last_row_reg[2]/P0001 ,
		_w4602_
	);
	LUT2 #(
		.INIT('h2)
	) name3644 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b0_last_row_reg[9]/P0001 ,
		_w4603_
	);
	LUT2 #(
		.INIT('h2)
	) name3645 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u1_b0_last_row_reg[10]/P0001 ,
		_w4604_
	);
	LUT2 #(
		.INIT('h2)
	) name3646 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b0_last_row_reg[1]/P0001 ,
		_w4605_
	);
	LUT2 #(
		.INIT('h2)
	) name3647 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b0_last_row_reg[5]/P0001 ,
		_w4606_
	);
	LUT2 #(
		.INIT('h1)
	) name3648 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		_w4607_
	);
	LUT2 #(
		.INIT('h4)
	) name3649 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b0_last_row_reg[4]/P0001 ,
		_w4608_
	);
	LUT2 #(
		.INIT('h1)
	) name3650 (
		_w4580_,
		_w4584_,
		_w4609_
	);
	LUT2 #(
		.INIT('h1)
	) name3651 (
		_w4585_,
		_w4589_,
		_w4610_
	);
	LUT2 #(
		.INIT('h1)
	) name3652 (
		_w4590_,
		_w4591_,
		_w4611_
	);
	LUT2 #(
		.INIT('h1)
	) name3653 (
		_w4592_,
		_w4593_,
		_w4612_
	);
	LUT2 #(
		.INIT('h1)
	) name3654 (
		_w4594_,
		_w4595_,
		_w4613_
	);
	LUT2 #(
		.INIT('h1)
	) name3655 (
		_w4596_,
		_w4597_,
		_w4614_
	);
	LUT2 #(
		.INIT('h1)
	) name3656 (
		_w4598_,
		_w4599_,
		_w4615_
	);
	LUT2 #(
		.INIT('h1)
	) name3657 (
		_w4600_,
		_w4601_,
		_w4616_
	);
	LUT2 #(
		.INIT('h1)
	) name3658 (
		_w4602_,
		_w4603_,
		_w4617_
	);
	LUT2 #(
		.INIT('h1)
	) name3659 (
		_w4604_,
		_w4605_,
		_w4618_
	);
	LUT2 #(
		.INIT('h4)
	) name3660 (
		_w4606_,
		_w4607_,
		_w4619_
	);
	LUT2 #(
		.INIT('h4)
	) name3661 (
		_w4608_,
		_w4619_,
		_w4620_
	);
	LUT2 #(
		.INIT('h8)
	) name3662 (
		_w4617_,
		_w4618_,
		_w4621_
	);
	LUT2 #(
		.INIT('h8)
	) name3663 (
		_w4615_,
		_w4616_,
		_w4622_
	);
	LUT2 #(
		.INIT('h8)
	) name3664 (
		_w4613_,
		_w4614_,
		_w4623_
	);
	LUT2 #(
		.INIT('h8)
	) name3665 (
		_w4611_,
		_w4612_,
		_w4624_
	);
	LUT2 #(
		.INIT('h8)
	) name3666 (
		_w4609_,
		_w4610_,
		_w4625_
	);
	LUT2 #(
		.INIT('h1)
	) name3667 (
		_w4583_,
		_w4588_,
		_w4626_
	);
	LUT2 #(
		.INIT('h8)
	) name3668 (
		_w4625_,
		_w4626_,
		_w4627_
	);
	LUT2 #(
		.INIT('h8)
	) name3669 (
		_w4623_,
		_w4624_,
		_w4628_
	);
	LUT2 #(
		.INIT('h8)
	) name3670 (
		_w4621_,
		_w4622_,
		_w4629_
	);
	LUT2 #(
		.INIT('h8)
	) name3671 (
		_w4620_,
		_w4629_,
		_w4630_
	);
	LUT2 #(
		.INIT('h8)
	) name3672 (
		_w4627_,
		_w4628_,
		_w4631_
	);
	LUT2 #(
		.INIT('h8)
	) name3673 (
		_w4630_,
		_w4631_,
		_w4632_
	);
	LUT2 #(
		.INIT('h2)
	) name3674 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b1_last_row_reg[11]/P0001 ,
		_w4633_
	);
	LUT2 #(
		.INIT('h2)
	) name3675 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b1_last_row_reg[2]/P0001 ,
		_w4634_
	);
	LUT2 #(
		.INIT('h2)
	) name3676 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u1_b1_last_row_reg[0]/P0001 ,
		_w4635_
	);
	LUT2 #(
		.INIT('h4)
	) name3677 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b1_last_row_reg[7]/P0001 ,
		_w4636_
	);
	LUT2 #(
		.INIT('h4)
	) name3678 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b1_last_row_reg[11]/P0001 ,
		_w4637_
	);
	LUT2 #(
		.INIT('h2)
	) name3679 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b1_last_row_reg[8]/P0001 ,
		_w4638_
	);
	LUT2 #(
		.INIT('h2)
	) name3680 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u1_b1_last_row_reg[10]/P0001 ,
		_w4639_
	);
	LUT2 #(
		.INIT('h2)
	) name3681 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b1_last_row_reg[4]/P0001 ,
		_w4640_
	);
	LUT2 #(
		.INIT('h4)
	) name3682 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u1_b1_last_row_reg[0]/P0001 ,
		_w4641_
	);
	LUT2 #(
		.INIT('h2)
	) name3683 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b1_last_row_reg[7]/P0001 ,
		_w4642_
	);
	LUT2 #(
		.INIT('h4)
	) name3684 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b1_last_row_reg[4]/P0001 ,
		_w4643_
	);
	LUT2 #(
		.INIT('h4)
	) name3685 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b1_last_row_reg[1]/P0001 ,
		_w4644_
	);
	LUT2 #(
		.INIT('h4)
	) name3686 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b1_last_row_reg[8]/P0001 ,
		_w4645_
	);
	LUT2 #(
		.INIT('h4)
	) name3687 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b1_last_row_reg[9]/P0001 ,
		_w4646_
	);
	LUT2 #(
		.INIT('h4)
	) name3688 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b1_last_row_reg[2]/P0001 ,
		_w4647_
	);
	LUT2 #(
		.INIT('h2)
	) name3689 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b1_last_row_reg[9]/P0001 ,
		_w4648_
	);
	LUT2 #(
		.INIT('h4)
	) name3690 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b1_last_row_reg[5]/P0001 ,
		_w4649_
	);
	LUT2 #(
		.INIT('h4)
	) name3691 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u1_b1_last_row_reg[10]/P0001 ,
		_w4650_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b1_last_row_reg[6]/P0001 ,
		_w4651_
	);
	LUT2 #(
		.INIT('h2)
	) name3693 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b1_last_row_reg[1]/P0001 ,
		_w4652_
	);
	LUT2 #(
		.INIT('h4)
	) name3694 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b1_last_row_reg[6]/P0001 ,
		_w4653_
	);
	LUT2 #(
		.INIT('h2)
	) name3695 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b1_last_row_reg[5]/P0001 ,
		_w4654_
	);
	LUT2 #(
		.INIT('h4)
	) name3696 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b1_last_row_reg[12]/P0001 ,
		_w4655_
	);
	LUT2 #(
		.INIT('h2)
	) name3697 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b1_last_row_reg[12]/P0001 ,
		_w4656_
	);
	LUT2 #(
		.INIT('h2)
	) name3698 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b1_last_row_reg[3]/P0001 ,
		_w4657_
	);
	LUT2 #(
		.INIT('h4)
	) name3699 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b1_last_row_reg[3]/P0001 ,
		_w4658_
	);
	LUT2 #(
		.INIT('h2)
	) name3700 (
		_w3049_,
		_w4633_,
		_w4659_
	);
	LUT2 #(
		.INIT('h1)
	) name3701 (
		_w4634_,
		_w4635_,
		_w4660_
	);
	LUT2 #(
		.INIT('h1)
	) name3702 (
		_w4636_,
		_w4637_,
		_w4661_
	);
	LUT2 #(
		.INIT('h1)
	) name3703 (
		_w4638_,
		_w4639_,
		_w4662_
	);
	LUT2 #(
		.INIT('h1)
	) name3704 (
		_w4640_,
		_w4641_,
		_w4663_
	);
	LUT2 #(
		.INIT('h1)
	) name3705 (
		_w4642_,
		_w4643_,
		_w4664_
	);
	LUT2 #(
		.INIT('h1)
	) name3706 (
		_w4644_,
		_w4645_,
		_w4665_
	);
	LUT2 #(
		.INIT('h1)
	) name3707 (
		_w4646_,
		_w4647_,
		_w4666_
	);
	LUT2 #(
		.INIT('h1)
	) name3708 (
		_w4648_,
		_w4649_,
		_w4667_
	);
	LUT2 #(
		.INIT('h1)
	) name3709 (
		_w4650_,
		_w4651_,
		_w4668_
	);
	LUT2 #(
		.INIT('h1)
	) name3710 (
		_w4652_,
		_w4653_,
		_w4669_
	);
	LUT2 #(
		.INIT('h1)
	) name3711 (
		_w4654_,
		_w4655_,
		_w4670_
	);
	LUT2 #(
		.INIT('h1)
	) name3712 (
		_w4656_,
		_w4657_,
		_w4671_
	);
	LUT2 #(
		.INIT('h4)
	) name3713 (
		_w4658_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h8)
	) name3714 (
		_w4669_,
		_w4670_,
		_w4673_
	);
	LUT2 #(
		.INIT('h8)
	) name3715 (
		_w4667_,
		_w4668_,
		_w4674_
	);
	LUT2 #(
		.INIT('h8)
	) name3716 (
		_w4665_,
		_w4666_,
		_w4675_
	);
	LUT2 #(
		.INIT('h8)
	) name3717 (
		_w4663_,
		_w4664_,
		_w4676_
	);
	LUT2 #(
		.INIT('h8)
	) name3718 (
		_w4661_,
		_w4662_,
		_w4677_
	);
	LUT2 #(
		.INIT('h8)
	) name3719 (
		_w4659_,
		_w4660_,
		_w4678_
	);
	LUT2 #(
		.INIT('h8)
	) name3720 (
		_w4677_,
		_w4678_,
		_w4679_
	);
	LUT2 #(
		.INIT('h8)
	) name3721 (
		_w4675_,
		_w4676_,
		_w4680_
	);
	LUT2 #(
		.INIT('h8)
	) name3722 (
		_w4673_,
		_w4674_,
		_w4681_
	);
	LUT2 #(
		.INIT('h8)
	) name3723 (
		_w4672_,
		_w4681_,
		_w4682_
	);
	LUT2 #(
		.INIT('h8)
	) name3724 (
		_w4679_,
		_w4680_,
		_w4683_
	);
	LUT2 #(
		.INIT('h8)
	) name3725 (
		_w4682_,
		_w4683_,
		_w4684_
	);
	LUT2 #(
		.INIT('h1)
	) name3726 (
		_w4527_,
		_w4579_,
		_w4685_
	);
	LUT2 #(
		.INIT('h1)
	) name3727 (
		_w4632_,
		_w4684_,
		_w4686_
	);
	LUT2 #(
		.INIT('h8)
	) name3728 (
		_w4685_,
		_w4686_,
		_w4687_
	);
	LUT2 #(
		.INIT('h1)
	) name3729 (
		_w1676_,
		_w4687_,
		_w4688_
	);
	LUT2 #(
		.INIT('h2)
	) name3730 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b2_last_row_reg[7]/P0001 ,
		_w4689_
	);
	LUT2 #(
		.INIT('h1)
	) name3731 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b2_last_row_reg[4]/P0001 ,
		_w4690_
	);
	LUT2 #(
		.INIT('h8)
	) name3732 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b2_last_row_reg[4]/P0001 ,
		_w4691_
	);
	LUT2 #(
		.INIT('h1)
	) name3733 (
		_w4690_,
		_w4691_,
		_w4692_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b2_last_row_reg[6]/P0001 ,
		_w4693_
	);
	LUT2 #(
		.INIT('h2)
	) name3735 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b2_last_row_reg[2]/P0001 ,
		_w4694_
	);
	LUT2 #(
		.INIT('h1)
	) name3736 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u0_b2_last_row_reg[0]/P0001 ,
		_w4695_
	);
	LUT2 #(
		.INIT('h8)
	) name3737 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u0_b2_last_row_reg[0]/P0001 ,
		_w4696_
	);
	LUT2 #(
		.INIT('h1)
	) name3738 (
		_w4695_,
		_w4696_,
		_w4697_
	);
	LUT2 #(
		.INIT('h4)
	) name3739 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b2_last_row_reg[6]/P0001 ,
		_w4698_
	);
	LUT2 #(
		.INIT('h4)
	) name3740 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b2_last_row_reg[7]/P0001 ,
		_w4699_
	);
	LUT2 #(
		.INIT('h4)
	) name3741 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b2_last_row_reg[3]/P0001 ,
		_w4700_
	);
	LUT2 #(
		.INIT('h2)
	) name3742 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b2_last_row_reg[1]/P0001 ,
		_w4701_
	);
	LUT2 #(
		.INIT('h2)
	) name3743 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u0_b2_last_row_reg[12]/P0001 ,
		_w4702_
	);
	LUT2 #(
		.INIT('h4)
	) name3744 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u0_b2_last_row_reg[12]/P0001 ,
		_w4703_
	);
	LUT2 #(
		.INIT('h4)
	) name3745 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b2_last_row_reg[5]/P0001 ,
		_w4704_
	);
	LUT2 #(
		.INIT('h2)
	) name3746 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u0_b2_last_row_reg[10]/P0001 ,
		_w4705_
	);
	LUT2 #(
		.INIT('h4)
	) name3747 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b2_last_row_reg[2]/P0001 ,
		_w4706_
	);
	LUT2 #(
		.INIT('h4)
	) name3748 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b2_last_row_reg[1]/P0001 ,
		_w4707_
	);
	LUT2 #(
		.INIT('h4)
	) name3749 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b2_last_row_reg[9]/P0001 ,
		_w4708_
	);
	LUT2 #(
		.INIT('h2)
	) name3750 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b2_last_row_reg[3]/P0001 ,
		_w4709_
	);
	LUT2 #(
		.INIT('h4)
	) name3751 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u0_b2_last_row_reg[10]/P0001 ,
		_w4710_
	);
	LUT2 #(
		.INIT('h2)
	) name3752 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b2_last_row_reg[9]/P0001 ,
		_w4711_
	);
	LUT2 #(
		.INIT('h4)
	) name3753 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b2_last_row_reg[8]/P0001 ,
		_w4712_
	);
	LUT2 #(
		.INIT('h2)
	) name3754 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b2_last_row_reg[8]/P0001 ,
		_w4713_
	);
	LUT2 #(
		.INIT('h2)
	) name3755 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b2_last_row_reg[11]/P0001 ,
		_w4714_
	);
	LUT2 #(
		.INIT('h4)
	) name3756 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b2_last_row_reg[11]/P0001 ,
		_w4715_
	);
	LUT2 #(
		.INIT('h2)
	) name3757 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b2_last_row_reg[5]/P0001 ,
		_w4716_
	);
	LUT2 #(
		.INIT('h2)
	) name3758 (
		_w3103_,
		_w4689_,
		_w4717_
	);
	LUT2 #(
		.INIT('h1)
	) name3759 (
		_w4693_,
		_w4694_,
		_w4718_
	);
	LUT2 #(
		.INIT('h1)
	) name3760 (
		_w4698_,
		_w4699_,
		_w4719_
	);
	LUT2 #(
		.INIT('h1)
	) name3761 (
		_w4700_,
		_w4701_,
		_w4720_
	);
	LUT2 #(
		.INIT('h1)
	) name3762 (
		_w4702_,
		_w4703_,
		_w4721_
	);
	LUT2 #(
		.INIT('h1)
	) name3763 (
		_w4704_,
		_w4705_,
		_w4722_
	);
	LUT2 #(
		.INIT('h1)
	) name3764 (
		_w4706_,
		_w4707_,
		_w4723_
	);
	LUT2 #(
		.INIT('h1)
	) name3765 (
		_w4708_,
		_w4709_,
		_w4724_
	);
	LUT2 #(
		.INIT('h1)
	) name3766 (
		_w4710_,
		_w4711_,
		_w4725_
	);
	LUT2 #(
		.INIT('h1)
	) name3767 (
		_w4712_,
		_w4713_,
		_w4726_
	);
	LUT2 #(
		.INIT('h1)
	) name3768 (
		_w4714_,
		_w4715_,
		_w4727_
	);
	LUT2 #(
		.INIT('h4)
	) name3769 (
		_w4716_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h8)
	) name3770 (
		_w4725_,
		_w4726_,
		_w4729_
	);
	LUT2 #(
		.INIT('h8)
	) name3771 (
		_w4723_,
		_w4724_,
		_w4730_
	);
	LUT2 #(
		.INIT('h8)
	) name3772 (
		_w4721_,
		_w4722_,
		_w4731_
	);
	LUT2 #(
		.INIT('h8)
	) name3773 (
		_w4719_,
		_w4720_,
		_w4732_
	);
	LUT2 #(
		.INIT('h8)
	) name3774 (
		_w4717_,
		_w4718_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name3775 (
		_w4692_,
		_w4697_,
		_w4734_
	);
	LUT2 #(
		.INIT('h8)
	) name3776 (
		_w4733_,
		_w4734_,
		_w4735_
	);
	LUT2 #(
		.INIT('h8)
	) name3777 (
		_w4731_,
		_w4732_,
		_w4736_
	);
	LUT2 #(
		.INIT('h8)
	) name3778 (
		_w4729_,
		_w4730_,
		_w4737_
	);
	LUT2 #(
		.INIT('h8)
	) name3779 (
		_w4728_,
		_w4737_,
		_w4738_
	);
	LUT2 #(
		.INIT('h8)
	) name3780 (
		_w4735_,
		_w4736_,
		_w4739_
	);
	LUT2 #(
		.INIT('h8)
	) name3781 (
		_w4738_,
		_w4739_,
		_w4740_
	);
	LUT2 #(
		.INIT('h4)
	) name3782 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b1_last_row_reg[1]/P0001 ,
		_w4741_
	);
	LUT2 #(
		.INIT('h2)
	) name3783 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b1_last_row_reg[9]/P0001 ,
		_w4742_
	);
	LUT2 #(
		.INIT('h2)
	) name3784 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b1_last_row_reg[4]/P0001 ,
		_w4743_
	);
	LUT2 #(
		.INIT('h2)
	) name3785 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b1_last_row_reg[5]/P0001 ,
		_w4744_
	);
	LUT2 #(
		.INIT('h4)
	) name3786 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b1_last_row_reg[9]/P0001 ,
		_w4745_
	);
	LUT2 #(
		.INIT('h2)
	) name3787 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u0_b1_last_row_reg[12]/P0001 ,
		_w4746_
	);
	LUT2 #(
		.INIT('h4)
	) name3788 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b1_last_row_reg[6]/P0001 ,
		_w4747_
	);
	LUT2 #(
		.INIT('h2)
	) name3789 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b1_last_row_reg[7]/P0001 ,
		_w4748_
	);
	LUT2 #(
		.INIT('h4)
	) name3790 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b1_last_row_reg[5]/P0001 ,
		_w4749_
	);
	LUT2 #(
		.INIT('h4)
	) name3791 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b1_last_row_reg[4]/P0001 ,
		_w4750_
	);
	LUT2 #(
		.INIT('h2)
	) name3792 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b1_last_row_reg[2]/P0001 ,
		_w4751_
	);
	LUT2 #(
		.INIT('h2)
	) name3793 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u0_b1_last_row_reg[10]/P0001 ,
		_w4752_
	);
	LUT2 #(
		.INIT('h4)
	) name3794 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b1_last_row_reg[2]/P0001 ,
		_w4753_
	);
	LUT2 #(
		.INIT('h4)
	) name3795 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b1_last_row_reg[8]/P0001 ,
		_w4754_
	);
	LUT2 #(
		.INIT('h2)
	) name3796 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u0_b1_last_row_reg[0]/P0001 ,
		_w4755_
	);
	LUT2 #(
		.INIT('h4)
	) name3797 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b1_last_row_reg[3]/P0001 ,
		_w4756_
	);
	LUT2 #(
		.INIT('h2)
	) name3798 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b1_last_row_reg[8]/P0001 ,
		_w4757_
	);
	LUT2 #(
		.INIT('h4)
	) name3799 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u0_b1_last_row_reg[10]/P0001 ,
		_w4758_
	);
	LUT2 #(
		.INIT('h4)
	) name3800 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u0_b1_last_row_reg[0]/P0001 ,
		_w4759_
	);
	LUT2 #(
		.INIT('h4)
	) name3801 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b1_last_row_reg[7]/P0001 ,
		_w4760_
	);
	LUT2 #(
		.INIT('h2)
	) name3802 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b1_last_row_reg[1]/P0001 ,
		_w4761_
	);
	LUT2 #(
		.INIT('h4)
	) name3803 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b1_last_row_reg[11]/P0001 ,
		_w4762_
	);
	LUT2 #(
		.INIT('h2)
	) name3804 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b1_last_row_reg[11]/P0001 ,
		_w4763_
	);
	LUT2 #(
		.INIT('h2)
	) name3805 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b1_last_row_reg[6]/P0001 ,
		_w4764_
	);
	LUT2 #(
		.INIT('h4)
	) name3806 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u0_b1_last_row_reg[12]/P0001 ,
		_w4765_
	);
	LUT2 #(
		.INIT('h2)
	) name3807 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b1_last_row_reg[3]/P0001 ,
		_w4766_
	);
	LUT2 #(
		.INIT('h2)
	) name3808 (
		_w3049_,
		_w4741_,
		_w4767_
	);
	LUT2 #(
		.INIT('h1)
	) name3809 (
		_w4742_,
		_w4743_,
		_w4768_
	);
	LUT2 #(
		.INIT('h1)
	) name3810 (
		_w4744_,
		_w4745_,
		_w4769_
	);
	LUT2 #(
		.INIT('h1)
	) name3811 (
		_w4746_,
		_w4747_,
		_w4770_
	);
	LUT2 #(
		.INIT('h1)
	) name3812 (
		_w4748_,
		_w4749_,
		_w4771_
	);
	LUT2 #(
		.INIT('h1)
	) name3813 (
		_w4750_,
		_w4751_,
		_w4772_
	);
	LUT2 #(
		.INIT('h1)
	) name3814 (
		_w4752_,
		_w4753_,
		_w4773_
	);
	LUT2 #(
		.INIT('h1)
	) name3815 (
		_w4754_,
		_w4755_,
		_w4774_
	);
	LUT2 #(
		.INIT('h1)
	) name3816 (
		_w4756_,
		_w4757_,
		_w4775_
	);
	LUT2 #(
		.INIT('h1)
	) name3817 (
		_w4758_,
		_w4759_,
		_w4776_
	);
	LUT2 #(
		.INIT('h1)
	) name3818 (
		_w4760_,
		_w4761_,
		_w4777_
	);
	LUT2 #(
		.INIT('h1)
	) name3819 (
		_w4762_,
		_w4763_,
		_w4778_
	);
	LUT2 #(
		.INIT('h1)
	) name3820 (
		_w4764_,
		_w4765_,
		_w4779_
	);
	LUT2 #(
		.INIT('h4)
	) name3821 (
		_w4766_,
		_w4779_,
		_w4780_
	);
	LUT2 #(
		.INIT('h8)
	) name3822 (
		_w4777_,
		_w4778_,
		_w4781_
	);
	LUT2 #(
		.INIT('h8)
	) name3823 (
		_w4775_,
		_w4776_,
		_w4782_
	);
	LUT2 #(
		.INIT('h8)
	) name3824 (
		_w4773_,
		_w4774_,
		_w4783_
	);
	LUT2 #(
		.INIT('h8)
	) name3825 (
		_w4771_,
		_w4772_,
		_w4784_
	);
	LUT2 #(
		.INIT('h8)
	) name3826 (
		_w4769_,
		_w4770_,
		_w4785_
	);
	LUT2 #(
		.INIT('h8)
	) name3827 (
		_w4767_,
		_w4768_,
		_w4786_
	);
	LUT2 #(
		.INIT('h8)
	) name3828 (
		_w4785_,
		_w4786_,
		_w4787_
	);
	LUT2 #(
		.INIT('h8)
	) name3829 (
		_w4783_,
		_w4784_,
		_w4788_
	);
	LUT2 #(
		.INIT('h8)
	) name3830 (
		_w4781_,
		_w4782_,
		_w4789_
	);
	LUT2 #(
		.INIT('h8)
	) name3831 (
		_w4780_,
		_w4789_,
		_w4790_
	);
	LUT2 #(
		.INIT('h8)
	) name3832 (
		_w4787_,
		_w4788_,
		_w4791_
	);
	LUT2 #(
		.INIT('h8)
	) name3833 (
		_w4790_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h4)
	) name3834 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b0_last_row_reg[5]/P0001 ,
		_w4793_
	);
	LUT2 #(
		.INIT('h4)
	) name3835 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b0_last_row_reg[8]/P0001 ,
		_w4794_
	);
	LUT2 #(
		.INIT('h4)
	) name3836 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b0_last_row_reg[4]/P0001 ,
		_w4795_
	);
	LUT2 #(
		.INIT('h2)
	) name3837 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b0_last_row_reg[7]/P0001 ,
		_w4796_
	);
	LUT2 #(
		.INIT('h2)
	) name3838 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b0_last_row_reg[1]/P0001 ,
		_w4797_
	);
	LUT2 #(
		.INIT('h2)
	) name3839 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b0_last_row_reg[8]/P0001 ,
		_w4798_
	);
	LUT2 #(
		.INIT('h4)
	) name3840 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b0_last_row_reg[11]/P0001 ,
		_w4799_
	);
	LUT2 #(
		.INIT('h2)
	) name3841 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b0_last_row_reg[3]/P0001 ,
		_w4800_
	);
	LUT2 #(
		.INIT('h2)
	) name3842 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b0_last_row_reg[4]/P0001 ,
		_w4801_
	);
	LUT2 #(
		.INIT('h2)
	) name3843 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b0_last_row_reg[9]/P0001 ,
		_w4802_
	);
	LUT2 #(
		.INIT('h4)
	) name3844 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b0_last_row_reg[7]/P0001 ,
		_w4803_
	);
	LUT2 #(
		.INIT('h4)
	) name3845 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b0_last_row_reg[3]/P0001 ,
		_w4804_
	);
	LUT2 #(
		.INIT('h4)
	) name3846 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b0_last_row_reg[1]/P0001 ,
		_w4805_
	);
	LUT2 #(
		.INIT('h2)
	) name3847 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u0_b0_last_row_reg[0]/P0001 ,
		_w4806_
	);
	LUT2 #(
		.INIT('h2)
	) name3848 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b0_last_row_reg[2]/P0001 ,
		_w4807_
	);
	LUT2 #(
		.INIT('h4)
	) name3849 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u0_b0_last_row_reg[10]/P0001 ,
		_w4808_
	);
	LUT2 #(
		.INIT('h2)
	) name3850 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b0_last_row_reg[6]/P0001 ,
		_w4809_
	);
	LUT2 #(
		.INIT('h4)
	) name3851 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b0_last_row_reg[2]/P0001 ,
		_w4810_
	);
	LUT2 #(
		.INIT('h4)
	) name3852 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b0_last_row_reg[9]/P0001 ,
		_w4811_
	);
	LUT2 #(
		.INIT('h2)
	) name3853 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u0_b0_last_row_reg[10]/P0001 ,
		_w4812_
	);
	LUT2 #(
		.INIT('h2)
	) name3854 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b0_last_row_reg[11]/P0001 ,
		_w4813_
	);
	LUT2 #(
		.INIT('h4)
	) name3855 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u0_b0_last_row_reg[0]/P0001 ,
		_w4814_
	);
	LUT2 #(
		.INIT('h4)
	) name3856 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b0_last_row_reg[6]/P0001 ,
		_w4815_
	);
	LUT2 #(
		.INIT('h2)
	) name3857 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u0_b0_last_row_reg[12]/P0001 ,
		_w4816_
	);
	LUT2 #(
		.INIT('h2)
	) name3858 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b0_last_row_reg[5]/P0001 ,
		_w4817_
	);
	LUT2 #(
		.INIT('h4)
	) name3859 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u0_b0_last_row_reg[12]/P0001 ,
		_w4818_
	);
	LUT2 #(
		.INIT('h2)
	) name3860 (
		_w4607_,
		_w4793_,
		_w4819_
	);
	LUT2 #(
		.INIT('h1)
	) name3861 (
		_w4794_,
		_w4795_,
		_w4820_
	);
	LUT2 #(
		.INIT('h1)
	) name3862 (
		_w4796_,
		_w4797_,
		_w4821_
	);
	LUT2 #(
		.INIT('h1)
	) name3863 (
		_w4798_,
		_w4799_,
		_w4822_
	);
	LUT2 #(
		.INIT('h1)
	) name3864 (
		_w4800_,
		_w4801_,
		_w4823_
	);
	LUT2 #(
		.INIT('h1)
	) name3865 (
		_w4802_,
		_w4803_,
		_w4824_
	);
	LUT2 #(
		.INIT('h1)
	) name3866 (
		_w4804_,
		_w4805_,
		_w4825_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w4806_,
		_w4807_,
		_w4826_
	);
	LUT2 #(
		.INIT('h1)
	) name3868 (
		_w4808_,
		_w4809_,
		_w4827_
	);
	LUT2 #(
		.INIT('h1)
	) name3869 (
		_w4810_,
		_w4811_,
		_w4828_
	);
	LUT2 #(
		.INIT('h1)
	) name3870 (
		_w4812_,
		_w4813_,
		_w4829_
	);
	LUT2 #(
		.INIT('h1)
	) name3871 (
		_w4814_,
		_w4815_,
		_w4830_
	);
	LUT2 #(
		.INIT('h1)
	) name3872 (
		_w4816_,
		_w4817_,
		_w4831_
	);
	LUT2 #(
		.INIT('h4)
	) name3873 (
		_w4818_,
		_w4831_,
		_w4832_
	);
	LUT2 #(
		.INIT('h8)
	) name3874 (
		_w4829_,
		_w4830_,
		_w4833_
	);
	LUT2 #(
		.INIT('h8)
	) name3875 (
		_w4827_,
		_w4828_,
		_w4834_
	);
	LUT2 #(
		.INIT('h8)
	) name3876 (
		_w4825_,
		_w4826_,
		_w4835_
	);
	LUT2 #(
		.INIT('h8)
	) name3877 (
		_w4823_,
		_w4824_,
		_w4836_
	);
	LUT2 #(
		.INIT('h8)
	) name3878 (
		_w4821_,
		_w4822_,
		_w4837_
	);
	LUT2 #(
		.INIT('h8)
	) name3879 (
		_w4819_,
		_w4820_,
		_w4838_
	);
	LUT2 #(
		.INIT('h8)
	) name3880 (
		_w4837_,
		_w4838_,
		_w4839_
	);
	LUT2 #(
		.INIT('h8)
	) name3881 (
		_w4835_,
		_w4836_,
		_w4840_
	);
	LUT2 #(
		.INIT('h8)
	) name3882 (
		_w4833_,
		_w4834_,
		_w4841_
	);
	LUT2 #(
		.INIT('h8)
	) name3883 (
		_w4832_,
		_w4841_,
		_w4842_
	);
	LUT2 #(
		.INIT('h8)
	) name3884 (
		_w4839_,
		_w4840_,
		_w4843_
	);
	LUT2 #(
		.INIT('h8)
	) name3885 (
		_w4842_,
		_w4843_,
		_w4844_
	);
	LUT2 #(
		.INIT('h2)
	) name3886 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b3_last_row_reg[6]/P0001 ,
		_w4845_
	);
	LUT2 #(
		.INIT('h1)
	) name3887 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b3_last_row_reg[4]/P0001 ,
		_w4846_
	);
	LUT2 #(
		.INIT('h8)
	) name3888 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b3_last_row_reg[4]/P0001 ,
		_w4847_
	);
	LUT2 #(
		.INIT('h1)
	) name3889 (
		_w4846_,
		_w4847_,
		_w4848_
	);
	LUT2 #(
		.INIT('h2)
	) name3890 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b3_last_row_reg[5]/P0001 ,
		_w4849_
	);
	LUT2 #(
		.INIT('h4)
	) name3891 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u0_b3_last_row_reg[10]/P0001 ,
		_w4850_
	);
	LUT2 #(
		.INIT('h2)
	) name3892 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b3_last_row_reg[2]/P0001 ,
		_w4851_
	);
	LUT2 #(
		.INIT('h4)
	) name3893 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b3_last_row_reg[8]/P0001 ,
		_w4852_
	);
	LUT2 #(
		.INIT('h4)
	) name3894 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b3_last_row_reg[7]/P0001 ,
		_w4853_
	);
	LUT2 #(
		.INIT('h2)
	) name3895 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b3_last_row_reg[9]/P0001 ,
		_w4854_
	);
	LUT2 #(
		.INIT('h4)
	) name3896 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b3_last_row_reg[1]/P0001 ,
		_w4855_
	);
	LUT2 #(
		.INIT('h2)
	) name3897 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u0_b3_last_row_reg[12]/P0001 ,
		_w4856_
	);
	LUT2 #(
		.INIT('h2)
	) name3898 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b3_last_row_reg[3]/P0001 ,
		_w4857_
	);
	LUT2 #(
		.INIT('h2)
	) name3899 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b3_last_row_reg[8]/P0001 ,
		_w4858_
	);
	LUT2 #(
		.INIT('h4)
	) name3900 (
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b3_last_row_reg[2]/P0001 ,
		_w4859_
	);
	LUT2 #(
		.INIT('h4)
	) name3901 (
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b3_last_row_reg[6]/P0001 ,
		_w4860_
	);
	LUT2 #(
		.INIT('h4)
	) name3902 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b3_last_row_reg[3]/P0001 ,
		_w4861_
	);
	LUT2 #(
		.INIT('h2)
	) name3903 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u0_b3_last_row_reg[10]/P0001 ,
		_w4862_
	);
	LUT2 #(
		.INIT('h4)
	) name3904 (
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b3_last_row_reg[5]/P0001 ,
		_w4863_
	);
	LUT2 #(
		.INIT('h4)
	) name3905 (
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b3_last_row_reg[9]/P0001 ,
		_w4864_
	);
	LUT2 #(
		.INIT('h4)
	) name3906 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b3_last_row_reg[11]/P0001 ,
		_w4865_
	);
	LUT2 #(
		.INIT('h2)
	) name3907 (
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b3_last_row_reg[7]/P0001 ,
		_w4866_
	);
	LUT2 #(
		.INIT('h2)
	) name3908 (
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b3_last_row_reg[1]/P0001 ,
		_w4867_
	);
	LUT2 #(
		.INIT('h4)
	) name3909 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u0_b3_last_row_reg[12]/P0001 ,
		_w4868_
	);
	LUT2 #(
		.INIT('h2)
	) name3910 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u0_b3_last_row_reg[0]/P0001 ,
		_w4869_
	);
	LUT2 #(
		.INIT('h2)
	) name3911 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b3_last_row_reg[11]/P0001 ,
		_w4870_
	);
	LUT2 #(
		.INIT('h4)
	) name3912 (
		\u1_row_adr_reg[0]/P0001 ,
		\u2_u0_b3_last_row_reg[0]/P0001 ,
		_w4871_
	);
	LUT2 #(
		.INIT('h2)
	) name3913 (
		_w3133_,
		_w4845_,
		_w4872_
	);
	LUT2 #(
		.INIT('h1)
	) name3914 (
		_w4849_,
		_w4850_,
		_w4873_
	);
	LUT2 #(
		.INIT('h1)
	) name3915 (
		_w4851_,
		_w4852_,
		_w4874_
	);
	LUT2 #(
		.INIT('h1)
	) name3916 (
		_w4853_,
		_w4854_,
		_w4875_
	);
	LUT2 #(
		.INIT('h1)
	) name3917 (
		_w4855_,
		_w4856_,
		_w4876_
	);
	LUT2 #(
		.INIT('h1)
	) name3918 (
		_w4857_,
		_w4858_,
		_w4877_
	);
	LUT2 #(
		.INIT('h1)
	) name3919 (
		_w4859_,
		_w4860_,
		_w4878_
	);
	LUT2 #(
		.INIT('h1)
	) name3920 (
		_w4861_,
		_w4862_,
		_w4879_
	);
	LUT2 #(
		.INIT('h1)
	) name3921 (
		_w4863_,
		_w4864_,
		_w4880_
	);
	LUT2 #(
		.INIT('h1)
	) name3922 (
		_w4865_,
		_w4866_,
		_w4881_
	);
	LUT2 #(
		.INIT('h1)
	) name3923 (
		_w4867_,
		_w4868_,
		_w4882_
	);
	LUT2 #(
		.INIT('h1)
	) name3924 (
		_w4869_,
		_w4870_,
		_w4883_
	);
	LUT2 #(
		.INIT('h4)
	) name3925 (
		_w4871_,
		_w4883_,
		_w4884_
	);
	LUT2 #(
		.INIT('h8)
	) name3926 (
		_w4881_,
		_w4882_,
		_w4885_
	);
	LUT2 #(
		.INIT('h8)
	) name3927 (
		_w4879_,
		_w4880_,
		_w4886_
	);
	LUT2 #(
		.INIT('h8)
	) name3928 (
		_w4877_,
		_w4878_,
		_w4887_
	);
	LUT2 #(
		.INIT('h8)
	) name3929 (
		_w4875_,
		_w4876_,
		_w4888_
	);
	LUT2 #(
		.INIT('h8)
	) name3930 (
		_w4873_,
		_w4874_,
		_w4889_
	);
	LUT2 #(
		.INIT('h4)
	) name3931 (
		_w4848_,
		_w4872_,
		_w4890_
	);
	LUT2 #(
		.INIT('h8)
	) name3932 (
		_w4889_,
		_w4890_,
		_w4891_
	);
	LUT2 #(
		.INIT('h8)
	) name3933 (
		_w4887_,
		_w4888_,
		_w4892_
	);
	LUT2 #(
		.INIT('h8)
	) name3934 (
		_w4885_,
		_w4886_,
		_w4893_
	);
	LUT2 #(
		.INIT('h8)
	) name3935 (
		_w4884_,
		_w4893_,
		_w4894_
	);
	LUT2 #(
		.INIT('h8)
	) name3936 (
		_w4891_,
		_w4892_,
		_w4895_
	);
	LUT2 #(
		.INIT('h8)
	) name3937 (
		_w4894_,
		_w4895_,
		_w4896_
	);
	LUT2 #(
		.INIT('h1)
	) name3938 (
		_w4740_,
		_w4792_,
		_w4897_
	);
	LUT2 #(
		.INIT('h1)
	) name3939 (
		_w4844_,
		_w4896_,
		_w4898_
	);
	LUT2 #(
		.INIT('h8)
	) name3940 (
		_w4897_,
		_w4898_,
		_w4899_
	);
	LUT2 #(
		.INIT('h2)
	) name3941 (
		_w1623_,
		_w4899_,
		_w4900_
	);
	LUT2 #(
		.INIT('h1)
	) name3942 (
		_w4688_,
		_w4900_,
		_w4901_
	);
	LUT2 #(
		.INIT('h8)
	) name3943 (
		_w2842_,
		_w3035_,
		_w4902_
	);
	LUT2 #(
		.INIT('h4)
	) name3944 (
		_w2818_,
		_w4902_,
		_w4903_
	);
	LUT2 #(
		.INIT('h8)
	) name3945 (
		_w2821_,
		_w4903_,
		_w4904_
	);
	LUT2 #(
		.INIT('h8)
	) name3946 (
		_w3032_,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('h8)
	) name3947 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1362_,
		_w4906_
	);
	LUT2 #(
		.INIT('h2)
	) name3948 (
		\u5_susp_sel_r_reg/NET0131 ,
		_w4906_,
		_w4907_
	);
	LUT2 #(
		.INIT('h8)
	) name3949 (
		_w1680_,
		_w1682_,
		_w4908_
	);
	LUT2 #(
		.INIT('h8)
	) name3950 (
		_w3178_,
		_w4908_,
		_w4909_
	);
	LUT2 #(
		.INIT('h1)
	) name3951 (
		_w4907_,
		_w4909_,
		_w4910_
	);
	LUT2 #(
		.INIT('h8)
	) name3952 (
		\u0_u1_csc_reg[1]/NET0131 ,
		_w3458_,
		_w4911_
	);
	LUT2 #(
		.INIT('h8)
	) name3953 (
		\u0_u0_csc_reg[1]/NET0131 ,
		_w3415_,
		_w4912_
	);
	LUT2 #(
		.INIT('h1)
	) name3954 (
		_w4911_,
		_w4912_,
		_w4913_
	);
	LUT2 #(
		.INIT('h8)
	) name3955 (
		\u0_u1_csc_reg[2]/NET0131 ,
		_w3458_,
		_w4914_
	);
	LUT2 #(
		.INIT('h8)
	) name3956 (
		\u0_u0_csc_reg[2]/NET0131 ,
		_w3415_,
		_w4915_
	);
	LUT2 #(
		.INIT('h1)
	) name3957 (
		_w4914_,
		_w4915_,
		_w4916_
	);
	LUT2 #(
		.INIT('h8)
	) name3958 (
		\u0_u1_csc_reg[3]/NET0131 ,
		_w3458_,
		_w4917_
	);
	LUT2 #(
		.INIT('h8)
	) name3959 (
		\u0_u0_csc_reg[3]/NET0131 ,
		_w3415_,
		_w4918_
	);
	LUT2 #(
		.INIT('h1)
	) name3960 (
		_w4917_,
		_w4918_,
		_w4919_
	);
	LUT2 #(
		.INIT('h1)
	) name3961 (
		\u4_ps_cnt_reg[3]/NET0131 ,
		_w4333_,
		_w4920_
	);
	LUT2 #(
		.INIT('h1)
	) name3962 (
		_w4334_,
		_w4920_,
		_w4921_
	);
	LUT2 #(
		.INIT('h4)
	) name3963 (
		_w4375_,
		_w4921_,
		_w4922_
	);
	LUT2 #(
		.INIT('h8)
	) name3964 (
		\u1_bank_adr_reg[0]/P0001 ,
		_w1062_,
		_w4923_
	);
	LUT2 #(
		.INIT('h8)
	) name3965 (
		\u1_acs_addr_reg[13]/P0001 ,
		_w1438_,
		_w4924_
	);
	LUT2 #(
		.INIT('h1)
	) name3966 (
		\wb_addr_i[15]_pad ,
		_w1442_,
		_w4925_
	);
	LUT2 #(
		.INIT('h4)
	) name3967 (
		\u1_sram_addr_reg[13]/P0001 ,
		_w1442_,
		_w4926_
	);
	LUT2 #(
		.INIT('h1)
	) name3968 (
		_w1058_,
		_w4925_,
		_w4927_
	);
	LUT2 #(
		.INIT('h4)
	) name3969 (
		_w4926_,
		_w4927_,
		_w4928_
	);
	LUT2 #(
		.INIT('h1)
	) name3970 (
		_w4923_,
		_w4924_,
		_w4929_
	);
	LUT2 #(
		.INIT('h4)
	) name3971 (
		_w4928_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('h8)
	) name3972 (
		\u1_bank_adr_reg[1]/P0001 ,
		_w1062_,
		_w4931_
	);
	LUT2 #(
		.INIT('h8)
	) name3973 (
		\u1_acs_addr_reg[14]/P0001 ,
		_w1438_,
		_w4932_
	);
	LUT2 #(
		.INIT('h1)
	) name3974 (
		\wb_addr_i[16]_pad ,
		_w1442_,
		_w4933_
	);
	LUT2 #(
		.INIT('h4)
	) name3975 (
		\u1_sram_addr_reg[14]/P0001 ,
		_w1442_,
		_w4934_
	);
	LUT2 #(
		.INIT('h1)
	) name3976 (
		_w1058_,
		_w4933_,
		_w4935_
	);
	LUT2 #(
		.INIT('h4)
	) name3977 (
		_w4934_,
		_w4935_,
		_w4936_
	);
	LUT2 #(
		.INIT('h1)
	) name3978 (
		_w4931_,
		_w4932_,
		_w4937_
	);
	LUT2 #(
		.INIT('h4)
	) name3979 (
		_w4936_,
		_w4937_,
		_w4938_
	);
	LUT2 #(
		.INIT('h8)
	) name3980 (
		\u1_col_adr_reg[9]/P0001 ,
		_w4316_,
		_w4939_
	);
	LUT2 #(
		.INIT('h2)
	) name3981 (
		_w3840_,
		_w4316_,
		_w4940_
	);
	LUT2 #(
		.INIT('h4)
	) name3982 (
		_w3977_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h1)
	) name3983 (
		_w4939_,
		_w4941_,
		_w4942_
	);
	LUT2 #(
		.INIT('h8)
	) name3984 (
		\u1_acs_addr_reg[16]/P0001 ,
		_w1438_,
		_w4943_
	);
	LUT2 #(
		.INIT('h1)
	) name3985 (
		\wb_addr_i[18]_pad ,
		_w1442_,
		_w4944_
	);
	LUT2 #(
		.INIT('h4)
	) name3986 (
		\u1_sram_addr_reg[16]/P0001 ,
		_w1442_,
		_w4945_
	);
	LUT2 #(
		.INIT('h1)
	) name3987 (
		_w1058_,
		_w4944_,
		_w4946_
	);
	LUT2 #(
		.INIT('h4)
	) name3988 (
		_w4945_,
		_w4946_,
		_w4947_
	);
	LUT2 #(
		.INIT('h1)
	) name3989 (
		_w4943_,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h8)
	) name3990 (
		\u1_acs_addr_reg[17]/P0001 ,
		_w1438_,
		_w4949_
	);
	LUT2 #(
		.INIT('h1)
	) name3991 (
		\wb_addr_i[19]_pad ,
		_w1442_,
		_w4950_
	);
	LUT2 #(
		.INIT('h4)
	) name3992 (
		\u1_sram_addr_reg[17]/P0001 ,
		_w1442_,
		_w4951_
	);
	LUT2 #(
		.INIT('h1)
	) name3993 (
		_w1058_,
		_w4950_,
		_w4952_
	);
	LUT2 #(
		.INIT('h4)
	) name3994 (
		_w4951_,
		_w4952_,
		_w4953_
	);
	LUT2 #(
		.INIT('h1)
	) name3995 (
		_w4949_,
		_w4953_,
		_w4954_
	);
	LUT2 #(
		.INIT('h8)
	) name3996 (
		\u1_acs_addr_reg[18]/P0001 ,
		_w1438_,
		_w4955_
	);
	LUT2 #(
		.INIT('h1)
	) name3997 (
		\wb_addr_i[20]_pad ,
		_w1442_,
		_w4956_
	);
	LUT2 #(
		.INIT('h4)
	) name3998 (
		\u1_sram_addr_reg[18]/P0001 ,
		_w1442_,
		_w4957_
	);
	LUT2 #(
		.INIT('h1)
	) name3999 (
		_w1058_,
		_w4956_,
		_w4958_
	);
	LUT2 #(
		.INIT('h4)
	) name4000 (
		_w4957_,
		_w4958_,
		_w4959_
	);
	LUT2 #(
		.INIT('h1)
	) name4001 (
		_w4955_,
		_w4959_,
		_w4960_
	);
	LUT2 #(
		.INIT('h8)
	) name4002 (
		\u1_acs_addr_reg[19]/P0001 ,
		_w1438_,
		_w4961_
	);
	LUT2 #(
		.INIT('h1)
	) name4003 (
		\wb_addr_i[21]_pad ,
		_w1442_,
		_w4962_
	);
	LUT2 #(
		.INIT('h4)
	) name4004 (
		\u1_sram_addr_reg[19]/P0001 ,
		_w1442_,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name4005 (
		_w1058_,
		_w4962_,
		_w4964_
	);
	LUT2 #(
		.INIT('h4)
	) name4006 (
		_w4963_,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h1)
	) name4007 (
		_w4961_,
		_w4965_,
		_w4966_
	);
	LUT2 #(
		.INIT('h8)
	) name4008 (
		\u1_acs_addr_reg[21]/P0001 ,
		_w1438_,
		_w4967_
	);
	LUT2 #(
		.INIT('h1)
	) name4009 (
		\wb_addr_i[23]_pad ,
		_w1442_,
		_w4968_
	);
	LUT2 #(
		.INIT('h4)
	) name4010 (
		\u1_sram_addr_reg[21]/P0001 ,
		_w1442_,
		_w4969_
	);
	LUT2 #(
		.INIT('h1)
	) name4011 (
		_w1058_,
		_w4968_,
		_w4970_
	);
	LUT2 #(
		.INIT('h4)
	) name4012 (
		_w4969_,
		_w4970_,
		_w4971_
	);
	LUT2 #(
		.INIT('h1)
	) name4013 (
		_w4967_,
		_w4971_,
		_w4972_
	);
	LUT2 #(
		.INIT('h8)
	) name4014 (
		\u1_acs_addr_reg[22]/P0001 ,
		_w1438_,
		_w4973_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		\wb_addr_i[24]_pad ,
		_w1442_,
		_w4974_
	);
	LUT2 #(
		.INIT('h4)
	) name4016 (
		\u1_sram_addr_reg[22]/P0001 ,
		_w1442_,
		_w4975_
	);
	LUT2 #(
		.INIT('h1)
	) name4017 (
		_w1058_,
		_w4974_,
		_w4976_
	);
	LUT2 #(
		.INIT('h4)
	) name4018 (
		_w4975_,
		_w4976_,
		_w4977_
	);
	LUT2 #(
		.INIT('h1)
	) name4019 (
		_w4973_,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h8)
	) name4020 (
		\u1_acs_addr_reg[23]/P0001 ,
		_w1438_,
		_w4979_
	);
	LUT2 #(
		.INIT('h1)
	) name4021 (
		\wb_addr_i[25]_pad ,
		_w1442_,
		_w4980_
	);
	LUT2 #(
		.INIT('h4)
	) name4022 (
		\u1_sram_addr_reg[23]/P0001 ,
		_w1442_,
		_w4981_
	);
	LUT2 #(
		.INIT('h1)
	) name4023 (
		_w1058_,
		_w4980_,
		_w4982_
	);
	LUT2 #(
		.INIT('h4)
	) name4024 (
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT2 #(
		.INIT('h1)
	) name4025 (
		_w4979_,
		_w4983_,
		_w4984_
	);
	LUT2 #(
		.INIT('h8)
	) name4026 (
		\u1_acs_addr_reg[15]/P0001 ,
		_w1438_,
		_w4985_
	);
	LUT2 #(
		.INIT('h1)
	) name4027 (
		\wb_addr_i[17]_pad ,
		_w1442_,
		_w4986_
	);
	LUT2 #(
		.INIT('h4)
	) name4028 (
		\u1_sram_addr_reg[15]/P0001 ,
		_w1442_,
		_w4987_
	);
	LUT2 #(
		.INIT('h1)
	) name4029 (
		_w1058_,
		_w4986_,
		_w4988_
	);
	LUT2 #(
		.INIT('h4)
	) name4030 (
		_w4987_,
		_w4988_,
		_w4989_
	);
	LUT2 #(
		.INIT('h1)
	) name4031 (
		_w4985_,
		_w4989_,
		_w4990_
	);
	LUT2 #(
		.INIT('h8)
	) name4032 (
		\u1_acs_addr_reg[20]/P0001 ,
		_w1438_,
		_w4991_
	);
	LUT2 #(
		.INIT('h1)
	) name4033 (
		\wb_addr_i[22]_pad ,
		_w1442_,
		_w4992_
	);
	LUT2 #(
		.INIT('h4)
	) name4034 (
		\u1_sram_addr_reg[20]/P0001 ,
		_w1442_,
		_w4993_
	);
	LUT2 #(
		.INIT('h1)
	) name4035 (
		_w1058_,
		_w4992_,
		_w4994_
	);
	LUT2 #(
		.INIT('h4)
	) name4036 (
		_w4993_,
		_w4994_,
		_w4995_
	);
	LUT2 #(
		.INIT('h1)
	) name4037 (
		_w4991_,
		_w4995_,
		_w4996_
	);
	LUT2 #(
		.INIT('h1)
	) name4038 (
		\u1_acs_addr_reg[8]/P0001 ,
		_w4007_,
		_w4997_
	);
	LUT2 #(
		.INIT('h1)
	) name4039 (
		_w4008_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h1)
	) name4040 (
		\u4_ps_cnt_reg[2]/NET0131 ,
		_w4332_,
		_w4999_
	);
	LUT2 #(
		.INIT('h1)
	) name4041 (
		_w4333_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('h4)
	) name4042 (
		_w4375_,
		_w5000_,
		_w5001_
	);
	LUT2 #(
		.INIT('h1)
	) name4043 (
		\u4_ps_cnt_reg[5]/NET0131 ,
		_w4335_,
		_w5002_
	);
	LUT2 #(
		.INIT('h1)
	) name4044 (
		_w4375_,
		_w4457_,
		_w5003_
	);
	LUT2 #(
		.INIT('h4)
	) name4045 (
		_w5002_,
		_w5003_,
		_w5004_
	);
	LUT2 #(
		.INIT('h1)
	) name4046 (
		\u4_ps_cnt_reg[6]/NET0131 ,
		_w4457_,
		_w5005_
	);
	LUT2 #(
		.INIT('h1)
	) name4047 (
		_w4375_,
		_w4458_,
		_w5006_
	);
	LUT2 #(
		.INIT('h4)
	) name4048 (
		_w5005_,
		_w5006_,
		_w5007_
	);
	LUT2 #(
		.INIT('h1)
	) name4049 (
		\u4_ps_cnt_reg[0]/NET0131 ,
		\u4_rfr_en_reg/NET0131 ,
		_w5008_
	);
	LUT2 #(
		.INIT('h1)
	) name4050 (
		_w4331_,
		_w5008_,
		_w5009_
	);
	LUT2 #(
		.INIT('h4)
	) name4051 (
		_w4375_,
		_w5009_,
		_w5010_
	);
	LUT2 #(
		.INIT('h1)
	) name4052 (
		\u4_ps_cnt_reg[1]/NET0131 ,
		_w4331_,
		_w5011_
	);
	LUT2 #(
		.INIT('h1)
	) name4053 (
		_w4332_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h4)
	) name4054 (
		_w4375_,
		_w5012_,
		_w5013_
	);
	LUT2 #(
		.INIT('h8)
	) name4055 (
		\u0_init_req_reg/NET0131 ,
		_w3178_,
		_w5014_
	);
	LUT2 #(
		.INIT('h1)
	) name4056 (
		\u1_acs_addr_reg[4]/P0001 ,
		_w4003_,
		_w5015_
	);
	LUT2 #(
		.INIT('h1)
	) name4057 (
		_w4004_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h8)
	) name4058 (
		\mem_ack_r_reg/P0001 ,
		_w1627_,
		_w5017_
	);
	LUT2 #(
		.INIT('h8)
	) name4059 (
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h2)
	) name4060 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		_w5017_,
		_w5019_
	);
	LUT2 #(
		.INIT('h2)
	) name4061 (
		_w4203_,
		_w5018_,
		_w5020_
	);
	LUT2 #(
		.INIT('h4)
	) name4062 (
		_w5019_,
		_w5020_,
		_w5021_
	);
	LUT2 #(
		.INIT('h1)
	) name4063 (
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		_w5017_,
		_w5022_
	);
	LUT2 #(
		.INIT('h4)
	) name4064 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		_w5017_,
		_w5023_
	);
	LUT2 #(
		.INIT('h2)
	) name4065 (
		_w4203_,
		_w5022_,
		_w5024_
	);
	LUT2 #(
		.INIT('h4)
	) name4066 (
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT2 #(
		.INIT('h1)
	) name4067 (
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		_w5017_,
		_w5026_
	);
	LUT2 #(
		.INIT('h4)
	) name4068 (
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		_w5017_,
		_w5027_
	);
	LUT2 #(
		.INIT('h2)
	) name4069 (
		_w4203_,
		_w5026_,
		_w5028_
	);
	LUT2 #(
		.INIT('h4)
	) name4070 (
		_w5027_,
		_w5028_,
		_w5029_
	);
	LUT2 #(
		.INIT('h1)
	) name4071 (
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		_w5017_,
		_w5030_
	);
	LUT2 #(
		.INIT('h4)
	) name4072 (
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		_w5017_,
		_w5031_
	);
	LUT2 #(
		.INIT('h2)
	) name4073 (
		_w4203_,
		_w5030_,
		_w5032_
	);
	LUT2 #(
		.INIT('h4)
	) name4074 (
		_w5031_,
		_w5032_,
		_w5033_
	);
	LUT2 #(
		.INIT('h8)
	) name4075 (
		\u2_u0_bank2_open_reg/NET0131 ,
		_w3103_,
		_w5034_
	);
	LUT2 #(
		.INIT('h8)
	) name4076 (
		\u2_u0_bank1_open_reg/NET0131 ,
		_w3049_,
		_w5035_
	);
	LUT2 #(
		.INIT('h8)
	) name4077 (
		\u2_u0_bank3_open_reg/NET0131 ,
		_w3133_,
		_w5036_
	);
	LUT2 #(
		.INIT('h8)
	) name4078 (
		\u2_u0_bank0_open_reg/NET0131 ,
		_w4607_,
		_w5037_
	);
	LUT2 #(
		.INIT('h1)
	) name4079 (
		_w5034_,
		_w5035_,
		_w5038_
	);
	LUT2 #(
		.INIT('h1)
	) name4080 (
		_w5036_,
		_w5037_,
		_w5039_
	);
	LUT2 #(
		.INIT('h8)
	) name4081 (
		_w5038_,
		_w5039_,
		_w5040_
	);
	LUT2 #(
		.INIT('h2)
	) name4082 (
		_w1623_,
		_w5040_,
		_w5041_
	);
	LUT2 #(
		.INIT('h8)
	) name4083 (
		\u2_u1_bank2_open_reg/NET0131 ,
		_w3103_,
		_w5042_
	);
	LUT2 #(
		.INIT('h8)
	) name4084 (
		\u2_u1_bank3_open_reg/NET0131 ,
		_w3133_,
		_w5043_
	);
	LUT2 #(
		.INIT('h8)
	) name4085 (
		\u2_u1_bank0_open_reg/NET0131 ,
		_w4607_,
		_w5044_
	);
	LUT2 #(
		.INIT('h8)
	) name4086 (
		\u2_u1_bank1_open_reg/NET0131 ,
		_w3049_,
		_w5045_
	);
	LUT2 #(
		.INIT('h1)
	) name4087 (
		_w5042_,
		_w5043_,
		_w5046_
	);
	LUT2 #(
		.INIT('h1)
	) name4088 (
		_w5044_,
		_w5045_,
		_w5047_
	);
	LUT2 #(
		.INIT('h8)
	) name4089 (
		_w5046_,
		_w5047_,
		_w5048_
	);
	LUT2 #(
		.INIT('h1)
	) name4090 (
		_w1676_,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h1)
	) name4091 (
		_w5041_,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('h8)
	) name4092 (
		\poc_o[3]_pad ,
		\u0_rst_r2_reg/NET0131 ,
		_w5051_
	);
	LUT2 #(
		.INIT('h8)
	) name4093 (
		\poc_o[2]_pad ,
		\u0_rst_r2_reg/NET0131 ,
		_w5052_
	);
	LUT2 #(
		.INIT('h8)
	) name4094 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		_w5053_
	);
	LUT2 #(
		.INIT('h1)
	) name4095 (
		\u0_u0_addr_r_reg[5]/P0001 ,
		\u0_u0_addr_r_reg[6]/P0001 ,
		_w5054_
	);
	LUT2 #(
		.INIT('h4)
	) name4096 (
		\u0_u0_addr_r_reg[3]/P0001 ,
		_w5054_,
		_w5055_
	);
	LUT2 #(
		.INIT('h8)
	) name4097 (
		_w5053_,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h4)
	) name4098 (
		\u0_u0_addr_r_reg[2]/P0001 ,
		_w5056_,
		_w5057_
	);
	LUT2 #(
		.INIT('h1)
	) name4099 (
		\u0_u0_csc_reg[0]/NET0131 ,
		_w5057_,
		_w5058_
	);
	LUT2 #(
		.INIT('h4)
	) name4100 (
		\wb_data_i[0]_pad ,
		_w5057_,
		_w5059_
	);
	LUT2 #(
		.INIT('h1)
	) name4101 (
		\u0_rst_r2_reg/NET0131 ,
		_w5058_,
		_w5060_
	);
	LUT2 #(
		.INIT('h4)
	) name4102 (
		_w5059_,
		_w5060_,
		_w5061_
	);
	LUT2 #(
		.INIT('h1)
	) name4103 (
		_w5051_,
		_w5052_,
		_w5062_
	);
	LUT2 #(
		.INIT('h4)
	) name4104 (
		_w5061_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h1)
	) name4105 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		_w5064_
	);
	LUT2 #(
		.INIT('h4)
	) name4106 (
		_w2072_,
		_w5064_,
		_w5065_
	);
	LUT2 #(
		.INIT('h8)
	) name4107 (
		\u7_mc_data_ir_reg[2]/P0001 ,
		_w4151_,
		_w5066_
	);
	LUT2 #(
		.INIT('h8)
	) name4108 (
		\u7_mc_data_ir_reg[10]/P0001 ,
		_w4153_,
		_w5067_
	);
	LUT2 #(
		.INIT('h8)
	) name4109 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[26]/P0001 ,
		_w5068_
	);
	LUT2 #(
		.INIT('h1)
	) name4110 (
		_w5066_,
		_w5068_,
		_w5069_
	);
	LUT2 #(
		.INIT('h4)
	) name4111 (
		_w5067_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h1)
	) name4112 (
		_w5064_,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h2)
	) name4113 (
		_w2269_,
		_w5071_,
		_w5072_
	);
	LUT2 #(
		.INIT('h4)
	) name4114 (
		_w5065_,
		_w5072_,
		_w5073_
	);
	LUT2 #(
		.INIT('h1)
	) name4115 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w5074_
	);
	LUT2 #(
		.INIT('h4)
	) name4116 (
		\wb_addr_i[3]_pad ,
		_w5074_,
		_w5075_
	);
	LUT2 #(
		.INIT('h8)
	) name4117 (
		\wb_addr_i[2]_pad ,
		_w5075_,
		_w5076_
	);
	LUT2 #(
		.INIT('h8)
	) name4118 (
		\wb_addr_i[4]_pad ,
		_w5076_,
		_w5077_
	);
	LUT2 #(
		.INIT('h8)
	) name4119 (
		\u0_u0_tms_reg[26]/P0001 ,
		_w5077_,
		_w5078_
	);
	LUT2 #(
		.INIT('h4)
	) name4120 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w5079_
	);
	LUT2 #(
		.INIT('h8)
	) name4121 (
		\wb_addr_i[3]_pad ,
		_w5074_,
		_w5080_
	);
	LUT2 #(
		.INIT('h8)
	) name4122 (
		_w5079_,
		_w5080_,
		_w5081_
	);
	LUT2 #(
		.INIT('h8)
	) name4123 (
		\u0_u1_csc_reg[26]/P0001 ,
		_w5081_,
		_w5082_
	);
	LUT2 #(
		.INIT('h8)
	) name4124 (
		_w5075_,
		_w5079_,
		_w5083_
	);
	LUT2 #(
		.INIT('h8)
	) name4125 (
		\u0_u0_csc_reg[26]/P0001 ,
		_w5083_,
		_w5084_
	);
	LUT2 #(
		.INIT('h8)
	) name4126 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w5085_
	);
	LUT2 #(
		.INIT('h8)
	) name4127 (
		_w5080_,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('h8)
	) name4128 (
		\u0_u1_tms_reg[26]/P0001 ,
		_w5086_,
		_w5087_
	);
	LUT2 #(
		.INIT('h1)
	) name4129 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w5088_
	);
	LUT2 #(
		.INIT('h8)
	) name4130 (
		_w5075_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h8)
	) name4131 (
		\u0_csr_r2_reg[2]/NET0131 ,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h4)
	) name4132 (
		\wb_addr_i[4]_pad ,
		_w5076_,
		_w5091_
	);
	LUT2 #(
		.INIT('h8)
	) name4133 (
		\poc_o[26]_pad ,
		_w5091_,
		_w5092_
	);
	LUT2 #(
		.INIT('h1)
	) name4134 (
		_w2269_,
		_w5082_,
		_w5093_
	);
	LUT2 #(
		.INIT('h1)
	) name4135 (
		_w5084_,
		_w5087_,
		_w5094_
	);
	LUT2 #(
		.INIT('h4)
	) name4136 (
		_w5090_,
		_w5094_,
		_w5095_
	);
	LUT2 #(
		.INIT('h4)
	) name4137 (
		_w5078_,
		_w5093_,
		_w5096_
	);
	LUT2 #(
		.INIT('h4)
	) name4138 (
		_w5092_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h8)
	) name4139 (
		_w5095_,
		_w5097_,
		_w5098_
	);
	LUT2 #(
		.INIT('h1)
	) name4140 (
		_w5073_,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h8)
	) name4141 (
		_w2018_,
		_w5064_,
		_w5100_
	);
	LUT2 #(
		.INIT('h8)
	) name4142 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[27]/P0001 ,
		_w5101_
	);
	LUT2 #(
		.INIT('h8)
	) name4143 (
		\u7_mc_data_ir_reg[3]/P0001 ,
		_w4151_,
		_w5102_
	);
	LUT2 #(
		.INIT('h8)
	) name4144 (
		\u7_mc_data_ir_reg[11]/P0001 ,
		_w4153_,
		_w5103_
	);
	LUT2 #(
		.INIT('h1)
	) name4145 (
		_w5064_,
		_w5101_,
		_w5104_
	);
	LUT2 #(
		.INIT('h4)
	) name4146 (
		_w5102_,
		_w5104_,
		_w5105_
	);
	LUT2 #(
		.INIT('h4)
	) name4147 (
		_w5103_,
		_w5105_,
		_w5106_
	);
	LUT2 #(
		.INIT('h1)
	) name4148 (
		_w5100_,
		_w5106_,
		_w5107_
	);
	LUT2 #(
		.INIT('h2)
	) name4149 (
		_w2269_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h8)
	) name4150 (
		\u0_u0_tms_reg[27]/P0001 ,
		_w5077_,
		_w5109_
	);
	LUT2 #(
		.INIT('h8)
	) name4151 (
		\u0_csr_r2_reg[3]/NET0131 ,
		_w5089_,
		_w5110_
	);
	LUT2 #(
		.INIT('h8)
	) name4152 (
		\u0_u0_csc_reg[27]/P0001 ,
		_w5083_,
		_w5111_
	);
	LUT2 #(
		.INIT('h8)
	) name4153 (
		\u0_u1_tms_reg[27]/P0001 ,
		_w5086_,
		_w5112_
	);
	LUT2 #(
		.INIT('h8)
	) name4154 (
		\u0_u1_csc_reg[27]/P0001 ,
		_w5081_,
		_w5113_
	);
	LUT2 #(
		.INIT('h8)
	) name4155 (
		\poc_o[27]_pad ,
		_w5091_,
		_w5114_
	);
	LUT2 #(
		.INIT('h1)
	) name4156 (
		_w2269_,
		_w5110_,
		_w5115_
	);
	LUT2 #(
		.INIT('h1)
	) name4157 (
		_w5111_,
		_w5112_,
		_w5116_
	);
	LUT2 #(
		.INIT('h4)
	) name4158 (
		_w5113_,
		_w5116_,
		_w5117_
	);
	LUT2 #(
		.INIT('h4)
	) name4159 (
		_w5109_,
		_w5115_,
		_w5118_
	);
	LUT2 #(
		.INIT('h4)
	) name4160 (
		_w5114_,
		_w5118_,
		_w5119_
	);
	LUT2 #(
		.INIT('h8)
	) name4161 (
		_w5117_,
		_w5119_,
		_w5120_
	);
	LUT2 #(
		.INIT('h1)
	) name4162 (
		_w5108_,
		_w5120_,
		_w5121_
	);
	LUT2 #(
		.INIT('h8)
	) name4163 (
		_w2032_,
		_w5064_,
		_w5122_
	);
	LUT2 #(
		.INIT('h8)
	) name4164 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[28]/P0001 ,
		_w5123_
	);
	LUT2 #(
		.INIT('h8)
	) name4165 (
		\u7_mc_data_ir_reg[4]/P0001 ,
		_w4151_,
		_w5124_
	);
	LUT2 #(
		.INIT('h8)
	) name4166 (
		\u7_mc_data_ir_reg[12]/P0001 ,
		_w4153_,
		_w5125_
	);
	LUT2 #(
		.INIT('h1)
	) name4167 (
		_w5064_,
		_w5123_,
		_w5126_
	);
	LUT2 #(
		.INIT('h4)
	) name4168 (
		_w5124_,
		_w5126_,
		_w5127_
	);
	LUT2 #(
		.INIT('h4)
	) name4169 (
		_w5125_,
		_w5127_,
		_w5128_
	);
	LUT2 #(
		.INIT('h1)
	) name4170 (
		_w5122_,
		_w5128_,
		_w5129_
	);
	LUT2 #(
		.INIT('h2)
	) name4171 (
		_w2269_,
		_w5129_,
		_w5130_
	);
	LUT2 #(
		.INIT('h8)
	) name4172 (
		\u0_u0_tms_reg[28]/P0001 ,
		_w5077_,
		_w5131_
	);
	LUT2 #(
		.INIT('h8)
	) name4173 (
		\u0_csr_r2_reg[4]/NET0131 ,
		_w5089_,
		_w5132_
	);
	LUT2 #(
		.INIT('h8)
	) name4174 (
		\u0_u0_csc_reg[28]/P0001 ,
		_w5083_,
		_w5133_
	);
	LUT2 #(
		.INIT('h8)
	) name4175 (
		\u0_u1_tms_reg[28]/P0001 ,
		_w5086_,
		_w5134_
	);
	LUT2 #(
		.INIT('h8)
	) name4176 (
		\u0_u1_csc_reg[28]/P0001 ,
		_w5081_,
		_w5135_
	);
	LUT2 #(
		.INIT('h8)
	) name4177 (
		\poc_o[28]_pad ,
		_w5091_,
		_w5136_
	);
	LUT2 #(
		.INIT('h1)
	) name4178 (
		_w2269_,
		_w5132_,
		_w5137_
	);
	LUT2 #(
		.INIT('h1)
	) name4179 (
		_w5133_,
		_w5134_,
		_w5138_
	);
	LUT2 #(
		.INIT('h4)
	) name4180 (
		_w5135_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h4)
	) name4181 (
		_w5131_,
		_w5137_,
		_w5140_
	);
	LUT2 #(
		.INIT('h4)
	) name4182 (
		_w5136_,
		_w5140_,
		_w5141_
	);
	LUT2 #(
		.INIT('h8)
	) name4183 (
		_w5139_,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('h1)
	) name4184 (
		_w5130_,
		_w5142_,
		_w5143_
	);
	LUT2 #(
		.INIT('h8)
	) name4185 (
		_w2008_,
		_w5064_,
		_w5144_
	);
	LUT2 #(
		.INIT('h8)
	) name4186 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[29]/P0001 ,
		_w5145_
	);
	LUT2 #(
		.INIT('h8)
	) name4187 (
		\u7_mc_data_ir_reg[5]/P0001 ,
		_w4151_,
		_w5146_
	);
	LUT2 #(
		.INIT('h8)
	) name4188 (
		\u7_mc_data_ir_reg[13]/P0001 ,
		_w4153_,
		_w5147_
	);
	LUT2 #(
		.INIT('h1)
	) name4189 (
		_w5064_,
		_w5145_,
		_w5148_
	);
	LUT2 #(
		.INIT('h4)
	) name4190 (
		_w5146_,
		_w5148_,
		_w5149_
	);
	LUT2 #(
		.INIT('h4)
	) name4191 (
		_w5147_,
		_w5149_,
		_w5150_
	);
	LUT2 #(
		.INIT('h1)
	) name4192 (
		_w5144_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h2)
	) name4193 (
		_w2269_,
		_w5151_,
		_w5152_
	);
	LUT2 #(
		.INIT('h8)
	) name4194 (
		\u0_u0_tms_reg[29]/P0001 ,
		_w5077_,
		_w5153_
	);
	LUT2 #(
		.INIT('h8)
	) name4195 (
		\u0_csr_r2_reg[5]/NET0131 ,
		_w5089_,
		_w5154_
	);
	LUT2 #(
		.INIT('h8)
	) name4196 (
		\u0_u0_csc_reg[29]/P0001 ,
		_w5083_,
		_w5155_
	);
	LUT2 #(
		.INIT('h8)
	) name4197 (
		\u0_u1_tms_reg[29]/P0001 ,
		_w5086_,
		_w5156_
	);
	LUT2 #(
		.INIT('h8)
	) name4198 (
		\u0_u1_csc_reg[29]/P0001 ,
		_w5081_,
		_w5157_
	);
	LUT2 #(
		.INIT('h8)
	) name4199 (
		\poc_o[29]_pad ,
		_w5091_,
		_w5158_
	);
	LUT2 #(
		.INIT('h1)
	) name4200 (
		_w2269_,
		_w5154_,
		_w5159_
	);
	LUT2 #(
		.INIT('h1)
	) name4201 (
		_w5155_,
		_w5156_,
		_w5160_
	);
	LUT2 #(
		.INIT('h4)
	) name4202 (
		_w5157_,
		_w5160_,
		_w5161_
	);
	LUT2 #(
		.INIT('h4)
	) name4203 (
		_w5153_,
		_w5159_,
		_w5162_
	);
	LUT2 #(
		.INIT('h4)
	) name4204 (
		_w5158_,
		_w5162_,
		_w5163_
	);
	LUT2 #(
		.INIT('h8)
	) name4205 (
		_w5161_,
		_w5163_,
		_w5164_
	);
	LUT2 #(
		.INIT('h1)
	) name4206 (
		_w5152_,
		_w5164_,
		_w5165_
	);
	LUT2 #(
		.INIT('h8)
	) name4207 (
		_w2055_,
		_w5064_,
		_w5166_
	);
	LUT2 #(
		.INIT('h8)
	) name4208 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[31]/P0001 ,
		_w5167_
	);
	LUT2 #(
		.INIT('h8)
	) name4209 (
		\u7_mc_data_ir_reg[7]/P0001 ,
		_w4151_,
		_w5168_
	);
	LUT2 #(
		.INIT('h8)
	) name4210 (
		\u7_mc_data_ir_reg[15]/P0001 ,
		_w4153_,
		_w5169_
	);
	LUT2 #(
		.INIT('h1)
	) name4211 (
		_w5064_,
		_w5167_,
		_w5170_
	);
	LUT2 #(
		.INIT('h4)
	) name4212 (
		_w5168_,
		_w5170_,
		_w5171_
	);
	LUT2 #(
		.INIT('h4)
	) name4213 (
		_w5169_,
		_w5171_,
		_w5172_
	);
	LUT2 #(
		.INIT('h1)
	) name4214 (
		_w5166_,
		_w5172_,
		_w5173_
	);
	LUT2 #(
		.INIT('h2)
	) name4215 (
		_w2269_,
		_w5173_,
		_w5174_
	);
	LUT2 #(
		.INIT('h8)
	) name4216 (
		\u0_u0_tms_reg[31]/P0001 ,
		_w5077_,
		_w5175_
	);
	LUT2 #(
		.INIT('h8)
	) name4217 (
		\u0_u0_csc_reg[31]/P0001 ,
		_w5083_,
		_w5176_
	);
	LUT2 #(
		.INIT('h8)
	) name4218 (
		\u0_u1_tms_reg[31]/P0001 ,
		_w5086_,
		_w5177_
	);
	LUT2 #(
		.INIT('h8)
	) name4219 (
		\u0_csr_r2_reg[7]/NET0131 ,
		_w5089_,
		_w5178_
	);
	LUT2 #(
		.INIT('h8)
	) name4220 (
		\u0_u1_csc_reg[31]/P0001 ,
		_w5081_,
		_w5179_
	);
	LUT2 #(
		.INIT('h8)
	) name4221 (
		\poc_o[31]_pad ,
		_w5091_,
		_w5180_
	);
	LUT2 #(
		.INIT('h1)
	) name4222 (
		_w2269_,
		_w5176_,
		_w5181_
	);
	LUT2 #(
		.INIT('h1)
	) name4223 (
		_w5177_,
		_w5178_,
		_w5182_
	);
	LUT2 #(
		.INIT('h4)
	) name4224 (
		_w5179_,
		_w5182_,
		_w5183_
	);
	LUT2 #(
		.INIT('h4)
	) name4225 (
		_w5175_,
		_w5181_,
		_w5184_
	);
	LUT2 #(
		.INIT('h4)
	) name4226 (
		_w5180_,
		_w5184_,
		_w5185_
	);
	LUT2 #(
		.INIT('h8)
	) name4227 (
		_w5183_,
		_w5185_,
		_w5186_
	);
	LUT2 #(
		.INIT('h1)
	) name4228 (
		_w5174_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('h8)
	) name4229 (
		\u0_u0_lmr_req_we_reg/NET0131 ,
		_w1620_,
		_w5188_
	);
	LUT2 #(
		.INIT('h8)
	) name4230 (
		\u0_u0_inited_reg/NET0131 ,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('h2)
	) name4231 (
		\u0_lmr_ack_r_reg/P0001 ,
		\u5_lmr_ack_reg/NET0131 ,
		_w5190_
	);
	LUT2 #(
		.INIT('h8)
	) name4232 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		_w5190_,
		_w5191_
	);
	LUT2 #(
		.INIT('h2)
	) name4233 (
		\u0_u0_lmr_req_reg/NET0131 ,
		_w5191_,
		_w5192_
	);
	LUT2 #(
		.INIT('h4)
	) name4234 (
		_w5188_,
		_w5192_,
		_w5193_
	);
	LUT2 #(
		.INIT('h1)
	) name4235 (
		_w5189_,
		_w5193_,
		_w5194_
	);
	LUT2 #(
		.INIT('h8)
	) name4236 (
		\u0_u1_lmr_req_we_reg/NET0131 ,
		_w1673_,
		_w5195_
	);
	LUT2 #(
		.INIT('h8)
	) name4237 (
		\u0_u1_inited_reg/NET0131 ,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h8)
	) name4238 (
		\u0_spec_req_cs_reg[1]/NET0131 ,
		_w5190_,
		_w5197_
	);
	LUT2 #(
		.INIT('h2)
	) name4239 (
		\u0_u1_lmr_req_reg/NET0131 ,
		_w5197_,
		_w5198_
	);
	LUT2 #(
		.INIT('h4)
	) name4240 (
		_w5195_,
		_w5198_,
		_w5199_
	);
	LUT2 #(
		.INIT('h1)
	) name4241 (
		_w5196_,
		_w5199_,
		_w5200_
	);
	LUT2 #(
		.INIT('h8)
	) name4242 (
		_w2001_,
		_w5064_,
		_w5201_
	);
	LUT2 #(
		.INIT('h8)
	) name4243 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[30]/P0001 ,
		_w5202_
	);
	LUT2 #(
		.INIT('h8)
	) name4244 (
		\u7_mc_data_ir_reg[6]/P0001 ,
		_w4151_,
		_w5203_
	);
	LUT2 #(
		.INIT('h8)
	) name4245 (
		\u7_mc_data_ir_reg[14]/P0001 ,
		_w4153_,
		_w5204_
	);
	LUT2 #(
		.INIT('h1)
	) name4246 (
		_w5064_,
		_w5202_,
		_w5205_
	);
	LUT2 #(
		.INIT('h4)
	) name4247 (
		_w5203_,
		_w5205_,
		_w5206_
	);
	LUT2 #(
		.INIT('h4)
	) name4248 (
		_w5204_,
		_w5206_,
		_w5207_
	);
	LUT2 #(
		.INIT('h1)
	) name4249 (
		_w5201_,
		_w5207_,
		_w5208_
	);
	LUT2 #(
		.INIT('h2)
	) name4250 (
		_w2269_,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('h8)
	) name4251 (
		\u0_u0_tms_reg[30]/P0001 ,
		_w5077_,
		_w5210_
	);
	LUT2 #(
		.INIT('h8)
	) name4252 (
		\u0_csr_r2_reg[6]/NET0131 ,
		_w5089_,
		_w5211_
	);
	LUT2 #(
		.INIT('h8)
	) name4253 (
		\u0_u0_csc_reg[30]/P0001 ,
		_w5083_,
		_w5212_
	);
	LUT2 #(
		.INIT('h8)
	) name4254 (
		\u0_u1_tms_reg[30]/P0001 ,
		_w5086_,
		_w5213_
	);
	LUT2 #(
		.INIT('h8)
	) name4255 (
		\u0_u1_csc_reg[30]/P0001 ,
		_w5081_,
		_w5214_
	);
	LUT2 #(
		.INIT('h8)
	) name4256 (
		\poc_o[30]_pad ,
		_w5091_,
		_w5215_
	);
	LUT2 #(
		.INIT('h1)
	) name4257 (
		_w2269_,
		_w5211_,
		_w5216_
	);
	LUT2 #(
		.INIT('h1)
	) name4258 (
		_w5212_,
		_w5213_,
		_w5217_
	);
	LUT2 #(
		.INIT('h4)
	) name4259 (
		_w5214_,
		_w5217_,
		_w5218_
	);
	LUT2 #(
		.INIT('h4)
	) name4260 (
		_w5210_,
		_w5216_,
		_w5219_
	);
	LUT2 #(
		.INIT('h4)
	) name4261 (
		_w5215_,
		_w5219_,
		_w5220_
	);
	LUT2 #(
		.INIT('h8)
	) name4262 (
		_w5218_,
		_w5220_,
		_w5221_
	);
	LUT2 #(
		.INIT('h1)
	) name4263 (
		_w5209_,
		_w5221_,
		_w5222_
	);
	LUT2 #(
		.INIT('h8)
	) name4264 (
		_w2048_,
		_w5064_,
		_w5223_
	);
	LUT2 #(
		.INIT('h8)
	) name4265 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[24]/P0001 ,
		_w5224_
	);
	LUT2 #(
		.INIT('h8)
	) name4266 (
		\u7_mc_data_ir_reg[8]/P0001 ,
		_w4153_,
		_w5225_
	);
	LUT2 #(
		.INIT('h8)
	) name4267 (
		\u7_mc_data_ir_reg[0]/P0001 ,
		_w4151_,
		_w5226_
	);
	LUT2 #(
		.INIT('h1)
	) name4268 (
		_w5064_,
		_w5224_,
		_w5227_
	);
	LUT2 #(
		.INIT('h4)
	) name4269 (
		_w5225_,
		_w5227_,
		_w5228_
	);
	LUT2 #(
		.INIT('h4)
	) name4270 (
		_w5226_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('h1)
	) name4271 (
		_w5223_,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h2)
	) name4272 (
		_w2269_,
		_w5230_,
		_w5231_
	);
	LUT2 #(
		.INIT('h8)
	) name4273 (
		\u0_u0_tms_reg[24]/P0001 ,
		_w5077_,
		_w5232_
	);
	LUT2 #(
		.INIT('h8)
	) name4274 (
		\u0_csr_r2_reg[0]/NET0131 ,
		_w5089_,
		_w5233_
	);
	LUT2 #(
		.INIT('h8)
	) name4275 (
		\u0_u0_csc_reg[24]/P0001 ,
		_w5083_,
		_w5234_
	);
	LUT2 #(
		.INIT('h8)
	) name4276 (
		\u0_u1_tms_reg[24]/P0001 ,
		_w5086_,
		_w5235_
	);
	LUT2 #(
		.INIT('h8)
	) name4277 (
		\u0_u1_csc_reg[24]/P0001 ,
		_w5081_,
		_w5236_
	);
	LUT2 #(
		.INIT('h8)
	) name4278 (
		\poc_o[24]_pad ,
		_w5091_,
		_w5237_
	);
	LUT2 #(
		.INIT('h1)
	) name4279 (
		_w2269_,
		_w5233_,
		_w5238_
	);
	LUT2 #(
		.INIT('h1)
	) name4280 (
		_w5234_,
		_w5235_,
		_w5239_
	);
	LUT2 #(
		.INIT('h4)
	) name4281 (
		_w5236_,
		_w5239_,
		_w5240_
	);
	LUT2 #(
		.INIT('h4)
	) name4282 (
		_w5232_,
		_w5238_,
		_w5241_
	);
	LUT2 #(
		.INIT('h4)
	) name4283 (
		_w5237_,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('h8)
	) name4284 (
		_w5240_,
		_w5242_,
		_w5243_
	);
	LUT2 #(
		.INIT('h1)
	) name4285 (
		_w5231_,
		_w5243_,
		_w5244_
	);
	LUT2 #(
		.INIT('h8)
	) name4286 (
		_w2025_,
		_w5064_,
		_w5245_
	);
	LUT2 #(
		.INIT('h8)
	) name4287 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[25]/P0001 ,
		_w5246_
	);
	LUT2 #(
		.INIT('h8)
	) name4288 (
		\u7_mc_data_ir_reg[9]/P0001 ,
		_w4153_,
		_w5247_
	);
	LUT2 #(
		.INIT('h8)
	) name4289 (
		\u7_mc_data_ir_reg[1]/P0001 ,
		_w4151_,
		_w5248_
	);
	LUT2 #(
		.INIT('h1)
	) name4290 (
		_w5064_,
		_w5246_,
		_w5249_
	);
	LUT2 #(
		.INIT('h4)
	) name4291 (
		_w5247_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h4)
	) name4292 (
		_w5248_,
		_w5250_,
		_w5251_
	);
	LUT2 #(
		.INIT('h1)
	) name4293 (
		_w5245_,
		_w5251_,
		_w5252_
	);
	LUT2 #(
		.INIT('h2)
	) name4294 (
		_w2269_,
		_w5252_,
		_w5253_
	);
	LUT2 #(
		.INIT('h8)
	) name4295 (
		\u0_u0_tms_reg[25]/P0001 ,
		_w5077_,
		_w5254_
	);
	LUT2 #(
		.INIT('h8)
	) name4296 (
		\u0_csr_r2_reg[1]/NET0131 ,
		_w5089_,
		_w5255_
	);
	LUT2 #(
		.INIT('h8)
	) name4297 (
		\u0_u0_csc_reg[25]/P0001 ,
		_w5083_,
		_w5256_
	);
	LUT2 #(
		.INIT('h8)
	) name4298 (
		\u0_u1_tms_reg[25]/P0001 ,
		_w5086_,
		_w5257_
	);
	LUT2 #(
		.INIT('h8)
	) name4299 (
		\u0_u1_csc_reg[25]/P0001 ,
		_w5081_,
		_w5258_
	);
	LUT2 #(
		.INIT('h8)
	) name4300 (
		\poc_o[25]_pad ,
		_w5091_,
		_w5259_
	);
	LUT2 #(
		.INIT('h1)
	) name4301 (
		_w2269_,
		_w5255_,
		_w5260_
	);
	LUT2 #(
		.INIT('h1)
	) name4302 (
		_w5256_,
		_w5257_,
		_w5261_
	);
	LUT2 #(
		.INIT('h4)
	) name4303 (
		_w5258_,
		_w5261_,
		_w5262_
	);
	LUT2 #(
		.INIT('h4)
	) name4304 (
		_w5254_,
		_w5260_,
		_w5263_
	);
	LUT2 #(
		.INIT('h4)
	) name4305 (
		_w5259_,
		_w5263_,
		_w5264_
	);
	LUT2 #(
		.INIT('h8)
	) name4306 (
		_w5262_,
		_w5264_,
		_w5265_
	);
	LUT2 #(
		.INIT('h1)
	) name4307 (
		_w5253_,
		_w5265_,
		_w5266_
	);
	LUT2 #(
		.INIT('h4)
	) name4308 (
		_w2248_,
		_w5064_,
		_w5267_
	);
	LUT2 #(
		.INIT('h4)
	) name4309 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[1]/P0001 ,
		_w5268_
	);
	LUT2 #(
		.INIT('h8)
	) name4310 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[1]/P0001 ,
		_w5269_
	);
	LUT2 #(
		.INIT('h1)
	) name4311 (
		_w5268_,
		_w5269_,
		_w5270_
	);
	LUT2 #(
		.INIT('h1)
	) name4312 (
		_w5064_,
		_w5270_,
		_w5271_
	);
	LUT2 #(
		.INIT('h2)
	) name4313 (
		_w2269_,
		_w5271_,
		_w5272_
	);
	LUT2 #(
		.INIT('h4)
	) name4314 (
		_w5267_,
		_w5272_,
		_w5273_
	);
	LUT2 #(
		.INIT('h8)
	) name4315 (
		\poc_o[1]_pad ,
		_w5091_,
		_w5274_
	);
	LUT2 #(
		.INIT('h8)
	) name4316 (
		\u0_u0_csc_reg[1]/NET0131 ,
		_w5083_,
		_w5275_
	);
	LUT2 #(
		.INIT('h8)
	) name4317 (
		\u0_u1_csc_reg[1]/NET0131 ,
		_w5081_,
		_w5276_
	);
	LUT2 #(
		.INIT('h8)
	) name4318 (
		_w5080_,
		_w5088_,
		_w5277_
	);
	LUT2 #(
		.INIT('h8)
	) name4319 (
		\u0_csc_mask_r_reg[1]/NET0131 ,
		_w5277_,
		_w5278_
	);
	LUT2 #(
		.INIT('h8)
	) name4320 (
		\u0_u1_tms_reg[1]/P0001 ,
		_w5086_,
		_w5279_
	);
	LUT2 #(
		.INIT('h8)
	) name4321 (
		mc_vpen_pad_o_pad,
		_w5089_,
		_w5280_
	);
	LUT2 #(
		.INIT('h8)
	) name4322 (
		\u0_u0_tms_reg[1]/P0001 ,
		_w5077_,
		_w5281_
	);
	LUT2 #(
		.INIT('h1)
	) name4323 (
		_w2269_,
		_w5275_,
		_w5282_
	);
	LUT2 #(
		.INIT('h1)
	) name4324 (
		_w5276_,
		_w5278_,
		_w5283_
	);
	LUT2 #(
		.INIT('h1)
	) name4325 (
		_w5279_,
		_w5280_,
		_w5284_
	);
	LUT2 #(
		.INIT('h8)
	) name4326 (
		_w5283_,
		_w5284_,
		_w5285_
	);
	LUT2 #(
		.INIT('h4)
	) name4327 (
		_w5274_,
		_w5282_,
		_w5286_
	);
	LUT2 #(
		.INIT('h4)
	) name4328 (
		_w5281_,
		_w5286_,
		_w5287_
	);
	LUT2 #(
		.INIT('h8)
	) name4329 (
		_w5285_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h1)
	) name4330 (
		_w5273_,
		_w5288_,
		_w5289_
	);
	LUT2 #(
		.INIT('h4)
	) name4331 (
		_w2231_,
		_w5064_,
		_w5290_
	);
	LUT2 #(
		.INIT('h4)
	) name4332 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[3]/P0001 ,
		_w5291_
	);
	LUT2 #(
		.INIT('h8)
	) name4333 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[3]/P0001 ,
		_w5292_
	);
	LUT2 #(
		.INIT('h1)
	) name4334 (
		_w5291_,
		_w5292_,
		_w5293_
	);
	LUT2 #(
		.INIT('h1)
	) name4335 (
		_w5064_,
		_w5293_,
		_w5294_
	);
	LUT2 #(
		.INIT('h2)
	) name4336 (
		_w2269_,
		_w5294_,
		_w5295_
	);
	LUT2 #(
		.INIT('h4)
	) name4337 (
		_w5290_,
		_w5295_,
		_w5296_
	);
	LUT2 #(
		.INIT('h8)
	) name4338 (
		\poc_o[3]_pad ,
		_w5091_,
		_w5297_
	);
	LUT2 #(
		.INIT('h8)
	) name4339 (
		\u0_u1_csc_reg[3]/NET0131 ,
		_w5081_,
		_w5298_
	);
	LUT2 #(
		.INIT('h8)
	) name4340 (
		\u0_csc_mask_r_reg[3]/NET0131 ,
		_w5277_,
		_w5299_
	);
	LUT2 #(
		.INIT('h8)
	) name4341 (
		\u0_u0_csc_reg[3]/NET0131 ,
		_w5083_,
		_w5300_
	);
	LUT2 #(
		.INIT('h8)
	) name4342 (
		\u0_u1_tms_reg[3]/P0001 ,
		_w5086_,
		_w5301_
	);
	LUT2 #(
		.INIT('h8)
	) name4343 (
		\u0_csr_r_reg[3]/NET0131 ,
		_w5089_,
		_w5302_
	);
	LUT2 #(
		.INIT('h8)
	) name4344 (
		\u0_u0_tms_reg[3]/P0001 ,
		_w5077_,
		_w5303_
	);
	LUT2 #(
		.INIT('h1)
	) name4345 (
		_w2269_,
		_w5298_,
		_w5304_
	);
	LUT2 #(
		.INIT('h1)
	) name4346 (
		_w5299_,
		_w5300_,
		_w5305_
	);
	LUT2 #(
		.INIT('h1)
	) name4347 (
		_w5301_,
		_w5302_,
		_w5306_
	);
	LUT2 #(
		.INIT('h8)
	) name4348 (
		_w5305_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('h4)
	) name4349 (
		_w5297_,
		_w5304_,
		_w5308_
	);
	LUT2 #(
		.INIT('h4)
	) name4350 (
		_w5303_,
		_w5308_,
		_w5309_
	);
	LUT2 #(
		.INIT('h8)
	) name4351 (
		_w5307_,
		_w5309_,
		_w5310_
	);
	LUT2 #(
		.INIT('h1)
	) name4352 (
		_w5296_,
		_w5310_,
		_w5311_
	);
	LUT2 #(
		.INIT('h4)
	) name4353 (
		_w2224_,
		_w5064_,
		_w5312_
	);
	LUT2 #(
		.INIT('h4)
	) name4354 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[5]/P0001 ,
		_w5313_
	);
	LUT2 #(
		.INIT('h8)
	) name4355 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[5]/P0001 ,
		_w5314_
	);
	LUT2 #(
		.INIT('h1)
	) name4356 (
		_w5313_,
		_w5314_,
		_w5315_
	);
	LUT2 #(
		.INIT('h1)
	) name4357 (
		_w5064_,
		_w5315_,
		_w5316_
	);
	LUT2 #(
		.INIT('h2)
	) name4358 (
		_w2269_,
		_w5316_,
		_w5317_
	);
	LUT2 #(
		.INIT('h4)
	) name4359 (
		_w5312_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h8)
	) name4360 (
		\u0_u0_tms_reg[5]/P0001 ,
		_w5077_,
		_w5319_
	);
	LUT2 #(
		.INIT('h8)
	) name4361 (
		\u0_u0_csc_reg[5]/P0001 ,
		_w5083_,
		_w5320_
	);
	LUT2 #(
		.INIT('h8)
	) name4362 (
		\u0_csc_mask_r_reg[5]/NET0131 ,
		_w5277_,
		_w5321_
	);
	LUT2 #(
		.INIT('h8)
	) name4363 (
		\u0_u1_tms_reg[5]/P0001 ,
		_w5086_,
		_w5322_
	);
	LUT2 #(
		.INIT('h8)
	) name4364 (
		\u0_u1_csc_reg[5]/P0001 ,
		_w5081_,
		_w5323_
	);
	LUT2 #(
		.INIT('h8)
	) name4365 (
		\u0_csr_r_reg[5]/NET0131 ,
		_w5089_,
		_w5324_
	);
	LUT2 #(
		.INIT('h8)
	) name4366 (
		\poc_o[5]_pad ,
		_w5091_,
		_w5325_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		_w2269_,
		_w5320_,
		_w5326_
	);
	LUT2 #(
		.INIT('h1)
	) name4368 (
		_w5321_,
		_w5322_,
		_w5327_
	);
	LUT2 #(
		.INIT('h1)
	) name4369 (
		_w5323_,
		_w5324_,
		_w5328_
	);
	LUT2 #(
		.INIT('h8)
	) name4370 (
		_w5327_,
		_w5328_,
		_w5329_
	);
	LUT2 #(
		.INIT('h4)
	) name4371 (
		_w5319_,
		_w5326_,
		_w5330_
	);
	LUT2 #(
		.INIT('h4)
	) name4372 (
		_w5325_,
		_w5330_,
		_w5331_
	);
	LUT2 #(
		.INIT('h8)
	) name4373 (
		_w5329_,
		_w5331_,
		_w5332_
	);
	LUT2 #(
		.INIT('h1)
	) name4374 (
		_w5318_,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('h4)
	) name4375 (
		_w1920_,
		_w5064_,
		_w5334_
	);
	LUT2 #(
		.INIT('h4)
	) name4376 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[1]/P0001 ,
		_w5335_
	);
	LUT2 #(
		.INIT('h8)
	) name4377 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[9]/P0001 ,
		_w5336_
	);
	LUT2 #(
		.INIT('h1)
	) name4378 (
		_w5335_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h1)
	) name4379 (
		_w5064_,
		_w5337_,
		_w5338_
	);
	LUT2 #(
		.INIT('h2)
	) name4380 (
		_w2269_,
		_w5338_,
		_w5339_
	);
	LUT2 #(
		.INIT('h4)
	) name4381 (
		_w5334_,
		_w5339_,
		_w5340_
	);
	LUT2 #(
		.INIT('h8)
	) name4382 (
		\u0_u0_tms_reg[9]/P0001 ,
		_w5077_,
		_w5341_
	);
	LUT2 #(
		.INIT('h8)
	) name4383 (
		\u0_csr_r_reg[9]/NET0131 ,
		_w5089_,
		_w5342_
	);
	LUT2 #(
		.INIT('h8)
	) name4384 (
		\u0_u1_csc_reg[9]/P0001 ,
		_w5081_,
		_w5343_
	);
	LUT2 #(
		.INIT('h8)
	) name4385 (
		\u0_u1_tms_reg[9]/P0001 ,
		_w5086_,
		_w5344_
	);
	LUT2 #(
		.INIT('h8)
	) name4386 (
		\u0_u0_csc_reg[9]/P0001 ,
		_w5083_,
		_w5345_
	);
	LUT2 #(
		.INIT('h8)
	) name4387 (
		\u0_csc_mask_r_reg[9]/NET0131 ,
		_w5277_,
		_w5346_
	);
	LUT2 #(
		.INIT('h8)
	) name4388 (
		\poc_o[9]_pad ,
		_w5091_,
		_w5347_
	);
	LUT2 #(
		.INIT('h1)
	) name4389 (
		_w2269_,
		_w5342_,
		_w5348_
	);
	LUT2 #(
		.INIT('h1)
	) name4390 (
		_w5343_,
		_w5344_,
		_w5349_
	);
	LUT2 #(
		.INIT('h1)
	) name4391 (
		_w5345_,
		_w5346_,
		_w5350_
	);
	LUT2 #(
		.INIT('h8)
	) name4392 (
		_w5349_,
		_w5350_,
		_w5351_
	);
	LUT2 #(
		.INIT('h4)
	) name4393 (
		_w5341_,
		_w5348_,
		_w5352_
	);
	LUT2 #(
		.INIT('h4)
	) name4394 (
		_w5347_,
		_w5352_,
		_w5353_
	);
	LUT2 #(
		.INIT('h8)
	) name4395 (
		_w5351_,
		_w5353_,
		_w5354_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		_w5340_,
		_w5354_,
		_w5355_
	);
	LUT2 #(
		.INIT('h4)
	) name4397 (
		_w2208_,
		_w5064_,
		_w5356_
	);
	LUT2 #(
		.INIT('h4)
	) name4398 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[6]/P0001 ,
		_w5357_
	);
	LUT2 #(
		.INIT('h8)
	) name4399 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[6]/P0001 ,
		_w5358_
	);
	LUT2 #(
		.INIT('h1)
	) name4400 (
		_w5357_,
		_w5358_,
		_w5359_
	);
	LUT2 #(
		.INIT('h1)
	) name4401 (
		_w5064_,
		_w5359_,
		_w5360_
	);
	LUT2 #(
		.INIT('h2)
	) name4402 (
		_w2269_,
		_w5360_,
		_w5361_
	);
	LUT2 #(
		.INIT('h4)
	) name4403 (
		_w5356_,
		_w5361_,
		_w5362_
	);
	LUT2 #(
		.INIT('h8)
	) name4404 (
		\u0_u0_tms_reg[6]/P0001 ,
		_w5077_,
		_w5363_
	);
	LUT2 #(
		.INIT('h8)
	) name4405 (
		\u0_u1_tms_reg[6]/P0001 ,
		_w5086_,
		_w5364_
	);
	LUT2 #(
		.INIT('h8)
	) name4406 (
		\u0_u0_csc_reg[6]/P0001 ,
		_w5083_,
		_w5365_
	);
	LUT2 #(
		.INIT('h8)
	) name4407 (
		\u0_u1_csc_reg[6]/P0001 ,
		_w5081_,
		_w5366_
	);
	LUT2 #(
		.INIT('h8)
	) name4408 (
		\u0_csc_mask_r_reg[6]/NET0131 ,
		_w5277_,
		_w5367_
	);
	LUT2 #(
		.INIT('h8)
	) name4409 (
		\u0_csr_r_reg[6]/NET0131 ,
		_w5089_,
		_w5368_
	);
	LUT2 #(
		.INIT('h8)
	) name4410 (
		\poc_o[6]_pad ,
		_w5091_,
		_w5369_
	);
	LUT2 #(
		.INIT('h1)
	) name4411 (
		_w2269_,
		_w5364_,
		_w5370_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		_w5365_,
		_w5366_,
		_w5371_
	);
	LUT2 #(
		.INIT('h1)
	) name4413 (
		_w5367_,
		_w5368_,
		_w5372_
	);
	LUT2 #(
		.INIT('h8)
	) name4414 (
		_w5371_,
		_w5372_,
		_w5373_
	);
	LUT2 #(
		.INIT('h4)
	) name4415 (
		_w5363_,
		_w5370_,
		_w5374_
	);
	LUT2 #(
		.INIT('h4)
	) name4416 (
		_w5369_,
		_w5374_,
		_w5375_
	);
	LUT2 #(
		.INIT('h8)
	) name4417 (
		_w5373_,
		_w5375_,
		_w5376_
	);
	LUT2 #(
		.INIT('h1)
	) name4418 (
		_w5362_,
		_w5376_,
		_w5377_
	);
	LUT2 #(
		.INIT('h4)
	) name4419 (
		_w2194_,
		_w5064_,
		_w5378_
	);
	LUT2 #(
		.INIT('h4)
	) name4420 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[4]/P0001 ,
		_w5379_
	);
	LUT2 #(
		.INIT('h8)
	) name4421 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[4]/P0001 ,
		_w5380_
	);
	LUT2 #(
		.INIT('h1)
	) name4422 (
		_w5379_,
		_w5380_,
		_w5381_
	);
	LUT2 #(
		.INIT('h1)
	) name4423 (
		_w5064_,
		_w5381_,
		_w5382_
	);
	LUT2 #(
		.INIT('h2)
	) name4424 (
		_w2269_,
		_w5382_,
		_w5383_
	);
	LUT2 #(
		.INIT('h4)
	) name4425 (
		_w5378_,
		_w5383_,
		_w5384_
	);
	LUT2 #(
		.INIT('h8)
	) name4426 (
		\u0_u0_tms_reg[4]/P0001 ,
		_w5077_,
		_w5385_
	);
	LUT2 #(
		.INIT('h8)
	) name4427 (
		\u0_u1_tms_reg[4]/P0001 ,
		_w5086_,
		_w5386_
	);
	LUT2 #(
		.INIT('h8)
	) name4428 (
		\u0_u0_csc_reg[4]/P0001 ,
		_w5083_,
		_w5387_
	);
	LUT2 #(
		.INIT('h8)
	) name4429 (
		\u0_u1_csc_reg[4]/P0001 ,
		_w5081_,
		_w5388_
	);
	LUT2 #(
		.INIT('h8)
	) name4430 (
		\u0_csc_mask_r_reg[4]/NET0131 ,
		_w5277_,
		_w5389_
	);
	LUT2 #(
		.INIT('h8)
	) name4431 (
		\u0_csr_r_reg[4]/NET0131 ,
		_w5089_,
		_w5390_
	);
	LUT2 #(
		.INIT('h8)
	) name4432 (
		\poc_o[4]_pad ,
		_w5091_,
		_w5391_
	);
	LUT2 #(
		.INIT('h1)
	) name4433 (
		_w2269_,
		_w5386_,
		_w5392_
	);
	LUT2 #(
		.INIT('h1)
	) name4434 (
		_w5387_,
		_w5388_,
		_w5393_
	);
	LUT2 #(
		.INIT('h1)
	) name4435 (
		_w5389_,
		_w5390_,
		_w5394_
	);
	LUT2 #(
		.INIT('h8)
	) name4436 (
		_w5393_,
		_w5394_,
		_w5395_
	);
	LUT2 #(
		.INIT('h4)
	) name4437 (
		_w5385_,
		_w5392_,
		_w5396_
	);
	LUT2 #(
		.INIT('h4)
	) name4438 (
		_w5391_,
		_w5396_,
		_w5397_
	);
	LUT2 #(
		.INIT('h8)
	) name4439 (
		_w5395_,
		_w5397_,
		_w5398_
	);
	LUT2 #(
		.INIT('h1)
	) name4440 (
		_w5384_,
		_w5398_,
		_w5399_
	);
	LUT2 #(
		.INIT('h8)
	) name4441 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1146_,
		_w5400_
	);
	LUT2 #(
		.INIT('h8)
	) name4442 (
		\u5_state_reg[45]/NET0131 ,
		_w2606_,
		_w5401_
	);
	LUT2 #(
		.INIT('h8)
	) name4443 (
		_w3075_,
		_w4388_,
		_w5402_
	);
	LUT2 #(
		.INIT('h8)
	) name4444 (
		_w3073_,
		_w5402_,
		_w5403_
	);
	LUT2 #(
		.INIT('h8)
	) name4445 (
		_w4386_,
		_w5403_,
		_w5404_
	);
	LUT2 #(
		.INIT('h8)
	) name4446 (
		_w964_,
		_w989_,
		_w5405_
	);
	LUT2 #(
		.INIT('h8)
	) name4447 (
		_w1257_,
		_w1340_,
		_w5406_
	);
	LUT2 #(
		.INIT('h8)
	) name4448 (
		_w5405_,
		_w5406_,
		_w5407_
	);
	LUT2 #(
		.INIT('h8)
	) name4449 (
		_w1336_,
		_w5407_,
		_w5408_
	);
	LUT2 #(
		.INIT('h8)
	) name4450 (
		_w5404_,
		_w5408_,
		_w5409_
	);
	LUT2 #(
		.INIT('h1)
	) name4451 (
		_w5401_,
		_w5409_,
		_w5410_
	);
	LUT2 #(
		.INIT('h1)
	) name4452 (
		\u1_acs_addr_reg[10]/P0001 ,
		_w4009_,
		_w5411_
	);
	LUT2 #(
		.INIT('h1)
	) name4453 (
		_w4010_,
		_w5411_,
		_w5412_
	);
	LUT2 #(
		.INIT('h8)
	) name4454 (
		\u0_init_ack_r_reg/P0001 ,
		_w1050_,
		_w5413_
	);
	LUT2 #(
		.INIT('h8)
	) name4455 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		_w5413_,
		_w5414_
	);
	LUT2 #(
		.INIT('h2)
	) name4456 (
		\u0_u0_init_req_reg/NET0131 ,
		_w5414_,
		_w5415_
	);
	LUT2 #(
		.INIT('h2)
	) name4457 (
		\u0_u0_init_req_we_reg/NET0131 ,
		\u0_u0_inited_reg/NET0131 ,
		_w5416_
	);
	LUT2 #(
		.INIT('h8)
	) name4458 (
		_w1621_,
		_w5416_,
		_w5417_
	);
	LUT2 #(
		.INIT('h1)
	) name4459 (
		_w5415_,
		_w5417_,
		_w5418_
	);
	LUT2 #(
		.INIT('h8)
	) name4460 (
		\u0_spec_req_cs_reg[1]/NET0131 ,
		_w5413_,
		_w5419_
	);
	LUT2 #(
		.INIT('h2)
	) name4461 (
		\u0_u1_init_req_reg/NET0131 ,
		_w5419_,
		_w5420_
	);
	LUT2 #(
		.INIT('h2)
	) name4462 (
		\u0_u1_init_req_we_reg/NET0131 ,
		\u0_u1_inited_reg/NET0131 ,
		_w5421_
	);
	LUT2 #(
		.INIT('h8)
	) name4463 (
		_w1674_,
		_w5421_,
		_w5422_
	);
	LUT2 #(
		.INIT('h1)
	) name4464 (
		_w5420_,
		_w5422_,
		_w5423_
	);
	LUT2 #(
		.INIT('h8)
	) name4465 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1272_,
		_w5424_
	);
	LUT2 #(
		.INIT('h8)
	) name4466 (
		_w2136_,
		_w5064_,
		_w5425_
	);
	LUT2 #(
		.INIT('h8)
	) name4467 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[16]/P0001 ,
		_w5426_
	);
	LUT2 #(
		.INIT('h8)
	) name4468 (
		\u7_mc_data_ir_reg[0]/P0001 ,
		_w4153_,
		_w5427_
	);
	LUT2 #(
		.INIT('h8)
	) name4469 (
		\u3_byte2_reg[0]/P0001 ,
		_w4151_,
		_w5428_
	);
	LUT2 #(
		.INIT('h1)
	) name4470 (
		_w5064_,
		_w5426_,
		_w5429_
	);
	LUT2 #(
		.INIT('h4)
	) name4471 (
		_w5427_,
		_w5429_,
		_w5430_
	);
	LUT2 #(
		.INIT('h4)
	) name4472 (
		_w5428_,
		_w5430_,
		_w5431_
	);
	LUT2 #(
		.INIT('h1)
	) name4473 (
		_w5425_,
		_w5431_,
		_w5432_
	);
	LUT2 #(
		.INIT('h2)
	) name4474 (
		_w2269_,
		_w5432_,
		_w5433_
	);
	LUT2 #(
		.INIT('h8)
	) name4475 (
		\u0_u0_tms_reg[16]/P0001 ,
		_w5077_,
		_w5434_
	);
	LUT2 #(
		.INIT('h8)
	) name4476 (
		\u0_u1_csc_reg[16]/P0001 ,
		_w5081_,
		_w5435_
	);
	LUT2 #(
		.INIT('h8)
	) name4477 (
		\u0_u1_tms_reg[16]/P0001 ,
		_w5086_,
		_w5436_
	);
	LUT2 #(
		.INIT('h8)
	) name4478 (
		\u0_u0_csc_reg[16]/P0001 ,
		_w5083_,
		_w5437_
	);
	LUT2 #(
		.INIT('h8)
	) name4479 (
		\poc_o[16]_pad ,
		_w5091_,
		_w5438_
	);
	LUT2 #(
		.INIT('h1)
	) name4480 (
		_w2269_,
		_w5435_,
		_w5439_
	);
	LUT2 #(
		.INIT('h1)
	) name4481 (
		_w5436_,
		_w5437_,
		_w5440_
	);
	LUT2 #(
		.INIT('h8)
	) name4482 (
		_w5439_,
		_w5440_,
		_w5441_
	);
	LUT2 #(
		.INIT('h1)
	) name4483 (
		_w5434_,
		_w5438_,
		_w5442_
	);
	LUT2 #(
		.INIT('h8)
	) name4484 (
		_w5441_,
		_w5442_,
		_w5443_
	);
	LUT2 #(
		.INIT('h1)
	) name4485 (
		_w5433_,
		_w5443_,
		_w5444_
	);
	LUT2 #(
		.INIT('h8)
	) name4486 (
		_w2096_,
		_w5064_,
		_w5445_
	);
	LUT2 #(
		.INIT('h8)
	) name4487 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[17]/P0001 ,
		_w5446_
	);
	LUT2 #(
		.INIT('h8)
	) name4488 (
		\u7_mc_data_ir_reg[1]/P0001 ,
		_w4153_,
		_w5447_
	);
	LUT2 #(
		.INIT('h8)
	) name4489 (
		\u3_byte2_reg[1]/P0001 ,
		_w4151_,
		_w5448_
	);
	LUT2 #(
		.INIT('h1)
	) name4490 (
		_w5064_,
		_w5446_,
		_w5449_
	);
	LUT2 #(
		.INIT('h4)
	) name4491 (
		_w5447_,
		_w5449_,
		_w5450_
	);
	LUT2 #(
		.INIT('h4)
	) name4492 (
		_w5448_,
		_w5450_,
		_w5451_
	);
	LUT2 #(
		.INIT('h1)
	) name4493 (
		_w5445_,
		_w5451_,
		_w5452_
	);
	LUT2 #(
		.INIT('h2)
	) name4494 (
		_w2269_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h8)
	) name4495 (
		\u0_u0_tms_reg[17]/P0001 ,
		_w5077_,
		_w5454_
	);
	LUT2 #(
		.INIT('h8)
	) name4496 (
		\u0_u1_csc_reg[17]/P0001 ,
		_w5081_,
		_w5455_
	);
	LUT2 #(
		.INIT('h8)
	) name4497 (
		\u0_u1_tms_reg[17]/P0001 ,
		_w5086_,
		_w5456_
	);
	LUT2 #(
		.INIT('h8)
	) name4498 (
		\u0_u0_csc_reg[17]/P0001 ,
		_w5083_,
		_w5457_
	);
	LUT2 #(
		.INIT('h8)
	) name4499 (
		\poc_o[17]_pad ,
		_w5091_,
		_w5458_
	);
	LUT2 #(
		.INIT('h1)
	) name4500 (
		_w2269_,
		_w5455_,
		_w5459_
	);
	LUT2 #(
		.INIT('h1)
	) name4501 (
		_w5456_,
		_w5457_,
		_w5460_
	);
	LUT2 #(
		.INIT('h8)
	) name4502 (
		_w5459_,
		_w5460_,
		_w5461_
	);
	LUT2 #(
		.INIT('h1)
	) name4503 (
		_w5454_,
		_w5458_,
		_w5462_
	);
	LUT2 #(
		.INIT('h8)
	) name4504 (
		_w5461_,
		_w5462_,
		_w5463_
	);
	LUT2 #(
		.INIT('h1)
	) name4505 (
		_w5453_,
		_w5463_,
		_w5464_
	);
	LUT2 #(
		.INIT('h8)
	) name4506 (
		_w2160_,
		_w5064_,
		_w5465_
	);
	LUT2 #(
		.INIT('h8)
	) name4507 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[18]/P0001 ,
		_w5466_
	);
	LUT2 #(
		.INIT('h8)
	) name4508 (
		\u7_mc_data_ir_reg[2]/P0001 ,
		_w4153_,
		_w5467_
	);
	LUT2 #(
		.INIT('h8)
	) name4509 (
		\u3_byte2_reg[2]/P0001 ,
		_w4151_,
		_w5468_
	);
	LUT2 #(
		.INIT('h1)
	) name4510 (
		_w5064_,
		_w5466_,
		_w5469_
	);
	LUT2 #(
		.INIT('h4)
	) name4511 (
		_w5467_,
		_w5469_,
		_w5470_
	);
	LUT2 #(
		.INIT('h4)
	) name4512 (
		_w5468_,
		_w5470_,
		_w5471_
	);
	LUT2 #(
		.INIT('h1)
	) name4513 (
		_w5465_,
		_w5471_,
		_w5472_
	);
	LUT2 #(
		.INIT('h2)
	) name4514 (
		_w2269_,
		_w5472_,
		_w5473_
	);
	LUT2 #(
		.INIT('h8)
	) name4515 (
		\u0_u0_tms_reg[18]/P0001 ,
		_w5077_,
		_w5474_
	);
	LUT2 #(
		.INIT('h8)
	) name4516 (
		\u0_u1_csc_reg[18]/P0001 ,
		_w5081_,
		_w5475_
	);
	LUT2 #(
		.INIT('h8)
	) name4517 (
		\u0_u1_tms_reg[18]/P0001 ,
		_w5086_,
		_w5476_
	);
	LUT2 #(
		.INIT('h8)
	) name4518 (
		\u0_u0_csc_reg[18]/P0001 ,
		_w5083_,
		_w5477_
	);
	LUT2 #(
		.INIT('h8)
	) name4519 (
		\poc_o[18]_pad ,
		_w5091_,
		_w5478_
	);
	LUT2 #(
		.INIT('h1)
	) name4520 (
		_w2269_,
		_w5475_,
		_w5479_
	);
	LUT2 #(
		.INIT('h1)
	) name4521 (
		_w5476_,
		_w5477_,
		_w5480_
	);
	LUT2 #(
		.INIT('h8)
	) name4522 (
		_w5479_,
		_w5480_,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name4523 (
		_w5474_,
		_w5478_,
		_w5482_
	);
	LUT2 #(
		.INIT('h8)
	) name4524 (
		_w5481_,
		_w5482_,
		_w5483_
	);
	LUT2 #(
		.INIT('h1)
	) name4525 (
		_w5473_,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h8)
	) name4526 (
		_w2113_,
		_w5064_,
		_w5485_
	);
	LUT2 #(
		.INIT('h8)
	) name4527 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[19]/P0001 ,
		_w5486_
	);
	LUT2 #(
		.INIT('h8)
	) name4528 (
		\u7_mc_data_ir_reg[3]/P0001 ,
		_w4153_,
		_w5487_
	);
	LUT2 #(
		.INIT('h8)
	) name4529 (
		\u3_byte2_reg[3]/P0001 ,
		_w4151_,
		_w5488_
	);
	LUT2 #(
		.INIT('h1)
	) name4530 (
		_w5064_,
		_w5486_,
		_w5489_
	);
	LUT2 #(
		.INIT('h4)
	) name4531 (
		_w5487_,
		_w5489_,
		_w5490_
	);
	LUT2 #(
		.INIT('h4)
	) name4532 (
		_w5488_,
		_w5490_,
		_w5491_
	);
	LUT2 #(
		.INIT('h1)
	) name4533 (
		_w5485_,
		_w5491_,
		_w5492_
	);
	LUT2 #(
		.INIT('h2)
	) name4534 (
		_w2269_,
		_w5492_,
		_w5493_
	);
	LUT2 #(
		.INIT('h8)
	) name4535 (
		\u0_u0_tms_reg[19]/P0001 ,
		_w5077_,
		_w5494_
	);
	LUT2 #(
		.INIT('h8)
	) name4536 (
		\u0_u1_csc_reg[19]/P0001 ,
		_w5081_,
		_w5495_
	);
	LUT2 #(
		.INIT('h8)
	) name4537 (
		\u0_u1_tms_reg[19]/P0001 ,
		_w5086_,
		_w5496_
	);
	LUT2 #(
		.INIT('h8)
	) name4538 (
		\u0_u0_csc_reg[19]/P0001 ,
		_w5083_,
		_w5497_
	);
	LUT2 #(
		.INIT('h8)
	) name4539 (
		\poc_o[19]_pad ,
		_w5091_,
		_w5498_
	);
	LUT2 #(
		.INIT('h1)
	) name4540 (
		_w2269_,
		_w5495_,
		_w5499_
	);
	LUT2 #(
		.INIT('h1)
	) name4541 (
		_w5496_,
		_w5497_,
		_w5500_
	);
	LUT2 #(
		.INIT('h8)
	) name4542 (
		_w5499_,
		_w5500_,
		_w5501_
	);
	LUT2 #(
		.INIT('h1)
	) name4543 (
		_w5494_,
		_w5498_,
		_w5502_
	);
	LUT2 #(
		.INIT('h8)
	) name4544 (
		_w5501_,
		_w5502_,
		_w5503_
	);
	LUT2 #(
		.INIT('h1)
	) name4545 (
		_w5493_,
		_w5503_,
		_w5504_
	);
	LUT2 #(
		.INIT('h8)
	) name4546 (
		_w2120_,
		_w5064_,
		_w5505_
	);
	LUT2 #(
		.INIT('h8)
	) name4547 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[20]/P0001 ,
		_w5506_
	);
	LUT2 #(
		.INIT('h8)
	) name4548 (
		\u7_mc_data_ir_reg[4]/P0001 ,
		_w4153_,
		_w5507_
	);
	LUT2 #(
		.INIT('h8)
	) name4549 (
		\u3_byte2_reg[4]/P0001 ,
		_w4151_,
		_w5508_
	);
	LUT2 #(
		.INIT('h1)
	) name4550 (
		_w5064_,
		_w5506_,
		_w5509_
	);
	LUT2 #(
		.INIT('h4)
	) name4551 (
		_w5507_,
		_w5509_,
		_w5510_
	);
	LUT2 #(
		.INIT('h4)
	) name4552 (
		_w5508_,
		_w5510_,
		_w5511_
	);
	LUT2 #(
		.INIT('h1)
	) name4553 (
		_w5505_,
		_w5511_,
		_w5512_
	);
	LUT2 #(
		.INIT('h2)
	) name4554 (
		_w2269_,
		_w5512_,
		_w5513_
	);
	LUT2 #(
		.INIT('h8)
	) name4555 (
		\u0_u0_tms_reg[20]/P0001 ,
		_w5077_,
		_w5514_
	);
	LUT2 #(
		.INIT('h8)
	) name4556 (
		\u0_u1_csc_reg[20]/P0001 ,
		_w5081_,
		_w5515_
	);
	LUT2 #(
		.INIT('h8)
	) name4557 (
		\u0_u1_tms_reg[20]/P0001 ,
		_w5086_,
		_w5516_
	);
	LUT2 #(
		.INIT('h8)
	) name4558 (
		\u0_u0_csc_reg[20]/P0001 ,
		_w5083_,
		_w5517_
	);
	LUT2 #(
		.INIT('h8)
	) name4559 (
		\poc_o[20]_pad ,
		_w5091_,
		_w5518_
	);
	LUT2 #(
		.INIT('h1)
	) name4560 (
		_w2269_,
		_w5515_,
		_w5519_
	);
	LUT2 #(
		.INIT('h1)
	) name4561 (
		_w5516_,
		_w5517_,
		_w5520_
	);
	LUT2 #(
		.INIT('h8)
	) name4562 (
		_w5519_,
		_w5520_,
		_w5521_
	);
	LUT2 #(
		.INIT('h1)
	) name4563 (
		_w5514_,
		_w5518_,
		_w5522_
	);
	LUT2 #(
		.INIT('h8)
	) name4564 (
		_w5521_,
		_w5522_,
		_w5523_
	);
	LUT2 #(
		.INIT('h1)
	) name4565 (
		_w5513_,
		_w5523_,
		_w5524_
	);
	LUT2 #(
		.INIT('h8)
	) name4566 (
		_w2106_,
		_w5064_,
		_w5525_
	);
	LUT2 #(
		.INIT('h8)
	) name4567 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[22]/P0001 ,
		_w5526_
	);
	LUT2 #(
		.INIT('h8)
	) name4568 (
		\u7_mc_data_ir_reg[6]/P0001 ,
		_w4153_,
		_w5527_
	);
	LUT2 #(
		.INIT('h8)
	) name4569 (
		\u3_byte2_reg[6]/P0001 ,
		_w4151_,
		_w5528_
	);
	LUT2 #(
		.INIT('h1)
	) name4570 (
		_w5064_,
		_w5526_,
		_w5529_
	);
	LUT2 #(
		.INIT('h4)
	) name4571 (
		_w5527_,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('h4)
	) name4572 (
		_w5528_,
		_w5530_,
		_w5531_
	);
	LUT2 #(
		.INIT('h1)
	) name4573 (
		_w5525_,
		_w5531_,
		_w5532_
	);
	LUT2 #(
		.INIT('h2)
	) name4574 (
		_w2269_,
		_w5532_,
		_w5533_
	);
	LUT2 #(
		.INIT('h8)
	) name4575 (
		\u0_u0_tms_reg[22]/P0001 ,
		_w5077_,
		_w5534_
	);
	LUT2 #(
		.INIT('h8)
	) name4576 (
		\u0_u1_csc_reg[22]/P0001 ,
		_w5081_,
		_w5535_
	);
	LUT2 #(
		.INIT('h8)
	) name4577 (
		\u0_u1_tms_reg[22]/P0001 ,
		_w5086_,
		_w5536_
	);
	LUT2 #(
		.INIT('h8)
	) name4578 (
		\u0_u0_csc_reg[22]/P0001 ,
		_w5083_,
		_w5537_
	);
	LUT2 #(
		.INIT('h8)
	) name4579 (
		\poc_o[22]_pad ,
		_w5091_,
		_w5538_
	);
	LUT2 #(
		.INIT('h1)
	) name4580 (
		_w2269_,
		_w5535_,
		_w5539_
	);
	LUT2 #(
		.INIT('h1)
	) name4581 (
		_w5536_,
		_w5537_,
		_w5540_
	);
	LUT2 #(
		.INIT('h8)
	) name4582 (
		_w5539_,
		_w5540_,
		_w5541_
	);
	LUT2 #(
		.INIT('h1)
	) name4583 (
		_w5534_,
		_w5538_,
		_w5542_
	);
	LUT2 #(
		.INIT('h8)
	) name4584 (
		_w5541_,
		_w5542_,
		_w5543_
	);
	LUT2 #(
		.INIT('h1)
	) name4585 (
		_w5533_,
		_w5543_,
		_w5544_
	);
	LUT2 #(
		.INIT('h8)
	) name4586 (
		_w2143_,
		_w5064_,
		_w5545_
	);
	LUT2 #(
		.INIT('h8)
	) name4587 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[23]/P0001 ,
		_w5546_
	);
	LUT2 #(
		.INIT('h8)
	) name4588 (
		\u7_mc_data_ir_reg[7]/P0001 ,
		_w4153_,
		_w5547_
	);
	LUT2 #(
		.INIT('h8)
	) name4589 (
		\u3_byte2_reg[7]/P0001 ,
		_w4151_,
		_w5548_
	);
	LUT2 #(
		.INIT('h1)
	) name4590 (
		_w5064_,
		_w5546_,
		_w5549_
	);
	LUT2 #(
		.INIT('h4)
	) name4591 (
		_w5547_,
		_w5549_,
		_w5550_
	);
	LUT2 #(
		.INIT('h4)
	) name4592 (
		_w5548_,
		_w5550_,
		_w5551_
	);
	LUT2 #(
		.INIT('h1)
	) name4593 (
		_w5545_,
		_w5551_,
		_w5552_
	);
	LUT2 #(
		.INIT('h2)
	) name4594 (
		_w2269_,
		_w5552_,
		_w5553_
	);
	LUT2 #(
		.INIT('h8)
	) name4595 (
		\u0_u0_tms_reg[23]/P0001 ,
		_w5077_,
		_w5554_
	);
	LUT2 #(
		.INIT('h8)
	) name4596 (
		\u0_u1_csc_reg[23]/P0001 ,
		_w5081_,
		_w5555_
	);
	LUT2 #(
		.INIT('h8)
	) name4597 (
		\u0_u1_tms_reg[23]/P0001 ,
		_w5086_,
		_w5556_
	);
	LUT2 #(
		.INIT('h8)
	) name4598 (
		\u0_u0_csc_reg[23]/P0001 ,
		_w5083_,
		_w5557_
	);
	LUT2 #(
		.INIT('h8)
	) name4599 (
		\poc_o[23]_pad ,
		_w5091_,
		_w5558_
	);
	LUT2 #(
		.INIT('h1)
	) name4600 (
		_w2269_,
		_w5555_,
		_w5559_
	);
	LUT2 #(
		.INIT('h1)
	) name4601 (
		_w5556_,
		_w5557_,
		_w5560_
	);
	LUT2 #(
		.INIT('h8)
	) name4602 (
		_w5559_,
		_w5560_,
		_w5561_
	);
	LUT2 #(
		.INIT('h1)
	) name4603 (
		_w5554_,
		_w5558_,
		_w5562_
	);
	LUT2 #(
		.INIT('h8)
	) name4604 (
		_w5561_,
		_w5562_,
		_w5563_
	);
	LUT2 #(
		.INIT('h1)
	) name4605 (
		_w5553_,
		_w5563_,
		_w5564_
	);
	LUT2 #(
		.INIT('h8)
	) name4606 (
		_w2089_,
		_w5064_,
		_w5565_
	);
	LUT2 #(
		.INIT('h8)
	) name4607 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[21]/P0001 ,
		_w5566_
	);
	LUT2 #(
		.INIT('h8)
	) name4608 (
		\u7_mc_data_ir_reg[5]/P0001 ,
		_w4153_,
		_w5567_
	);
	LUT2 #(
		.INIT('h8)
	) name4609 (
		\u3_byte2_reg[5]/P0001 ,
		_w4151_,
		_w5568_
	);
	LUT2 #(
		.INIT('h1)
	) name4610 (
		_w5064_,
		_w5566_,
		_w5569_
	);
	LUT2 #(
		.INIT('h4)
	) name4611 (
		_w5567_,
		_w5569_,
		_w5570_
	);
	LUT2 #(
		.INIT('h4)
	) name4612 (
		_w5568_,
		_w5570_,
		_w5571_
	);
	LUT2 #(
		.INIT('h1)
	) name4613 (
		_w5565_,
		_w5571_,
		_w5572_
	);
	LUT2 #(
		.INIT('h2)
	) name4614 (
		_w2269_,
		_w5572_,
		_w5573_
	);
	LUT2 #(
		.INIT('h8)
	) name4615 (
		\u0_u0_tms_reg[21]/P0001 ,
		_w5077_,
		_w5574_
	);
	LUT2 #(
		.INIT('h8)
	) name4616 (
		\u0_u1_csc_reg[21]/P0001 ,
		_w5081_,
		_w5575_
	);
	LUT2 #(
		.INIT('h8)
	) name4617 (
		\u0_u1_tms_reg[21]/P0001 ,
		_w5086_,
		_w5576_
	);
	LUT2 #(
		.INIT('h8)
	) name4618 (
		\u0_u0_csc_reg[21]/P0001 ,
		_w5083_,
		_w5577_
	);
	LUT2 #(
		.INIT('h8)
	) name4619 (
		\poc_o[21]_pad ,
		_w5091_,
		_w5578_
	);
	LUT2 #(
		.INIT('h1)
	) name4620 (
		_w2269_,
		_w5575_,
		_w5579_
	);
	LUT2 #(
		.INIT('h1)
	) name4621 (
		_w5576_,
		_w5577_,
		_w5580_
	);
	LUT2 #(
		.INIT('h8)
	) name4622 (
		_w5579_,
		_w5580_,
		_w5581_
	);
	LUT2 #(
		.INIT('h1)
	) name4623 (
		_w5574_,
		_w5578_,
		_w5582_
	);
	LUT2 #(
		.INIT('h8)
	) name4624 (
		_w5581_,
		_w5582_,
		_w5583_
	);
	LUT2 #(
		.INIT('h1)
	) name4625 (
		_w5573_,
		_w5583_,
		_w5584_
	);
	LUT2 #(
		.INIT('h4)
	) name4626 (
		_w1937_,
		_w5064_,
		_w5585_
	);
	LUT2 #(
		.INIT('h4)
	) name4627 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[3]/P0001 ,
		_w5586_
	);
	LUT2 #(
		.INIT('h8)
	) name4628 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[11]/P0001 ,
		_w5587_
	);
	LUT2 #(
		.INIT('h1)
	) name4629 (
		_w5586_,
		_w5587_,
		_w5588_
	);
	LUT2 #(
		.INIT('h1)
	) name4630 (
		_w5064_,
		_w5588_,
		_w5589_
	);
	LUT2 #(
		.INIT('h2)
	) name4631 (
		_w2269_,
		_w5589_,
		_w5590_
	);
	LUT2 #(
		.INIT('h4)
	) name4632 (
		_w5585_,
		_w5590_,
		_w5591_
	);
	LUT2 #(
		.INIT('h8)
	) name4633 (
		\u0_u0_tms_reg[11]/P0001 ,
		_w5077_,
		_w5592_
	);
	LUT2 #(
		.INIT('h8)
	) name4634 (
		\u0_u1_csc_reg[11]/P0001 ,
		_w5081_,
		_w5593_
	);
	LUT2 #(
		.INIT('h8)
	) name4635 (
		\u0_u1_tms_reg[11]/P0001 ,
		_w5086_,
		_w5594_
	);
	LUT2 #(
		.INIT('h8)
	) name4636 (
		\u0_u0_csc_reg[11]/P0001 ,
		_w5083_,
		_w5595_
	);
	LUT2 #(
		.INIT('h8)
	) name4637 (
		\poc_o[11]_pad ,
		_w5091_,
		_w5596_
	);
	LUT2 #(
		.INIT('h1)
	) name4638 (
		_w2269_,
		_w5593_,
		_w5597_
	);
	LUT2 #(
		.INIT('h1)
	) name4639 (
		_w5594_,
		_w5595_,
		_w5598_
	);
	LUT2 #(
		.INIT('h8)
	) name4640 (
		_w5597_,
		_w5598_,
		_w5599_
	);
	LUT2 #(
		.INIT('h1)
	) name4641 (
		_w5592_,
		_w5596_,
		_w5600_
	);
	LUT2 #(
		.INIT('h8)
	) name4642 (
		_w5599_,
		_w5600_,
		_w5601_
	);
	LUT2 #(
		.INIT('h1)
	) name4643 (
		_w5591_,
		_w5601_,
		_w5602_
	);
	LUT2 #(
		.INIT('h4)
	) name4644 (
		_w1944_,
		_w5064_,
		_w5603_
	);
	LUT2 #(
		.INIT('h4)
	) name4645 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[4]/P0001 ,
		_w5604_
	);
	LUT2 #(
		.INIT('h8)
	) name4646 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[12]/P0001 ,
		_w5605_
	);
	LUT2 #(
		.INIT('h1)
	) name4647 (
		_w5604_,
		_w5605_,
		_w5606_
	);
	LUT2 #(
		.INIT('h1)
	) name4648 (
		_w5064_,
		_w5606_,
		_w5607_
	);
	LUT2 #(
		.INIT('h2)
	) name4649 (
		_w2269_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('h4)
	) name4650 (
		_w5603_,
		_w5608_,
		_w5609_
	);
	LUT2 #(
		.INIT('h8)
	) name4651 (
		\u0_u0_tms_reg[12]/P0001 ,
		_w5077_,
		_w5610_
	);
	LUT2 #(
		.INIT('h8)
	) name4652 (
		\u0_u1_csc_reg[12]/P0001 ,
		_w5081_,
		_w5611_
	);
	LUT2 #(
		.INIT('h8)
	) name4653 (
		\u0_u1_tms_reg[12]/P0001 ,
		_w5086_,
		_w5612_
	);
	LUT2 #(
		.INIT('h8)
	) name4654 (
		\u0_u0_csc_reg[12]/P0001 ,
		_w5083_,
		_w5613_
	);
	LUT2 #(
		.INIT('h8)
	) name4655 (
		\poc_o[12]_pad ,
		_w5091_,
		_w5614_
	);
	LUT2 #(
		.INIT('h1)
	) name4656 (
		_w2269_,
		_w5611_,
		_w5615_
	);
	LUT2 #(
		.INIT('h1)
	) name4657 (
		_w5612_,
		_w5613_,
		_w5616_
	);
	LUT2 #(
		.INIT('h8)
	) name4658 (
		_w5615_,
		_w5616_,
		_w5617_
	);
	LUT2 #(
		.INIT('h1)
	) name4659 (
		_w5610_,
		_w5614_,
		_w5618_
	);
	LUT2 #(
		.INIT('h8)
	) name4660 (
		_w5617_,
		_w5618_,
		_w5619_
	);
	LUT2 #(
		.INIT('h1)
	) name4661 (
		_w5609_,
		_w5619_,
		_w5620_
	);
	LUT2 #(
		.INIT('h4)
	) name4662 (
		_w1930_,
		_w5064_,
		_w5621_
	);
	LUT2 #(
		.INIT('h4)
	) name4663 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[6]/P0001 ,
		_w5622_
	);
	LUT2 #(
		.INIT('h8)
	) name4664 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[14]/P0001 ,
		_w5623_
	);
	LUT2 #(
		.INIT('h1)
	) name4665 (
		_w5622_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h1)
	) name4666 (
		_w5064_,
		_w5624_,
		_w5625_
	);
	LUT2 #(
		.INIT('h2)
	) name4667 (
		_w2269_,
		_w5625_,
		_w5626_
	);
	LUT2 #(
		.INIT('h4)
	) name4668 (
		_w5621_,
		_w5626_,
		_w5627_
	);
	LUT2 #(
		.INIT('h8)
	) name4669 (
		\u0_u0_tms_reg[14]/P0001 ,
		_w5077_,
		_w5628_
	);
	LUT2 #(
		.INIT('h8)
	) name4670 (
		\u0_u1_csc_reg[14]/P0001 ,
		_w5081_,
		_w5629_
	);
	LUT2 #(
		.INIT('h8)
	) name4671 (
		\u0_u1_tms_reg[14]/P0001 ,
		_w5086_,
		_w5630_
	);
	LUT2 #(
		.INIT('h8)
	) name4672 (
		\u0_u0_csc_reg[14]/P0001 ,
		_w5083_,
		_w5631_
	);
	LUT2 #(
		.INIT('h8)
	) name4673 (
		\poc_o[14]_pad ,
		_w5091_,
		_w5632_
	);
	LUT2 #(
		.INIT('h1)
	) name4674 (
		_w2269_,
		_w5629_,
		_w5633_
	);
	LUT2 #(
		.INIT('h1)
	) name4675 (
		_w5630_,
		_w5631_,
		_w5634_
	);
	LUT2 #(
		.INIT('h8)
	) name4676 (
		_w5633_,
		_w5634_,
		_w5635_
	);
	LUT2 #(
		.INIT('h1)
	) name4677 (
		_w5628_,
		_w5632_,
		_w5636_
	);
	LUT2 #(
		.INIT('h8)
	) name4678 (
		_w5635_,
		_w5636_,
		_w5637_
	);
	LUT2 #(
		.INIT('h1)
	) name4679 (
		_w5627_,
		_w5637_,
		_w5638_
	);
	LUT2 #(
		.INIT('h4)
	) name4680 (
		_w1967_,
		_w5064_,
		_w5639_
	);
	LUT2 #(
		.INIT('h4)
	) name4681 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[7]/P0001 ,
		_w5640_
	);
	LUT2 #(
		.INIT('h8)
	) name4682 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[15]/P0001 ,
		_w5641_
	);
	LUT2 #(
		.INIT('h1)
	) name4683 (
		_w5640_,
		_w5641_,
		_w5642_
	);
	LUT2 #(
		.INIT('h1)
	) name4684 (
		_w5064_,
		_w5642_,
		_w5643_
	);
	LUT2 #(
		.INIT('h2)
	) name4685 (
		_w2269_,
		_w5643_,
		_w5644_
	);
	LUT2 #(
		.INIT('h4)
	) name4686 (
		_w5639_,
		_w5644_,
		_w5645_
	);
	LUT2 #(
		.INIT('h8)
	) name4687 (
		\u0_u0_tms_reg[15]/P0001 ,
		_w5077_,
		_w5646_
	);
	LUT2 #(
		.INIT('h8)
	) name4688 (
		\u0_u1_csc_reg[15]/P0001 ,
		_w5081_,
		_w5647_
	);
	LUT2 #(
		.INIT('h8)
	) name4689 (
		\u0_u1_tms_reg[15]/P0001 ,
		_w5086_,
		_w5648_
	);
	LUT2 #(
		.INIT('h8)
	) name4690 (
		\u0_u0_csc_reg[15]/P0001 ,
		_w5083_,
		_w5649_
	);
	LUT2 #(
		.INIT('h8)
	) name4691 (
		\poc_o[15]_pad ,
		_w5091_,
		_w5650_
	);
	LUT2 #(
		.INIT('h1)
	) name4692 (
		_w2269_,
		_w5647_,
		_w5651_
	);
	LUT2 #(
		.INIT('h1)
	) name4693 (
		_w5648_,
		_w5649_,
		_w5652_
	);
	LUT2 #(
		.INIT('h8)
	) name4694 (
		_w5651_,
		_w5652_,
		_w5653_
	);
	LUT2 #(
		.INIT('h1)
	) name4695 (
		_w5646_,
		_w5650_,
		_w5654_
	);
	LUT2 #(
		.INIT('h8)
	) name4696 (
		_w5653_,
		_w5654_,
		_w5655_
	);
	LUT2 #(
		.INIT('h1)
	) name4697 (
		_w5645_,
		_w5655_,
		_w5656_
	);
	LUT2 #(
		.INIT('h4)
	) name4698 (
		_w1913_,
		_w5064_,
		_w5657_
	);
	LUT2 #(
		.INIT('h4)
	) name4699 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[5]/P0001 ,
		_w5658_
	);
	LUT2 #(
		.INIT('h8)
	) name4700 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[13]/P0001 ,
		_w5659_
	);
	LUT2 #(
		.INIT('h1)
	) name4701 (
		_w5658_,
		_w5659_,
		_w5660_
	);
	LUT2 #(
		.INIT('h1)
	) name4702 (
		_w5064_,
		_w5660_,
		_w5661_
	);
	LUT2 #(
		.INIT('h2)
	) name4703 (
		_w2269_,
		_w5661_,
		_w5662_
	);
	LUT2 #(
		.INIT('h4)
	) name4704 (
		_w5657_,
		_w5662_,
		_w5663_
	);
	LUT2 #(
		.INIT('h8)
	) name4705 (
		\u0_u0_tms_reg[13]/P0001 ,
		_w5077_,
		_w5664_
	);
	LUT2 #(
		.INIT('h8)
	) name4706 (
		\u0_u1_csc_reg[13]/P0001 ,
		_w5081_,
		_w5665_
	);
	LUT2 #(
		.INIT('h8)
	) name4707 (
		\u0_u1_tms_reg[13]/P0001 ,
		_w5086_,
		_w5666_
	);
	LUT2 #(
		.INIT('h8)
	) name4708 (
		\u0_u0_csc_reg[13]/P0001 ,
		_w5083_,
		_w5667_
	);
	LUT2 #(
		.INIT('h8)
	) name4709 (
		\poc_o[13]_pad ,
		_w5091_,
		_w5668_
	);
	LUT2 #(
		.INIT('h1)
	) name4710 (
		_w2269_,
		_w5665_,
		_w5669_
	);
	LUT2 #(
		.INIT('h1)
	) name4711 (
		_w5666_,
		_w5667_,
		_w5670_
	);
	LUT2 #(
		.INIT('h8)
	) name4712 (
		_w5669_,
		_w5670_,
		_w5671_
	);
	LUT2 #(
		.INIT('h1)
	) name4713 (
		_w5664_,
		_w5668_,
		_w5672_
	);
	LUT2 #(
		.INIT('h8)
	) name4714 (
		_w5671_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w5663_,
		_w5673_,
		_w5674_
	);
	LUT2 #(
		.INIT('h1)
	) name4716 (
		\u0_u0_csc_reg[1]/NET0131 ,
		_w5057_,
		_w5675_
	);
	LUT2 #(
		.INIT('h4)
	) name4717 (
		\wb_data_i[1]_pad ,
		_w5057_,
		_w5676_
	);
	LUT2 #(
		.INIT('h1)
	) name4718 (
		\u0_rst_r2_reg/NET0131 ,
		_w5675_,
		_w5677_
	);
	LUT2 #(
		.INIT('h4)
	) name4719 (
		_w5676_,
		_w5677_,
		_w5678_
	);
	LUT2 #(
		.INIT('h1)
	) name4720 (
		_w5052_,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h1)
	) name4721 (
		\u0_u0_csc_reg[2]/NET0131 ,
		_w5057_,
		_w5680_
	);
	LUT2 #(
		.INIT('h4)
	) name4722 (
		\wb_data_i[2]_pad ,
		_w5057_,
		_w5681_
	);
	LUT2 #(
		.INIT('h1)
	) name4723 (
		\u0_rst_r2_reg/NET0131 ,
		_w5680_,
		_w5682_
	);
	LUT2 #(
		.INIT('h4)
	) name4724 (
		_w5681_,
		_w5682_,
		_w5683_
	);
	LUT2 #(
		.INIT('h1)
	) name4725 (
		_w5051_,
		_w5683_,
		_w5684_
	);
	LUT2 #(
		.INIT('h1)
	) name4726 (
		\u1_acs_addr_reg[6]/P0001 ,
		_w4005_,
		_w5685_
	);
	LUT2 #(
		.INIT('h1)
	) name4727 (
		_w4006_,
		_w5685_,
		_w5686_
	);
	LUT2 #(
		.INIT('h4)
	) name4728 (
		_w2177_,
		_w5064_,
		_w5687_
	);
	LUT2 #(
		.INIT('h4)
	) name4729 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[0]/P0001 ,
		_w5688_
	);
	LUT2 #(
		.INIT('h8)
	) name4730 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[0]/P0001 ,
		_w5689_
	);
	LUT2 #(
		.INIT('h1)
	) name4731 (
		_w5688_,
		_w5689_,
		_w5690_
	);
	LUT2 #(
		.INIT('h1)
	) name4732 (
		_w5064_,
		_w5690_,
		_w5691_
	);
	LUT2 #(
		.INIT('h2)
	) name4733 (
		_w2269_,
		_w5691_,
		_w5692_
	);
	LUT2 #(
		.INIT('h4)
	) name4734 (
		_w5687_,
		_w5692_,
		_w5693_
	);
	LUT2 #(
		.INIT('h8)
	) name4735 (
		\u0_u0_tms_reg[0]/P0001 ,
		_w5077_,
		_w5694_
	);
	LUT2 #(
		.INIT('h8)
	) name4736 (
		\u0_u1_tms_reg[0]/P0001 ,
		_w5086_,
		_w5695_
	);
	LUT2 #(
		.INIT('h8)
	) name4737 (
		\u0_u0_csc_reg[0]/NET0131 ,
		_w5083_,
		_w5696_
	);
	LUT2 #(
		.INIT('h8)
	) name4738 (
		\u0_csc_mask_r_reg[0]/NET0131 ,
		_w5277_,
		_w5697_
	);
	LUT2 #(
		.INIT('h8)
	) name4739 (
		\u0_u1_csc_reg[0]/NET0131 ,
		_w5081_,
		_w5698_
	);
	LUT2 #(
		.INIT('h8)
	) name4740 (
		\u0_csr_r_reg[0]/P0001 ,
		_w5089_,
		_w5699_
	);
	LUT2 #(
		.INIT('h8)
	) name4741 (
		\poc_o[0]_pad ,
		_w5091_,
		_w5700_
	);
	LUT2 #(
		.INIT('h1)
	) name4742 (
		_w2269_,
		_w5695_,
		_w5701_
	);
	LUT2 #(
		.INIT('h1)
	) name4743 (
		_w5696_,
		_w5697_,
		_w5702_
	);
	LUT2 #(
		.INIT('h1)
	) name4744 (
		_w5698_,
		_w5699_,
		_w5703_
	);
	LUT2 #(
		.INIT('h8)
	) name4745 (
		_w5702_,
		_w5703_,
		_w5704_
	);
	LUT2 #(
		.INIT('h4)
	) name4746 (
		_w5694_,
		_w5701_,
		_w5705_
	);
	LUT2 #(
		.INIT('h4)
	) name4747 (
		_w5700_,
		_w5705_,
		_w5706_
	);
	LUT2 #(
		.INIT('h8)
	) name4748 (
		_w5704_,
		_w5706_,
		_w5707_
	);
	LUT2 #(
		.INIT('h1)
	) name4749 (
		_w5693_,
		_w5707_,
		_w5708_
	);
	LUT2 #(
		.INIT('h4)
	) name4750 (
		_w1984_,
		_w5064_,
		_w5709_
	);
	LUT2 #(
		.INIT('h4)
	) name4751 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[2]/P0001 ,
		_w5710_
	);
	LUT2 #(
		.INIT('h8)
	) name4752 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[10]/P0001 ,
		_w5711_
	);
	LUT2 #(
		.INIT('h1)
	) name4753 (
		_w5710_,
		_w5711_,
		_w5712_
	);
	LUT2 #(
		.INIT('h1)
	) name4754 (
		_w5064_,
		_w5712_,
		_w5713_
	);
	LUT2 #(
		.INIT('h2)
	) name4755 (
		_w2269_,
		_w5713_,
		_w5714_
	);
	LUT2 #(
		.INIT('h4)
	) name4756 (
		_w5709_,
		_w5714_,
		_w5715_
	);
	LUT2 #(
		.INIT('h8)
	) name4757 (
		\u0_u0_tms_reg[10]/P0001 ,
		_w5077_,
		_w5716_
	);
	LUT2 #(
		.INIT('h8)
	) name4758 (
		\u0_u1_tms_reg[10]/P0001 ,
		_w5086_,
		_w5717_
	);
	LUT2 #(
		.INIT('h8)
	) name4759 (
		\u0_u0_csc_reg[10]/P0001 ,
		_w5083_,
		_w5718_
	);
	LUT2 #(
		.INIT('h8)
	) name4760 (
		\u0_csr_r_reg[10]/NET0131 ,
		_w5089_,
		_w5719_
	);
	LUT2 #(
		.INIT('h8)
	) name4761 (
		\u0_u1_csc_reg[10]/P0001 ,
		_w5081_,
		_w5720_
	);
	LUT2 #(
		.INIT('h8)
	) name4762 (
		\u0_csc_mask_r_reg[10]/NET0131 ,
		_w5277_,
		_w5721_
	);
	LUT2 #(
		.INIT('h8)
	) name4763 (
		\poc_o[10]_pad ,
		_w5091_,
		_w5722_
	);
	LUT2 #(
		.INIT('h1)
	) name4764 (
		_w2269_,
		_w5717_,
		_w5723_
	);
	LUT2 #(
		.INIT('h1)
	) name4765 (
		_w5718_,
		_w5719_,
		_w5724_
	);
	LUT2 #(
		.INIT('h1)
	) name4766 (
		_w5720_,
		_w5721_,
		_w5725_
	);
	LUT2 #(
		.INIT('h8)
	) name4767 (
		_w5724_,
		_w5725_,
		_w5726_
	);
	LUT2 #(
		.INIT('h4)
	) name4768 (
		_w5716_,
		_w5723_,
		_w5727_
	);
	LUT2 #(
		.INIT('h4)
	) name4769 (
		_w5722_,
		_w5727_,
		_w5728_
	);
	LUT2 #(
		.INIT('h8)
	) name4770 (
		_w5726_,
		_w5728_,
		_w5729_
	);
	LUT2 #(
		.INIT('h1)
	) name4771 (
		_w5715_,
		_w5729_,
		_w5730_
	);
	LUT2 #(
		.INIT('h4)
	) name4772 (
		_w2184_,
		_w5064_,
		_w5731_
	);
	LUT2 #(
		.INIT('h4)
	) name4773 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[2]/P0001 ,
		_w5732_
	);
	LUT2 #(
		.INIT('h8)
	) name4774 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[2]/P0001 ,
		_w5733_
	);
	LUT2 #(
		.INIT('h1)
	) name4775 (
		_w5732_,
		_w5733_,
		_w5734_
	);
	LUT2 #(
		.INIT('h1)
	) name4776 (
		_w5064_,
		_w5734_,
		_w5735_
	);
	LUT2 #(
		.INIT('h2)
	) name4777 (
		_w2269_,
		_w5735_,
		_w5736_
	);
	LUT2 #(
		.INIT('h4)
	) name4778 (
		_w5731_,
		_w5736_,
		_w5737_
	);
	LUT2 #(
		.INIT('h8)
	) name4779 (
		\u0_u0_tms_reg[2]/P0001 ,
		_w5077_,
		_w5738_
	);
	LUT2 #(
		.INIT('h8)
	) name4780 (
		\u0_u1_csc_reg[2]/NET0131 ,
		_w5081_,
		_w5739_
	);
	LUT2 #(
		.INIT('h8)
	) name4781 (
		\u0_csr_r_reg[2]/NET0131 ,
		_w5089_,
		_w5740_
	);
	LUT2 #(
		.INIT('h8)
	) name4782 (
		\u0_u0_csc_reg[2]/NET0131 ,
		_w5083_,
		_w5741_
	);
	LUT2 #(
		.INIT('h8)
	) name4783 (
		\u0_u1_tms_reg[2]/P0001 ,
		_w5086_,
		_w5742_
	);
	LUT2 #(
		.INIT('h8)
	) name4784 (
		\u0_csc_mask_r_reg[2]/NET0131 ,
		_w5277_,
		_w5743_
	);
	LUT2 #(
		.INIT('h8)
	) name4785 (
		\poc_o[2]_pad ,
		_w5091_,
		_w5744_
	);
	LUT2 #(
		.INIT('h1)
	) name4786 (
		_w2269_,
		_w5739_,
		_w5745_
	);
	LUT2 #(
		.INIT('h1)
	) name4787 (
		_w5740_,
		_w5741_,
		_w5746_
	);
	LUT2 #(
		.INIT('h1)
	) name4788 (
		_w5742_,
		_w5743_,
		_w5747_
	);
	LUT2 #(
		.INIT('h8)
	) name4789 (
		_w5746_,
		_w5747_,
		_w5748_
	);
	LUT2 #(
		.INIT('h4)
	) name4790 (
		_w5738_,
		_w5745_,
		_w5749_
	);
	LUT2 #(
		.INIT('h4)
	) name4791 (
		_w5744_,
		_w5749_,
		_w5750_
	);
	LUT2 #(
		.INIT('h8)
	) name4792 (
		_w5748_,
		_w5750_,
		_w5751_
	);
	LUT2 #(
		.INIT('h1)
	) name4793 (
		_w5737_,
		_w5751_,
		_w5752_
	);
	LUT2 #(
		.INIT('h4)
	) name4794 (
		_w2201_,
		_w5064_,
		_w5753_
	);
	LUT2 #(
		.INIT('h4)
	) name4795 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[7]/P0001 ,
		_w5754_
	);
	LUT2 #(
		.INIT('h8)
	) name4796 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[7]/P0001 ,
		_w5755_
	);
	LUT2 #(
		.INIT('h1)
	) name4797 (
		_w5754_,
		_w5755_,
		_w5756_
	);
	LUT2 #(
		.INIT('h1)
	) name4798 (
		_w5064_,
		_w5756_,
		_w5757_
	);
	LUT2 #(
		.INIT('h2)
	) name4799 (
		_w2269_,
		_w5757_,
		_w5758_
	);
	LUT2 #(
		.INIT('h4)
	) name4800 (
		_w5753_,
		_w5758_,
		_w5759_
	);
	LUT2 #(
		.INIT('h8)
	) name4801 (
		\u0_u0_tms_reg[7]/P0001 ,
		_w5077_,
		_w5760_
	);
	LUT2 #(
		.INIT('h8)
	) name4802 (
		\u0_u1_tms_reg[7]/P0001 ,
		_w5086_,
		_w5761_
	);
	LUT2 #(
		.INIT('h8)
	) name4803 (
		\u0_u0_csc_reg[7]/P0001 ,
		_w5083_,
		_w5762_
	);
	LUT2 #(
		.INIT('h8)
	) name4804 (
		\u0_csc_mask_r_reg[7]/NET0131 ,
		_w5277_,
		_w5763_
	);
	LUT2 #(
		.INIT('h8)
	) name4805 (
		\u0_u1_csc_reg[7]/P0001 ,
		_w5081_,
		_w5764_
	);
	LUT2 #(
		.INIT('h8)
	) name4806 (
		\u0_csr_r_reg[7]/NET0131 ,
		_w5089_,
		_w5765_
	);
	LUT2 #(
		.INIT('h8)
	) name4807 (
		\poc_o[7]_pad ,
		_w5091_,
		_w5766_
	);
	LUT2 #(
		.INIT('h1)
	) name4808 (
		_w2269_,
		_w5761_,
		_w5767_
	);
	LUT2 #(
		.INIT('h1)
	) name4809 (
		_w5762_,
		_w5763_,
		_w5768_
	);
	LUT2 #(
		.INIT('h1)
	) name4810 (
		_w5764_,
		_w5765_,
		_w5769_
	);
	LUT2 #(
		.INIT('h8)
	) name4811 (
		_w5768_,
		_w5769_,
		_w5770_
	);
	LUT2 #(
		.INIT('h4)
	) name4812 (
		_w5760_,
		_w5767_,
		_w5771_
	);
	LUT2 #(
		.INIT('h4)
	) name4813 (
		_w5766_,
		_w5771_,
		_w5772_
	);
	LUT2 #(
		.INIT('h8)
	) name4814 (
		_w5770_,
		_w5772_,
		_w5773_
	);
	LUT2 #(
		.INIT('h1)
	) name4815 (
		_w5759_,
		_w5773_,
		_w5774_
	);
	LUT2 #(
		.INIT('h4)
	) name4816 (
		_w1960_,
		_w5064_,
		_w5775_
	);
	LUT2 #(
		.INIT('h4)
	) name4817 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[0]/P0001 ,
		_w5776_
	);
	LUT2 #(
		.INIT('h8)
	) name4818 (
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[8]/P0001 ,
		_w5777_
	);
	LUT2 #(
		.INIT('h1)
	) name4819 (
		_w5776_,
		_w5777_,
		_w5778_
	);
	LUT2 #(
		.INIT('h1)
	) name4820 (
		_w5064_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('h2)
	) name4821 (
		_w2269_,
		_w5779_,
		_w5780_
	);
	LUT2 #(
		.INIT('h4)
	) name4822 (
		_w5775_,
		_w5780_,
		_w5781_
	);
	LUT2 #(
		.INIT('h8)
	) name4823 (
		\u0_u0_tms_reg[8]/P0001 ,
		_w5077_,
		_w5782_
	);
	LUT2 #(
		.INIT('h8)
	) name4824 (
		\u0_u1_tms_reg[8]/P0001 ,
		_w5086_,
		_w5783_
	);
	LUT2 #(
		.INIT('h8)
	) name4825 (
		\u0_u0_csc_reg[8]/P0001 ,
		_w5083_,
		_w5784_
	);
	LUT2 #(
		.INIT('h8)
	) name4826 (
		\u0_csr_r_reg[8]/NET0131 ,
		_w5089_,
		_w5785_
	);
	LUT2 #(
		.INIT('h8)
	) name4827 (
		\u0_u1_csc_reg[8]/P0001 ,
		_w5081_,
		_w5786_
	);
	LUT2 #(
		.INIT('h8)
	) name4828 (
		\u0_csc_mask_r_reg[8]/NET0131 ,
		_w5277_,
		_w5787_
	);
	LUT2 #(
		.INIT('h8)
	) name4829 (
		\poc_o[8]_pad ,
		_w5091_,
		_w5788_
	);
	LUT2 #(
		.INIT('h1)
	) name4830 (
		_w2269_,
		_w5783_,
		_w5789_
	);
	LUT2 #(
		.INIT('h1)
	) name4831 (
		_w5784_,
		_w5785_,
		_w5790_
	);
	LUT2 #(
		.INIT('h1)
	) name4832 (
		_w5786_,
		_w5787_,
		_w5791_
	);
	LUT2 #(
		.INIT('h8)
	) name4833 (
		_w5790_,
		_w5791_,
		_w5792_
	);
	LUT2 #(
		.INIT('h4)
	) name4834 (
		_w5782_,
		_w5789_,
		_w5793_
	);
	LUT2 #(
		.INIT('h4)
	) name4835 (
		_w5788_,
		_w5793_,
		_w5794_
	);
	LUT2 #(
		.INIT('h8)
	) name4836 (
		_w5792_,
		_w5794_,
		_w5795_
	);
	LUT2 #(
		.INIT('h1)
	) name4837 (
		_w5781_,
		_w5795_,
		_w5796_
	);
	LUT2 #(
		.INIT('h2)
	) name4838 (
		\u0_u0_csc_reg[5]/P0001 ,
		_w5057_,
		_w5797_
	);
	LUT2 #(
		.INIT('h8)
	) name4839 (
		\wb_data_i[5]_pad ,
		_w5057_,
		_w5798_
	);
	LUT2 #(
		.INIT('h1)
	) name4840 (
		_w5797_,
		_w5798_,
		_w5799_
	);
	LUT2 #(
		.INIT('h1)
	) name4841 (
		\u0_rst_r2_reg/NET0131 ,
		_w5799_,
		_w5800_
	);
	LUT2 #(
		.INIT('h8)
	) name4842 (
		\poc_o[1]_pad ,
		\u0_rst_r2_reg/NET0131 ,
		_w5801_
	);
	LUT2 #(
		.INIT('h1)
	) name4843 (
		_w5800_,
		_w5801_,
		_w5802_
	);
	LUT2 #(
		.INIT('h2)
	) name4844 (
		\u0_u0_csc_reg[4]/P0001 ,
		_w5057_,
		_w5803_
	);
	LUT2 #(
		.INIT('h8)
	) name4845 (
		\wb_data_i[4]_pad ,
		_w5057_,
		_w5804_
	);
	LUT2 #(
		.INIT('h1)
	) name4846 (
		_w5803_,
		_w5804_,
		_w5805_
	);
	LUT2 #(
		.INIT('h1)
	) name4847 (
		\u0_rst_r2_reg/NET0131 ,
		_w5805_,
		_w5806_
	);
	LUT2 #(
		.INIT('h8)
	) name4848 (
		\poc_o[0]_pad ,
		\u0_rst_r2_reg/NET0131 ,
		_w5807_
	);
	LUT2 #(
		.INIT('h1)
	) name4849 (
		_w5806_,
		_w5807_,
		_w5808_
	);
	LUT2 #(
		.INIT('h8)
	) name4850 (
		\u5_state_reg[45]/NET0131 ,
		_w2388_,
		_w5809_
	);
	LUT2 #(
		.INIT('h1)
	) name4851 (
		\u0_u0_csc_reg[11]/P0001 ,
		_w5057_,
		_w5810_
	);
	LUT2 #(
		.INIT('h4)
	) name4852 (
		\wb_data_i[11]_pad ,
		_w5057_,
		_w5811_
	);
	LUT2 #(
		.INIT('h1)
	) name4853 (
		\u0_rst_r2_reg/NET0131 ,
		_w5810_,
		_w5812_
	);
	LUT2 #(
		.INIT('h4)
	) name4854 (
		_w5811_,
		_w5812_,
		_w5813_
	);
	LUT2 #(
		.INIT('h1)
	) name4855 (
		\u0_u0_csc_reg[12]/P0001 ,
		_w5057_,
		_w5814_
	);
	LUT2 #(
		.INIT('h4)
	) name4856 (
		\wb_data_i[12]_pad ,
		_w5057_,
		_w5815_
	);
	LUT2 #(
		.INIT('h1)
	) name4857 (
		\u0_rst_r2_reg/NET0131 ,
		_w5814_,
		_w5816_
	);
	LUT2 #(
		.INIT('h4)
	) name4858 (
		_w5815_,
		_w5816_,
		_w5817_
	);
	LUT2 #(
		.INIT('h8)
	) name4859 (
		\u0_u0_addr_r_reg[3]/P0001 ,
		_w5054_,
		_w5818_
	);
	LUT2 #(
		.INIT('h8)
	) name4860 (
		_w5053_,
		_w5818_,
		_w5819_
	);
	LUT2 #(
		.INIT('h8)
	) name4861 (
		\u0_u0_addr_r_reg[2]/P0001 ,
		_w5819_,
		_w5820_
	);
	LUT2 #(
		.INIT('h1)
	) name4862 (
		\u0_u1_tms_reg[19]/P0001 ,
		_w5820_,
		_w5821_
	);
	LUT2 #(
		.INIT('h4)
	) name4863 (
		\wb_data_i[19]_pad ,
		_w5820_,
		_w5822_
	);
	LUT2 #(
		.INIT('h1)
	) name4864 (
		\u0_rst_r2_reg/NET0131 ,
		_w5821_,
		_w5823_
	);
	LUT2 #(
		.INIT('h4)
	) name4865 (
		_w5822_,
		_w5823_,
		_w5824_
	);
	LUT2 #(
		.INIT('h1)
	) name4866 (
		\u0_u0_csc_reg[13]/P0001 ,
		_w5057_,
		_w5825_
	);
	LUT2 #(
		.INIT('h4)
	) name4867 (
		\wb_data_i[13]_pad ,
		_w5057_,
		_w5826_
	);
	LUT2 #(
		.INIT('h1)
	) name4868 (
		\u0_rst_r2_reg/NET0131 ,
		_w5825_,
		_w5827_
	);
	LUT2 #(
		.INIT('h4)
	) name4869 (
		_w5826_,
		_w5827_,
		_w5828_
	);
	LUT2 #(
		.INIT('h1)
	) name4870 (
		\u0_u0_csc_reg[14]/P0001 ,
		_w5057_,
		_w5829_
	);
	LUT2 #(
		.INIT('h4)
	) name4871 (
		\wb_data_i[14]_pad ,
		_w5057_,
		_w5830_
	);
	LUT2 #(
		.INIT('h1)
	) name4872 (
		\u0_rst_r2_reg/NET0131 ,
		_w5829_,
		_w5831_
	);
	LUT2 #(
		.INIT('h4)
	) name4873 (
		_w5830_,
		_w5831_,
		_w5832_
	);
	LUT2 #(
		.INIT('h1)
	) name4874 (
		\u0_u0_csc_reg[16]/P0001 ,
		_w5057_,
		_w5833_
	);
	LUT2 #(
		.INIT('h4)
	) name4875 (
		\wb_data_i[16]_pad ,
		_w5057_,
		_w5834_
	);
	LUT2 #(
		.INIT('h1)
	) name4876 (
		\u0_rst_r2_reg/NET0131 ,
		_w5833_,
		_w5835_
	);
	LUT2 #(
		.INIT('h4)
	) name4877 (
		_w5834_,
		_w5835_,
		_w5836_
	);
	LUT2 #(
		.INIT('h1)
	) name4878 (
		\u0_u0_csc_reg[17]/P0001 ,
		_w5057_,
		_w5837_
	);
	LUT2 #(
		.INIT('h4)
	) name4879 (
		\wb_data_i[17]_pad ,
		_w5057_,
		_w5838_
	);
	LUT2 #(
		.INIT('h1)
	) name4880 (
		\u0_rst_r2_reg/NET0131 ,
		_w5837_,
		_w5839_
	);
	LUT2 #(
		.INIT('h4)
	) name4881 (
		_w5838_,
		_w5839_,
		_w5840_
	);
	LUT2 #(
		.INIT('h1)
	) name4882 (
		\u0_u0_csc_reg[20]/P0001 ,
		_w5057_,
		_w5841_
	);
	LUT2 #(
		.INIT('h4)
	) name4883 (
		\wb_data_i[20]_pad ,
		_w5057_,
		_w5842_
	);
	LUT2 #(
		.INIT('h1)
	) name4884 (
		\u0_rst_r2_reg/NET0131 ,
		_w5841_,
		_w5843_
	);
	LUT2 #(
		.INIT('h4)
	) name4885 (
		_w5842_,
		_w5843_,
		_w5844_
	);
	LUT2 #(
		.INIT('h1)
	) name4886 (
		\u0_u0_csc_reg[21]/P0001 ,
		_w5057_,
		_w5845_
	);
	LUT2 #(
		.INIT('h4)
	) name4887 (
		\wb_data_i[21]_pad ,
		_w5057_,
		_w5846_
	);
	LUT2 #(
		.INIT('h1)
	) name4888 (
		\u0_rst_r2_reg/NET0131 ,
		_w5845_,
		_w5847_
	);
	LUT2 #(
		.INIT('h4)
	) name4889 (
		_w5846_,
		_w5847_,
		_w5848_
	);
	LUT2 #(
		.INIT('h1)
	) name4890 (
		\u0_u0_csc_reg[22]/P0001 ,
		_w5057_,
		_w5849_
	);
	LUT2 #(
		.INIT('h4)
	) name4891 (
		\wb_data_i[22]_pad ,
		_w5057_,
		_w5850_
	);
	LUT2 #(
		.INIT('h1)
	) name4892 (
		\u0_rst_r2_reg/NET0131 ,
		_w5849_,
		_w5851_
	);
	LUT2 #(
		.INIT('h4)
	) name4893 (
		_w5850_,
		_w5851_,
		_w5852_
	);
	LUT2 #(
		.INIT('h1)
	) name4894 (
		\u0_u0_csc_reg[24]/P0001 ,
		_w5057_,
		_w5853_
	);
	LUT2 #(
		.INIT('h4)
	) name4895 (
		\wb_data_i[24]_pad ,
		_w5057_,
		_w5854_
	);
	LUT2 #(
		.INIT('h1)
	) name4896 (
		\u0_rst_r2_reg/NET0131 ,
		_w5853_,
		_w5855_
	);
	LUT2 #(
		.INIT('h4)
	) name4897 (
		_w5854_,
		_w5855_,
		_w5856_
	);
	LUT2 #(
		.INIT('h1)
	) name4898 (
		\u0_u0_csc_reg[26]/P0001 ,
		_w5057_,
		_w5857_
	);
	LUT2 #(
		.INIT('h4)
	) name4899 (
		\wb_data_i[26]_pad ,
		_w5057_,
		_w5858_
	);
	LUT2 #(
		.INIT('h1)
	) name4900 (
		\u0_rst_r2_reg/NET0131 ,
		_w5857_,
		_w5859_
	);
	LUT2 #(
		.INIT('h4)
	) name4901 (
		_w5858_,
		_w5859_,
		_w5860_
	);
	LUT2 #(
		.INIT('h1)
	) name4902 (
		\u0_u0_csc_reg[27]/P0001 ,
		_w5057_,
		_w5861_
	);
	LUT2 #(
		.INIT('h4)
	) name4903 (
		\wb_data_i[27]_pad ,
		_w5057_,
		_w5862_
	);
	LUT2 #(
		.INIT('h1)
	) name4904 (
		\u0_rst_r2_reg/NET0131 ,
		_w5861_,
		_w5863_
	);
	LUT2 #(
		.INIT('h4)
	) name4905 (
		_w5862_,
		_w5863_,
		_w5864_
	);
	LUT2 #(
		.INIT('h1)
	) name4906 (
		\u0_u0_csc_reg[28]/P0001 ,
		_w5057_,
		_w5865_
	);
	LUT2 #(
		.INIT('h4)
	) name4907 (
		\wb_data_i[28]_pad ,
		_w5057_,
		_w5866_
	);
	LUT2 #(
		.INIT('h1)
	) name4908 (
		\u0_rst_r2_reg/NET0131 ,
		_w5865_,
		_w5867_
	);
	LUT2 #(
		.INIT('h4)
	) name4909 (
		_w5866_,
		_w5867_,
		_w5868_
	);
	LUT2 #(
		.INIT('h1)
	) name4910 (
		\u0_u1_tms_reg[23]/P0001 ,
		_w5820_,
		_w5869_
	);
	LUT2 #(
		.INIT('h4)
	) name4911 (
		\wb_data_i[23]_pad ,
		_w5820_,
		_w5870_
	);
	LUT2 #(
		.INIT('h1)
	) name4912 (
		\u0_rst_r2_reg/NET0131 ,
		_w5869_,
		_w5871_
	);
	LUT2 #(
		.INIT('h4)
	) name4913 (
		_w5870_,
		_w5871_,
		_w5872_
	);
	LUT2 #(
		.INIT('h1)
	) name4914 (
		\u0_u0_csc_reg[30]/P0001 ,
		_w5057_,
		_w5873_
	);
	LUT2 #(
		.INIT('h4)
	) name4915 (
		\wb_data_i[30]_pad ,
		_w5057_,
		_w5874_
	);
	LUT2 #(
		.INIT('h1)
	) name4916 (
		\u0_rst_r2_reg/NET0131 ,
		_w5873_,
		_w5875_
	);
	LUT2 #(
		.INIT('h4)
	) name4917 (
		_w5874_,
		_w5875_,
		_w5876_
	);
	LUT2 #(
		.INIT('h1)
	) name4918 (
		\u0_u0_csc_reg[3]/NET0131 ,
		_w5057_,
		_w5877_
	);
	LUT2 #(
		.INIT('h4)
	) name4919 (
		\wb_data_i[3]_pad ,
		_w5057_,
		_w5878_
	);
	LUT2 #(
		.INIT('h1)
	) name4920 (
		\u0_rst_r2_reg/NET0131 ,
		_w5877_,
		_w5879_
	);
	LUT2 #(
		.INIT('h4)
	) name4921 (
		_w5878_,
		_w5879_,
		_w5880_
	);
	LUT2 #(
		.INIT('h1)
	) name4922 (
		\u0_u0_csc_reg[25]/P0001 ,
		_w5057_,
		_w5881_
	);
	LUT2 #(
		.INIT('h4)
	) name4923 (
		\wb_data_i[25]_pad ,
		_w5057_,
		_w5882_
	);
	LUT2 #(
		.INIT('h1)
	) name4924 (
		\u0_rst_r2_reg/NET0131 ,
		_w5881_,
		_w5883_
	);
	LUT2 #(
		.INIT('h4)
	) name4925 (
		_w5882_,
		_w5883_,
		_w5884_
	);
	LUT2 #(
		.INIT('h1)
	) name4926 (
		\u0_u1_tms_reg[17]/P0001 ,
		_w5820_,
		_w5885_
	);
	LUT2 #(
		.INIT('h4)
	) name4927 (
		\wb_data_i[17]_pad ,
		_w5820_,
		_w5886_
	);
	LUT2 #(
		.INIT('h1)
	) name4928 (
		\u0_rst_r2_reg/NET0131 ,
		_w5885_,
		_w5887_
	);
	LUT2 #(
		.INIT('h4)
	) name4929 (
		_w5886_,
		_w5887_,
		_w5888_
	);
	LUT2 #(
		.INIT('h1)
	) name4930 (
		\u0_u1_tms_reg[16]/P0001 ,
		_w5820_,
		_w5889_
	);
	LUT2 #(
		.INIT('h4)
	) name4931 (
		\wb_data_i[16]_pad ,
		_w5820_,
		_w5890_
	);
	LUT2 #(
		.INIT('h1)
	) name4932 (
		\u0_rst_r2_reg/NET0131 ,
		_w5889_,
		_w5891_
	);
	LUT2 #(
		.INIT('h4)
	) name4933 (
		_w5890_,
		_w5891_,
		_w5892_
	);
	LUT2 #(
		.INIT('h8)
	) name4934 (
		\u0_u0_addr_r_reg[2]/P0001 ,
		_w5056_,
		_w5893_
	);
	LUT2 #(
		.INIT('h8)
	) name4935 (
		\wb_data_i[0]_pad ,
		_w5893_,
		_w5894_
	);
	LUT2 #(
		.INIT('h2)
	) name4936 (
		\u0_u0_tms_reg[0]/P0001 ,
		_w5893_,
		_w5895_
	);
	LUT2 #(
		.INIT('h1)
	) name4937 (
		\u0_rst_r2_reg/NET0131 ,
		_w5894_,
		_w5896_
	);
	LUT2 #(
		.INIT('h4)
	) name4938 (
		_w5895_,
		_w5896_,
		_w5897_
	);
	LUT2 #(
		.INIT('h8)
	) name4939 (
		\wb_data_i[10]_pad ,
		_w5893_,
		_w5898_
	);
	LUT2 #(
		.INIT('h2)
	) name4940 (
		\u0_u0_tms_reg[10]/P0001 ,
		_w5893_,
		_w5899_
	);
	LUT2 #(
		.INIT('h1)
	) name4941 (
		\u0_rst_r2_reg/NET0131 ,
		_w5898_,
		_w5900_
	);
	LUT2 #(
		.INIT('h4)
	) name4942 (
		_w5899_,
		_w5900_,
		_w5901_
	);
	LUT2 #(
		.INIT('h8)
	) name4943 (
		\wb_data_i[11]_pad ,
		_w5893_,
		_w5902_
	);
	LUT2 #(
		.INIT('h2)
	) name4944 (
		\u0_u0_tms_reg[11]/P0001 ,
		_w5893_,
		_w5903_
	);
	LUT2 #(
		.INIT('h1)
	) name4945 (
		\u0_rst_r2_reg/NET0131 ,
		_w5902_,
		_w5904_
	);
	LUT2 #(
		.INIT('h4)
	) name4946 (
		_w5903_,
		_w5904_,
		_w5905_
	);
	LUT2 #(
		.INIT('h8)
	) name4947 (
		\wb_data_i[12]_pad ,
		_w5893_,
		_w5906_
	);
	LUT2 #(
		.INIT('h2)
	) name4948 (
		\u0_u0_tms_reg[12]/P0001 ,
		_w5893_,
		_w5907_
	);
	LUT2 #(
		.INIT('h1)
	) name4949 (
		\u0_rst_r2_reg/NET0131 ,
		_w5906_,
		_w5908_
	);
	LUT2 #(
		.INIT('h4)
	) name4950 (
		_w5907_,
		_w5908_,
		_w5909_
	);
	LUT2 #(
		.INIT('h8)
	) name4951 (
		\wb_data_i[14]_pad ,
		_w5893_,
		_w5910_
	);
	LUT2 #(
		.INIT('h2)
	) name4952 (
		\u0_u0_tms_reg[14]/P0001 ,
		_w5893_,
		_w5911_
	);
	LUT2 #(
		.INIT('h1)
	) name4953 (
		\u0_rst_r2_reg/NET0131 ,
		_w5910_,
		_w5912_
	);
	LUT2 #(
		.INIT('h4)
	) name4954 (
		_w5911_,
		_w5912_,
		_w5913_
	);
	LUT2 #(
		.INIT('h8)
	) name4955 (
		\wb_data_i[13]_pad ,
		_w5893_,
		_w5914_
	);
	LUT2 #(
		.INIT('h2)
	) name4956 (
		\u0_u0_tms_reg[13]/P0001 ,
		_w5893_,
		_w5915_
	);
	LUT2 #(
		.INIT('h1)
	) name4957 (
		\u0_rst_r2_reg/NET0131 ,
		_w5914_,
		_w5916_
	);
	LUT2 #(
		.INIT('h4)
	) name4958 (
		_w5915_,
		_w5916_,
		_w5917_
	);
	LUT2 #(
		.INIT('h8)
	) name4959 (
		\wb_data_i[15]_pad ,
		_w5893_,
		_w5918_
	);
	LUT2 #(
		.INIT('h2)
	) name4960 (
		\u0_u0_tms_reg[15]/P0001 ,
		_w5893_,
		_w5919_
	);
	LUT2 #(
		.INIT('h1)
	) name4961 (
		\u0_rst_r2_reg/NET0131 ,
		_w5918_,
		_w5920_
	);
	LUT2 #(
		.INIT('h4)
	) name4962 (
		_w5919_,
		_w5920_,
		_w5921_
	);
	LUT2 #(
		.INIT('h8)
	) name4963 (
		\wb_data_i[16]_pad ,
		_w5893_,
		_w5922_
	);
	LUT2 #(
		.INIT('h2)
	) name4964 (
		\u0_u0_tms_reg[16]/P0001 ,
		_w5893_,
		_w5923_
	);
	LUT2 #(
		.INIT('h1)
	) name4965 (
		\u0_rst_r2_reg/NET0131 ,
		_w5922_,
		_w5924_
	);
	LUT2 #(
		.INIT('h4)
	) name4966 (
		_w5923_,
		_w5924_,
		_w5925_
	);
	LUT2 #(
		.INIT('h8)
	) name4967 (
		\wb_data_i[17]_pad ,
		_w5893_,
		_w5926_
	);
	LUT2 #(
		.INIT('h2)
	) name4968 (
		\u0_u0_tms_reg[17]/P0001 ,
		_w5893_,
		_w5927_
	);
	LUT2 #(
		.INIT('h1)
	) name4969 (
		\u0_rst_r2_reg/NET0131 ,
		_w5926_,
		_w5928_
	);
	LUT2 #(
		.INIT('h4)
	) name4970 (
		_w5927_,
		_w5928_,
		_w5929_
	);
	LUT2 #(
		.INIT('h8)
	) name4971 (
		\wb_data_i[18]_pad ,
		_w5893_,
		_w5930_
	);
	LUT2 #(
		.INIT('h2)
	) name4972 (
		\u0_u0_tms_reg[18]/P0001 ,
		_w5893_,
		_w5931_
	);
	LUT2 #(
		.INIT('h1)
	) name4973 (
		\u0_rst_r2_reg/NET0131 ,
		_w5930_,
		_w5932_
	);
	LUT2 #(
		.INIT('h4)
	) name4974 (
		_w5931_,
		_w5932_,
		_w5933_
	);
	LUT2 #(
		.INIT('h8)
	) name4975 (
		\wb_data_i[19]_pad ,
		_w5893_,
		_w5934_
	);
	LUT2 #(
		.INIT('h2)
	) name4976 (
		\u0_u0_tms_reg[19]/P0001 ,
		_w5893_,
		_w5935_
	);
	LUT2 #(
		.INIT('h1)
	) name4977 (
		\u0_rst_r2_reg/NET0131 ,
		_w5934_,
		_w5936_
	);
	LUT2 #(
		.INIT('h4)
	) name4978 (
		_w5935_,
		_w5936_,
		_w5937_
	);
	LUT2 #(
		.INIT('h8)
	) name4979 (
		\wb_data_i[1]_pad ,
		_w5893_,
		_w5938_
	);
	LUT2 #(
		.INIT('h2)
	) name4980 (
		\u0_u0_tms_reg[1]/P0001 ,
		_w5893_,
		_w5939_
	);
	LUT2 #(
		.INIT('h1)
	) name4981 (
		\u0_rst_r2_reg/NET0131 ,
		_w5938_,
		_w5940_
	);
	LUT2 #(
		.INIT('h4)
	) name4982 (
		_w5939_,
		_w5940_,
		_w5941_
	);
	LUT2 #(
		.INIT('h8)
	) name4983 (
		\wb_data_i[21]_pad ,
		_w5893_,
		_w5942_
	);
	LUT2 #(
		.INIT('h2)
	) name4984 (
		\u0_u0_tms_reg[21]/P0001 ,
		_w5893_,
		_w5943_
	);
	LUT2 #(
		.INIT('h1)
	) name4985 (
		\u0_rst_r2_reg/NET0131 ,
		_w5942_,
		_w5944_
	);
	LUT2 #(
		.INIT('h4)
	) name4986 (
		_w5943_,
		_w5944_,
		_w5945_
	);
	LUT2 #(
		.INIT('h8)
	) name4987 (
		\wb_data_i[22]_pad ,
		_w5893_,
		_w5946_
	);
	LUT2 #(
		.INIT('h2)
	) name4988 (
		\u0_u0_tms_reg[22]/P0001 ,
		_w5893_,
		_w5947_
	);
	LUT2 #(
		.INIT('h1)
	) name4989 (
		\u0_rst_r2_reg/NET0131 ,
		_w5946_,
		_w5948_
	);
	LUT2 #(
		.INIT('h4)
	) name4990 (
		_w5947_,
		_w5948_,
		_w5949_
	);
	LUT2 #(
		.INIT('h8)
	) name4991 (
		\wb_data_i[23]_pad ,
		_w5893_,
		_w5950_
	);
	LUT2 #(
		.INIT('h2)
	) name4992 (
		\u0_u0_tms_reg[23]/P0001 ,
		_w5893_,
		_w5951_
	);
	LUT2 #(
		.INIT('h1)
	) name4993 (
		\u0_rst_r2_reg/NET0131 ,
		_w5950_,
		_w5952_
	);
	LUT2 #(
		.INIT('h4)
	) name4994 (
		_w5951_,
		_w5952_,
		_w5953_
	);
	LUT2 #(
		.INIT('h8)
	) name4995 (
		\wb_data_i[24]_pad ,
		_w5893_,
		_w5954_
	);
	LUT2 #(
		.INIT('h2)
	) name4996 (
		\u0_u0_tms_reg[24]/P0001 ,
		_w5893_,
		_w5955_
	);
	LUT2 #(
		.INIT('h1)
	) name4997 (
		\u0_rst_r2_reg/NET0131 ,
		_w5954_,
		_w5956_
	);
	LUT2 #(
		.INIT('h4)
	) name4998 (
		_w5955_,
		_w5956_,
		_w5957_
	);
	LUT2 #(
		.INIT('h8)
	) name4999 (
		\wb_data_i[25]_pad ,
		_w5893_,
		_w5958_
	);
	LUT2 #(
		.INIT('h2)
	) name5000 (
		\u0_u0_tms_reg[25]/P0001 ,
		_w5893_,
		_w5959_
	);
	LUT2 #(
		.INIT('h1)
	) name5001 (
		\u0_rst_r2_reg/NET0131 ,
		_w5958_,
		_w5960_
	);
	LUT2 #(
		.INIT('h4)
	) name5002 (
		_w5959_,
		_w5960_,
		_w5961_
	);
	LUT2 #(
		.INIT('h8)
	) name5003 (
		\wb_data_i[26]_pad ,
		_w5893_,
		_w5962_
	);
	LUT2 #(
		.INIT('h2)
	) name5004 (
		\u0_u0_tms_reg[26]/P0001 ,
		_w5893_,
		_w5963_
	);
	LUT2 #(
		.INIT('h1)
	) name5005 (
		\u0_rst_r2_reg/NET0131 ,
		_w5962_,
		_w5964_
	);
	LUT2 #(
		.INIT('h4)
	) name5006 (
		_w5963_,
		_w5964_,
		_w5965_
	);
	LUT2 #(
		.INIT('h8)
	) name5007 (
		\wb_data_i[27]_pad ,
		_w5893_,
		_w5966_
	);
	LUT2 #(
		.INIT('h2)
	) name5008 (
		\u0_u0_tms_reg[27]/P0001 ,
		_w5893_,
		_w5967_
	);
	LUT2 #(
		.INIT('h1)
	) name5009 (
		\u0_rst_r2_reg/NET0131 ,
		_w5966_,
		_w5968_
	);
	LUT2 #(
		.INIT('h4)
	) name5010 (
		_w5967_,
		_w5968_,
		_w5969_
	);
	LUT2 #(
		.INIT('h1)
	) name5011 (
		\u0_u1_tms_reg[22]/P0001 ,
		_w5820_,
		_w5970_
	);
	LUT2 #(
		.INIT('h4)
	) name5012 (
		\wb_data_i[22]_pad ,
		_w5820_,
		_w5971_
	);
	LUT2 #(
		.INIT('h1)
	) name5013 (
		\u0_rst_r2_reg/NET0131 ,
		_w5970_,
		_w5972_
	);
	LUT2 #(
		.INIT('h4)
	) name5014 (
		_w5971_,
		_w5972_,
		_w5973_
	);
	LUT2 #(
		.INIT('h8)
	) name5015 (
		\wb_data_i[28]_pad ,
		_w5893_,
		_w5974_
	);
	LUT2 #(
		.INIT('h2)
	) name5016 (
		\u0_u0_tms_reg[28]/P0001 ,
		_w5893_,
		_w5975_
	);
	LUT2 #(
		.INIT('h1)
	) name5017 (
		\u0_rst_r2_reg/NET0131 ,
		_w5974_,
		_w5976_
	);
	LUT2 #(
		.INIT('h4)
	) name5018 (
		_w5975_,
		_w5976_,
		_w5977_
	);
	LUT2 #(
		.INIT('h8)
	) name5019 (
		\wb_data_i[29]_pad ,
		_w5893_,
		_w5978_
	);
	LUT2 #(
		.INIT('h2)
	) name5020 (
		\u0_u0_tms_reg[29]/P0001 ,
		_w5893_,
		_w5979_
	);
	LUT2 #(
		.INIT('h1)
	) name5021 (
		\u0_rst_r2_reg/NET0131 ,
		_w5978_,
		_w5980_
	);
	LUT2 #(
		.INIT('h4)
	) name5022 (
		_w5979_,
		_w5980_,
		_w5981_
	);
	LUT2 #(
		.INIT('h8)
	) name5023 (
		\wb_data_i[2]_pad ,
		_w5893_,
		_w5982_
	);
	LUT2 #(
		.INIT('h2)
	) name5024 (
		\u0_u0_tms_reg[2]/P0001 ,
		_w5893_,
		_w5983_
	);
	LUT2 #(
		.INIT('h1)
	) name5025 (
		\u0_rst_r2_reg/NET0131 ,
		_w5982_,
		_w5984_
	);
	LUT2 #(
		.INIT('h4)
	) name5026 (
		_w5983_,
		_w5984_,
		_w5985_
	);
	LUT2 #(
		.INIT('h1)
	) name5027 (
		\u0_u0_csc_reg[15]/P0001 ,
		_w5057_,
		_w5986_
	);
	LUT2 #(
		.INIT('h4)
	) name5028 (
		\wb_data_i[15]_pad ,
		_w5057_,
		_w5987_
	);
	LUT2 #(
		.INIT('h1)
	) name5029 (
		\u0_rst_r2_reg/NET0131 ,
		_w5986_,
		_w5988_
	);
	LUT2 #(
		.INIT('h4)
	) name5030 (
		_w5987_,
		_w5988_,
		_w5989_
	);
	LUT2 #(
		.INIT('h8)
	) name5031 (
		\wb_data_i[30]_pad ,
		_w5893_,
		_w5990_
	);
	LUT2 #(
		.INIT('h2)
	) name5032 (
		\u0_u0_tms_reg[30]/P0001 ,
		_w5893_,
		_w5991_
	);
	LUT2 #(
		.INIT('h1)
	) name5033 (
		\u0_rst_r2_reg/NET0131 ,
		_w5990_,
		_w5992_
	);
	LUT2 #(
		.INIT('h4)
	) name5034 (
		_w5991_,
		_w5992_,
		_w5993_
	);
	LUT2 #(
		.INIT('h8)
	) name5035 (
		\wb_data_i[3]_pad ,
		_w5893_,
		_w5994_
	);
	LUT2 #(
		.INIT('h2)
	) name5036 (
		\u0_u0_tms_reg[3]/P0001 ,
		_w5893_,
		_w5995_
	);
	LUT2 #(
		.INIT('h1)
	) name5037 (
		\u0_rst_r2_reg/NET0131 ,
		_w5994_,
		_w5996_
	);
	LUT2 #(
		.INIT('h4)
	) name5038 (
		_w5995_,
		_w5996_,
		_w5997_
	);
	LUT2 #(
		.INIT('h8)
	) name5039 (
		\wb_data_i[4]_pad ,
		_w5893_,
		_w5998_
	);
	LUT2 #(
		.INIT('h2)
	) name5040 (
		\u0_u0_tms_reg[4]/P0001 ,
		_w5893_,
		_w5999_
	);
	LUT2 #(
		.INIT('h1)
	) name5041 (
		\u0_rst_r2_reg/NET0131 ,
		_w5998_,
		_w6000_
	);
	LUT2 #(
		.INIT('h4)
	) name5042 (
		_w5999_,
		_w6000_,
		_w6001_
	);
	LUT2 #(
		.INIT('h8)
	) name5043 (
		\wb_data_i[5]_pad ,
		_w5893_,
		_w6002_
	);
	LUT2 #(
		.INIT('h2)
	) name5044 (
		\u0_u0_tms_reg[5]/P0001 ,
		_w5893_,
		_w6003_
	);
	LUT2 #(
		.INIT('h1)
	) name5045 (
		\u0_rst_r2_reg/NET0131 ,
		_w6002_,
		_w6004_
	);
	LUT2 #(
		.INIT('h4)
	) name5046 (
		_w6003_,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h8)
	) name5047 (
		\wb_data_i[6]_pad ,
		_w5893_,
		_w6006_
	);
	LUT2 #(
		.INIT('h2)
	) name5048 (
		\u0_u0_tms_reg[6]/P0001 ,
		_w5893_,
		_w6007_
	);
	LUT2 #(
		.INIT('h1)
	) name5049 (
		\u0_rst_r2_reg/NET0131 ,
		_w6006_,
		_w6008_
	);
	LUT2 #(
		.INIT('h4)
	) name5050 (
		_w6007_,
		_w6008_,
		_w6009_
	);
	LUT2 #(
		.INIT('h8)
	) name5051 (
		\wb_data_i[7]_pad ,
		_w5893_,
		_w6010_
	);
	LUT2 #(
		.INIT('h2)
	) name5052 (
		\u0_u0_tms_reg[7]/P0001 ,
		_w5893_,
		_w6011_
	);
	LUT2 #(
		.INIT('h1)
	) name5053 (
		\u0_rst_r2_reg/NET0131 ,
		_w6010_,
		_w6012_
	);
	LUT2 #(
		.INIT('h4)
	) name5054 (
		_w6011_,
		_w6012_,
		_w6013_
	);
	LUT2 #(
		.INIT('h8)
	) name5055 (
		\wb_data_i[8]_pad ,
		_w5893_,
		_w6014_
	);
	LUT2 #(
		.INIT('h2)
	) name5056 (
		\u0_u0_tms_reg[8]/P0001 ,
		_w5893_,
		_w6015_
	);
	LUT2 #(
		.INIT('h1)
	) name5057 (
		\u0_rst_r2_reg/NET0131 ,
		_w6014_,
		_w6016_
	);
	LUT2 #(
		.INIT('h4)
	) name5058 (
		_w6015_,
		_w6016_,
		_w6017_
	);
	LUT2 #(
		.INIT('h8)
	) name5059 (
		\wb_data_i[9]_pad ,
		_w5893_,
		_w6018_
	);
	LUT2 #(
		.INIT('h2)
	) name5060 (
		\u0_u0_tms_reg[9]/P0001 ,
		_w5893_,
		_w6019_
	);
	LUT2 #(
		.INIT('h1)
	) name5061 (
		\u0_rst_r2_reg/NET0131 ,
		_w6018_,
		_w6020_
	);
	LUT2 #(
		.INIT('h4)
	) name5062 (
		_w6019_,
		_w6020_,
		_w6021_
	);
	LUT2 #(
		.INIT('h4)
	) name5063 (
		\u0_u0_addr_r_reg[2]/P0001 ,
		_w5819_,
		_w6022_
	);
	LUT2 #(
		.INIT('h1)
	) name5064 (
		\u0_u1_csc_reg[0]/NET0131 ,
		_w6022_,
		_w6023_
	);
	LUT2 #(
		.INIT('h4)
	) name5065 (
		\wb_data_i[0]_pad ,
		_w6022_,
		_w6024_
	);
	LUT2 #(
		.INIT('h1)
	) name5066 (
		\u0_rst_r2_reg/NET0131 ,
		_w6023_,
		_w6025_
	);
	LUT2 #(
		.INIT('h4)
	) name5067 (
		_w6024_,
		_w6025_,
		_w6026_
	);
	LUT2 #(
		.INIT('h1)
	) name5068 (
		\u0_u1_csc_reg[10]/P0001 ,
		_w6022_,
		_w6027_
	);
	LUT2 #(
		.INIT('h4)
	) name5069 (
		\wb_data_i[10]_pad ,
		_w6022_,
		_w6028_
	);
	LUT2 #(
		.INIT('h1)
	) name5070 (
		\u0_rst_r2_reg/NET0131 ,
		_w6027_,
		_w6029_
	);
	LUT2 #(
		.INIT('h4)
	) name5071 (
		_w6028_,
		_w6029_,
		_w6030_
	);
	LUT2 #(
		.INIT('h1)
	) name5072 (
		\u0_u1_csc_reg[11]/P0001 ,
		_w6022_,
		_w6031_
	);
	LUT2 #(
		.INIT('h4)
	) name5073 (
		\wb_data_i[11]_pad ,
		_w6022_,
		_w6032_
	);
	LUT2 #(
		.INIT('h1)
	) name5074 (
		\u0_rst_r2_reg/NET0131 ,
		_w6031_,
		_w6033_
	);
	LUT2 #(
		.INIT('h4)
	) name5075 (
		_w6032_,
		_w6033_,
		_w6034_
	);
	LUT2 #(
		.INIT('h1)
	) name5076 (
		\u0_u1_csc_reg[12]/P0001 ,
		_w6022_,
		_w6035_
	);
	LUT2 #(
		.INIT('h4)
	) name5077 (
		\wb_data_i[12]_pad ,
		_w6022_,
		_w6036_
	);
	LUT2 #(
		.INIT('h1)
	) name5078 (
		\u0_rst_r2_reg/NET0131 ,
		_w6035_,
		_w6037_
	);
	LUT2 #(
		.INIT('h4)
	) name5079 (
		_w6036_,
		_w6037_,
		_w6038_
	);
	LUT2 #(
		.INIT('h1)
	) name5080 (
		\u0_u1_csc_reg[13]/P0001 ,
		_w6022_,
		_w6039_
	);
	LUT2 #(
		.INIT('h4)
	) name5081 (
		\wb_data_i[13]_pad ,
		_w6022_,
		_w6040_
	);
	LUT2 #(
		.INIT('h1)
	) name5082 (
		\u0_rst_r2_reg/NET0131 ,
		_w6039_,
		_w6041_
	);
	LUT2 #(
		.INIT('h4)
	) name5083 (
		_w6040_,
		_w6041_,
		_w6042_
	);
	LUT2 #(
		.INIT('h1)
	) name5084 (
		\u0_u1_csc_reg[14]/P0001 ,
		_w6022_,
		_w6043_
	);
	LUT2 #(
		.INIT('h4)
	) name5085 (
		\wb_data_i[14]_pad ,
		_w6022_,
		_w6044_
	);
	LUT2 #(
		.INIT('h1)
	) name5086 (
		\u0_rst_r2_reg/NET0131 ,
		_w6043_,
		_w6045_
	);
	LUT2 #(
		.INIT('h4)
	) name5087 (
		_w6044_,
		_w6045_,
		_w6046_
	);
	LUT2 #(
		.INIT('h1)
	) name5088 (
		\u0_u1_csc_reg[15]/P0001 ,
		_w6022_,
		_w6047_
	);
	LUT2 #(
		.INIT('h4)
	) name5089 (
		\wb_data_i[15]_pad ,
		_w6022_,
		_w6048_
	);
	LUT2 #(
		.INIT('h1)
	) name5090 (
		\u0_rst_r2_reg/NET0131 ,
		_w6047_,
		_w6049_
	);
	LUT2 #(
		.INIT('h4)
	) name5091 (
		_w6048_,
		_w6049_,
		_w6050_
	);
	LUT2 #(
		.INIT('h1)
	) name5092 (
		\u0_u1_csc_reg[17]/P0001 ,
		_w6022_,
		_w6051_
	);
	LUT2 #(
		.INIT('h4)
	) name5093 (
		\wb_data_i[17]_pad ,
		_w6022_,
		_w6052_
	);
	LUT2 #(
		.INIT('h1)
	) name5094 (
		\u0_rst_r2_reg/NET0131 ,
		_w6051_,
		_w6053_
	);
	LUT2 #(
		.INIT('h4)
	) name5095 (
		_w6052_,
		_w6053_,
		_w6054_
	);
	LUT2 #(
		.INIT('h1)
	) name5096 (
		\u0_u1_csc_reg[18]/P0001 ,
		_w6022_,
		_w6055_
	);
	LUT2 #(
		.INIT('h4)
	) name5097 (
		\wb_data_i[18]_pad ,
		_w6022_,
		_w6056_
	);
	LUT2 #(
		.INIT('h1)
	) name5098 (
		\u0_rst_r2_reg/NET0131 ,
		_w6055_,
		_w6057_
	);
	LUT2 #(
		.INIT('h4)
	) name5099 (
		_w6056_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('h1)
	) name5100 (
		\u0_u1_csc_reg[19]/P0001 ,
		_w6022_,
		_w6059_
	);
	LUT2 #(
		.INIT('h4)
	) name5101 (
		\wb_data_i[19]_pad ,
		_w6022_,
		_w6060_
	);
	LUT2 #(
		.INIT('h1)
	) name5102 (
		\u0_rst_r2_reg/NET0131 ,
		_w6059_,
		_w6061_
	);
	LUT2 #(
		.INIT('h4)
	) name5103 (
		_w6060_,
		_w6061_,
		_w6062_
	);
	LUT2 #(
		.INIT('h1)
	) name5104 (
		\u0_u1_csc_reg[1]/NET0131 ,
		_w6022_,
		_w6063_
	);
	LUT2 #(
		.INIT('h4)
	) name5105 (
		\wb_data_i[1]_pad ,
		_w6022_,
		_w6064_
	);
	LUT2 #(
		.INIT('h1)
	) name5106 (
		\u0_rst_r2_reg/NET0131 ,
		_w6063_,
		_w6065_
	);
	LUT2 #(
		.INIT('h4)
	) name5107 (
		_w6064_,
		_w6065_,
		_w6066_
	);
	LUT2 #(
		.INIT('h1)
	) name5108 (
		\u0_u1_csc_reg[20]/P0001 ,
		_w6022_,
		_w6067_
	);
	LUT2 #(
		.INIT('h4)
	) name5109 (
		\wb_data_i[20]_pad ,
		_w6022_,
		_w6068_
	);
	LUT2 #(
		.INIT('h1)
	) name5110 (
		\u0_rst_r2_reg/NET0131 ,
		_w6067_,
		_w6069_
	);
	LUT2 #(
		.INIT('h4)
	) name5111 (
		_w6068_,
		_w6069_,
		_w6070_
	);
	LUT2 #(
		.INIT('h1)
	) name5112 (
		\u0_u0_csc_reg[29]/P0001 ,
		_w5057_,
		_w6071_
	);
	LUT2 #(
		.INIT('h4)
	) name5113 (
		\wb_data_i[29]_pad ,
		_w5057_,
		_w6072_
	);
	LUT2 #(
		.INIT('h1)
	) name5114 (
		\u0_rst_r2_reg/NET0131 ,
		_w6071_,
		_w6073_
	);
	LUT2 #(
		.INIT('h4)
	) name5115 (
		_w6072_,
		_w6073_,
		_w6074_
	);
	LUT2 #(
		.INIT('h1)
	) name5116 (
		\u0_u1_csc_reg[22]/P0001 ,
		_w6022_,
		_w6075_
	);
	LUT2 #(
		.INIT('h4)
	) name5117 (
		\wb_data_i[22]_pad ,
		_w6022_,
		_w6076_
	);
	LUT2 #(
		.INIT('h1)
	) name5118 (
		\u0_rst_r2_reg/NET0131 ,
		_w6075_,
		_w6077_
	);
	LUT2 #(
		.INIT('h4)
	) name5119 (
		_w6076_,
		_w6077_,
		_w6078_
	);
	LUT2 #(
		.INIT('h1)
	) name5120 (
		\u0_u1_csc_reg[23]/P0001 ,
		_w6022_,
		_w6079_
	);
	LUT2 #(
		.INIT('h4)
	) name5121 (
		\wb_data_i[23]_pad ,
		_w6022_,
		_w6080_
	);
	LUT2 #(
		.INIT('h1)
	) name5122 (
		\u0_rst_r2_reg/NET0131 ,
		_w6079_,
		_w6081_
	);
	LUT2 #(
		.INIT('h4)
	) name5123 (
		_w6080_,
		_w6081_,
		_w6082_
	);
	LUT2 #(
		.INIT('h1)
	) name5124 (
		\u0_u1_csc_reg[21]/P0001 ,
		_w6022_,
		_w6083_
	);
	LUT2 #(
		.INIT('h4)
	) name5125 (
		\wb_data_i[21]_pad ,
		_w6022_,
		_w6084_
	);
	LUT2 #(
		.INIT('h1)
	) name5126 (
		\u0_rst_r2_reg/NET0131 ,
		_w6083_,
		_w6085_
	);
	LUT2 #(
		.INIT('h4)
	) name5127 (
		_w6084_,
		_w6085_,
		_w6086_
	);
	LUT2 #(
		.INIT('h1)
	) name5128 (
		\u0_u1_csc_reg[24]/P0001 ,
		_w6022_,
		_w6087_
	);
	LUT2 #(
		.INIT('h4)
	) name5129 (
		\wb_data_i[24]_pad ,
		_w6022_,
		_w6088_
	);
	LUT2 #(
		.INIT('h1)
	) name5130 (
		\u0_rst_r2_reg/NET0131 ,
		_w6087_,
		_w6089_
	);
	LUT2 #(
		.INIT('h4)
	) name5131 (
		_w6088_,
		_w6089_,
		_w6090_
	);
	LUT2 #(
		.INIT('h1)
	) name5132 (
		\u0_u1_csc_reg[25]/P0001 ,
		_w6022_,
		_w6091_
	);
	LUT2 #(
		.INIT('h4)
	) name5133 (
		\wb_data_i[25]_pad ,
		_w6022_,
		_w6092_
	);
	LUT2 #(
		.INIT('h1)
	) name5134 (
		\u0_rst_r2_reg/NET0131 ,
		_w6091_,
		_w6093_
	);
	LUT2 #(
		.INIT('h4)
	) name5135 (
		_w6092_,
		_w6093_,
		_w6094_
	);
	LUT2 #(
		.INIT('h1)
	) name5136 (
		\u0_u1_csc_reg[26]/P0001 ,
		_w6022_,
		_w6095_
	);
	LUT2 #(
		.INIT('h4)
	) name5137 (
		\wb_data_i[26]_pad ,
		_w6022_,
		_w6096_
	);
	LUT2 #(
		.INIT('h1)
	) name5138 (
		\u0_rst_r2_reg/NET0131 ,
		_w6095_,
		_w6097_
	);
	LUT2 #(
		.INIT('h4)
	) name5139 (
		_w6096_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h1)
	) name5140 (
		\u0_u1_csc_reg[27]/P0001 ,
		_w6022_,
		_w6099_
	);
	LUT2 #(
		.INIT('h4)
	) name5141 (
		\wb_data_i[27]_pad ,
		_w6022_,
		_w6100_
	);
	LUT2 #(
		.INIT('h1)
	) name5142 (
		\u0_rst_r2_reg/NET0131 ,
		_w6099_,
		_w6101_
	);
	LUT2 #(
		.INIT('h4)
	) name5143 (
		_w6100_,
		_w6101_,
		_w6102_
	);
	LUT2 #(
		.INIT('h1)
	) name5144 (
		\u0_u1_csc_reg[28]/P0001 ,
		_w6022_,
		_w6103_
	);
	LUT2 #(
		.INIT('h4)
	) name5145 (
		\wb_data_i[28]_pad ,
		_w6022_,
		_w6104_
	);
	LUT2 #(
		.INIT('h1)
	) name5146 (
		\u0_rst_r2_reg/NET0131 ,
		_w6103_,
		_w6105_
	);
	LUT2 #(
		.INIT('h4)
	) name5147 (
		_w6104_,
		_w6105_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name5148 (
		\u0_u0_csc_reg[7]/P0001 ,
		_w5057_,
		_w6107_
	);
	LUT2 #(
		.INIT('h4)
	) name5149 (
		\wb_data_i[7]_pad ,
		_w5057_,
		_w6108_
	);
	LUT2 #(
		.INIT('h1)
	) name5150 (
		\u0_rst_r2_reg/NET0131 ,
		_w6107_,
		_w6109_
	);
	LUT2 #(
		.INIT('h4)
	) name5151 (
		_w6108_,
		_w6109_,
		_w6110_
	);
	LUT2 #(
		.INIT('h1)
	) name5152 (
		\u0_u1_csc_reg[29]/P0001 ,
		_w6022_,
		_w6111_
	);
	LUT2 #(
		.INIT('h4)
	) name5153 (
		\wb_data_i[29]_pad ,
		_w6022_,
		_w6112_
	);
	LUT2 #(
		.INIT('h1)
	) name5154 (
		\u0_rst_r2_reg/NET0131 ,
		_w6111_,
		_w6113_
	);
	LUT2 #(
		.INIT('h4)
	) name5155 (
		_w6112_,
		_w6113_,
		_w6114_
	);
	LUT2 #(
		.INIT('h1)
	) name5156 (
		\u0_u1_csc_reg[2]/NET0131 ,
		_w6022_,
		_w6115_
	);
	LUT2 #(
		.INIT('h4)
	) name5157 (
		\wb_data_i[2]_pad ,
		_w6022_,
		_w6116_
	);
	LUT2 #(
		.INIT('h1)
	) name5158 (
		\u0_rst_r2_reg/NET0131 ,
		_w6115_,
		_w6117_
	);
	LUT2 #(
		.INIT('h4)
	) name5159 (
		_w6116_,
		_w6117_,
		_w6118_
	);
	LUT2 #(
		.INIT('h1)
	) name5160 (
		\u0_u1_csc_reg[30]/P0001 ,
		_w6022_,
		_w6119_
	);
	LUT2 #(
		.INIT('h4)
	) name5161 (
		\wb_data_i[30]_pad ,
		_w6022_,
		_w6120_
	);
	LUT2 #(
		.INIT('h1)
	) name5162 (
		\u0_rst_r2_reg/NET0131 ,
		_w6119_,
		_w6121_
	);
	LUT2 #(
		.INIT('h4)
	) name5163 (
		_w6120_,
		_w6121_,
		_w6122_
	);
	LUT2 #(
		.INIT('h1)
	) name5164 (
		\u0_u1_csc_reg[31]/P0001 ,
		_w6022_,
		_w6123_
	);
	LUT2 #(
		.INIT('h4)
	) name5165 (
		\wb_data_i[31]_pad ,
		_w6022_,
		_w6124_
	);
	LUT2 #(
		.INIT('h1)
	) name5166 (
		\u0_rst_r2_reg/NET0131 ,
		_w6123_,
		_w6125_
	);
	LUT2 #(
		.INIT('h4)
	) name5167 (
		_w6124_,
		_w6125_,
		_w6126_
	);
	LUT2 #(
		.INIT('h1)
	) name5168 (
		\u0_u1_csc_reg[4]/P0001 ,
		_w6022_,
		_w6127_
	);
	LUT2 #(
		.INIT('h4)
	) name5169 (
		\wb_data_i[4]_pad ,
		_w6022_,
		_w6128_
	);
	LUT2 #(
		.INIT('h1)
	) name5170 (
		\u0_rst_r2_reg/NET0131 ,
		_w6127_,
		_w6129_
	);
	LUT2 #(
		.INIT('h4)
	) name5171 (
		_w6128_,
		_w6129_,
		_w6130_
	);
	LUT2 #(
		.INIT('h1)
	) name5172 (
		\u0_u1_csc_reg[3]/NET0131 ,
		_w6022_,
		_w6131_
	);
	LUT2 #(
		.INIT('h4)
	) name5173 (
		\wb_data_i[3]_pad ,
		_w6022_,
		_w6132_
	);
	LUT2 #(
		.INIT('h1)
	) name5174 (
		\u0_rst_r2_reg/NET0131 ,
		_w6131_,
		_w6133_
	);
	LUT2 #(
		.INIT('h4)
	) name5175 (
		_w6132_,
		_w6133_,
		_w6134_
	);
	LUT2 #(
		.INIT('h1)
	) name5176 (
		\u0_u1_csc_reg[5]/P0001 ,
		_w6022_,
		_w6135_
	);
	LUT2 #(
		.INIT('h4)
	) name5177 (
		\wb_data_i[5]_pad ,
		_w6022_,
		_w6136_
	);
	LUT2 #(
		.INIT('h1)
	) name5178 (
		\u0_rst_r2_reg/NET0131 ,
		_w6135_,
		_w6137_
	);
	LUT2 #(
		.INIT('h4)
	) name5179 (
		_w6136_,
		_w6137_,
		_w6138_
	);
	LUT2 #(
		.INIT('h1)
	) name5180 (
		\u0_u1_csc_reg[6]/P0001 ,
		_w6022_,
		_w6139_
	);
	LUT2 #(
		.INIT('h4)
	) name5181 (
		\wb_data_i[6]_pad ,
		_w6022_,
		_w6140_
	);
	LUT2 #(
		.INIT('h1)
	) name5182 (
		\u0_rst_r2_reg/NET0131 ,
		_w6139_,
		_w6141_
	);
	LUT2 #(
		.INIT('h4)
	) name5183 (
		_w6140_,
		_w6141_,
		_w6142_
	);
	LUT2 #(
		.INIT('h1)
	) name5184 (
		\u0_u0_csc_reg[8]/P0001 ,
		_w5057_,
		_w6143_
	);
	LUT2 #(
		.INIT('h4)
	) name5185 (
		\wb_data_i[8]_pad ,
		_w5057_,
		_w6144_
	);
	LUT2 #(
		.INIT('h1)
	) name5186 (
		\u0_rst_r2_reg/NET0131 ,
		_w6143_,
		_w6145_
	);
	LUT2 #(
		.INIT('h4)
	) name5187 (
		_w6144_,
		_w6145_,
		_w6146_
	);
	LUT2 #(
		.INIT('h1)
	) name5188 (
		\u0_u1_csc_reg[8]/P0001 ,
		_w6022_,
		_w6147_
	);
	LUT2 #(
		.INIT('h4)
	) name5189 (
		\wb_data_i[8]_pad ,
		_w6022_,
		_w6148_
	);
	LUT2 #(
		.INIT('h1)
	) name5190 (
		\u0_rst_r2_reg/NET0131 ,
		_w6147_,
		_w6149_
	);
	LUT2 #(
		.INIT('h4)
	) name5191 (
		_w6148_,
		_w6149_,
		_w6150_
	);
	LUT2 #(
		.INIT('h1)
	) name5192 (
		\u0_u1_csc_reg[7]/P0001 ,
		_w6022_,
		_w6151_
	);
	LUT2 #(
		.INIT('h4)
	) name5193 (
		\wb_data_i[7]_pad ,
		_w6022_,
		_w6152_
	);
	LUT2 #(
		.INIT('h1)
	) name5194 (
		\u0_rst_r2_reg/NET0131 ,
		_w6151_,
		_w6153_
	);
	LUT2 #(
		.INIT('h4)
	) name5195 (
		_w6152_,
		_w6153_,
		_w6154_
	);
	LUT2 #(
		.INIT('h1)
	) name5196 (
		\u0_u1_csc_reg[9]/P0001 ,
		_w6022_,
		_w6155_
	);
	LUT2 #(
		.INIT('h4)
	) name5197 (
		\wb_data_i[9]_pad ,
		_w6022_,
		_w6156_
	);
	LUT2 #(
		.INIT('h1)
	) name5198 (
		\u0_rst_r2_reg/NET0131 ,
		_w6155_,
		_w6157_
	);
	LUT2 #(
		.INIT('h4)
	) name5199 (
		_w6156_,
		_w6157_,
		_w6158_
	);
	LUT2 #(
		.INIT('h1)
	) name5200 (
		\u0_u1_tms_reg[0]/P0001 ,
		_w5820_,
		_w6159_
	);
	LUT2 #(
		.INIT('h4)
	) name5201 (
		\wb_data_i[0]_pad ,
		_w5820_,
		_w6160_
	);
	LUT2 #(
		.INIT('h1)
	) name5202 (
		\u0_rst_r2_reg/NET0131 ,
		_w6159_,
		_w6161_
	);
	LUT2 #(
		.INIT('h4)
	) name5203 (
		_w6160_,
		_w6161_,
		_w6162_
	);
	LUT2 #(
		.INIT('h1)
	) name5204 (
		\u0_u1_tms_reg[30]/P0001 ,
		_w5820_,
		_w6163_
	);
	LUT2 #(
		.INIT('h4)
	) name5205 (
		\wb_data_i[30]_pad ,
		_w5820_,
		_w6164_
	);
	LUT2 #(
		.INIT('h1)
	) name5206 (
		\u0_rst_r2_reg/NET0131 ,
		_w6163_,
		_w6165_
	);
	LUT2 #(
		.INIT('h4)
	) name5207 (
		_w6164_,
		_w6165_,
		_w6166_
	);
	LUT2 #(
		.INIT('h1)
	) name5208 (
		\u0_u1_tms_reg[10]/P0001 ,
		_w5820_,
		_w6167_
	);
	LUT2 #(
		.INIT('h4)
	) name5209 (
		\wb_data_i[10]_pad ,
		_w5820_,
		_w6168_
	);
	LUT2 #(
		.INIT('h1)
	) name5210 (
		\u0_rst_r2_reg/NET0131 ,
		_w6167_,
		_w6169_
	);
	LUT2 #(
		.INIT('h4)
	) name5211 (
		_w6168_,
		_w6169_,
		_w6170_
	);
	LUT2 #(
		.INIT('h1)
	) name5212 (
		\u0_u1_tms_reg[11]/P0001 ,
		_w5820_,
		_w6171_
	);
	LUT2 #(
		.INIT('h4)
	) name5213 (
		\wb_data_i[11]_pad ,
		_w5820_,
		_w6172_
	);
	LUT2 #(
		.INIT('h1)
	) name5214 (
		\u0_rst_r2_reg/NET0131 ,
		_w6171_,
		_w6173_
	);
	LUT2 #(
		.INIT('h4)
	) name5215 (
		_w6172_,
		_w6173_,
		_w6174_
	);
	LUT2 #(
		.INIT('h1)
	) name5216 (
		\u0_u1_tms_reg[12]/P0001 ,
		_w5820_,
		_w6175_
	);
	LUT2 #(
		.INIT('h4)
	) name5217 (
		\wb_data_i[12]_pad ,
		_w5820_,
		_w6176_
	);
	LUT2 #(
		.INIT('h1)
	) name5218 (
		\u0_rst_r2_reg/NET0131 ,
		_w6175_,
		_w6177_
	);
	LUT2 #(
		.INIT('h4)
	) name5219 (
		_w6176_,
		_w6177_,
		_w6178_
	);
	LUT2 #(
		.INIT('h1)
	) name5220 (
		\u0_u1_tms_reg[13]/P0001 ,
		_w5820_,
		_w6179_
	);
	LUT2 #(
		.INIT('h4)
	) name5221 (
		\wb_data_i[13]_pad ,
		_w5820_,
		_w6180_
	);
	LUT2 #(
		.INIT('h1)
	) name5222 (
		\u0_rst_r2_reg/NET0131 ,
		_w6179_,
		_w6181_
	);
	LUT2 #(
		.INIT('h4)
	) name5223 (
		_w6180_,
		_w6181_,
		_w6182_
	);
	LUT2 #(
		.INIT('h1)
	) name5224 (
		\u0_u1_tms_reg[14]/P0001 ,
		_w5820_,
		_w6183_
	);
	LUT2 #(
		.INIT('h4)
	) name5225 (
		\wb_data_i[14]_pad ,
		_w5820_,
		_w6184_
	);
	LUT2 #(
		.INIT('h1)
	) name5226 (
		\u0_rst_r2_reg/NET0131 ,
		_w6183_,
		_w6185_
	);
	LUT2 #(
		.INIT('h4)
	) name5227 (
		_w6184_,
		_w6185_,
		_w6186_
	);
	LUT2 #(
		.INIT('h1)
	) name5228 (
		\u0_u1_tms_reg[15]/P0001 ,
		_w5820_,
		_w6187_
	);
	LUT2 #(
		.INIT('h4)
	) name5229 (
		\wb_data_i[15]_pad ,
		_w5820_,
		_w6188_
	);
	LUT2 #(
		.INIT('h1)
	) name5230 (
		\u0_rst_r2_reg/NET0131 ,
		_w6187_,
		_w6189_
	);
	LUT2 #(
		.INIT('h4)
	) name5231 (
		_w6188_,
		_w6189_,
		_w6190_
	);
	LUT2 #(
		.INIT('h1)
	) name5232 (
		\u0_u1_tms_reg[18]/P0001 ,
		_w5820_,
		_w6191_
	);
	LUT2 #(
		.INIT('h4)
	) name5233 (
		\wb_data_i[18]_pad ,
		_w5820_,
		_w6192_
	);
	LUT2 #(
		.INIT('h1)
	) name5234 (
		\u0_rst_r2_reg/NET0131 ,
		_w6191_,
		_w6193_
	);
	LUT2 #(
		.INIT('h4)
	) name5235 (
		_w6192_,
		_w6193_,
		_w6194_
	);
	LUT2 #(
		.INIT('h1)
	) name5236 (
		\u0_u1_tms_reg[20]/P0001 ,
		_w5820_,
		_w6195_
	);
	LUT2 #(
		.INIT('h4)
	) name5237 (
		\wb_data_i[20]_pad ,
		_w5820_,
		_w6196_
	);
	LUT2 #(
		.INIT('h1)
	) name5238 (
		\u0_rst_r2_reg/NET0131 ,
		_w6195_,
		_w6197_
	);
	LUT2 #(
		.INIT('h4)
	) name5239 (
		_w6196_,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h1)
	) name5240 (
		\u0_u1_tms_reg[21]/P0001 ,
		_w5820_,
		_w6199_
	);
	LUT2 #(
		.INIT('h4)
	) name5241 (
		\wb_data_i[21]_pad ,
		_w5820_,
		_w6200_
	);
	LUT2 #(
		.INIT('h1)
	) name5242 (
		\u0_rst_r2_reg/NET0131 ,
		_w6199_,
		_w6201_
	);
	LUT2 #(
		.INIT('h4)
	) name5243 (
		_w6200_,
		_w6201_,
		_w6202_
	);
	LUT2 #(
		.INIT('h1)
	) name5244 (
		\u0_u1_tms_reg[24]/P0001 ,
		_w5820_,
		_w6203_
	);
	LUT2 #(
		.INIT('h4)
	) name5245 (
		\wb_data_i[24]_pad ,
		_w5820_,
		_w6204_
	);
	LUT2 #(
		.INIT('h1)
	) name5246 (
		\u0_rst_r2_reg/NET0131 ,
		_w6203_,
		_w6205_
	);
	LUT2 #(
		.INIT('h4)
	) name5247 (
		_w6204_,
		_w6205_,
		_w6206_
	);
	LUT2 #(
		.INIT('h1)
	) name5248 (
		\u0_u1_tms_reg[25]/P0001 ,
		_w5820_,
		_w6207_
	);
	LUT2 #(
		.INIT('h4)
	) name5249 (
		\wb_data_i[25]_pad ,
		_w5820_,
		_w6208_
	);
	LUT2 #(
		.INIT('h1)
	) name5250 (
		\u0_rst_r2_reg/NET0131 ,
		_w6207_,
		_w6209_
	);
	LUT2 #(
		.INIT('h4)
	) name5251 (
		_w6208_,
		_w6209_,
		_w6210_
	);
	LUT2 #(
		.INIT('h1)
	) name5252 (
		\u0_u1_tms_reg[27]/P0001 ,
		_w5820_,
		_w6211_
	);
	LUT2 #(
		.INIT('h4)
	) name5253 (
		\wb_data_i[27]_pad ,
		_w5820_,
		_w6212_
	);
	LUT2 #(
		.INIT('h1)
	) name5254 (
		\u0_rst_r2_reg/NET0131 ,
		_w6211_,
		_w6213_
	);
	LUT2 #(
		.INIT('h4)
	) name5255 (
		_w6212_,
		_w6213_,
		_w6214_
	);
	LUT2 #(
		.INIT('h1)
	) name5256 (
		\u0_u1_tms_reg[2]/P0001 ,
		_w5820_,
		_w6215_
	);
	LUT2 #(
		.INIT('h4)
	) name5257 (
		\wb_data_i[2]_pad ,
		_w5820_,
		_w6216_
	);
	LUT2 #(
		.INIT('h1)
	) name5258 (
		\u0_rst_r2_reg/NET0131 ,
		_w6215_,
		_w6217_
	);
	LUT2 #(
		.INIT('h4)
	) name5259 (
		_w6216_,
		_w6217_,
		_w6218_
	);
	LUT2 #(
		.INIT('h1)
	) name5260 (
		\u0_u1_tms_reg[31]/P0001 ,
		_w5820_,
		_w6219_
	);
	LUT2 #(
		.INIT('h4)
	) name5261 (
		\wb_data_i[31]_pad ,
		_w5820_,
		_w6220_
	);
	LUT2 #(
		.INIT('h1)
	) name5262 (
		\u0_rst_r2_reg/NET0131 ,
		_w6219_,
		_w6221_
	);
	LUT2 #(
		.INIT('h4)
	) name5263 (
		_w6220_,
		_w6221_,
		_w6222_
	);
	LUT2 #(
		.INIT('h1)
	) name5264 (
		\u0_u0_csc_reg[23]/P0001 ,
		_w5057_,
		_w6223_
	);
	LUT2 #(
		.INIT('h4)
	) name5265 (
		\wb_data_i[23]_pad ,
		_w5057_,
		_w6224_
	);
	LUT2 #(
		.INIT('h1)
	) name5266 (
		\u0_rst_r2_reg/NET0131 ,
		_w6223_,
		_w6225_
	);
	LUT2 #(
		.INIT('h4)
	) name5267 (
		_w6224_,
		_w6225_,
		_w6226_
	);
	LUT2 #(
		.INIT('h1)
	) name5268 (
		\u0_u1_tms_reg[3]/P0001 ,
		_w5820_,
		_w6227_
	);
	LUT2 #(
		.INIT('h4)
	) name5269 (
		\wb_data_i[3]_pad ,
		_w5820_,
		_w6228_
	);
	LUT2 #(
		.INIT('h1)
	) name5270 (
		\u0_rst_r2_reg/NET0131 ,
		_w6227_,
		_w6229_
	);
	LUT2 #(
		.INIT('h4)
	) name5271 (
		_w6228_,
		_w6229_,
		_w6230_
	);
	LUT2 #(
		.INIT('h1)
	) name5272 (
		\u0_u1_tms_reg[5]/P0001 ,
		_w5820_,
		_w6231_
	);
	LUT2 #(
		.INIT('h4)
	) name5273 (
		\wb_data_i[5]_pad ,
		_w5820_,
		_w6232_
	);
	LUT2 #(
		.INIT('h1)
	) name5274 (
		\u0_rst_r2_reg/NET0131 ,
		_w6231_,
		_w6233_
	);
	LUT2 #(
		.INIT('h4)
	) name5275 (
		_w6232_,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h1)
	) name5276 (
		\u0_u1_tms_reg[8]/P0001 ,
		_w5820_,
		_w6235_
	);
	LUT2 #(
		.INIT('h4)
	) name5277 (
		\wb_data_i[8]_pad ,
		_w5820_,
		_w6236_
	);
	LUT2 #(
		.INIT('h1)
	) name5278 (
		\u0_rst_r2_reg/NET0131 ,
		_w6235_,
		_w6237_
	);
	LUT2 #(
		.INIT('h4)
	) name5279 (
		_w6236_,
		_w6237_,
		_w6238_
	);
	LUT2 #(
		.INIT('h1)
	) name5280 (
		\u0_u1_tms_reg[9]/P0001 ,
		_w5820_,
		_w6239_
	);
	LUT2 #(
		.INIT('h4)
	) name5281 (
		\wb_data_i[9]_pad ,
		_w5820_,
		_w6240_
	);
	LUT2 #(
		.INIT('h1)
	) name5282 (
		\u0_rst_r2_reg/NET0131 ,
		_w6239_,
		_w6241_
	);
	LUT2 #(
		.INIT('h4)
	) name5283 (
		_w6240_,
		_w6241_,
		_w6242_
	);
	LUT2 #(
		.INIT('h8)
	) name5284 (
		\wb_data_i[20]_pad ,
		_w5893_,
		_w6243_
	);
	LUT2 #(
		.INIT('h2)
	) name5285 (
		\u0_u0_tms_reg[20]/P0001 ,
		_w5893_,
		_w6244_
	);
	LUT2 #(
		.INIT('h1)
	) name5286 (
		\u0_rst_r2_reg/NET0131 ,
		_w6243_,
		_w6245_
	);
	LUT2 #(
		.INIT('h4)
	) name5287 (
		_w6244_,
		_w6245_,
		_w6246_
	);
	LUT2 #(
		.INIT('h1)
	) name5288 (
		\u0_u1_tms_reg[1]/P0001 ,
		_w5820_,
		_w6247_
	);
	LUT2 #(
		.INIT('h4)
	) name5289 (
		\wb_data_i[1]_pad ,
		_w5820_,
		_w6248_
	);
	LUT2 #(
		.INIT('h1)
	) name5290 (
		\u0_rst_r2_reg/NET0131 ,
		_w6247_,
		_w6249_
	);
	LUT2 #(
		.INIT('h4)
	) name5291 (
		_w6248_,
		_w6249_,
		_w6250_
	);
	LUT2 #(
		.INIT('h1)
	) name5292 (
		\u0_u1_tms_reg[6]/P0001 ,
		_w5820_,
		_w6251_
	);
	LUT2 #(
		.INIT('h4)
	) name5293 (
		\wb_data_i[6]_pad ,
		_w5820_,
		_w6252_
	);
	LUT2 #(
		.INIT('h1)
	) name5294 (
		\u0_rst_r2_reg/NET0131 ,
		_w6251_,
		_w6253_
	);
	LUT2 #(
		.INIT('h4)
	) name5295 (
		_w6252_,
		_w6253_,
		_w6254_
	);
	LUT2 #(
		.INIT('h1)
	) name5296 (
		\u0_u1_tms_reg[29]/P0001 ,
		_w5820_,
		_w6255_
	);
	LUT2 #(
		.INIT('h4)
	) name5297 (
		\wb_data_i[29]_pad ,
		_w5820_,
		_w6256_
	);
	LUT2 #(
		.INIT('h1)
	) name5298 (
		\u0_rst_r2_reg/NET0131 ,
		_w6255_,
		_w6257_
	);
	LUT2 #(
		.INIT('h4)
	) name5299 (
		_w6256_,
		_w6257_,
		_w6258_
	);
	LUT2 #(
		.INIT('h1)
	) name5300 (
		\u0_u1_tms_reg[28]/P0001 ,
		_w5820_,
		_w6259_
	);
	LUT2 #(
		.INIT('h4)
	) name5301 (
		\wb_data_i[28]_pad ,
		_w5820_,
		_w6260_
	);
	LUT2 #(
		.INIT('h1)
	) name5302 (
		\u0_rst_r2_reg/NET0131 ,
		_w6259_,
		_w6261_
	);
	LUT2 #(
		.INIT('h4)
	) name5303 (
		_w6260_,
		_w6261_,
		_w6262_
	);
	LUT2 #(
		.INIT('h1)
	) name5304 (
		\u0_u1_tms_reg[4]/P0001 ,
		_w5820_,
		_w6263_
	);
	LUT2 #(
		.INIT('h4)
	) name5305 (
		\wb_data_i[4]_pad ,
		_w5820_,
		_w6264_
	);
	LUT2 #(
		.INIT('h1)
	) name5306 (
		\u0_rst_r2_reg/NET0131 ,
		_w6263_,
		_w6265_
	);
	LUT2 #(
		.INIT('h4)
	) name5307 (
		_w6264_,
		_w6265_,
		_w6266_
	);
	LUT2 #(
		.INIT('h1)
	) name5308 (
		\u0_u0_csc_reg[10]/P0001 ,
		_w5057_,
		_w6267_
	);
	LUT2 #(
		.INIT('h4)
	) name5309 (
		\wb_data_i[10]_pad ,
		_w5057_,
		_w6268_
	);
	LUT2 #(
		.INIT('h1)
	) name5310 (
		\u0_rst_r2_reg/NET0131 ,
		_w6267_,
		_w6269_
	);
	LUT2 #(
		.INIT('h4)
	) name5311 (
		_w6268_,
		_w6269_,
		_w6270_
	);
	LUT2 #(
		.INIT('h1)
	) name5312 (
		\u0_u1_tms_reg[26]/P0001 ,
		_w5820_,
		_w6271_
	);
	LUT2 #(
		.INIT('h4)
	) name5313 (
		\wb_data_i[26]_pad ,
		_w5820_,
		_w6272_
	);
	LUT2 #(
		.INIT('h1)
	) name5314 (
		\u0_rst_r2_reg/NET0131 ,
		_w6271_,
		_w6273_
	);
	LUT2 #(
		.INIT('h4)
	) name5315 (
		_w6272_,
		_w6273_,
		_w6274_
	);
	LUT2 #(
		.INIT('h1)
	) name5316 (
		\u0_u1_csc_reg[16]/P0001 ,
		_w6022_,
		_w6275_
	);
	LUT2 #(
		.INIT('h4)
	) name5317 (
		\wb_data_i[16]_pad ,
		_w6022_,
		_w6276_
	);
	LUT2 #(
		.INIT('h1)
	) name5318 (
		\u0_rst_r2_reg/NET0131 ,
		_w6275_,
		_w6277_
	);
	LUT2 #(
		.INIT('h4)
	) name5319 (
		_w6276_,
		_w6277_,
		_w6278_
	);
	LUT2 #(
		.INIT('h1)
	) name5320 (
		\u0_u0_csc_reg[18]/P0001 ,
		_w5057_,
		_w6279_
	);
	LUT2 #(
		.INIT('h4)
	) name5321 (
		\wb_data_i[18]_pad ,
		_w5057_,
		_w6280_
	);
	LUT2 #(
		.INIT('h1)
	) name5322 (
		\u0_rst_r2_reg/NET0131 ,
		_w6279_,
		_w6281_
	);
	LUT2 #(
		.INIT('h4)
	) name5323 (
		_w6280_,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h1)
	) name5324 (
		\u0_u0_csc_reg[31]/P0001 ,
		_w5057_,
		_w6283_
	);
	LUT2 #(
		.INIT('h4)
	) name5325 (
		\wb_data_i[31]_pad ,
		_w5057_,
		_w6284_
	);
	LUT2 #(
		.INIT('h1)
	) name5326 (
		\u0_rst_r2_reg/NET0131 ,
		_w6283_,
		_w6285_
	);
	LUT2 #(
		.INIT('h4)
	) name5327 (
		_w6284_,
		_w6285_,
		_w6286_
	);
	LUT2 #(
		.INIT('h8)
	) name5328 (
		\wb_data_i[31]_pad ,
		_w5893_,
		_w6287_
	);
	LUT2 #(
		.INIT('h2)
	) name5329 (
		\u0_u0_tms_reg[31]/P0001 ,
		_w5893_,
		_w6288_
	);
	LUT2 #(
		.INIT('h1)
	) name5330 (
		\u0_rst_r2_reg/NET0131 ,
		_w6287_,
		_w6289_
	);
	LUT2 #(
		.INIT('h4)
	) name5331 (
		_w6288_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h1)
	) name5332 (
		\u0_u1_tms_reg[7]/P0001 ,
		_w5820_,
		_w6291_
	);
	LUT2 #(
		.INIT('h4)
	) name5333 (
		\wb_data_i[7]_pad ,
		_w5820_,
		_w6292_
	);
	LUT2 #(
		.INIT('h1)
	) name5334 (
		\u0_rst_r2_reg/NET0131 ,
		_w6291_,
		_w6293_
	);
	LUT2 #(
		.INIT('h4)
	) name5335 (
		_w6292_,
		_w6293_,
		_w6294_
	);
	LUT2 #(
		.INIT('h1)
	) name5336 (
		\u0_u0_csc_reg[19]/P0001 ,
		_w5057_,
		_w6295_
	);
	LUT2 #(
		.INIT('h4)
	) name5337 (
		\wb_data_i[19]_pad ,
		_w5057_,
		_w6296_
	);
	LUT2 #(
		.INIT('h1)
	) name5338 (
		\u0_rst_r2_reg/NET0131 ,
		_w6295_,
		_w6297_
	);
	LUT2 #(
		.INIT('h4)
	) name5339 (
		_w6296_,
		_w6297_,
		_w6298_
	);
	LUT2 #(
		.INIT('h1)
	) name5340 (
		\u0_u0_csc_reg[6]/P0001 ,
		_w5057_,
		_w6299_
	);
	LUT2 #(
		.INIT('h4)
	) name5341 (
		\wb_data_i[6]_pad ,
		_w5057_,
		_w6300_
	);
	LUT2 #(
		.INIT('h1)
	) name5342 (
		\u0_rst_r2_reg/NET0131 ,
		_w6299_,
		_w6301_
	);
	LUT2 #(
		.INIT('h4)
	) name5343 (
		_w6300_,
		_w6301_,
		_w6302_
	);
	LUT2 #(
		.INIT('h1)
	) name5344 (
		\u0_u0_csc_reg[9]/P0001 ,
		_w5057_,
		_w6303_
	);
	LUT2 #(
		.INIT('h4)
	) name5345 (
		\wb_data_i[9]_pad ,
		_w5057_,
		_w6304_
	);
	LUT2 #(
		.INIT('h1)
	) name5346 (
		\u0_rst_r2_reg/NET0131 ,
		_w6303_,
		_w6305_
	);
	LUT2 #(
		.INIT('h4)
	) name5347 (
		_w6304_,
		_w6305_,
		_w6306_
	);
	LUT2 #(
		.INIT('h1)
	) name5348 (
		\u1_acs_addr_reg[3]/P0001 ,
		_w4002_,
		_w6307_
	);
	LUT2 #(
		.INIT('h1)
	) name5349 (
		_w4003_,
		_w6307_,
		_w6308_
	);
	LUT2 #(
		.INIT('h1)
	) name5350 (
		\u0_u1_inited_reg/NET0131 ,
		_w5419_,
		_w6309_
	);
	LUT2 #(
		.INIT('h1)
	) name5351 (
		\u0_u0_inited_reg/NET0131 ,
		_w5414_,
		_w6310_
	);
	LUT2 #(
		.INIT('h1)
	) name5352 (
		_w4398_,
		_w5190_,
		_w6311_
	);
	LUT2 #(
		.INIT('h4)
	) name5353 (
		_w5413_,
		_w6311_,
		_w6312_
	);
	LUT2 #(
		.INIT('h8)
	) name5354 (
		_w1378_,
		_w2269_,
		_w6313_
	);
	LUT2 #(
		.INIT('h1)
	) name5355 (
		\u6_read_go_r_reg/NET0131 ,
		_w6313_,
		_w6314_
	);
	LUT2 #(
		.INIT('h2)
	) name5356 (
		_w1381_,
		_w6314_,
		_w6315_
	);
	LUT2 #(
		.INIT('h1)
	) name5357 (
		\u1_acs_addr_reg[9]/P0001 ,
		_w4008_,
		_w6316_
	);
	LUT2 #(
		.INIT('h1)
	) name5358 (
		_w4009_,
		_w6316_,
		_w6317_
	);
	LUT2 #(
		.INIT('h2)
	) name5359 (
		\wb_data_i[11]_pad ,
		\wb_data_i[13]_pad ,
		_w6318_
	);
	LUT2 #(
		.INIT('h4)
	) name5360 (
		\wb_data_i[11]_pad ,
		\wb_data_i[13]_pad ,
		_w6319_
	);
	LUT2 #(
		.INIT('h1)
	) name5361 (
		_w6318_,
		_w6319_,
		_w6320_
	);
	LUT2 #(
		.INIT('h1)
	) name5362 (
		\wb_data_i[15]_pad ,
		\wb_data_i[8]_pad ,
		_w6321_
	);
	LUT2 #(
		.INIT('h8)
	) name5363 (
		\wb_data_i[15]_pad ,
		\wb_data_i[8]_pad ,
		_w6322_
	);
	LUT2 #(
		.INIT('h1)
	) name5364 (
		_w6321_,
		_w6322_,
		_w6323_
	);
	LUT2 #(
		.INIT('h8)
	) name5365 (
		\wb_data_i[9]_pad ,
		_w6323_,
		_w6324_
	);
	LUT2 #(
		.INIT('h1)
	) name5366 (
		\wb_data_i[9]_pad ,
		_w6323_,
		_w6325_
	);
	LUT2 #(
		.INIT('h1)
	) name5367 (
		_w6324_,
		_w6325_,
		_w6326_
	);
	LUT2 #(
		.INIT('h2)
	) name5368 (
		\wb_data_i[10]_pad ,
		\wb_data_i[12]_pad ,
		_w6327_
	);
	LUT2 #(
		.INIT('h4)
	) name5369 (
		\wb_data_i[10]_pad ,
		\wb_data_i[12]_pad ,
		_w6328_
	);
	LUT2 #(
		.INIT('h1)
	) name5370 (
		_w6327_,
		_w6328_,
		_w6329_
	);
	LUT2 #(
		.INIT('h8)
	) name5371 (
		\wb_data_i[14]_pad ,
		_w6329_,
		_w6330_
	);
	LUT2 #(
		.INIT('h1)
	) name5372 (
		\wb_data_i[14]_pad ,
		_w6329_,
		_w6331_
	);
	LUT2 #(
		.INIT('h1)
	) name5373 (
		_w6330_,
		_w6331_,
		_w6332_
	);
	LUT2 #(
		.INIT('h2)
	) name5374 (
		_w6326_,
		_w6332_,
		_w6333_
	);
	LUT2 #(
		.INIT('h4)
	) name5375 (
		_w6326_,
		_w6332_,
		_w6334_
	);
	LUT2 #(
		.INIT('h1)
	) name5376 (
		_w6333_,
		_w6334_,
		_w6335_
	);
	LUT2 #(
		.INIT('h8)
	) name5377 (
		_w6320_,
		_w6335_,
		_w6336_
	);
	LUT2 #(
		.INIT('h1)
	) name5378 (
		_w6320_,
		_w6335_,
		_w6337_
	);
	LUT2 #(
		.INIT('h1)
	) name5379 (
		_w6336_,
		_w6337_,
		_w6338_
	);
	LUT2 #(
		.INIT('h2)
	) name5380 (
		\wb_data_i[1]_pad ,
		\wb_data_i[6]_pad ,
		_w6339_
	);
	LUT2 #(
		.INIT('h4)
	) name5381 (
		\wb_data_i[1]_pad ,
		\wb_data_i[6]_pad ,
		_w6340_
	);
	LUT2 #(
		.INIT('h1)
	) name5382 (
		_w6339_,
		_w6340_,
		_w6341_
	);
	LUT2 #(
		.INIT('h1)
	) name5383 (
		\wb_data_i[2]_pad ,
		\wb_data_i[4]_pad ,
		_w6342_
	);
	LUT2 #(
		.INIT('h8)
	) name5384 (
		\wb_data_i[2]_pad ,
		\wb_data_i[4]_pad ,
		_w6343_
	);
	LUT2 #(
		.INIT('h1)
	) name5385 (
		_w6342_,
		_w6343_,
		_w6344_
	);
	LUT2 #(
		.INIT('h8)
	) name5386 (
		\wb_data_i[5]_pad ,
		_w6344_,
		_w6345_
	);
	LUT2 #(
		.INIT('h1)
	) name5387 (
		\wb_data_i[5]_pad ,
		_w6344_,
		_w6346_
	);
	LUT2 #(
		.INIT('h1)
	) name5388 (
		_w6345_,
		_w6346_,
		_w6347_
	);
	LUT2 #(
		.INIT('h2)
	) name5389 (
		\wb_data_i[0]_pad ,
		\wb_data_i[7]_pad ,
		_w6348_
	);
	LUT2 #(
		.INIT('h4)
	) name5390 (
		\wb_data_i[0]_pad ,
		\wb_data_i[7]_pad ,
		_w6349_
	);
	LUT2 #(
		.INIT('h1)
	) name5391 (
		_w6348_,
		_w6349_,
		_w6350_
	);
	LUT2 #(
		.INIT('h8)
	) name5392 (
		\wb_data_i[3]_pad ,
		_w6350_,
		_w6351_
	);
	LUT2 #(
		.INIT('h1)
	) name5393 (
		\wb_data_i[3]_pad ,
		_w6350_,
		_w6352_
	);
	LUT2 #(
		.INIT('h1)
	) name5394 (
		_w6351_,
		_w6352_,
		_w6353_
	);
	LUT2 #(
		.INIT('h2)
	) name5395 (
		_w6347_,
		_w6353_,
		_w6354_
	);
	LUT2 #(
		.INIT('h4)
	) name5396 (
		_w6347_,
		_w6353_,
		_w6355_
	);
	LUT2 #(
		.INIT('h1)
	) name5397 (
		_w6354_,
		_w6355_,
		_w6356_
	);
	LUT2 #(
		.INIT('h8)
	) name5398 (
		_w6341_,
		_w6356_,
		_w6357_
	);
	LUT2 #(
		.INIT('h1)
	) name5399 (
		_w6341_,
		_w6356_,
		_w6358_
	);
	LUT2 #(
		.INIT('h1)
	) name5400 (
		_w6357_,
		_w6358_,
		_w6359_
	);
	LUT2 #(
		.INIT('h2)
	) name5401 (
		\wb_data_i[27]_pad ,
		\wb_data_i[29]_pad ,
		_w6360_
	);
	LUT2 #(
		.INIT('h4)
	) name5402 (
		\wb_data_i[27]_pad ,
		\wb_data_i[29]_pad ,
		_w6361_
	);
	LUT2 #(
		.INIT('h1)
	) name5403 (
		_w6360_,
		_w6361_,
		_w6362_
	);
	LUT2 #(
		.INIT('h1)
	) name5404 (
		\wb_data_i[24]_pad ,
		\wb_data_i[31]_pad ,
		_w6363_
	);
	LUT2 #(
		.INIT('h8)
	) name5405 (
		\wb_data_i[24]_pad ,
		\wb_data_i[31]_pad ,
		_w6364_
	);
	LUT2 #(
		.INIT('h1)
	) name5406 (
		_w6363_,
		_w6364_,
		_w6365_
	);
	LUT2 #(
		.INIT('h8)
	) name5407 (
		\wb_data_i[30]_pad ,
		_w6365_,
		_w6366_
	);
	LUT2 #(
		.INIT('h1)
	) name5408 (
		\wb_data_i[30]_pad ,
		_w6365_,
		_w6367_
	);
	LUT2 #(
		.INIT('h1)
	) name5409 (
		_w6366_,
		_w6367_,
		_w6368_
	);
	LUT2 #(
		.INIT('h2)
	) name5410 (
		\wb_data_i[26]_pad ,
		\wb_data_i[28]_pad ,
		_w6369_
	);
	LUT2 #(
		.INIT('h4)
	) name5411 (
		\wb_data_i[26]_pad ,
		\wb_data_i[28]_pad ,
		_w6370_
	);
	LUT2 #(
		.INIT('h1)
	) name5412 (
		_w6369_,
		_w6370_,
		_w6371_
	);
	LUT2 #(
		.INIT('h8)
	) name5413 (
		\wb_data_i[25]_pad ,
		_w6371_,
		_w6372_
	);
	LUT2 #(
		.INIT('h1)
	) name5414 (
		\wb_data_i[25]_pad ,
		_w6371_,
		_w6373_
	);
	LUT2 #(
		.INIT('h1)
	) name5415 (
		_w6372_,
		_w6373_,
		_w6374_
	);
	LUT2 #(
		.INIT('h2)
	) name5416 (
		_w6368_,
		_w6374_,
		_w6375_
	);
	LUT2 #(
		.INIT('h4)
	) name5417 (
		_w6368_,
		_w6374_,
		_w6376_
	);
	LUT2 #(
		.INIT('h1)
	) name5418 (
		_w6375_,
		_w6376_,
		_w6377_
	);
	LUT2 #(
		.INIT('h8)
	) name5419 (
		_w6362_,
		_w6377_,
		_w6378_
	);
	LUT2 #(
		.INIT('h1)
	) name5420 (
		_w6362_,
		_w6377_,
		_w6379_
	);
	LUT2 #(
		.INIT('h1)
	) name5421 (
		_w6378_,
		_w6379_,
		_w6380_
	);
	LUT2 #(
		.INIT('h2)
	) name5422 (
		\wb_data_i[17]_pad ,
		\wb_data_i[22]_pad ,
		_w6381_
	);
	LUT2 #(
		.INIT('h4)
	) name5423 (
		\wb_data_i[17]_pad ,
		\wb_data_i[22]_pad ,
		_w6382_
	);
	LUT2 #(
		.INIT('h1)
	) name5424 (
		_w6381_,
		_w6382_,
		_w6383_
	);
	LUT2 #(
		.INIT('h1)
	) name5425 (
		\wb_data_i[16]_pad ,
		\wb_data_i[23]_pad ,
		_w6384_
	);
	LUT2 #(
		.INIT('h8)
	) name5426 (
		\wb_data_i[16]_pad ,
		\wb_data_i[23]_pad ,
		_w6385_
	);
	LUT2 #(
		.INIT('h1)
	) name5427 (
		_w6384_,
		_w6385_,
		_w6386_
	);
	LUT2 #(
		.INIT('h8)
	) name5428 (
		\wb_data_i[21]_pad ,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h1)
	) name5429 (
		\wb_data_i[21]_pad ,
		_w6386_,
		_w6388_
	);
	LUT2 #(
		.INIT('h1)
	) name5430 (
		_w6387_,
		_w6388_,
		_w6389_
	);
	LUT2 #(
		.INIT('h2)
	) name5431 (
		\wb_data_i[18]_pad ,
		\wb_data_i[20]_pad ,
		_w6390_
	);
	LUT2 #(
		.INIT('h4)
	) name5432 (
		\wb_data_i[18]_pad ,
		\wb_data_i[20]_pad ,
		_w6391_
	);
	LUT2 #(
		.INIT('h1)
	) name5433 (
		_w6390_,
		_w6391_,
		_w6392_
	);
	LUT2 #(
		.INIT('h8)
	) name5434 (
		\wb_data_i[19]_pad ,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h1)
	) name5435 (
		\wb_data_i[19]_pad ,
		_w6392_,
		_w6394_
	);
	LUT2 #(
		.INIT('h1)
	) name5436 (
		_w6393_,
		_w6394_,
		_w6395_
	);
	LUT2 #(
		.INIT('h2)
	) name5437 (
		_w6389_,
		_w6395_,
		_w6396_
	);
	LUT2 #(
		.INIT('h4)
	) name5438 (
		_w6389_,
		_w6395_,
		_w6397_
	);
	LUT2 #(
		.INIT('h1)
	) name5439 (
		_w6396_,
		_w6397_,
		_w6398_
	);
	LUT2 #(
		.INIT('h8)
	) name5440 (
		_w6383_,
		_w6398_,
		_w6399_
	);
	LUT2 #(
		.INIT('h1)
	) name5441 (
		_w6383_,
		_w6398_,
		_w6400_
	);
	LUT2 #(
		.INIT('h1)
	) name5442 (
		_w6399_,
		_w6400_,
		_w6401_
	);
	LUT2 #(
		.INIT('h8)
	) name5443 (
		_w1870_,
		_w2269_,
		_w6402_
	);
	LUT2 #(
		.INIT('h1)
	) name5444 (
		\u6_write_go_r_reg/NET0131 ,
		_w6402_,
		_w6403_
	);
	LUT2 #(
		.INIT('h2)
	) name5445 (
		wb_cyc_i_pad,
		_w6403_,
		_w6404_
	);
	LUT2 #(
		.INIT('h1)
	) name5446 (
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_sreq_cs_le_reg/NET0131 ,
		_w6405_
	);
	LUT2 #(
		.INIT('h1)
	) name5447 (
		\u0_init_req_reg/NET0131 ,
		\u0_u0_lmr_req_reg/NET0131 ,
		_w6406_
	);
	LUT2 #(
		.INIT('h2)
	) name5448 (
		\u0_init_req_reg/NET0131 ,
		\u0_u0_init_req_reg/NET0131 ,
		_w6407_
	);
	LUT2 #(
		.INIT('h2)
	) name5449 (
		\u0_sreq_cs_le_reg/NET0131 ,
		_w6406_,
		_w6408_
	);
	LUT2 #(
		.INIT('h4)
	) name5450 (
		_w6407_,
		_w6408_,
		_w6409_
	);
	LUT2 #(
		.INIT('h1)
	) name5451 (
		\u0_init_req_reg/NET0131 ,
		\u0_u1_lmr_req_reg/NET0131 ,
		_w6410_
	);
	LUT2 #(
		.INIT('h2)
	) name5452 (
		\u0_init_req_reg/NET0131 ,
		\u0_u1_init_req_reg/NET0131 ,
		_w6411_
	);
	LUT2 #(
		.INIT('h1)
	) name5453 (
		_w6410_,
		_w6411_,
		_w6412_
	);
	LUT2 #(
		.INIT('h2)
	) name5454 (
		\u0_sreq_cs_le_reg/NET0131 ,
		_w6412_,
		_w6413_
	);
	LUT2 #(
		.INIT('h1)
	) name5455 (
		_w6405_,
		_w6409_,
		_w6414_
	);
	LUT2 #(
		.INIT('h4)
	) name5456 (
		_w6413_,
		_w6414_,
		_w6415_
	);
	LUT2 #(
		.INIT('h1)
	) name5457 (
		\u1_acs_addr_reg[2]/P0001 ,
		_w4001_,
		_w6416_
	);
	LUT2 #(
		.INIT('h1)
	) name5458 (
		_w4002_,
		_w6416_,
		_w6417_
	);
	LUT2 #(
		.INIT('h1)
	) name5459 (
		\u1_acs_addr_reg[5]/P0001 ,
		_w4004_,
		_w6418_
	);
	LUT2 #(
		.INIT('h1)
	) name5460 (
		_w4005_,
		_w6418_,
		_w6419_
	);
	LUT2 #(
		.INIT('h1)
	) name5461 (
		suspended_o_pad,
		\u0_csr_r_reg[2]/NET0131 ,
		_w6420_
	);
	LUT2 #(
		.INIT('h4)
	) name5462 (
		\u0_rf_we_reg/NET0131 ,
		_w1047_,
		_w6421_
	);
	LUT2 #(
		.INIT('h8)
	) name5463 (
		_w2273_,
		_w6421_,
		_w6422_
	);
	LUT2 #(
		.INIT('h8)
	) name5464 (
		\u5_lookup_ready1_reg/NET0131 ,
		_w1046_,
		_w6423_
	);
	LUT2 #(
		.INIT('h2)
	) name5465 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		_w6424_
	);
	LUT2 #(
		.INIT('h4)
	) name5466 (
		\u0_u0_addr_r_reg[4]/P0001 ,
		_w6424_,
		_w6425_
	);
	LUT2 #(
		.INIT('h8)
	) name5467 (
		_w5055_,
		_w6425_,
		_w6426_
	);
	LUT2 #(
		.INIT('h8)
	) name5468 (
		_w5818_,
		_w6425_,
		_w6427_
	);
	LUT2 #(
		.INIT('h2)
	) name5469 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_sreq_cs_le_reg/NET0131 ,
		_w6428_
	);
	LUT2 #(
		.INIT('h1)
	) name5470 (
		_w6409_,
		_w6428_,
		_w6429_
	);
	LUT2 #(
		.INIT('h1)
	) name5471 (
		\mem_ack_r_reg/P0001 ,
		\u0_csc_reg[1]/NET0131 ,
		_w6430_
	);
	LUT2 #(
		.INIT('h8)
	) name5472 (
		_w5064_,
		_w6430_,
		_w6431_
	);
	LUT2 #(
		.INIT('h1)
	) name5473 (
		_w1621_,
		_w1674_,
		_w6432_
	);
	LUT2 #(
		.INIT('h2)
	) name5474 (
		\u6_wr_hold_reg/NET0131 ,
		_w1046_,
		_w6433_
	);
	LUT2 #(
		.INIT('h1)
	) name5475 (
		_w1047_,
		_w6433_,
		_w6434_
	);
	LUT2 #(
		.INIT('h1)
	) name5476 (
		\u1_acs_addr_reg[0]/P0001 ,
		\u1_acs_addr_reg[1]/P0001 ,
		_w6435_
	);
	LUT2 #(
		.INIT('h1)
	) name5477 (
		_w4001_,
		_w6435_,
		_w6436_
	);
	LUT2 #(
		.INIT('h8)
	) name5478 (
		\u6_rmw_en_reg/NET0131 ,
		wb_cyc_i_pad,
		_w6437_
	);
	LUT2 #(
		.INIT('h1)
	) name5479 (
		wb_ack_o_pad,
		_w6437_,
		_w6438_
	);
	LUT2 #(
		.INIT('h2)
	) name5480 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_mc_le_reg/NET0131 ,
		_w6439_
	);
	LUT2 #(
		.INIT('h8)
	) name5481 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_mc_le_reg/NET0131 ,
		_w6440_
	);
	LUT2 #(
		.INIT('h1)
	) name5482 (
		_w6439_,
		_w6440_,
		_w6441_
	);
	LUT2 #(
		.INIT('h1)
	) name5483 (
		\u0_u0_lmr_req_reg/NET0131 ,
		\u0_u1_lmr_req_reg/NET0131 ,
		_w6442_
	);
	LUT2 #(
		.INIT('h1)
	) name5484 (
		\u0_u0_init_req_reg/NET0131 ,
		\u0_u1_init_req_reg/NET0131 ,
		_w6443_
	);
	LUT2 #(
		.INIT('h1)
	) name5485 (
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[54]/NET0131 ,
		_w6444_
	);
	LUT2 #(
		.INIT('h8)
	) name5486 (
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[54]/NET0131 ,
		_w6445_
	);
	LUT2 #(
		.INIT('h1)
	) name5487 (
		_w6444_,
		_w6445_,
		_w6446_
	);
	LUT2 #(
		.INIT('h1)
	) name5488 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[54]/NET0131 ,
		_w6447_
	);
	LUT2 #(
		.INIT('h8)
	) name5489 (
		_w1665_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h8)
	) name5490 (
		_w1742_,
		_w6448_,
		_w6449_
	);
	LUT2 #(
		.INIT('h4)
	) name5491 (
		\u5_state_reg[1]/NET0131 ,
		_w2778_,
		_w6450_
	);
	LUT2 #(
		.INIT('h1)
	) name5492 (
		_w6449_,
		_w6450_,
		_w6451_
	);
	LUT2 #(
		.INIT('h2)
	) name5493 (
		_w6446_,
		_w6451_,
		_w6452_
	);
	LUT2 #(
		.INIT('h1)
	) name5494 (
		\u5_state_reg[46]/NET0131 ,
		_w1132_,
		_w6453_
	);
	LUT2 #(
		.INIT('h4)
	) name5495 (
		_w1147_,
		_w6453_,
		_w6454_
	);
	LUT2 #(
		.INIT('h2)
	) name5496 (
		\u5_state_reg[46]/NET0131 ,
		_w1142_,
		_w6455_
	);
	LUT2 #(
		.INIT('h2)
	) name5497 (
		_w1225_,
		_w6455_,
		_w6456_
	);
	LUT2 #(
		.INIT('h4)
	) name5498 (
		_w6454_,
		_w6456_,
		_w6457_
	);
	LUT2 #(
		.INIT('h8)
	) name5499 (
		_w1280_,
		_w6457_,
		_w6458_
	);
	LUT2 #(
		.INIT('h1)
	) name5500 (
		_w1110_,
		_w1313_,
		_w6459_
	);
	LUT2 #(
		.INIT('h2)
	) name5501 (
		_w968_,
		_w6459_,
		_w6460_
	);
	LUT2 #(
		.INIT('h1)
	) name5502 (
		_w1235_,
		_w1265_,
		_w6461_
	);
	LUT2 #(
		.INIT('h2)
	) name5503 (
		_w1152_,
		_w6461_,
		_w6462_
	);
	LUT2 #(
		.INIT('h1)
	) name5504 (
		_w6460_,
		_w6462_,
		_w6463_
	);
	LUT2 #(
		.INIT('h8)
	) name5505 (
		_w1029_,
		_w1142_,
		_w6464_
	);
	LUT2 #(
		.INIT('h8)
	) name5506 (
		_w3053_,
		_w6464_,
		_w6465_
	);
	LUT2 #(
		.INIT('h4)
	) name5507 (
		_w6463_,
		_w6465_,
		_w6466_
	);
	LUT2 #(
		.INIT('h1)
	) name5508 (
		_w6458_,
		_w6466_,
		_w6467_
	);
	LUT2 #(
		.INIT('h2)
	) name5509 (
		_w1134_,
		_w6467_,
		_w6468_
	);
	LUT2 #(
		.INIT('h2)
	) name5510 (
		_w1133_,
		_w1258_,
		_w6469_
	);
	LUT2 #(
		.INIT('h1)
	) name5511 (
		_w1145_,
		_w1149_,
		_w6470_
	);
	LUT2 #(
		.INIT('h2)
	) name5512 (
		_w986_,
		_w6470_,
		_w6471_
	);
	LUT2 #(
		.INIT('h1)
	) name5513 (
		_w6469_,
		_w6471_,
		_w6472_
	);
	LUT2 #(
		.INIT('h8)
	) name5514 (
		_w968_,
		_w1142_,
		_w6473_
	);
	LUT2 #(
		.INIT('h8)
	) name5515 (
		_w1335_,
		_w6473_,
		_w6474_
	);
	LUT2 #(
		.INIT('h4)
	) name5516 (
		_w6472_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h1)
	) name5517 (
		_w6468_,
		_w6475_,
		_w6476_
	);
	LUT2 #(
		.INIT('h2)
	) name5518 (
		_w1340_,
		_w6476_,
		_w6477_
	);
	LUT2 #(
		.INIT('h1)
	) name5519 (
		_w1243_,
		_w1291_,
		_w6478_
	);
	LUT2 #(
		.INIT('h4)
	) name5520 (
		\u5_state_reg[0]/NET0131 ,
		_w964_,
		_w6479_
	);
	LUT2 #(
		.INIT('h4)
	) name5521 (
		_w6478_,
		_w6479_,
		_w6480_
	);
	LUT2 #(
		.INIT('h8)
	) name5522 (
		_w1337_,
		_w6480_,
		_w6481_
	);
	LUT2 #(
		.INIT('h1)
	) name5523 (
		_w6477_,
		_w6481_,
		_w6482_
	);
	LUT2 #(
		.INIT('h2)
	) name5524 (
		_w5404_,
		_w6446_,
		_w6483_
	);
	LUT2 #(
		.INIT('h4)
	) name5525 (
		_w6482_,
		_w6483_,
		_w6484_
	);
	LUT2 #(
		.INIT('h1)
	) name5526 (
		_w6452_,
		_w6484_,
		_w6485_
	);
	LUT2 #(
		.INIT('h1)
	) name5527 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[10]/NET0131 ,
		_w6486_
	);
	LUT2 #(
		.INIT('h2)
	) name5528 (
		_w1364_,
		_w6486_,
		_w6487_
	);
	LUT2 #(
		.INIT('h4)
	) name5529 (
		\u5_tmr_done_reg/NET0131 ,
		_w1246_,
		_w6488_
	);
	LUT2 #(
		.INIT('h1)
	) name5530 (
		_w6487_,
		_w6488_,
		_w6489_
	);
	LUT2 #(
		.INIT('h8)
	) name5531 (
		\u5_tmr_done_reg/NET0131 ,
		_w1295_,
		_w6490_
	);
	LUT2 #(
		.INIT('h4)
	) name5532 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1358_,
		_w6491_
	);
	LUT2 #(
		.INIT('h1)
	) name5533 (
		_w6490_,
		_w6491_,
		_w6492_
	);
	LUT2 #(
		.INIT('h4)
	) name5534 (
		\u5_tmr_done_reg/NET0131 ,
		_w1131_,
		_w6493_
	);
	LUT2 #(
		.INIT('h1)
	) name5535 (
		_w4450_,
		_w6493_,
		_w6494_
	);
	LUT2 #(
		.INIT('h4)
	) name5536 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1076_,
		_w6495_
	);
	LUT2 #(
		.INIT('h1)
	) name5537 (
		_w1263_,
		_w6495_,
		_w6496_
	);
	LUT2 #(
		.INIT('h2)
	) name5538 (
		\u5_state_reg[26]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w6497_
	);
	LUT2 #(
		.INIT('h1)
	) name5539 (
		_w2795_,
		_w6497_,
		_w6498_
	);
	LUT2 #(
		.INIT('h2)
	) name5540 (
		_w1131_,
		_w6498_,
		_w6499_
	);
	LUT2 #(
		.INIT('h4)
	) name5541 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1395_,
		_w6500_
	);
	LUT2 #(
		.INIT('h1)
	) name5542 (
		_w6499_,
		_w6500_,
		_w6501_
	);
	LUT2 #(
		.INIT('h1)
	) name5543 (
		\u5_state_reg[38]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w6502_
	);
	LUT2 #(
		.INIT('h8)
	) name5544 (
		\u5_tmr2_done_reg/NET0131 ,
		_w2365_,
		_w6503_
	);
	LUT2 #(
		.INIT('h1)
	) name5545 (
		_w6502_,
		_w6503_,
		_w6504_
	);
	LUT2 #(
		.INIT('h8)
	) name5546 (
		_w1292_,
		_w6504_,
		_w6505_
	);
	LUT2 #(
		.INIT('h8)
	) name5547 (
		_w1438_,
		_w1664_,
		_w6506_
	);
	LUT2 #(
		.INIT('h2)
	) name5548 (
		\u5_state_reg[36]/NET0131 ,
		_w2426_,
		_w6507_
	);
	LUT2 #(
		.INIT('h1)
	) name5549 (
		_w6506_,
		_w6507_,
		_w6508_
	);
	LUT2 #(
		.INIT('h2)
	) name5550 (
		_w1679_,
		_w6508_,
		_w6509_
	);
	LUT2 #(
		.INIT('h8)
	) name5551 (
		\u5_state_reg[36]/NET0131 ,
		_w2618_,
		_w6510_
	);
	LUT2 #(
		.INIT('h1)
	) name5552 (
		_w6509_,
		_w6510_,
		_w6511_
	);
	LUT2 #(
		.INIT('h2)
	) name5553 (
		_w1685_,
		_w6511_,
		_w6512_
	);
	LUT2 #(
		.INIT('h4)
	) name5554 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1397_,
		_w6513_
	);
	LUT2 #(
		.INIT('h2)
	) name5555 (
		\u5_state_reg[13]/NET0131 ,
		_w2671_,
		_w6514_
	);
	LUT2 #(
		.INIT('h1)
	) name5556 (
		_w1419_,
		_w6514_,
		_w6515_
	);
	LUT2 #(
		.INIT('h2)
	) name5557 (
		_w1253_,
		_w6515_,
		_w6516_
	);
	LUT2 #(
		.INIT('h1)
	) name5558 (
		_w1384_,
		_w6516_,
		_w6517_
	);
	LUT2 #(
		.INIT('h4)
	) name5559 (
		_w6513_,
		_w6517_,
		_w6518_
	);
	LUT2 #(
		.INIT('h8)
	) name5560 (
		_w3178_,
		_w4215_,
		_w6519_
	);
	LUT2 #(
		.INIT('h4)
	) name5561 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1070_,
		_w6520_
	);
	LUT2 #(
		.INIT('h1)
	) name5562 (
		_w6519_,
		_w6520_,
		_w6521_
	);
	LUT2 #(
		.INIT('h1)
	) name5563 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[28]/NET0131 ,
		_w6522_
	);
	LUT2 #(
		.INIT('h2)
	) name5564 (
		_w1214_,
		_w6522_,
		_w6523_
	);
	LUT2 #(
		.INIT('h8)
	) name5565 (
		\u5_state_reg[28]/NET0131 ,
		_w2646_,
		_w6524_
	);
	LUT2 #(
		.INIT('h1)
	) name5566 (
		_w6523_,
		_w6524_,
		_w6525_
	);
	LUT2 #(
		.INIT('h1)
	) name5567 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[30]/NET0131 ,
		_w6526_
	);
	LUT2 #(
		.INIT('h2)
	) name5568 (
		_w1358_,
		_w6526_,
		_w6527_
	);
	LUT2 #(
		.INIT('h4)
	) name5569 (
		\u5_resume_req_r_reg/NET0131 ,
		_w1206_,
		_w6528_
	);
	LUT2 #(
		.INIT('h1)
	) name5570 (
		_w6527_,
		_w6528_,
		_w6529_
	);
	LUT2 #(
		.INIT('h1)
	) name5571 (
		\u5_state_reg[33]/NET0131 ,
		_w2421_,
		_w6530_
	);
	LUT2 #(
		.INIT('h2)
	) name5572 (
		_w2428_,
		_w6530_,
		_w6531_
	);
	LUT2 #(
		.INIT('h4)
	) name5573 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1214_,
		_w6532_
	);
	LUT2 #(
		.INIT('h1)
	) name5574 (
		_w4909_,
		_w6532_,
		_w6533_
	);
	LUT2 #(
		.INIT('h8)
	) name5575 (
		\u5_state_reg[32]/NET0131 ,
		_w2968_,
		_w6534_
	);
	LUT2 #(
		.INIT('h1)
	) name5576 (
		_w1290_,
		_w6534_,
		_w6535_
	);
	LUT2 #(
		.INIT('h4)
	) name5577 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1217_,
		_w6536_
	);
	LUT2 #(
		.INIT('h2)
	) name5578 (
		\u5_state_reg[4]/NET0131 ,
		_w2426_,
		_w6537_
	);
	LUT2 #(
		.INIT('h4)
	) name5579 (
		\u2_row_same_reg/P0001 ,
		_w2679_,
		_w6538_
	);
	LUT2 #(
		.INIT('h8)
	) name5580 (
		_w2678_,
		_w6538_,
		_w6539_
	);
	LUT2 #(
		.INIT('h1)
	) name5581 (
		_w6537_,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h2)
	) name5582 (
		_w1679_,
		_w6540_,
		_w6541_
	);
	LUT2 #(
		.INIT('h8)
	) name5583 (
		\u5_state_reg[4]/NET0131 ,
		_w2618_,
		_w6542_
	);
	LUT2 #(
		.INIT('h1)
	) name5584 (
		_w6541_,
		_w6542_,
		_w6543_
	);
	LUT2 #(
		.INIT('h8)
	) name5585 (
		_w1283_,
		_w1683_,
		_w6544_
	);
	LUT2 #(
		.INIT('h4)
	) name5586 (
		_w6543_,
		_w6544_,
		_w6545_
	);
	LUT2 #(
		.INIT('h1)
	) name5587 (
		_w1747_,
		_w6536_,
		_w6546_
	);
	LUT2 #(
		.INIT('h4)
	) name5588 (
		_w6545_,
		_w6546_,
		_w6547_
	);
	LUT2 #(
		.INIT('h1)
	) name5589 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[23]/NET0131 ,
		_w6548_
	);
	LUT2 #(
		.INIT('h2)
	) name5590 (
		_w1076_,
		_w6548_,
		_w6549_
	);
	LUT2 #(
		.INIT('h8)
	) name5591 (
		\u5_state_reg[23]/NET0131 ,
		_w2968_,
		_w6550_
	);
	LUT2 #(
		.INIT('h1)
	) name5592 (
		_w6549_,
		_w6550_,
		_w6551_
	);
	LUT2 #(
		.INIT('h8)
	) name5593 (
		wb_cyc_i_pad,
		_w1379_,
		_w6552_
	);
	LUT2 #(
		.INIT('h8)
	) name5594 (
		\u5_state_reg[44]/NET0131 ,
		_w2611_,
		_w6553_
	);
	LUT2 #(
		.INIT('h1)
	) name5595 (
		_w1150_,
		_w6553_,
		_w6554_
	);
	LUT2 #(
		.INIT('h8)
	) name5596 (
		\u6_read_go_r1_reg/NET0131 ,
		wb_cyc_i_pad,
		_w6555_
	);
	LUT2 #(
		.INIT('h1)
	) name5597 (
		\u5_state_reg[39]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w6556_
	);
	LUT2 #(
		.INIT('h2)
	) name5598 (
		_w1227_,
		_w6556_,
		_w6557_
	);
	LUT2 #(
		.INIT('h8)
	) name5599 (
		_w1254_,
		_w1305_,
		_w6558_
	);
	LUT2 #(
		.INIT('h1)
	) name5600 (
		_w6557_,
		_w6558_,
		_w6559_
	);
	LUT2 #(
		.INIT('h2)
	) name5601 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1244_,
		_w6560_
	);
	LUT2 #(
		.INIT('h1)
	) name5602 (
		_w1690_,
		_w6560_,
		_w6561_
	);
	LUT2 #(
		.INIT('h4)
	) name5603 (
		_w2411_,
		_w2414_,
		_w6562_
	);
	LUT2 #(
		.INIT('h2)
	) name5604 (
		_w1106_,
		_w6562_,
		_w6563_
	);
	LUT2 #(
		.INIT('h2)
	) name5605 (
		_w1865_,
		_w6563_,
		_w6564_
	);
	LUT2 #(
		.INIT('h8)
	) name5606 (
		_w3051_,
		_w4607_,
		_w6565_
	);
	LUT2 #(
		.INIT('h8)
	) name5607 (
		_w3098_,
		_w4607_,
		_w6566_
	);
	LUT2 #(
		.INIT('h2)
	) name5608 (
		\u2_u0_bank0_open_reg/NET0131 ,
		_w6566_,
		_w6567_
	);
	LUT2 #(
		.INIT('h8)
	) name5609 (
		_w3092_,
		_w6567_,
		_w6568_
	);
	LUT2 #(
		.INIT('h1)
	) name5610 (
		_w6565_,
		_w6568_,
		_w6569_
	);
	LUT2 #(
		.INIT('h8)
	) name5611 (
		_w3109_,
		_w4607_,
		_w6570_
	);
	LUT2 #(
		.INIT('h8)
	) name5612 (
		_w3113_,
		_w4607_,
		_w6571_
	);
	LUT2 #(
		.INIT('h2)
	) name5613 (
		\u2_u1_bank0_open_reg/NET0131 ,
		_w6571_,
		_w6572_
	);
	LUT2 #(
		.INIT('h8)
	) name5614 (
		_w3112_,
		_w6572_,
		_w6573_
	);
	LUT2 #(
		.INIT('h1)
	) name5615 (
		_w6570_,
		_w6573_,
		_w6574_
	);
	LUT2 #(
		.INIT('h4)
	) name5616 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1390_,
		_w6575_
	);
	LUT2 #(
		.INIT('h8)
	) name5617 (
		\u5_tmr_done_reg/NET0131 ,
		_w1080_,
		_w6576_
	);
	LUT2 #(
		.INIT('h1)
	) name5618 (
		_w6575_,
		_w6576_,
		_w6577_
	);
	LUT2 #(
		.INIT('h1)
	) name5619 (
		_w1087_,
		_w1688_,
		_w6578_
	);
	LUT2 #(
		.INIT('h4)
	) name5620 (
		\u5_state_reg[12]/NET0131 ,
		_w1654_,
		_w6579_
	);
	LUT2 #(
		.INIT('h2)
	) name5621 (
		_w2725_,
		_w6579_,
		_w6580_
	);
	LUT2 #(
		.INIT('h2)
	) name5622 (
		\u5_state_reg[12]/NET0131 ,
		_w2338_,
		_w6581_
	);
	LUT2 #(
		.INIT('h4)
	) name5623 (
		_w1875_,
		_w6581_,
		_w6582_
	);
	LUT2 #(
		.INIT('h1)
	) name5624 (
		_w2340_,
		_w6582_,
		_w6583_
	);
	LUT2 #(
		.INIT('h2)
	) name5625 (
		_w1224_,
		_w6583_,
		_w6584_
	);
	LUT2 #(
		.INIT('h1)
	) name5626 (
		_w6580_,
		_w6584_,
		_w6585_
	);
	LUT2 #(
		.INIT('h1)
	) name5627 (
		_w1200_,
		_w3859_,
		_w6586_
	);
	LUT2 #(
		.INIT('h8)
	) name5628 (
		_w1139_,
		_w1873_,
		_w6587_
	);
	LUT2 #(
		.INIT('h8)
	) name5629 (
		_w1241_,
		_w1629_,
		_w6588_
	);
	LUT2 #(
		.INIT('h1)
	) name5630 (
		_w6587_,
		_w6588_,
		_w6589_
	);
	LUT2 #(
		.INIT('h2)
	) name5631 (
		_w1627_,
		_w6589_,
		_w6590_
	);
	LUT2 #(
		.INIT('h8)
	) name5632 (
		\u3_u0_wr_adr_reg[1]/NET0131 ,
		_w1044_,
		_w6591_
	);
	LUT2 #(
		.INIT('h2)
	) name5633 (
		\u3_u0_wr_adr_reg[0]/NET0131 ,
		_w1044_,
		_w6592_
	);
	LUT2 #(
		.INIT('h1)
	) name5634 (
		_w6591_,
		_w6592_,
		_w6593_
	);
	LUT2 #(
		.INIT('h2)
	) name5635 (
		_w4203_,
		_w6593_,
		_w6594_
	);
	LUT2 #(
		.INIT('h2)
	) name5636 (
		\u7_mc_dqm_r_reg[0]/P0001 ,
		_w1046_,
		_w6595_
	);
	LUT2 #(
		.INIT('h8)
	) name5637 (
		\wb_sel_i[0]_pad ,
		_w1046_,
		_w6596_
	);
	LUT2 #(
		.INIT('h1)
	) name5638 (
		_w6595_,
		_w6596_,
		_w6597_
	);
	LUT2 #(
		.INIT('h2)
	) name5639 (
		\u7_mc_dqm_r_reg[1]/P0001 ,
		_w1046_,
		_w6598_
	);
	LUT2 #(
		.INIT('h8)
	) name5640 (
		\wb_sel_i[1]_pad ,
		_w1046_,
		_w6599_
	);
	LUT2 #(
		.INIT('h1)
	) name5641 (
		_w6598_,
		_w6599_,
		_w6600_
	);
	LUT2 #(
		.INIT('h2)
	) name5642 (
		\u7_mc_dqm_r_reg[2]/P0001 ,
		_w1046_,
		_w6601_
	);
	LUT2 #(
		.INIT('h8)
	) name5643 (
		\wb_sel_i[2]_pad ,
		_w1046_,
		_w6602_
	);
	LUT2 #(
		.INIT('h1)
	) name5644 (
		_w6601_,
		_w6602_,
		_w6603_
	);
	LUT2 #(
		.INIT('h2)
	) name5645 (
		\u7_mc_dqm_r_reg[3]/P0001 ,
		_w1046_,
		_w6604_
	);
	LUT2 #(
		.INIT('h8)
	) name5646 (
		\wb_sel_i[3]_pad ,
		_w1046_,
		_w6605_
	);
	LUT2 #(
		.INIT('h1)
	) name5647 (
		_w6604_,
		_w6605_,
		_w6606_
	);
	LUT2 #(
		.INIT('h8)
	) name5648 (
		\u5_cmd_del_reg[0]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w6607_
	);
	LUT2 #(
		.INIT('h1)
	) name5649 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1771_,
		_w6608_
	);
	LUT2 #(
		.INIT('h1)
	) name5650 (
		_w6607_,
		_w6608_,
		_w6609_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g22/_0_  = _w1045_ ;
	assign \g23/_0_  = _w1044_ ;
	assign \g25_dup61718/_2_  = _w1049_ ;
	assign \g43466/_0_  = _w1449_ ;
	assign \g43467/_0_  = _w1463_ ;
	assign \g43468/_0_  = _w1475_ ;
	assign \g43469/_0_  = _w1487_ ;
	assign \g43470/_0_  = _w1501_ ;
	assign \g43471/_0_  = _w1515_ ;
	assign \g43472/_0_  = _w1529_ ;
	assign \g43473/_0_  = _w1543_ ;
	assign \g43474/_0_  = _w1557_ ;
	assign \g43475/_0_  = _w1571_ ;
	assign \g43476/_0_  = _w1585_ ;
	assign \g43477/_0_  = _w1599_ ;
	assign \g43478/_0_  = _w1613_ ;
	assign \g43512/_0_  = _w1740_ ;
	assign \g43513/_0_  = _w1741_ ;
	assign \g43544/_3_  = _w1771_ ;
	assign \g43545/_0_  = _w1774_ ;
	assign \g43554/_0_  = _w1862_ ;
	assign \g43555/_0_  = _w2276_ ;
	assign \g43557/_0_  = _w1737_ ;
	assign \g43558/_0_  = _w2319_ ;
	assign \g43571/_2_  = _w2351_ ;
	assign \g43632/_0_  = _w2382_ ;
	assign \g43633/_0_  = _w2392_ ;
	assign \g43635/_0_  = _w2401_ ;
	assign \g43636/_0_  = _w2408_ ;
	assign \g43637/_0_  = _w2410_ ;
	assign \g43638/_0_  = _w2434_ ;
	assign \g43639/_0_  = _w2443_ ;
	assign \g43640/_0_  = _w2452_ ;
	assign \g43642/_0_  = _w1307_ ;
	assign \g43662/_0_  = _w2457_ ;
	assign \g43663/_0_  = _w2459_ ;
	assign \g43664/_0_  = _w2461_ ;
	assign \g43665/_0_  = _w2463_ ;
	assign \g43668/_0_  = _w2495_ ;
	assign \g43670/_0_  = _w2508_ ;
	assign \g43671/_0_  = _w2513_ ;
	assign \g43673/_0_  = _w2557_ ;
	assign \g43674/_0_  = _w2600_ ;
	assign \g43692/_0_  = _w2604_ ;
	assign \g43695/_0_  = _w2610_ ;
	assign \g43696/_0_  = _w2613_ ;
	assign \g43697/_0_  = _w2621_ ;
	assign \g43698/_0_  = _w2631_ ;
	assign \g43700/_0_  = _w2642_ ;
	assign \g43701/_0_  = _w2648_ ;
	assign \g43703/_0_  = _w2658_ ;
	assign \g43705/_0_  = _w2668_ ;
	assign \g43707/_0_  = _w2676_ ;
	assign \g43708/_0_  = _w2691_ ;
	assign \g43710/_0_  = _w2699_ ;
	assign \g43717/_0_  = _w2702_ ;
	assign \g43719/_0_  = _w2704_ ;
	assign \g43720/_0_  = _w2708_ ;
	assign \g43721/_0_  = _w2721_ ;
	assign \g43722/_1_  = _w2728_ ;
	assign \g43723/_0_  = _w2737_ ;
	assign \g43725/_0_  = _w2743_ ;
	assign \g43729/_0_  = _w2744_ ;
	assign \g43731/_0_  = _w2747_ ;
	assign \g43734/_0_  = _w2752_ ;
	assign \g43735/_0_  = _w2755_ ;
	assign \g43737/_0_  = _w2756_ ;
	assign \g43744/_0_  = _w2759_ ;
	assign \g43747/_0_  = _w2762_ ;
	assign \g43760/_2_  = _w2766_ ;
	assign \g43770/_1_  = _w2776_ ;
	assign \g43775/_2_  = _w2780_ ;
	assign \g43780/_2_  = _w2791_ ;
	assign \g43786/_0_  = _w2793_ ;
	assign \g43787/_1_  = _w2800_ ;
	assign \g43847/_0_  = _w2809_ ;
	assign \g43848/_1_  = _w2813_ ;
	assign \g43858/_1_  = _w2817_ ;
	assign \g43891/_3_  = _w2857_ ;
	assign \g43895/_0_  = _w2885_ ;
	assign \g43934/_0_  = _w2904_ ;
	assign \g43936/_3_  = _w2926_ ;
	assign \g43954/_3_  = _w2938_ ;
	assign \g43961/_0_  = _w2966_ ;
	assign \g44016/_1_  = _w2969_ ;
	assign \g44067/_0_  = _w2979_ ;
	assign \g44094/_0_  = _w2989_ ;
	assign \g44096/_0_  = _w3005_ ;
	assign \g44104/_0_  = _w3020_ ;
	assign \g44122/_0_  = _w3030_ ;
	assign \g44172/_0_  = _w2935_ ;
	assign \g44209/_0_  = _w3048_ ;
	assign \g44219/_0_  = _w3102_ ;
	assign \g44220/_0_  = _w3108_ ;
	assign \g44222/_0_  = _w3117_ ;
	assign \g44223/_0_  = _w3122_ ;
	assign \g44241/_2_  = _w3132_ ;
	assign \g44252/_0_  = _w3138_ ;
	assign \g44253/_0_  = _w3143_ ;
	assign \g44255/_2_  = _w3153_ ;
	assign \g44263/_2_  = _w3167_ ;
	assign \g44470/_0_  = _w3177_ ;
	assign \g44538/_0_  = _w3210_ ;
	assign \g44539/_0_  = _w3216_ ;
	assign \g44540/_0_  = _w3222_ ;
	assign \g44541/_0_  = _w3228_ ;
	assign \g44542/_0_  = _w3234_ ;
	assign \g44543/_0_  = _w3240_ ;
	assign \g44544/_0_  = _w3246_ ;
	assign \g44545/_0_  = _w3252_ ;
	assign \g44546/_0_  = _w3258_ ;
	assign \g44547/_0_  = _w3264_ ;
	assign \g44548/_0_  = _w3270_ ;
	assign \g44549/_0_  = _w3276_ ;
	assign \g44550/_0_  = _w3282_ ;
	assign \g44551/_0_  = _w3288_ ;
	assign \g44552/_0_  = _w3294_ ;
	assign \g44553/_0_  = _w3300_ ;
	assign \g44554/_0_  = _w3306_ ;
	assign \g44555/_0_  = _w3312_ ;
	assign \g44556/_0_  = _w3318_ ;
	assign \g44557/_0_  = _w3324_ ;
	assign \g44558/_0_  = _w3330_ ;
	assign \g44559/_0_  = _w3336_ ;
	assign \g44560/_0_  = _w3342_ ;
	assign \g44561/_0_  = _w3348_ ;
	assign \g44562/_0_  = _w3354_ ;
	assign \g44563/_0_  = _w3360_ ;
	assign \g44564/_0_  = _w3366_ ;
	assign \g44565/_0_  = _w3372_ ;
	assign \g44566/_0_  = _w3463_ ;
	assign \g44567/_0_  = _w3469_ ;
	assign \g44568/_0_  = _w3475_ ;
	assign \g44569/_0_  = _w3481_ ;
	assign \g44570/_0_  = _w3487_ ;
	assign \g44571/_0_  = _w3493_ ;
	assign \g44572/_0_  = _w3499_ ;
	assign \g44573/_0_  = _w3505_ ;
	assign \g44574/_0_  = _w3511_ ;
	assign \g44575/_0_  = _w3517_ ;
	assign \g44576/_0_  = _w3523_ ;
	assign \g44577/_0_  = _w3529_ ;
	assign \g44578/_0_  = _w3535_ ;
	assign \g44579/_0_  = _w3541_ ;
	assign \g44580/_0_  = _w3547_ ;
	assign \g44581/_0_  = _w3553_ ;
	assign \g44582/_0_  = _w3559_ ;
	assign \g44583/_0_  = _w3565_ ;
	assign \g44584/_0_  = _w3571_ ;
	assign \g44585/_0_  = _w3577_ ;
	assign \g44586/_0_  = _w3583_ ;
	assign \g44588/_0_  = _w3589_ ;
	assign \g44589/_0_  = _w3595_ ;
	assign \g44590/_0_  = _w3601_ ;
	assign \g44591/_0_  = _w3607_ ;
	assign \g44592/_0_  = _w3613_ ;
	assign \g44593/_0_  = _w3619_ ;
	assign \g44594/_0_  = _w3625_ ;
	assign \g44595/_0_  = _w3638_ ;
	assign \g44596/_0_  = _w3649_ ;
	assign \g44636/_2_  = _w3659_ ;
	assign \g44646/_0_  = _w3667_ ;
	assign \g44647/_0_  = _w3673_ ;
	assign \g44648/_0_  = _w3679_ ;
	assign \g44649/_0_  = _w3685_ ;
	assign \g44650/_0_  = _w3691_ ;
	assign \g44651/_0_  = _w3698_ ;
	assign \g44652/_0_  = _w3703_ ;
	assign \g44653/_0_  = _w3708_ ;
	assign \g44654/_0_  = _w3713_ ;
	assign \g44655/_0_  = _w3718_ ;
	assign \g44656/_0_  = _w3723_ ;
	assign \g44657/_0_  = _w3728_ ;
	assign \g44665/_0_  = _w3731_ ;
	assign \g44666/_0_  = _w3737_ ;
	assign \g44667/_0_  = _w3743_ ;
	assign \g44668/_0_  = _w3749_ ;
	assign \g44752/_0_  = _w3759_ ;
	assign \g44753/_0_  = _w3766_ ;
	assign \g44873/_0_  = _w1432_ ;
	assign \g44939/_0_  = _w3774_ ;
	assign \g44942/_0_  = _w3779_ ;
	assign \g44945/_0_  = _w3785_ ;
	assign \g45023/_2_  = _w3795_ ;
	assign \g45090/_0_  = _w3660_ ;
	assign \g45141/_0_  = _w3804_ ;
	assign \g45147/_3_  = _w3813_ ;
	assign \g45155/_0_  = _w3823_ ;
	assign \g45190/_0_  = _w3825_ ;
	assign \g45195/_2_  = _w3835_ ;
	assign \g45199/_2_  = _w3846_ ;
	assign \g45201/_2_  = _w3856_ ;
	assign \g45324/_0_  = _w3868_ ;
	assign \g45334/_2_  = _w3879_ ;
	assign \g45336/_0_  = _w3811_ ;
	assign \g45388/_0_  = _w3885_ ;
	assign \g45391/_0_  = _w3904_ ;
	assign \g45413/_2_  = _w3914_ ;
	assign \g45530/_0_  = _w3922_ ;
	assign \g45532/_0_  = _w3929_ ;
	assign \g45533/_0_  = _w3940_ ;
	assign \g45534/_0_  = _w3950_ ;
	assign \g45739/_2_  = _w3961_ ;
	assign \g45743/_2_  = _w3972_ ;
	assign \g45767/_0_  = _w4000_ ;
	assign \g45782/_0_  = _w4013_ ;
	assign \g45830/_3_  = _w4039_ ;
	assign \g45834/_3_  = _w4061_ ;
	assign \g45835/_3_  = _w4071_ ;
	assign \g45836/_3_  = _w4085_ ;
	assign \g45837/_3_  = _w4094_ ;
	assign \g45839/_3_  = _w4103_ ;
	assign \g45840/_3_  = _w4112_ ;
	assign \g45841/_3_  = _w4121_ ;
	assign \g45842/_3_  = _w4130_ ;
	assign \g45843/_3_  = _w4138_ ;
	assign \g45844/_3_  = _w4141_ ;
	assign \g45845/_3_  = _w4144_ ;
	assign \g46191/_0_  = _w1640_ ;
	assign \g46193/_3_  = _w4150_ ;
	assign \g46256/_3_  = _w4160_ ;
	assign \g46257/_3_  = _w4166_ ;
	assign \g46258/_3_  = _w4172_ ;
	assign \g46259/_3_  = _w4178_ ;
	assign \g46260/_3_  = _w4184_ ;
	assign \g46261/_3_  = _w4190_ ;
	assign \g46262/_3_  = _w4196_ ;
	assign \g46263/_3_  = _w4202_ ;
	assign \g46278/_0_  = _w4206_ ;
	assign \g46292/_0_  = _w4210_ ;
	assign \g46293/_0_  = _w4214_ ;
	assign \g46312/_0_  = _w4223_ ;
	assign \g46367/_2_  = _w4234_ ;
	assign \g46370/_2_  = _w4243_ ;
	assign \g46380/_2_  = _w4254_ ;
	assign \g46386/_2_  = _w4265_ ;
	assign \g46388/_2_  = _w4276_ ;
	assign \g46392/_2_  = _w4287_ ;
	assign \g46395/_2_  = _w4298_ ;
	assign \g46399/_2_  = _w4307_ ;
	assign \g46420/_0_  = _w4309_ ;
	assign \g46446/_0_  = _w4313_ ;
	assign \g46493/_0_  = _w4321_ ;
	assign \g46510/_0_  = _w4323_ ;
	assign \g46669/_2_  = _w4330_ ;
	assign \g46691/_0_  = _w4377_ ;
	assign \g46708/_0_  = _w4382_ ;
	assign \g46721/_00_  = _w4403_ ;
	assign \g46776/_0_  = _w4406_ ;
	assign \g46777/_0_  = _w4410_ ;
	assign \g46778/_0_  = _w4414_ ;
	assign \g46779/_0_  = _w4418_ ;
	assign \g46780/_0_  = _w4422_ ;
	assign \g46782/_0_  = _w4426_ ;
	assign \g46784/_0_  = _w4430_ ;
	assign \g46932/_0_  = _w4439_ ;
	assign \g47112/_0_  = _w4446_ ;
	assign \g47124/_0_  = _w4449_ ;
	assign \g47265/_0_  = _w4456_ ;
	assign \g47270/_0_  = _w4462_ ;
	assign \g47275/_0_  = _w4469_ ;
	assign \g47300/_1_  = _w4208_ ;
	assign \g47305/_1_  = _w4212_ ;
	assign \g47338/_0_  = _w4472_ ;
	assign \g47339/_0_  = _w4475_ ;
	assign \g47352/_0_  = _w4901_ ;
	assign \g47699/_3_  = _w4905_ ;
	assign \g47711/_0_  = _w4910_ ;
	assign \g47719/_3_  = _w4913_ ;
	assign \g47721/_3_  = _w4916_ ;
	assign \g47723/_3_  = _w4919_ ;
	assign \g47853/_0_  = _w4922_ ;
	assign \g48094/_0_  = _w4930_ ;
	assign \g48095/_0_  = _w4938_ ;
	assign \g48177/_2_  = _w4942_ ;
	assign \g48194/_0_  = _w4444_ ;
	assign \g48369/_2_  = _w4948_ ;
	assign \g48371/_2_  = _w4954_ ;
	assign \g48373/_2_  = _w4960_ ;
	assign \g48375/_2_  = _w4966_ ;
	assign \g48377/_2_  = _w4972_ ;
	assign \g48379/_2_  = _w4978_ ;
	assign \g48381/_2_  = _w4984_ ;
	assign \g48383/_2_  = _w4990_ ;
	assign \g48385/_2_  = _w4996_ ;
	assign \g48535/_0_  = _w4998_ ;
	assign \g48569/_0_  = _w5001_ ;
	assign \g48570/_0_  = _w5004_ ;
	assign \g48571/_0_  = _w5007_ ;
	assign \g48836/_0_  = _w5010_ ;
	assign \g48843/_0_  = _w5013_ ;
	assign \g49187/_3_  = _w4011_ ;
	assign \g49375/_2_  = _w5014_ ;
	assign \g49633/_0_  = _w5016_ ;
	assign \g49788/_1_  = _w3118_ ;
	assign \g49800/_1_  = _w3110_ ;
	assign \g49802/_1_  = _w3139_ ;
	assign \g49806/_1_  = _w3052_ ;
	assign \g49853/_1_  = _w3134_ ;
	assign \g49883/_0_  = _w5021_ ;
	assign \g49884/_0_  = _w5025_ ;
	assign \g49885/_0_  = _w5029_ ;
	assign \g49886/_0_  = _w5033_ ;
	assign \g49976/_1_  = _w3104_ ;
	assign \g50038/_0_  = _w5050_ ;
	assign \g50082/_0_  = _w5063_ ;
	assign \g50083/_0_  = _w4375_ ;
	assign \g50167/_3_  = _w5099_ ;
	assign \g50168/_3_  = _w5121_ ;
	assign \g50169/_3_  = _w5143_ ;
	assign \g50170/_3_  = _w5165_ ;
	assign \g50171/_3_  = _w5187_ ;
	assign \g50177/_0_  = _w5194_ ;
	assign \g50190/_0_  = _w5200_ ;
	assign \g50236/_0_  = _w3415_ ;
	assign \g50251/_3_  = _w5222_ ;
	assign \g50256/_0_  = _w3457_ ;
	assign \g50318/_3_  = _w5244_ ;
	assign \g50319/_3_  = _w5266_ ;
	assign \g50350/_3_  = _w5289_ ;
	assign \g50351/_3_  = _w5311_ ;
	assign \g50352/_3_  = _w5333_ ;
	assign \g50353/_3_  = _w5355_ ;
	assign \g50354/_3_  = _w5377_ ;
	assign \g50355/_3_  = _w5399_ ;
	assign \g50361/_2_  = _w5400_ ;
	assign \g50366/_0_  = _w5410_ ;
	assign \g50393/_0_  = _w5412_ ;
	assign \g50552/_1_  = _w1784_ ;
	assign \g51108/_0_  = _w5418_ ;
	assign \g51160/_0_  = _w5423_ ;
	assign \g51290/_1_  = _w5424_ ;
	assign \g51327/_3_  = _w5444_ ;
	assign \g51328/_3_  = _w5464_ ;
	assign \g51329/_3_  = _w5484_ ;
	assign \g51330/_3_  = _w5504_ ;
	assign \g51331/_3_  = _w5524_ ;
	assign \g51332/_3_  = _w5544_ ;
	assign \g51333/_3_  = _w5564_ ;
	assign \g51334/_3_  = _w5584_ ;
	assign \g51339/_3_  = _w5602_ ;
	assign \g51340/_3_  = _w5620_ ;
	assign \g51341/_3_  = _w5638_ ;
	assign \g51342/_3_  = _w5656_ ;
	assign \g51343/_3_  = _w5674_ ;
	assign \g51346/_0_  = _w5679_ ;
	assign \g51347/_0_  = _w5684_ ;
	assign \g51348/_0_  = _w5686_ ;
	assign \g51381/_3_  = _w5708_ ;
	assign \g51382/_3_  = _w5730_ ;
	assign \g51383/_3_  = _w5752_ ;
	assign \g51386/_3_  = _w5774_ ;
	assign \g51387/_3_  = _w5796_ ;
	assign \g51405/_3_  = _w5802_ ;
	assign \g51410/_3_  = _w5808_ ;
	assign \g51883/_0_  = _w5809_ ;
	assign \g51916/_0_  = _w4367_ ;
	assign \g51947/_0_  = _w5813_ ;
	assign \g51948/_0_  = _w5817_ ;
	assign \g51949/_0_  = _w5824_ ;
	assign \g51950/_0_  = _w5828_ ;
	assign \g51951/_0_  = _w5832_ ;
	assign \g51952/_0_  = _w5836_ ;
	assign \g51953/_0_  = _w5840_ ;
	assign \g51954/_0_  = _w5844_ ;
	assign \g51955/_0_  = _w5848_ ;
	assign \g51956/_0_  = _w5852_ ;
	assign \g51957/_0_  = _w5856_ ;
	assign \g51958/_0_  = _w5860_ ;
	assign \g51959/_0_  = _w5864_ ;
	assign \g51960/_0_  = _w5868_ ;
	assign \g51961/_0_  = _w5872_ ;
	assign \g51962/_0_  = _w5876_ ;
	assign \g51963/_0_  = _w5880_ ;
	assign \g51964/_0_  = _w5884_ ;
	assign \g51965/_0_  = _w5888_ ;
	assign \g51967/_0_  = _w5892_ ;
	assign \g51968/_0_  = _w5897_ ;
	assign \g51969/_0_  = _w5901_ ;
	assign \g51970/_0_  = _w5905_ ;
	assign \g51971/_0_  = _w5909_ ;
	assign \g51972/_0_  = _w5913_ ;
	assign \g51973/_0_  = _w5917_ ;
	assign \g51974/_0_  = _w5921_ ;
	assign \g51975/_0_  = _w5925_ ;
	assign \g51976/_0_  = _w5929_ ;
	assign \g51977/_0_  = _w5933_ ;
	assign \g51978/_0_  = _w5937_ ;
	assign \g51979/_0_  = _w5941_ ;
	assign \g51980/_0_  = _w5945_ ;
	assign \g51981/_0_  = _w5949_ ;
	assign \g51982/_0_  = _w5953_ ;
	assign \g51983/_0_  = _w5957_ ;
	assign \g51984/_0_  = _w5961_ ;
	assign \g51985/_0_  = _w5965_ ;
	assign \g51986/_0_  = _w5969_ ;
	assign \g51987/_0_  = _w5973_ ;
	assign \g51988/_0_  = _w5977_ ;
	assign \g51989/_0_  = _w5981_ ;
	assign \g51990/_0_  = _w5985_ ;
	assign \g51991/_0_  = _w5989_ ;
	assign \g51992/_0_  = _w5993_ ;
	assign \g51993/_0_  = _w5997_ ;
	assign \g51994/_0_  = _w6001_ ;
	assign \g51995/_0_  = _w6005_ ;
	assign \g51996/_0_  = _w6009_ ;
	assign \g51997/_0_  = _w6013_ ;
	assign \g51998/_0_  = _w6017_ ;
	assign \g51999/_0_  = _w6021_ ;
	assign \g52000/_0_  = _w6026_ ;
	assign \g52001/_0_  = _w6030_ ;
	assign \g52002/_0_  = _w6034_ ;
	assign \g52003/_0_  = _w6038_ ;
	assign \g52004/_0_  = _w6042_ ;
	assign \g52005/_0_  = _w6046_ ;
	assign \g52006/_0_  = _w6050_ ;
	assign \g52007/_0_  = _w6054_ ;
	assign \g52008/_0_  = _w6058_ ;
	assign \g52009/_0_  = _w6062_ ;
	assign \g52010/_0_  = _w6066_ ;
	assign \g52011/_0_  = _w6070_ ;
	assign \g52012/_0_  = _w6074_ ;
	assign \g52013/_0_  = _w6078_ ;
	assign \g52014/_0_  = _w6082_ ;
	assign \g52015/_0_  = _w6086_ ;
	assign \g52016/_0_  = _w6090_ ;
	assign \g52017/_0_  = _w6094_ ;
	assign \g52018/_0_  = _w6098_ ;
	assign \g52019/_0_  = _w6102_ ;
	assign \g52020/_0_  = _w6106_ ;
	assign \g52021/_0_  = _w6110_ ;
	assign \g52022/_0_  = _w6114_ ;
	assign \g52023/_0_  = _w6118_ ;
	assign \g52024/_0_  = _w6122_ ;
	assign \g52025/_0_  = _w6126_ ;
	assign \g52026/_0_  = _w6130_ ;
	assign \g52027/_0_  = _w6134_ ;
	assign \g52028/_0_  = _w6138_ ;
	assign \g52029/_0_  = _w6142_ ;
	assign \g52030/_0_  = _w6146_ ;
	assign \g52031/_0_  = _w6150_ ;
	assign \g52032/_0_  = _w6154_ ;
	assign \g52033/_0_  = _w6158_ ;
	assign \g52034/_0_  = _w6162_ ;
	assign \g52035/_0_  = _w6166_ ;
	assign \g52036/_0_  = _w6170_ ;
	assign \g52037/_0_  = _w6174_ ;
	assign \g52038/_0_  = _w6178_ ;
	assign \g52039/_0_  = _w6182_ ;
	assign \g52040/_0_  = _w6186_ ;
	assign \g52041/_0_  = _w6190_ ;
	assign \g52042/_0_  = _w6194_ ;
	assign \g52043/_0_  = _w6198_ ;
	assign \g52044/_0_  = _w6202_ ;
	assign \g52045/_0_  = _w6206_ ;
	assign \g52046/_0_  = _w6210_ ;
	assign \g52047/_0_  = _w6214_ ;
	assign \g52049/_0_  = _w6218_ ;
	assign \g52050/_0_  = _w6222_ ;
	assign \g52051/_0_  = _w6226_ ;
	assign \g52052/_0_  = _w6230_ ;
	assign \g52053/_0_  = _w6234_ ;
	assign \g52054/_0_  = _w6238_ ;
	assign \g52055/_0_  = _w6242_ ;
	assign \g52056/_0_  = _w6246_ ;
	assign \g52057/_0_  = _w6250_ ;
	assign \g52058/_0_  = _w6254_ ;
	assign \g52061/_0_  = _w6258_ ;
	assign \g52065/_0_  = _w6262_ ;
	assign \g52066/_0_  = _w6266_ ;
	assign \g52067/_0_  = _w6270_ ;
	assign \g52068/_0_  = _w6274_ ;
	assign \g52069/_0_  = _w6278_ ;
	assign \g52070/_0_  = _w6282_ ;
	assign \g52071/_0_  = _w6286_ ;
	assign \g52073/_0_  = _w6290_ ;
	assign \g52074/_0_  = _w6294_ ;
	assign \g52075/_0_  = _w6298_ ;
	assign \g52082/_0_  = _w6302_ ;
	assign \g52083/_0_  = _w6306_ ;
	assign \g52158/_0_  = _w6308_ ;
	assign \g52201/_0_  = _w6309_ ;
	assign \g52202/_0_  = _w6310_ ;
	assign \g52346/_0_  = _w1827_ ;
	assign \g52351/_0_  = _w6312_ ;
	assign \g52390/_0_  = _w6315_ ;
	assign \g52847/_0_  = _w2806_ ;
	assign \g52854/_0_  = _w6317_ ;
	assign \g52968/_0_  = _w6338_ ;
	assign \g52969/_0_  = _w6359_ ;
	assign \g52970/_0_  = _w6380_ ;
	assign \g52971/_0_  = _w6401_ ;
	assign \g52984/_0_  = _w6404_ ;
	assign \g52994/_0_  = _w4466_ ;
	assign \g53019/_0_  = _w5893_ ;
	assign \g53030/_0_  = _w5820_ ;
	assign \g53094/_1_  = _w5057_ ;
	assign \g53106/_0_  = _w6022_ ;
	assign \g53150/_0_  = _w6415_ ;
	assign \g53256/_0_  = _w6417_ ;
	assign \g53297/_0_  = _w6419_ ;
	assign \g53345/_0_  = _w6420_ ;
	assign \g53359/_0_  = _w6422_ ;
	assign \g53375/_0_  = _w6423_ ;
	assign \g53474/_1__syn_2  = _w6426_ ;
	assign \g53475/_2_  = _w6427_ ;
	assign \g53593/_0_  = _w6429_ ;
	assign \g53643/_1_  = _w6431_ ;
	assign \g53655/_0_  = _w1050_ ;
	assign \g53710/_0_  = _w6432_ ;
	assign \g53786/_0_  = _w6434_ ;
	assign \g53837/_0_  = _w6436_ ;
	assign \g53888/_1_  = _w4431_ ;
	assign \g53909/_0_  = _w1196_ ;
	assign \g54253/_2_  = _w6438_ ;
	assign \g54394/_3_  = _w4316_ ;
	assign \g54413/_0_  = _w6441_ ;
	assign \g55420/_0_  = _w6442_ ;
	assign \g55587/_0_  = _w6443_ ;
	assign \g55852/_0_  = \u5_mc_le_reg/NET0131 ;
	assign \g57020/_0_  = \u1_acs_addr_reg[0]/P0001 ;
	assign \g59450/_0_  = _w6485_ ;
	assign \g59488/_2_  = _w1325_ ;
	assign \g59752/_0_  = _w6489_ ;
	assign \g59786/_0_  = _w6492_ ;
	assign \g59854/_0_  = _w6494_ ;
	assign \g59878/_0_  = _w6496_ ;
	assign \g59902/_0_  = _w6501_ ;
	assign \g59924/_0_  = _w6505_ ;
	assign \g59947/_0_  = _w6512_ ;
	assign \g59972/_0_  = _w6518_ ;
	assign \g59996/_0_  = _w6521_ ;
	assign \g60017/_0_  = _w6525_ ;
	assign \g60040/_0_  = _w6529_ ;
	assign \g60064/_0_  = _w6531_ ;
	assign \g60095/_0_  = _w6533_ ;
	assign \g60119/_0_  = _w6535_ ;
	assign \g60145/_1_  = _w6547_ ;
	assign \g60165/_0_  = _w6551_ ;
	assign \g60407/_2_  = _w1382_ ;
	assign \g60408/_0_  = _w6552_ ;
	assign \g60613/_2_  = _w6554_ ;
	assign \g60649/_0_  = _w1896_ ;
	assign \g60771/_0_  = _w6555_ ;
	assign \g60908/_1_  = _w6559_ ;
	assign \g60911/_0_  = _w6561_ ;
	assign \g60977/_0_  = _w3201_ ;
	assign \g61/_0_  = _w1198_ ;
	assign \g61002/_0_  = _w6564_ ;
	assign \g61308/_0_  = _w6569_ ;
	assign \g61312/_1_  = _w6565_ ;
	assign \g61314/_0_  = _w6574_ ;
	assign \g61319/_1_  = _w6570_ ;
	assign \g61342/_1_  = _w1328_ ;
	assign \g61360/_0_  = _w6577_ ;
	assign \g61377/_0_  = _w6578_ ;
	assign \g61423/_1_  = _w1629_ ;
	assign \g61426/_0_  = _w1628_ ;
	assign \g61479/_1_  = _w6585_ ;
	assign \g61523/_1_  = _w6586_ ;
	assign \g61558/_1_  = _w2822_ ;
	assign \g61652/_0_  = _w6590_ ;
	assign \g61866/_0_  = _w6594_ ;
	assign \g61868/_1_  = _w6592_ ;
	assign \g61887/_0_  = _w1653_ ;
	assign \u7_mc_dqm_r_reg[0]/P0001_reg_syn_3  = _w6597_ ;
	assign \u7_mc_dqm_r_reg[1]/P0001_reg_syn_3  = _w6600_ ;
	assign \u7_mc_dqm_r_reg[2]/P0001_reg_syn_3  = _w6603_ ;
	assign \u7_mc_dqm_r_reg[3]/P0001_reg_syn_3  = _w6606_ ;
	assign \u7_mc_we__reg/_05_  = _w6609_ ;
endmodule;