module top( \P1_B_reg/NET0131  , \P1_IR_reg[0]/NET0131  , \P1_IR_reg[10]/NET0131  , \P1_IR_reg[11]/NET0131  , \P1_IR_reg[12]/NET0131  , \P1_IR_reg[13]/NET0131  , \P1_IR_reg[14]/NET0131  , \P1_IR_reg[15]/NET0131  , \P1_IR_reg[16]/NET0131  , \P1_IR_reg[17]/NET0131  , \P1_IR_reg[18]/NET0131  , \P1_IR_reg[19]/NET0131  , \P1_IR_reg[1]/NET0131  , \P1_IR_reg[20]/NET0131  , \P1_IR_reg[21]/NET0131  , \P1_IR_reg[22]/NET0131  , \P1_IR_reg[23]/NET0131  , \P1_IR_reg[24]/NET0131  , \P1_IR_reg[25]/NET0131  , \P1_IR_reg[26]/NET0131  , \P1_IR_reg[27]/NET0131  , \P1_IR_reg[28]/NET0131  , \P1_IR_reg[29]/NET0131  , \P1_IR_reg[2]/NET0131  , \P1_IR_reg[30]/NET0131  , \P1_IR_reg[31]/NET0131  , \P1_IR_reg[3]/NET0131  , \P1_IR_reg[4]/NET0131  , \P1_IR_reg[5]/NET0131  , \P1_IR_reg[6]/NET0131  , \P1_IR_reg[7]/NET0131  , \P1_IR_reg[8]/NET0131  , \P1_IR_reg[9]/NET0131  , \P1_addr_reg[0]/NET0131  , \P1_addr_reg[10]/NET0131  , \P1_addr_reg[11]/NET0131  , \P1_addr_reg[12]/NET0131  , \P1_addr_reg[13]/NET0131  , \P1_addr_reg[14]/NET0131  , \P1_addr_reg[15]/NET0131  , \P1_addr_reg[16]/NET0131  , \P1_addr_reg[17]/NET0131  , \P1_addr_reg[18]/NET0131  , \P1_addr_reg[19]/NET0131  , \P1_addr_reg[1]/NET0131  , \P1_addr_reg[2]/NET0131  , \P1_addr_reg[3]/NET0131  , \P1_addr_reg[4]/NET0131  , \P1_addr_reg[5]/NET0131  , \P1_addr_reg[6]/NET0131  , \P1_addr_reg[7]/NET0131  , \P1_addr_reg[8]/NET0131  , \P1_addr_reg[9]/NET0131  , \P1_d_reg[0]/NET0131  , \P1_d_reg[1]/NET0131  , \P1_datao_reg[0]/NET0131  , \P1_datao_reg[10]/NET0131  , \P1_datao_reg[11]/NET0131  , \P1_datao_reg[12]/NET0131  , \P1_datao_reg[13]/NET0131  , \P1_datao_reg[14]/NET0131  , \P1_datao_reg[15]/NET0131  , \P1_datao_reg[16]/NET0131  , \P1_datao_reg[17]/NET0131  , \P1_datao_reg[18]/NET0131  , \P1_datao_reg[19]/NET0131  , \P1_datao_reg[1]/NET0131  , \P1_datao_reg[20]/NET0131  , \P1_datao_reg[21]/NET0131  , \P1_datao_reg[22]/NET0131  , \P1_datao_reg[23]/NET0131  , \P1_datao_reg[24]/NET0131  , \P1_datao_reg[25]/NET0131  , \P1_datao_reg[26]/NET0131  , \P1_datao_reg[27]/NET0131  , \P1_datao_reg[28]/NET0131  , \P1_datao_reg[29]/NET0131  , \P1_datao_reg[2]/NET0131  , \P1_datao_reg[30]/NET0131  , \P1_datao_reg[31]/NET0131  , \P1_datao_reg[3]/NET0131  , \P1_datao_reg[4]/NET0131  , \P1_datao_reg[5]/NET0131  , \P1_datao_reg[6]/NET0131  , \P1_datao_reg[7]/NET0131  , \P1_datao_reg[8]/NET0131  , \P1_datao_reg[9]/NET0131  , \P1_rd_reg/NET0131  , \P1_reg0_reg[0]/NET0131  , \P1_reg0_reg[10]/NET0131  , \P1_reg0_reg[11]/NET0131  , \P1_reg0_reg[12]/NET0131  , \P1_reg0_reg[13]/NET0131  , \P1_reg0_reg[14]/NET0131  , \P1_reg0_reg[15]/NET0131  , \P1_reg0_reg[16]/NET0131  , \P1_reg0_reg[17]/NET0131  , \P1_reg0_reg[18]/NET0131  , \P1_reg0_reg[19]/NET0131  , \P1_reg0_reg[1]/NET0131  , \P1_reg0_reg[20]/NET0131  , \P1_reg0_reg[21]/NET0131  , \P1_reg0_reg[22]/NET0131  , \P1_reg0_reg[23]/NET0131  , \P1_reg0_reg[24]/NET0131  , \P1_reg0_reg[25]/NET0131  , \P1_reg0_reg[26]/NET0131  , \P1_reg0_reg[27]/NET0131  , \P1_reg0_reg[28]/NET0131  , \P1_reg0_reg[29]/NET0131  , \P1_reg0_reg[2]/NET0131  , \P1_reg0_reg[30]/NET0131  , \P1_reg0_reg[31]/NET0131  , \P1_reg0_reg[3]/NET0131  , \P1_reg0_reg[4]/NET0131  , \P1_reg0_reg[5]/NET0131  , \P1_reg0_reg[6]/NET0131  , \P1_reg0_reg[7]/NET0131  , \P1_reg0_reg[8]/NET0131  , \P1_reg0_reg[9]/NET0131  , \P1_reg1_reg[0]/NET0131  , \P1_reg1_reg[10]/NET0131  , \P1_reg1_reg[11]/NET0131  , \P1_reg1_reg[12]/NET0131  , \P1_reg1_reg[13]/NET0131  , \P1_reg1_reg[14]/NET0131  , \P1_reg1_reg[15]/NET0131  , \P1_reg1_reg[16]/NET0131  , \P1_reg1_reg[17]/NET0131  , \P1_reg1_reg[18]/NET0131  , \P1_reg1_reg[19]/NET0131  , \P1_reg1_reg[1]/NET0131  , \P1_reg1_reg[20]/NET0131  , \P1_reg1_reg[21]/NET0131  , \P1_reg1_reg[22]/NET0131  , \P1_reg1_reg[23]/NET0131  , \P1_reg1_reg[24]/NET0131  , \P1_reg1_reg[25]/NET0131  , \P1_reg1_reg[26]/NET0131  , \P1_reg1_reg[27]/NET0131  , \P1_reg1_reg[28]/NET0131  , \P1_reg1_reg[29]/NET0131  , \P1_reg1_reg[2]/NET0131  , \P1_reg1_reg[30]/NET0131  , \P1_reg1_reg[31]/NET0131  , \P1_reg1_reg[3]/NET0131  , \P1_reg1_reg[4]/NET0131  , \P1_reg1_reg[5]/NET0131  , \P1_reg1_reg[6]/NET0131  , \P1_reg1_reg[7]/NET0131  , \P1_reg1_reg[8]/NET0131  , \P1_reg1_reg[9]/NET0131  , \P1_reg2_reg[0]/NET0131  , \P1_reg2_reg[10]/NET0131  , \P1_reg2_reg[11]/NET0131  , \P1_reg2_reg[12]/NET0131  , \P1_reg2_reg[13]/NET0131  , \P1_reg2_reg[14]/NET0131  , \P1_reg2_reg[15]/NET0131  , \P1_reg2_reg[16]/NET0131  , \P1_reg2_reg[17]/NET0131  , \P1_reg2_reg[18]/NET0131  , \P1_reg2_reg[19]/NET0131  , \P1_reg2_reg[1]/NET0131  , \P1_reg2_reg[20]/NET0131  , \P1_reg2_reg[21]/NET0131  , \P1_reg2_reg[22]/NET0131  , \P1_reg2_reg[23]/NET0131  , \P1_reg2_reg[24]/NET0131  , \P1_reg2_reg[25]/NET0131  , \P1_reg2_reg[26]/NET0131  , \P1_reg2_reg[27]/NET0131  , \P1_reg2_reg[28]/NET0131  , \P1_reg2_reg[29]/NET0131  , \P1_reg2_reg[2]/NET0131  , \P1_reg2_reg[30]/NET0131  , \P1_reg2_reg[31]/NET0131  , \P1_reg2_reg[3]/NET0131  , \P1_reg2_reg[4]/NET0131  , \P1_reg2_reg[5]/NET0131  , \P1_reg2_reg[6]/NET0131  , \P1_reg2_reg[7]/NET0131  , \P1_reg2_reg[8]/NET0131  , \P1_reg2_reg[9]/NET0131  , \P1_reg3_reg[0]/NET0131  , \P1_reg3_reg[10]/NET0131  , \P1_reg3_reg[11]/NET0131  , \P1_reg3_reg[12]/NET0131  , \P1_reg3_reg[13]/NET0131  , \P1_reg3_reg[14]/NET0131  , \P1_reg3_reg[15]/NET0131  , \P1_reg3_reg[16]/NET0131  , \P1_reg3_reg[17]/NET0131  , \P1_reg3_reg[18]/NET0131  , \P1_reg3_reg[19]/NET0131  , \P1_reg3_reg[1]/NET0131  , \P1_reg3_reg[20]/NET0131  , \P1_reg3_reg[21]/NET0131  , \P1_reg3_reg[22]/NET0131  , \P1_reg3_reg[23]/NET0131  , \P1_reg3_reg[24]/NET0131  , \P1_reg3_reg[25]/NET0131  , \P1_reg3_reg[26]/NET0131  , \P1_reg3_reg[27]/NET0131  , \P1_reg3_reg[28]/NET0131  , \P1_reg3_reg[2]/NET0131  , \P1_reg3_reg[3]/NET0131  , \P1_reg3_reg[4]/NET0131  , \P1_reg3_reg[5]/NET0131  , \P1_reg3_reg[6]/NET0131  , \P1_reg3_reg[7]/NET0131  , \P1_reg3_reg[8]/NET0131  , \P1_reg3_reg[9]/NET0131  , \P1_state_reg[0]/NET0131  , \P1_wr_reg/NET0131  , \P2_B_reg/NET0131  , \P2_IR_reg[0]/NET0131  , \P2_IR_reg[10]/NET0131  , \P2_IR_reg[11]/NET0131  , \P2_IR_reg[12]/NET0131  , \P2_IR_reg[13]/NET0131  , \P2_IR_reg[14]/NET0131  , \P2_IR_reg[15]/NET0131  , \P2_IR_reg[16]/NET0131  , \P2_IR_reg[17]/NET0131  , \P2_IR_reg[18]/NET0131  , \P2_IR_reg[19]/NET0131  , \P2_IR_reg[1]/NET0131  , \P2_IR_reg[20]/NET0131  , \P2_IR_reg[21]/NET0131  , \P2_IR_reg[22]/NET0131  , \P2_IR_reg[23]/NET0131  , \P2_IR_reg[24]/NET0131  , \P2_IR_reg[25]/NET0131  , \P2_IR_reg[26]/NET0131  , \P2_IR_reg[27]/NET0131  , \P2_IR_reg[28]/NET0131  , \P2_IR_reg[29]/NET0131  , \P2_IR_reg[2]/NET0131  , \P2_IR_reg[30]/NET0131  , \P2_IR_reg[31]/NET0131  , \P2_IR_reg[3]/NET0131  , \P2_IR_reg[4]/NET0131  , \P2_IR_reg[5]/NET0131  , \P2_IR_reg[6]/NET0131  , \P2_IR_reg[7]/NET0131  , \P2_IR_reg[8]/NET0131  , \P2_IR_reg[9]/NET0131  , \P2_addr_reg[0]/NET0131  , \P2_addr_reg[10]/NET0131  , \P2_addr_reg[11]/NET0131  , \P2_addr_reg[12]/NET0131  , \P2_addr_reg[13]/NET0131  , \P2_addr_reg[14]/NET0131  , \P2_addr_reg[15]/NET0131  , \P2_addr_reg[16]/NET0131  , \P2_addr_reg[17]/NET0131  , \P2_addr_reg[18]/NET0131  , \P2_addr_reg[19]/NET0131  , \P2_addr_reg[1]/NET0131  , \P2_addr_reg[2]/NET0131  , \P2_addr_reg[3]/NET0131  , \P2_addr_reg[4]/NET0131  , \P2_addr_reg[5]/NET0131  , \P2_addr_reg[6]/NET0131  , \P2_addr_reg[7]/NET0131  , \P2_addr_reg[8]/NET0131  , \P2_addr_reg[9]/NET0131  , \P2_d_reg[0]/NET0131  , \P2_d_reg[1]/NET0131  , \P2_datao_reg[0]/NET0131  , \P2_datao_reg[10]/NET0131  , \P2_datao_reg[11]/NET0131  , \P2_datao_reg[12]/NET0131  , \P2_datao_reg[13]/NET0131  , \P2_datao_reg[14]/NET0131  , \P2_datao_reg[15]/NET0131  , \P2_datao_reg[16]/NET0131  , \P2_datao_reg[17]/NET0131  , \P2_datao_reg[18]/NET0131  , \P2_datao_reg[19]/NET0131  , \P2_datao_reg[1]/NET0131  , \P2_datao_reg[20]/NET0131  , \P2_datao_reg[21]/NET0131  , \P2_datao_reg[22]/NET0131  , \P2_datao_reg[23]/NET0131  , \P2_datao_reg[24]/NET0131  , \P2_datao_reg[25]/NET0131  , \P2_datao_reg[26]/NET0131  , \P2_datao_reg[27]/NET0131  , \P2_datao_reg[28]/NET0131  , \P2_datao_reg[29]/NET0131  , \P2_datao_reg[2]/NET0131  , \P2_datao_reg[30]/NET0131  , \P2_datao_reg[31]/NET0131  , \P2_datao_reg[3]/NET0131  , \P2_datao_reg[4]/NET0131  , \P2_datao_reg[5]/NET0131  , \P2_datao_reg[6]/NET0131  , \P2_datao_reg[7]/NET0131  , \P2_datao_reg[8]/NET0131  , \P2_datao_reg[9]/NET0131  , \P2_rd_reg/NET0131  , \P2_reg0_reg[0]/NET0131  , \P2_reg0_reg[10]/NET0131  , \P2_reg0_reg[11]/NET0131  , \P2_reg0_reg[12]/NET0131  , \P2_reg0_reg[13]/NET0131  , \P2_reg0_reg[14]/NET0131  , \P2_reg0_reg[15]/NET0131  , \P2_reg0_reg[16]/NET0131  , \P2_reg0_reg[17]/NET0131  , \P2_reg0_reg[18]/NET0131  , \P2_reg0_reg[19]/NET0131  , \P2_reg0_reg[1]/NET0131  , \P2_reg0_reg[20]/NET0131  , \P2_reg0_reg[21]/NET0131  , \P2_reg0_reg[22]/NET0131  , \P2_reg0_reg[23]/NET0131  , \P2_reg0_reg[24]/NET0131  , \P2_reg0_reg[25]/NET0131  , \P2_reg0_reg[26]/NET0131  , \P2_reg0_reg[27]/NET0131  , \P2_reg0_reg[28]/NET0131  , \P2_reg0_reg[29]/NET0131  , \P2_reg0_reg[2]/NET0131  , \P2_reg0_reg[30]/NET0131  , \P2_reg0_reg[31]/NET0131  , \P2_reg0_reg[3]/NET0131  , \P2_reg0_reg[4]/NET0131  , \P2_reg0_reg[5]/NET0131  , \P2_reg0_reg[6]/NET0131  , \P2_reg0_reg[7]/NET0131  , \P2_reg0_reg[8]/NET0131  , \P2_reg0_reg[9]/NET0131  , \P2_reg1_reg[0]/NET0131  , \P2_reg1_reg[10]/NET0131  , \P2_reg1_reg[11]/NET0131  , \P2_reg1_reg[12]/NET0131  , \P2_reg1_reg[13]/NET0131  , \P2_reg1_reg[14]/NET0131  , \P2_reg1_reg[15]/NET0131  , \P2_reg1_reg[16]/NET0131  , \P2_reg1_reg[17]/NET0131  , \P2_reg1_reg[18]/NET0131  , \P2_reg1_reg[19]/NET0131  , \P2_reg1_reg[1]/NET0131  , \P2_reg1_reg[20]/NET0131  , \P2_reg1_reg[21]/NET0131  , \P2_reg1_reg[22]/NET0131  , \P2_reg1_reg[23]/NET0131  , \P2_reg1_reg[24]/NET0131  , \P2_reg1_reg[25]/NET0131  , \P2_reg1_reg[26]/NET0131  , \P2_reg1_reg[27]/NET0131  , \P2_reg1_reg[28]/NET0131  , \P2_reg1_reg[29]/NET0131  , \P2_reg1_reg[2]/NET0131  , \P2_reg1_reg[30]/NET0131  , \P2_reg1_reg[31]/NET0131  , \P2_reg1_reg[3]/NET0131  , \P2_reg1_reg[4]/NET0131  , \P2_reg1_reg[5]/NET0131  , \P2_reg1_reg[6]/NET0131  , \P2_reg1_reg[7]/NET0131  , \P2_reg1_reg[8]/NET0131  , \P2_reg1_reg[9]/NET0131  , \P2_reg2_reg[0]/NET0131  , \P2_reg2_reg[10]/NET0131  , \P2_reg2_reg[11]/NET0131  , \P2_reg2_reg[12]/NET0131  , \P2_reg2_reg[13]/NET0131  , \P2_reg2_reg[14]/NET0131  , \P2_reg2_reg[15]/NET0131  , \P2_reg2_reg[16]/NET0131  , \P2_reg2_reg[17]/NET0131  , \P2_reg2_reg[18]/NET0131  , \P2_reg2_reg[19]/NET0131  , \P2_reg2_reg[1]/NET0131  , \P2_reg2_reg[20]/NET0131  , \P2_reg2_reg[21]/NET0131  , \P2_reg2_reg[22]/NET0131  , \P2_reg2_reg[23]/NET0131  , \P2_reg2_reg[24]/NET0131  , \P2_reg2_reg[25]/NET0131  , \P2_reg2_reg[26]/NET0131  , \P2_reg2_reg[27]/NET0131  , \P2_reg2_reg[28]/NET0131  , \P2_reg2_reg[29]/NET0131  , \P2_reg2_reg[2]/NET0131  , \P2_reg2_reg[30]/NET0131  , \P2_reg2_reg[31]/NET0131  , \P2_reg2_reg[3]/NET0131  , \P2_reg2_reg[4]/NET0131  , \P2_reg2_reg[5]/NET0131  , \P2_reg2_reg[6]/NET0131  , \P2_reg2_reg[7]/NET0131  , \P2_reg2_reg[8]/NET0131  , \P2_reg2_reg[9]/NET0131  , \P2_reg3_reg[0]/NET0131  , \P2_reg3_reg[10]/NET0131  , \P2_reg3_reg[11]/NET0131  , \P2_reg3_reg[12]/NET0131  , \P2_reg3_reg[13]/NET0131  , \P2_reg3_reg[14]/NET0131  , \P2_reg3_reg[15]/NET0131  , \P2_reg3_reg[16]/NET0131  , \P2_reg3_reg[17]/NET0131  , \P2_reg3_reg[18]/NET0131  , \P2_reg3_reg[19]/NET0131  , \P2_reg3_reg[1]/NET0131  , \P2_reg3_reg[20]/NET0131  , \P2_reg3_reg[21]/NET0131  , \P2_reg3_reg[22]/NET0131  , \P2_reg3_reg[23]/NET0131  , \P2_reg3_reg[24]/NET0131  , \P2_reg3_reg[25]/NET0131  , \P2_reg3_reg[26]/NET0131  , \P2_reg3_reg[27]/NET0131  , \P2_reg3_reg[28]/NET0131  , \P2_reg3_reg[2]/NET0131  , \P2_reg3_reg[3]/NET0131  , \P2_reg3_reg[4]/NET0131  , \P2_reg3_reg[5]/NET0131  , \P2_reg3_reg[6]/NET0131  , \P2_reg3_reg[7]/NET0131  , \P2_reg3_reg[8]/NET0131  , \P2_reg3_reg[9]/NET0131  , \P2_wr_reg/NET0131  , \P3_B_reg/NET0131  , \P3_IR_reg[0]/NET0131  , \P3_IR_reg[10]/NET0131  , \P3_IR_reg[11]/NET0131  , \P3_IR_reg[12]/NET0131  , \P3_IR_reg[13]/NET0131  , \P3_IR_reg[14]/NET0131  , \P3_IR_reg[15]/NET0131  , \P3_IR_reg[16]/NET0131  , \P3_IR_reg[17]/NET0131  , \P3_IR_reg[18]/NET0131  , \P3_IR_reg[19]/NET0131  , \P3_IR_reg[1]/NET0131  , \P3_IR_reg[20]/NET0131  , \P3_IR_reg[21]/NET0131  , \P3_IR_reg[22]/NET0131  , \P3_IR_reg[23]/NET0131  , \P3_IR_reg[24]/NET0131  , \P3_IR_reg[25]/NET0131  , \P3_IR_reg[26]/NET0131  , \P3_IR_reg[27]/NET0131  , \P3_IR_reg[28]/NET0131  , \P3_IR_reg[29]/NET0131  , \P3_IR_reg[2]/NET0131  , \P3_IR_reg[30]/NET0131  , \P3_IR_reg[31]/NET0131  , \P3_IR_reg[3]/NET0131  , \P3_IR_reg[4]/NET0131  , \P3_IR_reg[5]/NET0131  , \P3_IR_reg[6]/NET0131  , \P3_IR_reg[7]/NET0131  , \P3_IR_reg[8]/NET0131  , \P3_IR_reg[9]/NET0131  , \P3_addr_reg[0]/NET0131  , \P3_addr_reg[10]/NET0131  , \P3_addr_reg[11]/NET0131  , \P3_addr_reg[12]/NET0131  , \P3_addr_reg[13]/NET0131  , \P3_addr_reg[14]/NET0131  , \P3_addr_reg[15]/NET0131  , \P3_addr_reg[16]/NET0131  , \P3_addr_reg[17]/NET0131  , \P3_addr_reg[18]/NET0131  , \P3_addr_reg[19]/NET0131  , \P3_addr_reg[1]/NET0131  , \P3_addr_reg[2]/NET0131  , \P3_addr_reg[3]/NET0131  , \P3_addr_reg[4]/NET0131  , \P3_addr_reg[5]/NET0131  , \P3_addr_reg[6]/NET0131  , \P3_addr_reg[7]/NET0131  , \P3_addr_reg[8]/NET0131  , \P3_addr_reg[9]/NET0131  , \P3_d_reg[0]/NET0131  , \P3_d_reg[1]/NET0131  , \P3_rd_reg/NET0131  , \P3_reg0_reg[0]/NET0131  , \P3_reg0_reg[10]/NET0131  , \P3_reg0_reg[11]/NET0131  , \P3_reg0_reg[12]/NET0131  , \P3_reg0_reg[13]/NET0131  , \P3_reg0_reg[14]/NET0131  , \P3_reg0_reg[15]/NET0131  , \P3_reg0_reg[16]/NET0131  , \P3_reg0_reg[17]/NET0131  , \P3_reg0_reg[18]/NET0131  , \P3_reg0_reg[19]/NET0131  , \P3_reg0_reg[1]/NET0131  , \P3_reg0_reg[20]/NET0131  , \P3_reg0_reg[21]/NET0131  , \P3_reg0_reg[22]/NET0131  , \P3_reg0_reg[23]/NET0131  , \P3_reg0_reg[24]/NET0131  , \P3_reg0_reg[25]/NET0131  , \P3_reg0_reg[26]/NET0131  , \P3_reg0_reg[27]/NET0131  , \P3_reg0_reg[28]/NET0131  , \P3_reg0_reg[29]/NET0131  , \P3_reg0_reg[2]/NET0131  , \P3_reg0_reg[30]/NET0131  , \P3_reg0_reg[31]/NET0131  , \P3_reg0_reg[3]/NET0131  , \P3_reg0_reg[4]/NET0131  , \P3_reg0_reg[5]/NET0131  , \P3_reg0_reg[6]/NET0131  , \P3_reg0_reg[7]/NET0131  , \P3_reg0_reg[8]/NET0131  , \P3_reg0_reg[9]/NET0131  , \P3_reg1_reg[0]/NET0131  , \P3_reg1_reg[10]/NET0131  , \P3_reg1_reg[11]/NET0131  , \P3_reg1_reg[12]/NET0131  , \P3_reg1_reg[13]/NET0131  , \P3_reg1_reg[14]/NET0131  , \P3_reg1_reg[15]/NET0131  , \P3_reg1_reg[16]/NET0131  , \P3_reg1_reg[17]/NET0131  , \P3_reg1_reg[18]/NET0131  , \P3_reg1_reg[19]/NET0131  , \P3_reg1_reg[1]/NET0131  , \P3_reg1_reg[20]/NET0131  , \P3_reg1_reg[21]/NET0131  , \P3_reg1_reg[22]/NET0131  , \P3_reg1_reg[23]/NET0131  , \P3_reg1_reg[24]/NET0131  , \P3_reg1_reg[25]/NET0131  , \P3_reg1_reg[26]/NET0131  , \P3_reg1_reg[27]/NET0131  , \P3_reg1_reg[28]/NET0131  , \P3_reg1_reg[29]/NET0131  , \P3_reg1_reg[2]/NET0131  , \P3_reg1_reg[30]/NET0131  , \P3_reg1_reg[31]/NET0131  , \P3_reg1_reg[3]/NET0131  , \P3_reg1_reg[4]/NET0131  , \P3_reg1_reg[5]/NET0131  , \P3_reg1_reg[6]/NET0131  , \P3_reg1_reg[7]/NET0131  , \P3_reg1_reg[8]/NET0131  , \P3_reg1_reg[9]/NET0131  , \P3_reg2_reg[0]/NET0131  , \P3_reg2_reg[10]/NET0131  , \P3_reg2_reg[11]/NET0131  , \P3_reg2_reg[12]/NET0131  , \P3_reg2_reg[13]/NET0131  , \P3_reg2_reg[14]/NET0131  , \P3_reg2_reg[15]/NET0131  , \P3_reg2_reg[16]/NET0131  , \P3_reg2_reg[17]/NET0131  , \P3_reg2_reg[18]/NET0131  , \P3_reg2_reg[19]/NET0131  , \P3_reg2_reg[1]/NET0131  , \P3_reg2_reg[20]/NET0131  , \P3_reg2_reg[21]/NET0131  , \P3_reg2_reg[22]/NET0131  , \P3_reg2_reg[23]/NET0131  , \P3_reg2_reg[24]/NET0131  , \P3_reg2_reg[25]/NET0131  , \P3_reg2_reg[26]/NET0131  , \P3_reg2_reg[27]/NET0131  , \P3_reg2_reg[28]/NET0131  , \P3_reg2_reg[29]/NET0131  , \P3_reg2_reg[2]/NET0131  , \P3_reg2_reg[30]/NET0131  , \P3_reg2_reg[31]/NET0131  , \P3_reg2_reg[3]/NET0131  , \P3_reg2_reg[4]/NET0131  , \P3_reg2_reg[5]/NET0131  , \P3_reg2_reg[6]/NET0131  , \P3_reg2_reg[7]/NET0131  , \P3_reg2_reg[8]/NET0131  , \P3_reg2_reg[9]/NET0131  , \P3_reg3_reg[0]/NET0131  , \P3_reg3_reg[10]/NET0131  , \P3_reg3_reg[11]/NET0131  , \P3_reg3_reg[12]/NET0131  , \P3_reg3_reg[13]/NET0131  , \P3_reg3_reg[14]/NET0131  , \P3_reg3_reg[15]/NET0131  , \P3_reg3_reg[16]/NET0131  , \P3_reg3_reg[17]/NET0131  , \P3_reg3_reg[18]/NET0131  , \P3_reg3_reg[19]/NET0131  , \P3_reg3_reg[1]/NET0131  , \P3_reg3_reg[20]/NET0131  , \P3_reg3_reg[21]/NET0131  , \P3_reg3_reg[22]/NET0131  , \P3_reg3_reg[23]/NET0131  , \P3_reg3_reg[24]/NET0131  , \P3_reg3_reg[25]/NET0131  , \P3_reg3_reg[26]/NET0131  , \P3_reg3_reg[27]/NET0131  , \P3_reg3_reg[28]/NET0131  , \P3_reg3_reg[2]/NET0131  , \P3_reg3_reg[3]/NET0131  , \P3_reg3_reg[4]/NET0131  , \P3_reg3_reg[5]/NET0131  , \P3_reg3_reg[6]/NET0131  , \P3_reg3_reg[7]/NET0131  , \P3_reg3_reg[8]/NET0131  , \P3_reg3_reg[9]/NET0131  , \P3_wr_reg/NET0131  , \si[0]_pad  , \si[10]_pad  , \si[11]_pad  , \si[12]_pad  , \si[13]_pad  , \si[14]_pad  , \si[15]_pad  , \si[16]_pad  , \si[17]_pad  , \si[18]_pad  , \si[19]_pad  , \si[1]_pad  , \si[20]_pad  , \si[21]_pad  , \si[22]_pad  , \si[23]_pad  , \si[24]_pad  , \si[25]_pad  , \si[26]_pad  , \si[27]_pad  , \si[28]_pad  , \si[29]_pad  , \si[2]_pad  , \si[30]_pad  , \si[31]_pad  , \si[3]_pad  , \si[4]_pad  , \si[5]_pad  , \si[6]_pad  , \si[7]_pad  , \si[8]_pad  , \si[9]_pad  , \P1_state_reg[0]/NET0131_syn_2  , \_al_n0  , \_al_n1  , \g106254/_0_  , \g106255/_0_  , \g106267/_0_  , \g106268/_0_  , \g106269/_0_  , \g106270/_0_  , \g106271/_0_  , \g106272/_0_  , \g106288/_0_  , \g106289/_0_  , \g106290/_0_  , \g106291/_0_  , \g106292/_0_  , \g106293/_0_  , \g106294/_0_  , \g106295/_0_  , \g106296/_0_  , \g106297/_0_  , \g106352/_0_  , \g106356/_0_  , \g106359/_0_  , \g106360/_0_  , \g106361/_0_  , \g106362/_0_  , \g106363/_0_  , \g106364/_0_  , \g106365/_0_  , \g106406/_0_  , \g106407/_0_  , \g106408/_0_  , \g106410/_0_  , \g106411/_0_  , \g106412/_0_  , \g106413/_0_  , \g106414/_0_  , \g106417/_0_  , \g106418/_0_  , \g106419/_0_  , \g106420/_0_  , \g106421/_0_  , \g106422/_0_  , \g106423/_0_  , \g106424/_0_  , \g106425/_0_  , \g106426/_0_  , \g106427/_0_  , \g106428/_0_  , \g106430/_0_  , \g106431/_0_  , \g106432/_0_  , \g106433/_0_  , \g106434/_0_  , \g106436/_0_  , \g106437/_0_  , \g106438/_0_  , \g106439/_0_  , \g106440/_0_  , \g106441/_0_  , \g106442/_0_  , \g106443/_0_  , \g106444/_0_  , \g106445/_0_  , \g106446/_0_  , \g106447/_0_  , \g106448/_0_  , \g106530/_0_  , \g106531/_0_  , \g106532/_0_  , \g106533/_0_  , \g106534/_0_  , \g106554/_0_  , \g106556/_0_  , \g106557/_0_  , \g106559/_0_  , \g106560/_0_  , \g106561/_0_  , \g106562/_0_  , \g106563/_0_  , \g106564/_0_  , \g106565/_0_  , \g106566/_0_  , \g106567/_0_  , \g106568/_0_  , \g106569/_0_  , \g106570/_0_  , \g106571/_0_  , \g106572/_0_  , \g106633/_0_  , \g106634/_0_  , \g106640/_0_  , \g106654/_0_  , \g106655/_0_  , \g106679/_0_  , \g106682/_0_  , \g106684/_0_  , \g106687/_0_  , \g106690/_0_  , \g106691/_0_  , \g106692/_0_  , \g106693/_0_  , \g106694/_0_  , \g106695/_0_  , \g106696/_0_  , \g106697/_0_  , \g106698/_0_  , \g106699/_0_  , \g106700/_0_  , \g106701/_0_  , \g106702/_0_  , \g106703/_0_  , \g106704/_0_  , \g106705/_0_  , \g106706/_0_  , \g106707/_0_  , \g106708/_0_  , \g106710/_0_  , \g106711/_0_  , \g106712/_0_  , \g106713/_0_  , \g106714/_0_  , \g106715/_0_  , \g106716/_0_  , \g106717/_0_  , \g106718/_0_  , \g106719/_0_  , \g106720/_0_  , \g106721/_0_  , \g106722/_0_  , \g106723/_0_  , \g106724/_0_  , \g106725/_0_  , \g106726/_0_  , \g106727/_0_  , \g106728/_0_  , \g106729/_0_  , \g106830/_0_  , \g106836/_0_  , \g106837/_0_  , \g106838/_0_  , \g106843/_0_  , \g106850/_0_  , \g106851/_0_  , \g106852/_0_  , \g106853/_0_  , \g106854/_0_  , \g106899/_0_  , \g106901/_0_  , \g106902/_0_  , \g106903/_0_  , \g106904/_0_  , \g106905/_0_  , \g106906/_0_  , \g106907/_0_  , \g106908/_0_  , \g106909/_0_  , \g106910/_0_  , \g106911/_0_  , \g106912/_0_  , \g106913/_0_  , \g106914/_0_  , \g106915/_0_  , \g106916/_0_  , \g106917/_0_  , \g106918/_0_  , \g106919/_0_  , \g106920/_0_  , \g106921/_0_  , \g106922/_0_  , \g106923/_0_  , \g106924/_0_  , \g106925/_0_  , \g106994/_0_  , \g106995/_0_  , \g106996/_0_  , \g106997/_0_  , \g106998/_0_  , \g106999/_0_  , \g107002/_0_  , \g107007/_0_  , \g107008/_0_  , \g107038/_0_  , \g107041/_0_  , \g107048/_0_  , \g107091/_0_  , \g107093/_0_  , \g107094/_0_  , \g107096/_0_  , \g107097/_0_  , \g107098/_0_  , \g107099/_0_  , \g107100/_0_  , \g107101/_0_  , \g107102/_0_  , \g107103/_0_  , \g107104/_0_  , \g107105/_0_  , \g107106/_0_  , \g107107/_0_  , \g107108/_0_  , \g107109/_0_  , \g107110/_0_  , \g107111/_0_  , \g107112/_0_  , \g107113/_0_  , \g107114/_0_  , \g107115/_0_  , \g107116/_0_  , \g107117/_0_  , \g107118/_0_  , \g107119/_0_  , \g107120/_0_  , \g107121/_0_  , \g107122/_0_  , \g107123/_0_  , \g107124/_0_  , \g107125/_0_  , \g107126/_0_  , \g107127/_0_  , \g107128/_0_  , \g107129/_0_  , \g107130/_0_  , \g107131/_0_  , \g107132/_0_  , \g107133/_0_  , \g107134/_0_  , \g107135/_0_  , \g107136/_0_  , \g107137/_0_  , \g107138/_0_  , \g107248/_0_  , \g107252/_0_  , \g107254/_0_  , \g107255/_0_  , \g107280/_0_  , \g107281/_0_  , \g107282/_0_  , \g107370/_0_  , \g107371/_0_  , \g107372/_0_  , \g107373/_0_  , \g107374/_0_  , \g107375/_0_  , \g107376/_0_  , \g107377/_0_  , \g107378/_0_  , \g107379/_0_  , \g107380/_0_  , \g107381/_0_  , \g107382/_0_  , \g107383/_0_  , \g107384/_0_  , \g107385/_0_  , \g107386/_0_  , \g107387/_0_  , \g107388/_0_  , \g107389/_0_  , \g107390/_0_  , \g107391/_0_  , \g107488/_0_  , \g107489/_0_  , \g107490/_0_  , \g107491/_0_  , \g107492/_0_  , \g107493/_0_  , \g107500/_0_  , \g107615/_0_  , \g107623/_0_  , \g107624/_0_  , \g107625/_0_  , \g107626/_0_  , \g107627/_0_  , \g107628/_0_  , \g107629/_0_  , \g107630/_0_  , \g107631/_0_  , \g107632/_0_  , \g107634/_0_  , \g107637/_0_  , \g107638/_0_  , \g107639/_0_  , \g107640/_0_  , \g107641/_0_  , \g107642/_0_  , \g107643/_0_  , \g107644/_0_  , \g107645/_0_  , \g107646/_0_  , \g107647/_0_  , \g107650/_0_  , \g107651/_0_  , \g107652/_0_  , \g107653/_0_  , \g107654/_0_  , \g107655/_0_  , \g107656/_0_  , \g107743/_0_  , \g107787/_0_  , \g107954/_0_  , \g107955/_0_  , \g107956/_0_  , \g107957/_0_  , \g107958/_0_  , \g107959/_0_  , \g107960/_0_  , \g107961/_0_  , \g107962/_0_  , \g107963/_0_  , \g107964/_0_  , \g107965/_0_  , \g107966/_0_  , \g107967/_0_  , \g108118/_0_  , \g108125/_0_  , \g108169/_0_  , \g108269/_0_  , \g108270/_0_  , \g108319/_0_  , \g108320/_0_  , \g108321/_0_  , \g108322/_0_  , \g108323/_0_  , \g108324/_0_  , \g108326/_0_  , \g108327/_0_  , \g108328/_0_  , \g108329/_0_  , \g108330/_0_  , \g108334/_0_  , \g108335/_0_  , \g108468/_0_  , \g108538/_0_  , \g108801/_0_  , \g108812/_0_  , \g108813/_0_  , \g108814/_0_  , \g108815/_0_  , \g108817/_0_  , \g108818/_0_  , \g108819/_0_  , \g108822/_0_  , \g109052/_0_  , \g109053/_0_  , \g109401/_0_  , \g109402/_0_  , \g109403/_0_  , \g109410/_0_  , \g109411/_0_  , \g109415/_0_  , \g109420/_0_  , \g109425/_0_  , \g109693/_0_  , \g110116/_0_  , \g110117/_0_  , \g110905/_0_  , \g110906/_0_  , \g110907/_0_  , \g111086/_0_  , \g111094/_0_  , \g112422/_0_  , \g112423/_0_  , \g112424/_0_  , \g112425/_0_  , \g112426/_0_  , \g112427/_0_  , \g113647/_0_  , \g113648/_0_  , \g113649/_0_  , \g113650/_0_  , \g113651/_0_  , \g114133/_0_  , \g117884/_0_  , \g117885/_0_  , \g117886/_0_  , \g117895/_3_  , \g117896/_3_  , \g117897/_0_  , \g117898/_0_  , \g117899/_0_  , \g117900/_3_  , \g120982/_0_  , \g120983/_0_  , \g120984/_0_  , \g120985/_0_  , \g120986/_0_  , \g120987/_0_  , \g120988/_3_  , \g120989/_0_  , \g120990/_0_  , \g120991/_0_  , \g120992/_0_  , \g120993/_0_  , \g120994/_0_  , \g120995/_0_  , \g120996/_3_  , \g120997/_0_  , \g120998/_0_  , \g120999/_0_  , \g121000/_0_  , \g121001/_0_  , \g121002/_3_  , \g121003/_0_  , \g121004/_0_  , \g121005/_3_  , \g121006/_0_  , \g121007/_0_  , \g121008/_0_  , \g121029/_0_  , \g121030/_3_  , \g121032/_3_  , \g121033/_3_  , \g121034/_3_  , \g121035/_3_  , \g121036/_3_  , \g121037/_3_  , \g121038/_3_  , \g121039/_3_  , \g121040/_3_  , \g121041/_3_  , \g121042/_3_  , \g121043/_3_  , \g121044/_3_  , \g121045/_3_  , \g121046/_3_  , \g121047/_3_  , \g121048/_3_  , \g121049/_3_  , \g121050/_3_  , \g121051/_0_  , \g121052/_3_  , \g121053/_3_  , \g121054/_3_  , \g121055/_3_  , \g121056/_3_  , \g121057/_3_  , \g121058/_3_  , \g121060/_3_  , \g121061/_3_  , \g121062/_3_  , \g121063/_3_  , \g121064/_3_  , \g121065/_3_  , \g121066/_3_  , \g121067/_3_  , \g121068/_3_  , \g121069/_3_  , \g121070/_3_  , \g121071/_3_  , \g121072/_3_  , \g121073/_3_  , \g121074/_3_  , \g121075/_3_  , \g121076/_3_  , \g121077/_3_  , \g121078/_3_  , \g121079/_3_  , \g121080/_0_  , \g121081/_3_  , \g121082/_0_  , \g121083/_3_  , \g121084/_3_  , \g121085/_3_  , \g121086/_3_  , \g121087/_3_  , \g121626/_0_  , \g121633/_0_  , \g121669/_0_  , \g122948/_0_  , \g122949/_0_  , \g122951/_0_  , \g122952/_0_  , \g122953/_0_  , \g122954/_0_  , \g122955/_0_  , \g122956/_0_  , \g122957/_0_  , \g122958/_0_  , \g122959/_0_  , \g122960/_0_  , \g122963/_0_  , \g122965/_0_  , \g122967/_0_  , \g122968/_0_  , \g122972/_0_  , \g122973/_0_  , \g122974/_0_  , \g122975/_0_  , \g122976/_0_  , \g122977/_0_  , \g122978/_0_  , \g122979/_0_  , \g122980/_0_  , \g122981/_0_  , \g122982/_0_  , \g122983/_0_  , \g122984/_0_  , \g122985/_0_  , \g122986/_0_  , \g122987/_0_  , \g122988/_0_  , \g122989/_0_  , \g122990/_0_  , \g122991/_0_  , \g122997/_0_  , \g122998/_0_  , \g122999/_0_  , \g123000/_0_  , \g123740/_0_  , \g123811/_0_  , \g123812/_0_  , \g123813/_0_  , \g123814/_0_  , \g123815/_0_  , \g123816/_0_  , \g123817/_0_  , \g123818/_0_  , \g123819/_0_  , \g123820/_0_  , \g123821/_0_  , \g123822/_0_  , \g123823/_0_  , \g123824/_0_  , \g123825/_0_  , \g123826/_0_  , \g123827/_0_  , \g123828/_0_  , \g123829/_0_  , \g123830/_0_  , \g123853/u3_syn_4  , \g123854/u3_syn_4  , \g123871/_0_  , \g124519/_0_  , \g124554/_0_  , \g124798/_0_  , \g124897/_0_  , \g125133/_0_  , \g125231/_0_  , \g125318/u3_syn_4  , \g125495/u3_syn_4  , \g126480/_0_  , \g126501/_0_  , \g127137/_0_  , \g127147/_0_  , \g127163/_0_  , \g127173/_0_  , \g127202/_0_  , \g127211/_0_  , \g127223/_0_  , \g127234/_0_  , \g127241/_0_  , \g127251/_0_  , \g127257/_0_  , \g127262/_0_  , \g127271/_0_  , \g127285/_0_  , \g127292/_0_  , \g127302/_0_  , \g127313/_0_  , \g127324/_0_  , \g127334/_0_  , \g127348/_0_  , \g127366/_0_  , \g127396/_0_  , \g127405/_0_  , \g127411/_0_  , \g127427/_0_  , \g127439/_0_  , \g127464/_0_  , \g127893/_0_  , \g128290/_0_  , \g128431/_0_  , \g128477/_0_  , \g128501/_0_  , \g128540/_0_  , \g128566/_0_  , \g128575/_0_  , \g128586/_0_  , \g128594/_1_  , \g128631/_0_  , \g128648/_0_  , \g128698/_0_  , \g131281/_1_  , \g140384/_0_  , \g140411/_0_  , \g140627/_0_  , \g140741/_0_  , \g140774/_0_  , \g140804/_0_  , \g140955/_0_  , \g140986/_0_  , \g141163/_0_  , \g141237/_0_  , \g141301/_0_  , \g141328/_0_  , \g141367/_0_  , \g141441/_0_  , \g141474/_0_  , \g141548/_0_  , \g141640/_0_  , \g141838/_0_  , \g141844/_0_  , \g141853/_0_  , \g141855/_0_  , \g141860/_0_  , \g141896/_0_  , \g141915/_0_  , \g141952/_0_  , \g142033/_0_  , \g142046/_0_  , \g29/_0_  , \g33/_0_  , \g53/_0_  , \g71/_0_  , \g90/_0_  , rd_pad , \so[0]_pad  , \so[10]_pad  , \so[11]_pad  , \so[12]_pad  , \so[13]_pad  , \so[14]_pad  , \so[15]_pad  , \so[16]_pad  , \so[17]_pad  , \so[18]_pad  , \so[19]_pad  , \so[1]_pad  , \so[2]_pad  , \so[3]_pad  , \so[4]_pad  , \so[5]_pad  , \so[6]_pad  , \so[7]_pad  , \so[8]_pad  , \so[9]_pad  , wr_pad );
  input \P1_B_reg/NET0131  ;
  input \P1_IR_reg[0]/NET0131  ;
  input \P1_IR_reg[10]/NET0131  ;
  input \P1_IR_reg[11]/NET0131  ;
  input \P1_IR_reg[12]/NET0131  ;
  input \P1_IR_reg[13]/NET0131  ;
  input \P1_IR_reg[14]/NET0131  ;
  input \P1_IR_reg[15]/NET0131  ;
  input \P1_IR_reg[16]/NET0131  ;
  input \P1_IR_reg[17]/NET0131  ;
  input \P1_IR_reg[18]/NET0131  ;
  input \P1_IR_reg[19]/NET0131  ;
  input \P1_IR_reg[1]/NET0131  ;
  input \P1_IR_reg[20]/NET0131  ;
  input \P1_IR_reg[21]/NET0131  ;
  input \P1_IR_reg[22]/NET0131  ;
  input \P1_IR_reg[23]/NET0131  ;
  input \P1_IR_reg[24]/NET0131  ;
  input \P1_IR_reg[25]/NET0131  ;
  input \P1_IR_reg[26]/NET0131  ;
  input \P1_IR_reg[27]/NET0131  ;
  input \P1_IR_reg[28]/NET0131  ;
  input \P1_IR_reg[29]/NET0131  ;
  input \P1_IR_reg[2]/NET0131  ;
  input \P1_IR_reg[30]/NET0131  ;
  input \P1_IR_reg[31]/NET0131  ;
  input \P1_IR_reg[3]/NET0131  ;
  input \P1_IR_reg[4]/NET0131  ;
  input \P1_IR_reg[5]/NET0131  ;
  input \P1_IR_reg[6]/NET0131  ;
  input \P1_IR_reg[7]/NET0131  ;
  input \P1_IR_reg[8]/NET0131  ;
  input \P1_IR_reg[9]/NET0131  ;
  input \P1_addr_reg[0]/NET0131  ;
  input \P1_addr_reg[10]/NET0131  ;
  input \P1_addr_reg[11]/NET0131  ;
  input \P1_addr_reg[12]/NET0131  ;
  input \P1_addr_reg[13]/NET0131  ;
  input \P1_addr_reg[14]/NET0131  ;
  input \P1_addr_reg[15]/NET0131  ;
  input \P1_addr_reg[16]/NET0131  ;
  input \P1_addr_reg[17]/NET0131  ;
  input \P1_addr_reg[18]/NET0131  ;
  input \P1_addr_reg[19]/NET0131  ;
  input \P1_addr_reg[1]/NET0131  ;
  input \P1_addr_reg[2]/NET0131  ;
  input \P1_addr_reg[3]/NET0131  ;
  input \P1_addr_reg[4]/NET0131  ;
  input \P1_addr_reg[5]/NET0131  ;
  input \P1_addr_reg[6]/NET0131  ;
  input \P1_addr_reg[7]/NET0131  ;
  input \P1_addr_reg[8]/NET0131  ;
  input \P1_addr_reg[9]/NET0131  ;
  input \P1_d_reg[0]/NET0131  ;
  input \P1_d_reg[1]/NET0131  ;
  input \P1_datao_reg[0]/NET0131  ;
  input \P1_datao_reg[10]/NET0131  ;
  input \P1_datao_reg[11]/NET0131  ;
  input \P1_datao_reg[12]/NET0131  ;
  input \P1_datao_reg[13]/NET0131  ;
  input \P1_datao_reg[14]/NET0131  ;
  input \P1_datao_reg[15]/NET0131  ;
  input \P1_datao_reg[16]/NET0131  ;
  input \P1_datao_reg[17]/NET0131  ;
  input \P1_datao_reg[18]/NET0131  ;
  input \P1_datao_reg[19]/NET0131  ;
  input \P1_datao_reg[1]/NET0131  ;
  input \P1_datao_reg[20]/NET0131  ;
  input \P1_datao_reg[21]/NET0131  ;
  input \P1_datao_reg[22]/NET0131  ;
  input \P1_datao_reg[23]/NET0131  ;
  input \P1_datao_reg[24]/NET0131  ;
  input \P1_datao_reg[25]/NET0131  ;
  input \P1_datao_reg[26]/NET0131  ;
  input \P1_datao_reg[27]/NET0131  ;
  input \P1_datao_reg[28]/NET0131  ;
  input \P1_datao_reg[29]/NET0131  ;
  input \P1_datao_reg[2]/NET0131  ;
  input \P1_datao_reg[30]/NET0131  ;
  input \P1_datao_reg[31]/NET0131  ;
  input \P1_datao_reg[3]/NET0131  ;
  input \P1_datao_reg[4]/NET0131  ;
  input \P1_datao_reg[5]/NET0131  ;
  input \P1_datao_reg[6]/NET0131  ;
  input \P1_datao_reg[7]/NET0131  ;
  input \P1_datao_reg[8]/NET0131  ;
  input \P1_datao_reg[9]/NET0131  ;
  input \P1_rd_reg/NET0131  ;
  input \P1_reg0_reg[0]/NET0131  ;
  input \P1_reg0_reg[10]/NET0131  ;
  input \P1_reg0_reg[11]/NET0131  ;
  input \P1_reg0_reg[12]/NET0131  ;
  input \P1_reg0_reg[13]/NET0131  ;
  input \P1_reg0_reg[14]/NET0131  ;
  input \P1_reg0_reg[15]/NET0131  ;
  input \P1_reg0_reg[16]/NET0131  ;
  input \P1_reg0_reg[17]/NET0131  ;
  input \P1_reg0_reg[18]/NET0131  ;
  input \P1_reg0_reg[19]/NET0131  ;
  input \P1_reg0_reg[1]/NET0131  ;
  input \P1_reg0_reg[20]/NET0131  ;
  input \P1_reg0_reg[21]/NET0131  ;
  input \P1_reg0_reg[22]/NET0131  ;
  input \P1_reg0_reg[23]/NET0131  ;
  input \P1_reg0_reg[24]/NET0131  ;
  input \P1_reg0_reg[25]/NET0131  ;
  input \P1_reg0_reg[26]/NET0131  ;
  input \P1_reg0_reg[27]/NET0131  ;
  input \P1_reg0_reg[28]/NET0131  ;
  input \P1_reg0_reg[29]/NET0131  ;
  input \P1_reg0_reg[2]/NET0131  ;
  input \P1_reg0_reg[30]/NET0131  ;
  input \P1_reg0_reg[31]/NET0131  ;
  input \P1_reg0_reg[3]/NET0131  ;
  input \P1_reg0_reg[4]/NET0131  ;
  input \P1_reg0_reg[5]/NET0131  ;
  input \P1_reg0_reg[6]/NET0131  ;
  input \P1_reg0_reg[7]/NET0131  ;
  input \P1_reg0_reg[8]/NET0131  ;
  input \P1_reg0_reg[9]/NET0131  ;
  input \P1_reg1_reg[0]/NET0131  ;
  input \P1_reg1_reg[10]/NET0131  ;
  input \P1_reg1_reg[11]/NET0131  ;
  input \P1_reg1_reg[12]/NET0131  ;
  input \P1_reg1_reg[13]/NET0131  ;
  input \P1_reg1_reg[14]/NET0131  ;
  input \P1_reg1_reg[15]/NET0131  ;
  input \P1_reg1_reg[16]/NET0131  ;
  input \P1_reg1_reg[17]/NET0131  ;
  input \P1_reg1_reg[18]/NET0131  ;
  input \P1_reg1_reg[19]/NET0131  ;
  input \P1_reg1_reg[1]/NET0131  ;
  input \P1_reg1_reg[20]/NET0131  ;
  input \P1_reg1_reg[21]/NET0131  ;
  input \P1_reg1_reg[22]/NET0131  ;
  input \P1_reg1_reg[23]/NET0131  ;
  input \P1_reg1_reg[24]/NET0131  ;
  input \P1_reg1_reg[25]/NET0131  ;
  input \P1_reg1_reg[26]/NET0131  ;
  input \P1_reg1_reg[27]/NET0131  ;
  input \P1_reg1_reg[28]/NET0131  ;
  input \P1_reg1_reg[29]/NET0131  ;
  input \P1_reg1_reg[2]/NET0131  ;
  input \P1_reg1_reg[30]/NET0131  ;
  input \P1_reg1_reg[31]/NET0131  ;
  input \P1_reg1_reg[3]/NET0131  ;
  input \P1_reg1_reg[4]/NET0131  ;
  input \P1_reg1_reg[5]/NET0131  ;
  input \P1_reg1_reg[6]/NET0131  ;
  input \P1_reg1_reg[7]/NET0131  ;
  input \P1_reg1_reg[8]/NET0131  ;
  input \P1_reg1_reg[9]/NET0131  ;
  input \P1_reg2_reg[0]/NET0131  ;
  input \P1_reg2_reg[10]/NET0131  ;
  input \P1_reg2_reg[11]/NET0131  ;
  input \P1_reg2_reg[12]/NET0131  ;
  input \P1_reg2_reg[13]/NET0131  ;
  input \P1_reg2_reg[14]/NET0131  ;
  input \P1_reg2_reg[15]/NET0131  ;
  input \P1_reg2_reg[16]/NET0131  ;
  input \P1_reg2_reg[17]/NET0131  ;
  input \P1_reg2_reg[18]/NET0131  ;
  input \P1_reg2_reg[19]/NET0131  ;
  input \P1_reg2_reg[1]/NET0131  ;
  input \P1_reg2_reg[20]/NET0131  ;
  input \P1_reg2_reg[21]/NET0131  ;
  input \P1_reg2_reg[22]/NET0131  ;
  input \P1_reg2_reg[23]/NET0131  ;
  input \P1_reg2_reg[24]/NET0131  ;
  input \P1_reg2_reg[25]/NET0131  ;
  input \P1_reg2_reg[26]/NET0131  ;
  input \P1_reg2_reg[27]/NET0131  ;
  input \P1_reg2_reg[28]/NET0131  ;
  input \P1_reg2_reg[29]/NET0131  ;
  input \P1_reg2_reg[2]/NET0131  ;
  input \P1_reg2_reg[30]/NET0131  ;
  input \P1_reg2_reg[31]/NET0131  ;
  input \P1_reg2_reg[3]/NET0131  ;
  input \P1_reg2_reg[4]/NET0131  ;
  input \P1_reg2_reg[5]/NET0131  ;
  input \P1_reg2_reg[6]/NET0131  ;
  input \P1_reg2_reg[7]/NET0131  ;
  input \P1_reg2_reg[8]/NET0131  ;
  input \P1_reg2_reg[9]/NET0131  ;
  input \P1_reg3_reg[0]/NET0131  ;
  input \P1_reg3_reg[10]/NET0131  ;
  input \P1_reg3_reg[11]/NET0131  ;
  input \P1_reg3_reg[12]/NET0131  ;
  input \P1_reg3_reg[13]/NET0131  ;
  input \P1_reg3_reg[14]/NET0131  ;
  input \P1_reg3_reg[15]/NET0131  ;
  input \P1_reg3_reg[16]/NET0131  ;
  input \P1_reg3_reg[17]/NET0131  ;
  input \P1_reg3_reg[18]/NET0131  ;
  input \P1_reg3_reg[19]/NET0131  ;
  input \P1_reg3_reg[1]/NET0131  ;
  input \P1_reg3_reg[20]/NET0131  ;
  input \P1_reg3_reg[21]/NET0131  ;
  input \P1_reg3_reg[22]/NET0131  ;
  input \P1_reg3_reg[23]/NET0131  ;
  input \P1_reg3_reg[24]/NET0131  ;
  input \P1_reg3_reg[25]/NET0131  ;
  input \P1_reg3_reg[26]/NET0131  ;
  input \P1_reg3_reg[27]/NET0131  ;
  input \P1_reg3_reg[28]/NET0131  ;
  input \P1_reg3_reg[2]/NET0131  ;
  input \P1_reg3_reg[3]/NET0131  ;
  input \P1_reg3_reg[4]/NET0131  ;
  input \P1_reg3_reg[5]/NET0131  ;
  input \P1_reg3_reg[6]/NET0131  ;
  input \P1_reg3_reg[7]/NET0131  ;
  input \P1_reg3_reg[8]/NET0131  ;
  input \P1_reg3_reg[9]/NET0131  ;
  input \P1_state_reg[0]/NET0131  ;
  input \P1_wr_reg/NET0131  ;
  input \P2_B_reg/NET0131  ;
  input \P2_IR_reg[0]/NET0131  ;
  input \P2_IR_reg[10]/NET0131  ;
  input \P2_IR_reg[11]/NET0131  ;
  input \P2_IR_reg[12]/NET0131  ;
  input \P2_IR_reg[13]/NET0131  ;
  input \P2_IR_reg[14]/NET0131  ;
  input \P2_IR_reg[15]/NET0131  ;
  input \P2_IR_reg[16]/NET0131  ;
  input \P2_IR_reg[17]/NET0131  ;
  input \P2_IR_reg[18]/NET0131  ;
  input \P2_IR_reg[19]/NET0131  ;
  input \P2_IR_reg[1]/NET0131  ;
  input \P2_IR_reg[20]/NET0131  ;
  input \P2_IR_reg[21]/NET0131  ;
  input \P2_IR_reg[22]/NET0131  ;
  input \P2_IR_reg[23]/NET0131  ;
  input \P2_IR_reg[24]/NET0131  ;
  input \P2_IR_reg[25]/NET0131  ;
  input \P2_IR_reg[26]/NET0131  ;
  input \P2_IR_reg[27]/NET0131  ;
  input \P2_IR_reg[28]/NET0131  ;
  input \P2_IR_reg[29]/NET0131  ;
  input \P2_IR_reg[2]/NET0131  ;
  input \P2_IR_reg[30]/NET0131  ;
  input \P2_IR_reg[31]/NET0131  ;
  input \P2_IR_reg[3]/NET0131  ;
  input \P2_IR_reg[4]/NET0131  ;
  input \P2_IR_reg[5]/NET0131  ;
  input \P2_IR_reg[6]/NET0131  ;
  input \P2_IR_reg[7]/NET0131  ;
  input \P2_IR_reg[8]/NET0131  ;
  input \P2_IR_reg[9]/NET0131  ;
  input \P2_addr_reg[0]/NET0131  ;
  input \P2_addr_reg[10]/NET0131  ;
  input \P2_addr_reg[11]/NET0131  ;
  input \P2_addr_reg[12]/NET0131  ;
  input \P2_addr_reg[13]/NET0131  ;
  input \P2_addr_reg[14]/NET0131  ;
  input \P2_addr_reg[15]/NET0131  ;
  input \P2_addr_reg[16]/NET0131  ;
  input \P2_addr_reg[17]/NET0131  ;
  input \P2_addr_reg[18]/NET0131  ;
  input \P2_addr_reg[19]/NET0131  ;
  input \P2_addr_reg[1]/NET0131  ;
  input \P2_addr_reg[2]/NET0131  ;
  input \P2_addr_reg[3]/NET0131  ;
  input \P2_addr_reg[4]/NET0131  ;
  input \P2_addr_reg[5]/NET0131  ;
  input \P2_addr_reg[6]/NET0131  ;
  input \P2_addr_reg[7]/NET0131  ;
  input \P2_addr_reg[8]/NET0131  ;
  input \P2_addr_reg[9]/NET0131  ;
  input \P2_d_reg[0]/NET0131  ;
  input \P2_d_reg[1]/NET0131  ;
  input \P2_datao_reg[0]/NET0131  ;
  input \P2_datao_reg[10]/NET0131  ;
  input \P2_datao_reg[11]/NET0131  ;
  input \P2_datao_reg[12]/NET0131  ;
  input \P2_datao_reg[13]/NET0131  ;
  input \P2_datao_reg[14]/NET0131  ;
  input \P2_datao_reg[15]/NET0131  ;
  input \P2_datao_reg[16]/NET0131  ;
  input \P2_datao_reg[17]/NET0131  ;
  input \P2_datao_reg[18]/NET0131  ;
  input \P2_datao_reg[19]/NET0131  ;
  input \P2_datao_reg[1]/NET0131  ;
  input \P2_datao_reg[20]/NET0131  ;
  input \P2_datao_reg[21]/NET0131  ;
  input \P2_datao_reg[22]/NET0131  ;
  input \P2_datao_reg[23]/NET0131  ;
  input \P2_datao_reg[24]/NET0131  ;
  input \P2_datao_reg[25]/NET0131  ;
  input \P2_datao_reg[26]/NET0131  ;
  input \P2_datao_reg[27]/NET0131  ;
  input \P2_datao_reg[28]/NET0131  ;
  input \P2_datao_reg[29]/NET0131  ;
  input \P2_datao_reg[2]/NET0131  ;
  input \P2_datao_reg[30]/NET0131  ;
  input \P2_datao_reg[31]/NET0131  ;
  input \P2_datao_reg[3]/NET0131  ;
  input \P2_datao_reg[4]/NET0131  ;
  input \P2_datao_reg[5]/NET0131  ;
  input \P2_datao_reg[6]/NET0131  ;
  input \P2_datao_reg[7]/NET0131  ;
  input \P2_datao_reg[8]/NET0131  ;
  input \P2_datao_reg[9]/NET0131  ;
  input \P2_rd_reg/NET0131  ;
  input \P2_reg0_reg[0]/NET0131  ;
  input \P2_reg0_reg[10]/NET0131  ;
  input \P2_reg0_reg[11]/NET0131  ;
  input \P2_reg0_reg[12]/NET0131  ;
  input \P2_reg0_reg[13]/NET0131  ;
  input \P2_reg0_reg[14]/NET0131  ;
  input \P2_reg0_reg[15]/NET0131  ;
  input \P2_reg0_reg[16]/NET0131  ;
  input \P2_reg0_reg[17]/NET0131  ;
  input \P2_reg0_reg[18]/NET0131  ;
  input \P2_reg0_reg[19]/NET0131  ;
  input \P2_reg0_reg[1]/NET0131  ;
  input \P2_reg0_reg[20]/NET0131  ;
  input \P2_reg0_reg[21]/NET0131  ;
  input \P2_reg0_reg[22]/NET0131  ;
  input \P2_reg0_reg[23]/NET0131  ;
  input \P2_reg0_reg[24]/NET0131  ;
  input \P2_reg0_reg[25]/NET0131  ;
  input \P2_reg0_reg[26]/NET0131  ;
  input \P2_reg0_reg[27]/NET0131  ;
  input \P2_reg0_reg[28]/NET0131  ;
  input \P2_reg0_reg[29]/NET0131  ;
  input \P2_reg0_reg[2]/NET0131  ;
  input \P2_reg0_reg[30]/NET0131  ;
  input \P2_reg0_reg[31]/NET0131  ;
  input \P2_reg0_reg[3]/NET0131  ;
  input \P2_reg0_reg[4]/NET0131  ;
  input \P2_reg0_reg[5]/NET0131  ;
  input \P2_reg0_reg[6]/NET0131  ;
  input \P2_reg0_reg[7]/NET0131  ;
  input \P2_reg0_reg[8]/NET0131  ;
  input \P2_reg0_reg[9]/NET0131  ;
  input \P2_reg1_reg[0]/NET0131  ;
  input \P2_reg1_reg[10]/NET0131  ;
  input \P2_reg1_reg[11]/NET0131  ;
  input \P2_reg1_reg[12]/NET0131  ;
  input \P2_reg1_reg[13]/NET0131  ;
  input \P2_reg1_reg[14]/NET0131  ;
  input \P2_reg1_reg[15]/NET0131  ;
  input \P2_reg1_reg[16]/NET0131  ;
  input \P2_reg1_reg[17]/NET0131  ;
  input \P2_reg1_reg[18]/NET0131  ;
  input \P2_reg1_reg[19]/NET0131  ;
  input \P2_reg1_reg[1]/NET0131  ;
  input \P2_reg1_reg[20]/NET0131  ;
  input \P2_reg1_reg[21]/NET0131  ;
  input \P2_reg1_reg[22]/NET0131  ;
  input \P2_reg1_reg[23]/NET0131  ;
  input \P2_reg1_reg[24]/NET0131  ;
  input \P2_reg1_reg[25]/NET0131  ;
  input \P2_reg1_reg[26]/NET0131  ;
  input \P2_reg1_reg[27]/NET0131  ;
  input \P2_reg1_reg[28]/NET0131  ;
  input \P2_reg1_reg[29]/NET0131  ;
  input \P2_reg1_reg[2]/NET0131  ;
  input \P2_reg1_reg[30]/NET0131  ;
  input \P2_reg1_reg[31]/NET0131  ;
  input \P2_reg1_reg[3]/NET0131  ;
  input \P2_reg1_reg[4]/NET0131  ;
  input \P2_reg1_reg[5]/NET0131  ;
  input \P2_reg1_reg[6]/NET0131  ;
  input \P2_reg1_reg[7]/NET0131  ;
  input \P2_reg1_reg[8]/NET0131  ;
  input \P2_reg1_reg[9]/NET0131  ;
  input \P2_reg2_reg[0]/NET0131  ;
  input \P2_reg2_reg[10]/NET0131  ;
  input \P2_reg2_reg[11]/NET0131  ;
  input \P2_reg2_reg[12]/NET0131  ;
  input \P2_reg2_reg[13]/NET0131  ;
  input \P2_reg2_reg[14]/NET0131  ;
  input \P2_reg2_reg[15]/NET0131  ;
  input \P2_reg2_reg[16]/NET0131  ;
  input \P2_reg2_reg[17]/NET0131  ;
  input \P2_reg2_reg[18]/NET0131  ;
  input \P2_reg2_reg[19]/NET0131  ;
  input \P2_reg2_reg[1]/NET0131  ;
  input \P2_reg2_reg[20]/NET0131  ;
  input \P2_reg2_reg[21]/NET0131  ;
  input \P2_reg2_reg[22]/NET0131  ;
  input \P2_reg2_reg[23]/NET0131  ;
  input \P2_reg2_reg[24]/NET0131  ;
  input \P2_reg2_reg[25]/NET0131  ;
  input \P2_reg2_reg[26]/NET0131  ;
  input \P2_reg2_reg[27]/NET0131  ;
  input \P2_reg2_reg[28]/NET0131  ;
  input \P2_reg2_reg[29]/NET0131  ;
  input \P2_reg2_reg[2]/NET0131  ;
  input \P2_reg2_reg[30]/NET0131  ;
  input \P2_reg2_reg[31]/NET0131  ;
  input \P2_reg2_reg[3]/NET0131  ;
  input \P2_reg2_reg[4]/NET0131  ;
  input \P2_reg2_reg[5]/NET0131  ;
  input \P2_reg2_reg[6]/NET0131  ;
  input \P2_reg2_reg[7]/NET0131  ;
  input \P2_reg2_reg[8]/NET0131  ;
  input \P2_reg2_reg[9]/NET0131  ;
  input \P2_reg3_reg[0]/NET0131  ;
  input \P2_reg3_reg[10]/NET0131  ;
  input \P2_reg3_reg[11]/NET0131  ;
  input \P2_reg3_reg[12]/NET0131  ;
  input \P2_reg3_reg[13]/NET0131  ;
  input \P2_reg3_reg[14]/NET0131  ;
  input \P2_reg3_reg[15]/NET0131  ;
  input \P2_reg3_reg[16]/NET0131  ;
  input \P2_reg3_reg[17]/NET0131  ;
  input \P2_reg3_reg[18]/NET0131  ;
  input \P2_reg3_reg[19]/NET0131  ;
  input \P2_reg3_reg[1]/NET0131  ;
  input \P2_reg3_reg[20]/NET0131  ;
  input \P2_reg3_reg[21]/NET0131  ;
  input \P2_reg3_reg[22]/NET0131  ;
  input \P2_reg3_reg[23]/NET0131  ;
  input \P2_reg3_reg[24]/NET0131  ;
  input \P2_reg3_reg[25]/NET0131  ;
  input \P2_reg3_reg[26]/NET0131  ;
  input \P2_reg3_reg[27]/NET0131  ;
  input \P2_reg3_reg[28]/NET0131  ;
  input \P2_reg3_reg[2]/NET0131  ;
  input \P2_reg3_reg[3]/NET0131  ;
  input \P2_reg3_reg[4]/NET0131  ;
  input \P2_reg3_reg[5]/NET0131  ;
  input \P2_reg3_reg[6]/NET0131  ;
  input \P2_reg3_reg[7]/NET0131  ;
  input \P2_reg3_reg[8]/NET0131  ;
  input \P2_reg3_reg[9]/NET0131  ;
  input \P2_wr_reg/NET0131  ;
  input \P3_B_reg/NET0131  ;
  input \P3_IR_reg[0]/NET0131  ;
  input \P3_IR_reg[10]/NET0131  ;
  input \P3_IR_reg[11]/NET0131  ;
  input \P3_IR_reg[12]/NET0131  ;
  input \P3_IR_reg[13]/NET0131  ;
  input \P3_IR_reg[14]/NET0131  ;
  input \P3_IR_reg[15]/NET0131  ;
  input \P3_IR_reg[16]/NET0131  ;
  input \P3_IR_reg[17]/NET0131  ;
  input \P3_IR_reg[18]/NET0131  ;
  input \P3_IR_reg[19]/NET0131  ;
  input \P3_IR_reg[1]/NET0131  ;
  input \P3_IR_reg[20]/NET0131  ;
  input \P3_IR_reg[21]/NET0131  ;
  input \P3_IR_reg[22]/NET0131  ;
  input \P3_IR_reg[23]/NET0131  ;
  input \P3_IR_reg[24]/NET0131  ;
  input \P3_IR_reg[25]/NET0131  ;
  input \P3_IR_reg[26]/NET0131  ;
  input \P3_IR_reg[27]/NET0131  ;
  input \P3_IR_reg[28]/NET0131  ;
  input \P3_IR_reg[29]/NET0131  ;
  input \P3_IR_reg[2]/NET0131  ;
  input \P3_IR_reg[30]/NET0131  ;
  input \P3_IR_reg[31]/NET0131  ;
  input \P3_IR_reg[3]/NET0131  ;
  input \P3_IR_reg[4]/NET0131  ;
  input \P3_IR_reg[5]/NET0131  ;
  input \P3_IR_reg[6]/NET0131  ;
  input \P3_IR_reg[7]/NET0131  ;
  input \P3_IR_reg[8]/NET0131  ;
  input \P3_IR_reg[9]/NET0131  ;
  input \P3_addr_reg[0]/NET0131  ;
  input \P3_addr_reg[10]/NET0131  ;
  input \P3_addr_reg[11]/NET0131  ;
  input \P3_addr_reg[12]/NET0131  ;
  input \P3_addr_reg[13]/NET0131  ;
  input \P3_addr_reg[14]/NET0131  ;
  input \P3_addr_reg[15]/NET0131  ;
  input \P3_addr_reg[16]/NET0131  ;
  input \P3_addr_reg[17]/NET0131  ;
  input \P3_addr_reg[18]/NET0131  ;
  input \P3_addr_reg[19]/NET0131  ;
  input \P3_addr_reg[1]/NET0131  ;
  input \P3_addr_reg[2]/NET0131  ;
  input \P3_addr_reg[3]/NET0131  ;
  input \P3_addr_reg[4]/NET0131  ;
  input \P3_addr_reg[5]/NET0131  ;
  input \P3_addr_reg[6]/NET0131  ;
  input \P3_addr_reg[7]/NET0131  ;
  input \P3_addr_reg[8]/NET0131  ;
  input \P3_addr_reg[9]/NET0131  ;
  input \P3_d_reg[0]/NET0131  ;
  input \P3_d_reg[1]/NET0131  ;
  input \P3_rd_reg/NET0131  ;
  input \P3_reg0_reg[0]/NET0131  ;
  input \P3_reg0_reg[10]/NET0131  ;
  input \P3_reg0_reg[11]/NET0131  ;
  input \P3_reg0_reg[12]/NET0131  ;
  input \P3_reg0_reg[13]/NET0131  ;
  input \P3_reg0_reg[14]/NET0131  ;
  input \P3_reg0_reg[15]/NET0131  ;
  input \P3_reg0_reg[16]/NET0131  ;
  input \P3_reg0_reg[17]/NET0131  ;
  input \P3_reg0_reg[18]/NET0131  ;
  input \P3_reg0_reg[19]/NET0131  ;
  input \P3_reg0_reg[1]/NET0131  ;
  input \P3_reg0_reg[20]/NET0131  ;
  input \P3_reg0_reg[21]/NET0131  ;
  input \P3_reg0_reg[22]/NET0131  ;
  input \P3_reg0_reg[23]/NET0131  ;
  input \P3_reg0_reg[24]/NET0131  ;
  input \P3_reg0_reg[25]/NET0131  ;
  input \P3_reg0_reg[26]/NET0131  ;
  input \P3_reg0_reg[27]/NET0131  ;
  input \P3_reg0_reg[28]/NET0131  ;
  input \P3_reg0_reg[29]/NET0131  ;
  input \P3_reg0_reg[2]/NET0131  ;
  input \P3_reg0_reg[30]/NET0131  ;
  input \P3_reg0_reg[31]/NET0131  ;
  input \P3_reg0_reg[3]/NET0131  ;
  input \P3_reg0_reg[4]/NET0131  ;
  input \P3_reg0_reg[5]/NET0131  ;
  input \P3_reg0_reg[6]/NET0131  ;
  input \P3_reg0_reg[7]/NET0131  ;
  input \P3_reg0_reg[8]/NET0131  ;
  input \P3_reg0_reg[9]/NET0131  ;
  input \P3_reg1_reg[0]/NET0131  ;
  input \P3_reg1_reg[10]/NET0131  ;
  input \P3_reg1_reg[11]/NET0131  ;
  input \P3_reg1_reg[12]/NET0131  ;
  input \P3_reg1_reg[13]/NET0131  ;
  input \P3_reg1_reg[14]/NET0131  ;
  input \P3_reg1_reg[15]/NET0131  ;
  input \P3_reg1_reg[16]/NET0131  ;
  input \P3_reg1_reg[17]/NET0131  ;
  input \P3_reg1_reg[18]/NET0131  ;
  input \P3_reg1_reg[19]/NET0131  ;
  input \P3_reg1_reg[1]/NET0131  ;
  input \P3_reg1_reg[20]/NET0131  ;
  input \P3_reg1_reg[21]/NET0131  ;
  input \P3_reg1_reg[22]/NET0131  ;
  input \P3_reg1_reg[23]/NET0131  ;
  input \P3_reg1_reg[24]/NET0131  ;
  input \P3_reg1_reg[25]/NET0131  ;
  input \P3_reg1_reg[26]/NET0131  ;
  input \P3_reg1_reg[27]/NET0131  ;
  input \P3_reg1_reg[28]/NET0131  ;
  input \P3_reg1_reg[29]/NET0131  ;
  input \P3_reg1_reg[2]/NET0131  ;
  input \P3_reg1_reg[30]/NET0131  ;
  input \P3_reg1_reg[31]/NET0131  ;
  input \P3_reg1_reg[3]/NET0131  ;
  input \P3_reg1_reg[4]/NET0131  ;
  input \P3_reg1_reg[5]/NET0131  ;
  input \P3_reg1_reg[6]/NET0131  ;
  input \P3_reg1_reg[7]/NET0131  ;
  input \P3_reg1_reg[8]/NET0131  ;
  input \P3_reg1_reg[9]/NET0131  ;
  input \P3_reg2_reg[0]/NET0131  ;
  input \P3_reg2_reg[10]/NET0131  ;
  input \P3_reg2_reg[11]/NET0131  ;
  input \P3_reg2_reg[12]/NET0131  ;
  input \P3_reg2_reg[13]/NET0131  ;
  input \P3_reg2_reg[14]/NET0131  ;
  input \P3_reg2_reg[15]/NET0131  ;
  input \P3_reg2_reg[16]/NET0131  ;
  input \P3_reg2_reg[17]/NET0131  ;
  input \P3_reg2_reg[18]/NET0131  ;
  input \P3_reg2_reg[19]/NET0131  ;
  input \P3_reg2_reg[1]/NET0131  ;
  input \P3_reg2_reg[20]/NET0131  ;
  input \P3_reg2_reg[21]/NET0131  ;
  input \P3_reg2_reg[22]/NET0131  ;
  input \P3_reg2_reg[23]/NET0131  ;
  input \P3_reg2_reg[24]/NET0131  ;
  input \P3_reg2_reg[25]/NET0131  ;
  input \P3_reg2_reg[26]/NET0131  ;
  input \P3_reg2_reg[27]/NET0131  ;
  input \P3_reg2_reg[28]/NET0131  ;
  input \P3_reg2_reg[29]/NET0131  ;
  input \P3_reg2_reg[2]/NET0131  ;
  input \P3_reg2_reg[30]/NET0131  ;
  input \P3_reg2_reg[31]/NET0131  ;
  input \P3_reg2_reg[3]/NET0131  ;
  input \P3_reg2_reg[4]/NET0131  ;
  input \P3_reg2_reg[5]/NET0131  ;
  input \P3_reg2_reg[6]/NET0131  ;
  input \P3_reg2_reg[7]/NET0131  ;
  input \P3_reg2_reg[8]/NET0131  ;
  input \P3_reg2_reg[9]/NET0131  ;
  input \P3_reg3_reg[0]/NET0131  ;
  input \P3_reg3_reg[10]/NET0131  ;
  input \P3_reg3_reg[11]/NET0131  ;
  input \P3_reg3_reg[12]/NET0131  ;
  input \P3_reg3_reg[13]/NET0131  ;
  input \P3_reg3_reg[14]/NET0131  ;
  input \P3_reg3_reg[15]/NET0131  ;
  input \P3_reg3_reg[16]/NET0131  ;
  input \P3_reg3_reg[17]/NET0131  ;
  input \P3_reg3_reg[18]/NET0131  ;
  input \P3_reg3_reg[19]/NET0131  ;
  input \P3_reg3_reg[1]/NET0131  ;
  input \P3_reg3_reg[20]/NET0131  ;
  input \P3_reg3_reg[21]/NET0131  ;
  input \P3_reg3_reg[22]/NET0131  ;
  input \P3_reg3_reg[23]/NET0131  ;
  input \P3_reg3_reg[24]/NET0131  ;
  input \P3_reg3_reg[25]/NET0131  ;
  input \P3_reg3_reg[26]/NET0131  ;
  input \P3_reg3_reg[27]/NET0131  ;
  input \P3_reg3_reg[28]/NET0131  ;
  input \P3_reg3_reg[2]/NET0131  ;
  input \P3_reg3_reg[3]/NET0131  ;
  input \P3_reg3_reg[4]/NET0131  ;
  input \P3_reg3_reg[5]/NET0131  ;
  input \P3_reg3_reg[6]/NET0131  ;
  input \P3_reg3_reg[7]/NET0131  ;
  input \P3_reg3_reg[8]/NET0131  ;
  input \P3_reg3_reg[9]/NET0131  ;
  input \P3_wr_reg/NET0131  ;
  input \si[0]_pad  ;
  input \si[10]_pad  ;
  input \si[11]_pad  ;
  input \si[12]_pad  ;
  input \si[13]_pad  ;
  input \si[14]_pad  ;
  input \si[15]_pad  ;
  input \si[16]_pad  ;
  input \si[17]_pad  ;
  input \si[18]_pad  ;
  input \si[19]_pad  ;
  input \si[1]_pad  ;
  input \si[20]_pad  ;
  input \si[21]_pad  ;
  input \si[22]_pad  ;
  input \si[23]_pad  ;
  input \si[24]_pad  ;
  input \si[25]_pad  ;
  input \si[26]_pad  ;
  input \si[27]_pad  ;
  input \si[28]_pad  ;
  input \si[29]_pad  ;
  input \si[2]_pad  ;
  input \si[30]_pad  ;
  input \si[31]_pad  ;
  input \si[3]_pad  ;
  input \si[4]_pad  ;
  input \si[5]_pad  ;
  input \si[6]_pad  ;
  input \si[7]_pad  ;
  input \si[8]_pad  ;
  input \si[9]_pad  ;
  output \P1_state_reg[0]/NET0131_syn_2  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g106254/_0_  ;
  output \g106255/_0_  ;
  output \g106267/_0_  ;
  output \g106268/_0_  ;
  output \g106269/_0_  ;
  output \g106270/_0_  ;
  output \g106271/_0_  ;
  output \g106272/_0_  ;
  output \g106288/_0_  ;
  output \g106289/_0_  ;
  output \g106290/_0_  ;
  output \g106291/_0_  ;
  output \g106292/_0_  ;
  output \g106293/_0_  ;
  output \g106294/_0_  ;
  output \g106295/_0_  ;
  output \g106296/_0_  ;
  output \g106297/_0_  ;
  output \g106352/_0_  ;
  output \g106356/_0_  ;
  output \g106359/_0_  ;
  output \g106360/_0_  ;
  output \g106361/_0_  ;
  output \g106362/_0_  ;
  output \g106363/_0_  ;
  output \g106364/_0_  ;
  output \g106365/_0_  ;
  output \g106406/_0_  ;
  output \g106407/_0_  ;
  output \g106408/_0_  ;
  output \g106410/_0_  ;
  output \g106411/_0_  ;
  output \g106412/_0_  ;
  output \g106413/_0_  ;
  output \g106414/_0_  ;
  output \g106417/_0_  ;
  output \g106418/_0_  ;
  output \g106419/_0_  ;
  output \g106420/_0_  ;
  output \g106421/_0_  ;
  output \g106422/_0_  ;
  output \g106423/_0_  ;
  output \g106424/_0_  ;
  output \g106425/_0_  ;
  output \g106426/_0_  ;
  output \g106427/_0_  ;
  output \g106428/_0_  ;
  output \g106430/_0_  ;
  output \g106431/_0_  ;
  output \g106432/_0_  ;
  output \g106433/_0_  ;
  output \g106434/_0_  ;
  output \g106436/_0_  ;
  output \g106437/_0_  ;
  output \g106438/_0_  ;
  output \g106439/_0_  ;
  output \g106440/_0_  ;
  output \g106441/_0_  ;
  output \g106442/_0_  ;
  output \g106443/_0_  ;
  output \g106444/_0_  ;
  output \g106445/_0_  ;
  output \g106446/_0_  ;
  output \g106447/_0_  ;
  output \g106448/_0_  ;
  output \g106530/_0_  ;
  output \g106531/_0_  ;
  output \g106532/_0_  ;
  output \g106533/_0_  ;
  output \g106534/_0_  ;
  output \g106554/_0_  ;
  output \g106556/_0_  ;
  output \g106557/_0_  ;
  output \g106559/_0_  ;
  output \g106560/_0_  ;
  output \g106561/_0_  ;
  output \g106562/_0_  ;
  output \g106563/_0_  ;
  output \g106564/_0_  ;
  output \g106565/_0_  ;
  output \g106566/_0_  ;
  output \g106567/_0_  ;
  output \g106568/_0_  ;
  output \g106569/_0_  ;
  output \g106570/_0_  ;
  output \g106571/_0_  ;
  output \g106572/_0_  ;
  output \g106633/_0_  ;
  output \g106634/_0_  ;
  output \g106640/_0_  ;
  output \g106654/_0_  ;
  output \g106655/_0_  ;
  output \g106679/_0_  ;
  output \g106682/_0_  ;
  output \g106684/_0_  ;
  output \g106687/_0_  ;
  output \g106690/_0_  ;
  output \g106691/_0_  ;
  output \g106692/_0_  ;
  output \g106693/_0_  ;
  output \g106694/_0_  ;
  output \g106695/_0_  ;
  output \g106696/_0_  ;
  output \g106697/_0_  ;
  output \g106698/_0_  ;
  output \g106699/_0_  ;
  output \g106700/_0_  ;
  output \g106701/_0_  ;
  output \g106702/_0_  ;
  output \g106703/_0_  ;
  output \g106704/_0_  ;
  output \g106705/_0_  ;
  output \g106706/_0_  ;
  output \g106707/_0_  ;
  output \g106708/_0_  ;
  output \g106710/_0_  ;
  output \g106711/_0_  ;
  output \g106712/_0_  ;
  output \g106713/_0_  ;
  output \g106714/_0_  ;
  output \g106715/_0_  ;
  output \g106716/_0_  ;
  output \g106717/_0_  ;
  output \g106718/_0_  ;
  output \g106719/_0_  ;
  output \g106720/_0_  ;
  output \g106721/_0_  ;
  output \g106722/_0_  ;
  output \g106723/_0_  ;
  output \g106724/_0_  ;
  output \g106725/_0_  ;
  output \g106726/_0_  ;
  output \g106727/_0_  ;
  output \g106728/_0_  ;
  output \g106729/_0_  ;
  output \g106830/_0_  ;
  output \g106836/_0_  ;
  output \g106837/_0_  ;
  output \g106838/_0_  ;
  output \g106843/_0_  ;
  output \g106850/_0_  ;
  output \g106851/_0_  ;
  output \g106852/_0_  ;
  output \g106853/_0_  ;
  output \g106854/_0_  ;
  output \g106899/_0_  ;
  output \g106901/_0_  ;
  output \g106902/_0_  ;
  output \g106903/_0_  ;
  output \g106904/_0_  ;
  output \g106905/_0_  ;
  output \g106906/_0_  ;
  output \g106907/_0_  ;
  output \g106908/_0_  ;
  output \g106909/_0_  ;
  output \g106910/_0_  ;
  output \g106911/_0_  ;
  output \g106912/_0_  ;
  output \g106913/_0_  ;
  output \g106914/_0_  ;
  output \g106915/_0_  ;
  output \g106916/_0_  ;
  output \g106917/_0_  ;
  output \g106918/_0_  ;
  output \g106919/_0_  ;
  output \g106920/_0_  ;
  output \g106921/_0_  ;
  output \g106922/_0_  ;
  output \g106923/_0_  ;
  output \g106924/_0_  ;
  output \g106925/_0_  ;
  output \g106994/_0_  ;
  output \g106995/_0_  ;
  output \g106996/_0_  ;
  output \g106997/_0_  ;
  output \g106998/_0_  ;
  output \g106999/_0_  ;
  output \g107002/_0_  ;
  output \g107007/_0_  ;
  output \g107008/_0_  ;
  output \g107038/_0_  ;
  output \g107041/_0_  ;
  output \g107048/_0_  ;
  output \g107091/_0_  ;
  output \g107093/_0_  ;
  output \g107094/_0_  ;
  output \g107096/_0_  ;
  output \g107097/_0_  ;
  output \g107098/_0_  ;
  output \g107099/_0_  ;
  output \g107100/_0_  ;
  output \g107101/_0_  ;
  output \g107102/_0_  ;
  output \g107103/_0_  ;
  output \g107104/_0_  ;
  output \g107105/_0_  ;
  output \g107106/_0_  ;
  output \g107107/_0_  ;
  output \g107108/_0_  ;
  output \g107109/_0_  ;
  output \g107110/_0_  ;
  output \g107111/_0_  ;
  output \g107112/_0_  ;
  output \g107113/_0_  ;
  output \g107114/_0_  ;
  output \g107115/_0_  ;
  output \g107116/_0_  ;
  output \g107117/_0_  ;
  output \g107118/_0_  ;
  output \g107119/_0_  ;
  output \g107120/_0_  ;
  output \g107121/_0_  ;
  output \g107122/_0_  ;
  output \g107123/_0_  ;
  output \g107124/_0_  ;
  output \g107125/_0_  ;
  output \g107126/_0_  ;
  output \g107127/_0_  ;
  output \g107128/_0_  ;
  output \g107129/_0_  ;
  output \g107130/_0_  ;
  output \g107131/_0_  ;
  output \g107132/_0_  ;
  output \g107133/_0_  ;
  output \g107134/_0_  ;
  output \g107135/_0_  ;
  output \g107136/_0_  ;
  output \g107137/_0_  ;
  output \g107138/_0_  ;
  output \g107248/_0_  ;
  output \g107252/_0_  ;
  output \g107254/_0_  ;
  output \g107255/_0_  ;
  output \g107280/_0_  ;
  output \g107281/_0_  ;
  output \g107282/_0_  ;
  output \g107370/_0_  ;
  output \g107371/_0_  ;
  output \g107372/_0_  ;
  output \g107373/_0_  ;
  output \g107374/_0_  ;
  output \g107375/_0_  ;
  output \g107376/_0_  ;
  output \g107377/_0_  ;
  output \g107378/_0_  ;
  output \g107379/_0_  ;
  output \g107380/_0_  ;
  output \g107381/_0_  ;
  output \g107382/_0_  ;
  output \g107383/_0_  ;
  output \g107384/_0_  ;
  output \g107385/_0_  ;
  output \g107386/_0_  ;
  output \g107387/_0_  ;
  output \g107388/_0_  ;
  output \g107389/_0_  ;
  output \g107390/_0_  ;
  output \g107391/_0_  ;
  output \g107488/_0_  ;
  output \g107489/_0_  ;
  output \g107490/_0_  ;
  output \g107491/_0_  ;
  output \g107492/_0_  ;
  output \g107493/_0_  ;
  output \g107500/_0_  ;
  output \g107615/_0_  ;
  output \g107623/_0_  ;
  output \g107624/_0_  ;
  output \g107625/_0_  ;
  output \g107626/_0_  ;
  output \g107627/_0_  ;
  output \g107628/_0_  ;
  output \g107629/_0_  ;
  output \g107630/_0_  ;
  output \g107631/_0_  ;
  output \g107632/_0_  ;
  output \g107634/_0_  ;
  output \g107637/_0_  ;
  output \g107638/_0_  ;
  output \g107639/_0_  ;
  output \g107640/_0_  ;
  output \g107641/_0_  ;
  output \g107642/_0_  ;
  output \g107643/_0_  ;
  output \g107644/_0_  ;
  output \g107645/_0_  ;
  output \g107646/_0_  ;
  output \g107647/_0_  ;
  output \g107650/_0_  ;
  output \g107651/_0_  ;
  output \g107652/_0_  ;
  output \g107653/_0_  ;
  output \g107654/_0_  ;
  output \g107655/_0_  ;
  output \g107656/_0_  ;
  output \g107743/_0_  ;
  output \g107787/_0_  ;
  output \g107954/_0_  ;
  output \g107955/_0_  ;
  output \g107956/_0_  ;
  output \g107957/_0_  ;
  output \g107958/_0_  ;
  output \g107959/_0_  ;
  output \g107960/_0_  ;
  output \g107961/_0_  ;
  output \g107962/_0_  ;
  output \g107963/_0_  ;
  output \g107964/_0_  ;
  output \g107965/_0_  ;
  output \g107966/_0_  ;
  output \g107967/_0_  ;
  output \g108118/_0_  ;
  output \g108125/_0_  ;
  output \g108169/_0_  ;
  output \g108269/_0_  ;
  output \g108270/_0_  ;
  output \g108319/_0_  ;
  output \g108320/_0_  ;
  output \g108321/_0_  ;
  output \g108322/_0_  ;
  output \g108323/_0_  ;
  output \g108324/_0_  ;
  output \g108326/_0_  ;
  output \g108327/_0_  ;
  output \g108328/_0_  ;
  output \g108329/_0_  ;
  output \g108330/_0_  ;
  output \g108334/_0_  ;
  output \g108335/_0_  ;
  output \g108468/_0_  ;
  output \g108538/_0_  ;
  output \g108801/_0_  ;
  output \g108812/_0_  ;
  output \g108813/_0_  ;
  output \g108814/_0_  ;
  output \g108815/_0_  ;
  output \g108817/_0_  ;
  output \g108818/_0_  ;
  output \g108819/_0_  ;
  output \g108822/_0_  ;
  output \g109052/_0_  ;
  output \g109053/_0_  ;
  output \g109401/_0_  ;
  output \g109402/_0_  ;
  output \g109403/_0_  ;
  output \g109410/_0_  ;
  output \g109411/_0_  ;
  output \g109415/_0_  ;
  output \g109420/_0_  ;
  output \g109425/_0_  ;
  output \g109693/_0_  ;
  output \g110116/_0_  ;
  output \g110117/_0_  ;
  output \g110905/_0_  ;
  output \g110906/_0_  ;
  output \g110907/_0_  ;
  output \g111086/_0_  ;
  output \g111094/_0_  ;
  output \g112422/_0_  ;
  output \g112423/_0_  ;
  output \g112424/_0_  ;
  output \g112425/_0_  ;
  output \g112426/_0_  ;
  output \g112427/_0_  ;
  output \g113647/_0_  ;
  output \g113648/_0_  ;
  output \g113649/_0_  ;
  output \g113650/_0_  ;
  output \g113651/_0_  ;
  output \g114133/_0_  ;
  output \g117884/_0_  ;
  output \g117885/_0_  ;
  output \g117886/_0_  ;
  output \g117895/_3_  ;
  output \g117896/_3_  ;
  output \g117897/_0_  ;
  output \g117898/_0_  ;
  output \g117899/_0_  ;
  output \g117900/_3_  ;
  output \g120982/_0_  ;
  output \g120983/_0_  ;
  output \g120984/_0_  ;
  output \g120985/_0_  ;
  output \g120986/_0_  ;
  output \g120987/_0_  ;
  output \g120988/_3_  ;
  output \g120989/_0_  ;
  output \g120990/_0_  ;
  output \g120991/_0_  ;
  output \g120992/_0_  ;
  output \g120993/_0_  ;
  output \g120994/_0_  ;
  output \g120995/_0_  ;
  output \g120996/_3_  ;
  output \g120997/_0_  ;
  output \g120998/_0_  ;
  output \g120999/_0_  ;
  output \g121000/_0_  ;
  output \g121001/_0_  ;
  output \g121002/_3_  ;
  output \g121003/_0_  ;
  output \g121004/_0_  ;
  output \g121005/_3_  ;
  output \g121006/_0_  ;
  output \g121007/_0_  ;
  output \g121008/_0_  ;
  output \g121029/_0_  ;
  output \g121030/_3_  ;
  output \g121032/_3_  ;
  output \g121033/_3_  ;
  output \g121034/_3_  ;
  output \g121035/_3_  ;
  output \g121036/_3_  ;
  output \g121037/_3_  ;
  output \g121038/_3_  ;
  output \g121039/_3_  ;
  output \g121040/_3_  ;
  output \g121041/_3_  ;
  output \g121042/_3_  ;
  output \g121043/_3_  ;
  output \g121044/_3_  ;
  output \g121045/_3_  ;
  output \g121046/_3_  ;
  output \g121047/_3_  ;
  output \g121048/_3_  ;
  output \g121049/_3_  ;
  output \g121050/_3_  ;
  output \g121051/_0_  ;
  output \g121052/_3_  ;
  output \g121053/_3_  ;
  output \g121054/_3_  ;
  output \g121055/_3_  ;
  output \g121056/_3_  ;
  output \g121057/_3_  ;
  output \g121058/_3_  ;
  output \g121060/_3_  ;
  output \g121061/_3_  ;
  output \g121062/_3_  ;
  output \g121063/_3_  ;
  output \g121064/_3_  ;
  output \g121065/_3_  ;
  output \g121066/_3_  ;
  output \g121067/_3_  ;
  output \g121068/_3_  ;
  output \g121069/_3_  ;
  output \g121070/_3_  ;
  output \g121071/_3_  ;
  output \g121072/_3_  ;
  output \g121073/_3_  ;
  output \g121074/_3_  ;
  output \g121075/_3_  ;
  output \g121076/_3_  ;
  output \g121077/_3_  ;
  output \g121078/_3_  ;
  output \g121079/_3_  ;
  output \g121080/_0_  ;
  output \g121081/_3_  ;
  output \g121082/_0_  ;
  output \g121083/_3_  ;
  output \g121084/_3_  ;
  output \g121085/_3_  ;
  output \g121086/_3_  ;
  output \g121087/_3_  ;
  output \g121626/_0_  ;
  output \g121633/_0_  ;
  output \g121669/_0_  ;
  output \g122948/_0_  ;
  output \g122949/_0_  ;
  output \g122951/_0_  ;
  output \g122952/_0_  ;
  output \g122953/_0_  ;
  output \g122954/_0_  ;
  output \g122955/_0_  ;
  output \g122956/_0_  ;
  output \g122957/_0_  ;
  output \g122958/_0_  ;
  output \g122959/_0_  ;
  output \g122960/_0_  ;
  output \g122963/_0_  ;
  output \g122965/_0_  ;
  output \g122967/_0_  ;
  output \g122968/_0_  ;
  output \g122972/_0_  ;
  output \g122973/_0_  ;
  output \g122974/_0_  ;
  output \g122975/_0_  ;
  output \g122976/_0_  ;
  output \g122977/_0_  ;
  output \g122978/_0_  ;
  output \g122979/_0_  ;
  output \g122980/_0_  ;
  output \g122981/_0_  ;
  output \g122982/_0_  ;
  output \g122983/_0_  ;
  output \g122984/_0_  ;
  output \g122985/_0_  ;
  output \g122986/_0_  ;
  output \g122987/_0_  ;
  output \g122988/_0_  ;
  output \g122989/_0_  ;
  output \g122990/_0_  ;
  output \g122991/_0_  ;
  output \g122997/_0_  ;
  output \g122998/_0_  ;
  output \g122999/_0_  ;
  output \g123000/_0_  ;
  output \g123740/_0_  ;
  output \g123811/_0_  ;
  output \g123812/_0_  ;
  output \g123813/_0_  ;
  output \g123814/_0_  ;
  output \g123815/_0_  ;
  output \g123816/_0_  ;
  output \g123817/_0_  ;
  output \g123818/_0_  ;
  output \g123819/_0_  ;
  output \g123820/_0_  ;
  output \g123821/_0_  ;
  output \g123822/_0_  ;
  output \g123823/_0_  ;
  output \g123824/_0_  ;
  output \g123825/_0_  ;
  output \g123826/_0_  ;
  output \g123827/_0_  ;
  output \g123828/_0_  ;
  output \g123829/_0_  ;
  output \g123830/_0_  ;
  output \g123853/u3_syn_4  ;
  output \g123854/u3_syn_4  ;
  output \g123871/_0_  ;
  output \g124519/_0_  ;
  output \g124554/_0_  ;
  output \g124798/_0_  ;
  output \g124897/_0_  ;
  output \g125133/_0_  ;
  output \g125231/_0_  ;
  output \g125318/u3_syn_4  ;
  output \g125495/u3_syn_4  ;
  output \g126480/_0_  ;
  output \g126501/_0_  ;
  output \g127137/_0_  ;
  output \g127147/_0_  ;
  output \g127163/_0_  ;
  output \g127173/_0_  ;
  output \g127202/_0_  ;
  output \g127211/_0_  ;
  output \g127223/_0_  ;
  output \g127234/_0_  ;
  output \g127241/_0_  ;
  output \g127251/_0_  ;
  output \g127257/_0_  ;
  output \g127262/_0_  ;
  output \g127271/_0_  ;
  output \g127285/_0_  ;
  output \g127292/_0_  ;
  output \g127302/_0_  ;
  output \g127313/_0_  ;
  output \g127324/_0_  ;
  output \g127334/_0_  ;
  output \g127348/_0_  ;
  output \g127366/_0_  ;
  output \g127396/_0_  ;
  output \g127405/_0_  ;
  output \g127411/_0_  ;
  output \g127427/_0_  ;
  output \g127439/_0_  ;
  output \g127464/_0_  ;
  output \g127893/_0_  ;
  output \g128290/_0_  ;
  output \g128431/_0_  ;
  output \g128477/_0_  ;
  output \g128501/_0_  ;
  output \g128540/_0_  ;
  output \g128566/_0_  ;
  output \g128575/_0_  ;
  output \g128586/_0_  ;
  output \g128594/_1_  ;
  output \g128631/_0_  ;
  output \g128648/_0_  ;
  output \g128698/_0_  ;
  output \g131281/_1_  ;
  output \g140384/_0_  ;
  output \g140411/_0_  ;
  output \g140627/_0_  ;
  output \g140741/_0_  ;
  output \g140774/_0_  ;
  output \g140804/_0_  ;
  output \g140955/_0_  ;
  output \g140986/_0_  ;
  output \g141163/_0_  ;
  output \g141237/_0_  ;
  output \g141301/_0_  ;
  output \g141328/_0_  ;
  output \g141367/_0_  ;
  output \g141441/_0_  ;
  output \g141474/_0_  ;
  output \g141548/_0_  ;
  output \g141640/_0_  ;
  output \g141838/_0_  ;
  output \g141844/_0_  ;
  output \g141853/_0_  ;
  output \g141855/_0_  ;
  output \g141860/_0_  ;
  output \g141896/_0_  ;
  output \g141915/_0_  ;
  output \g141952/_0_  ;
  output \g142033/_0_  ;
  output \g142046/_0_  ;
  output \g29/_0_  ;
  output \g33/_0_  ;
  output \g53/_0_  ;
  output \g71/_0_  ;
  output \g90/_0_  ;
  output rd_pad ;
  output \so[0]_pad  ;
  output \so[10]_pad  ;
  output \so[11]_pad  ;
  output \so[12]_pad  ;
  output \so[13]_pad  ;
  output \so[14]_pad  ;
  output \so[15]_pad  ;
  output \so[16]_pad  ;
  output \so[17]_pad  ;
  output \so[18]_pad  ;
  output \so[19]_pad  ;
  output \so[1]_pad  ;
  output \so[2]_pad  ;
  output \so[3]_pad  ;
  output \so[4]_pad  ;
  output \so[5]_pad  ;
  output \so[6]_pad  ;
  output \so[7]_pad  ;
  output \so[8]_pad  ;
  output \so[9]_pad  ;
  output wr_pad ;
  wire n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 ;
  assign n644 = ~\P3_IR_reg[0]/NET0131  & ~\P3_IR_reg[1]/NET0131  ;
  assign n645 = ~\P3_IR_reg[2]/NET0131  & ~\P3_IR_reg[3]/NET0131  ;
  assign n646 = n644 & n645 ;
  assign n647 = ~\P3_IR_reg[4]/NET0131  & n646 ;
  assign n648 = ~\P3_IR_reg[5]/NET0131  & n647 ;
  assign n650 = ~\P3_IR_reg[6]/NET0131  & ~\P3_IR_reg[7]/NET0131  ;
  assign n649 = ~\P3_IR_reg[8]/NET0131  & ~\P3_IR_reg[9]/NET0131  ;
  assign n651 = ~\P3_IR_reg[10]/NET0131  & n649 ;
  assign n652 = n650 & n651 ;
  assign n653 = n648 & n652 ;
  assign n654 = ~\P3_IR_reg[12]/NET0131  & ~\P3_IR_reg[13]/NET0131  ;
  assign n655 = ~\P3_IR_reg[11]/NET0131  & ~\P3_IR_reg[14]/NET0131  ;
  assign n656 = n654 & n655 ;
  assign n657 = n653 & n656 ;
  assign n658 = ~\P3_IR_reg[15]/NET0131  & n657 ;
  assign n659 = ~\P3_IR_reg[17]/NET0131  & ~\P3_IR_reg[18]/NET0131  ;
  assign n660 = ~\P3_IR_reg[16]/NET0131  & n659 ;
  assign n661 = n658 & n660 ;
  assign n662 = \P3_IR_reg[31]/NET0131  & ~n661 ;
  assign n663 = ~\P3_IR_reg[20]/NET0131  & ~\P3_IR_reg[21]/NET0131  ;
  assign n664 = ~\P3_IR_reg[19]/NET0131  & n663 ;
  assign n665 = ~\P3_IR_reg[22]/NET0131  & n664 ;
  assign n666 = \P3_IR_reg[31]/NET0131  & ~n665 ;
  assign n667 = ~n662 & ~n666 ;
  assign n668 = \P3_IR_reg[23]/NET0131  & ~n667 ;
  assign n669 = ~\P3_IR_reg[23]/NET0131  & n667 ;
  assign n670 = ~n668 & ~n669 ;
  assign n716 = ~\P3_IR_reg[24]/NET0131  & ~\P3_IR_reg[25]/NET0131  ;
  assign n717 = ~\P3_IR_reg[26]/NET0131  & n716 ;
  assign n715 = ~\P3_IR_reg[22]/NET0131  & ~\P3_IR_reg[23]/NET0131  ;
  assign n718 = n664 & n715 ;
  assign n719 = n717 & n718 ;
  assign n720 = n661 & n719 ;
  assign n721 = \P3_IR_reg[31]/NET0131  & ~n720 ;
  assign n722 = \P3_IR_reg[27]/NET0131  & n721 ;
  assign n723 = ~\P3_IR_reg[27]/NET0131  & ~n721 ;
  assign n724 = ~n722 & ~n723 ;
  assign n671 = ~\P3_IR_reg[10]/NET0131  & ~\P3_IR_reg[11]/NET0131  ;
  assign n672 = ~\P3_IR_reg[5]/NET0131  & n650 ;
  assign n673 = n649 & n672 ;
  assign n674 = n647 & n673 ;
  assign n675 = n671 & n674 ;
  assign n679 = ~\P3_IR_reg[14]/NET0131  & ~\P3_IR_reg[15]/NET0131  ;
  assign n680 = ~\P3_IR_reg[16]/NET0131  & n679 ;
  assign n689 = ~\P3_IR_reg[13]/NET0131  & n680 ;
  assign n678 = ~\P3_IR_reg[19]/NET0131  & n659 ;
  assign n702 = ~\P3_IR_reg[12]/NET0131  & n678 ;
  assign n703 = n689 & n702 ;
  assign n704 = n675 & n703 ;
  assign n725 = n663 & n715 ;
  assign n726 = n704 & n725 ;
  assign n727 = \P3_IR_reg[31]/NET0131  & ~n726 ;
  assign n728 = ~\P3_IR_reg[27]/NET0131  & n717 ;
  assign n729 = \P3_IR_reg[31]/NET0131  & ~n728 ;
  assign n730 = ~n727 & ~n729 ;
  assign n731 = \P3_IR_reg[28]/NET0131  & ~n730 ;
  assign n732 = ~\P3_IR_reg[28]/NET0131  & n730 ;
  assign n733 = ~n731 & ~n732 ;
  assign n734 = ~n724 & n733 ;
  assign n676 = n654 & n675 ;
  assign n677 = \P3_IR_reg[31]/NET0131  & ~n676 ;
  assign n681 = n663 & n678 ;
  assign n682 = n680 & n681 ;
  assign n683 = \P3_IR_reg[31]/NET0131  & ~n682 ;
  assign n684 = ~n677 & ~n683 ;
  assign n685 = \P3_IR_reg[22]/NET0131  & ~n684 ;
  assign n686 = ~\P3_IR_reg[22]/NET0131  & n684 ;
  assign n687 = ~n685 & ~n686 ;
  assign n690 = ~\P3_IR_reg[8]/NET0131  & n672 ;
  assign n691 = n647 & n690 ;
  assign n692 = ~\P3_IR_reg[12]/NET0131  & ~\P3_IR_reg[9]/NET0131  ;
  assign n693 = n671 & n692 ;
  assign n694 = n691 & n693 ;
  assign n695 = n689 & n694 ;
  assign n696 = ~\P3_IR_reg[20]/NET0131  & n678 ;
  assign n697 = n695 & n696 ;
  assign n698 = \P3_IR_reg[31]/NET0131  & ~n697 ;
  assign n699 = \P3_IR_reg[21]/NET0131  & n698 ;
  assign n700 = ~\P3_IR_reg[21]/NET0131  & ~n698 ;
  assign n701 = ~n699 & ~n700 ;
  assign n735 = n687 & ~n701 ;
  assign n705 = \P3_IR_reg[31]/NET0131  & ~n704 ;
  assign n706 = \P3_IR_reg[20]/NET0131  & n705 ;
  assign n707 = ~\P3_IR_reg[20]/NET0131  & ~n705 ;
  assign n708 = ~n706 & ~n707 ;
  assign n736 = n670 & ~n708 ;
  assign n737 = n735 & n736 ;
  assign n738 = ~n734 & n737 ;
  assign n688 = n670 & n687 ;
  assign n711 = n687 & n701 ;
  assign n712 = n670 & n708 ;
  assign n713 = ~n711 & ~n712 ;
  assign n714 = ~n688 & ~n713 ;
  assign n709 = ~n701 & ~n708 ;
  assign n710 = n688 & ~n709 ;
  assign n753 = ~\P3_IR_reg[24]/NET0131  & ~n727 ;
  assign n754 = \P3_IR_reg[24]/NET0131  & n727 ;
  assign n755 = ~n753 & ~n754 ;
  assign n739 = ~\P3_IR_reg[24]/NET0131  & n678 ;
  assign n740 = n725 & n739 ;
  assign n741 = n695 & n740 ;
  assign n742 = \P3_IR_reg[31]/NET0131  & ~n741 ;
  assign n743 = \P3_IR_reg[25]/NET0131  & ~n742 ;
  assign n744 = ~\P3_IR_reg[25]/NET0131  & n742 ;
  assign n745 = ~n743 & ~n744 ;
  assign n746 = n715 & n716 ;
  assign n747 = n682 & n746 ;
  assign n748 = n676 & n747 ;
  assign n749 = \P3_IR_reg[31]/NET0131  & ~n748 ;
  assign n750 = ~\P3_IR_reg[26]/NET0131  & ~n749 ;
  assign n751 = \P3_IR_reg[26]/NET0131  & n749 ;
  assign n752 = ~n750 & ~n751 ;
  assign n756 = ~n745 & n752 ;
  assign n757 = n755 & n756 ;
  assign n758 = n711 & ~n757 ;
  assign n759 = ~n710 & n758 ;
  assign n760 = ~n714 & n759 ;
  assign n761 = ~n738 & n760 ;
  assign n762 = ~n670 & ~n761 ;
  assign n763 = \P1_state_reg[0]/NET0131  & ~n762 ;
  assign n764 = \P3_B_reg/NET0131  & ~n763 ;
  assign n765 = \P1_state_reg[0]/NET0131  & n670 ;
  assign n887 = ~\P3_IR_reg[27]/NET0131  & ~\P3_IR_reg[28]/NET0131  ;
  assign n888 = ~\P3_IR_reg[26]/NET0131  & n887 ;
  assign n889 = ~\P3_IR_reg[25]/NET0131  & n888 ;
  assign n890 = \P3_IR_reg[31]/NET0131  & ~n889 ;
  assign n891 = ~n742 & ~n890 ;
  assign n892 = \P3_IR_reg[29]/NET0131  & ~n891 ;
  assign n893 = ~\P3_IR_reg[29]/NET0131  & n891 ;
  assign n894 = ~n892 & ~n893 ;
  assign n895 = ~\P3_IR_reg[29]/NET0131  & n888 ;
  assign n896 = \P3_IR_reg[31]/NET0131  & ~n895 ;
  assign n897 = ~n749 & ~n896 ;
  assign n898 = \P3_IR_reg[30]/NET0131  & ~n897 ;
  assign n899 = ~\P3_IR_reg[30]/NET0131  & n897 ;
  assign n900 = ~n898 & ~n899 ;
  assign n907 = n894 & n900 ;
  assign n908 = ~\P3_reg3_reg[3]/NET0131  & ~\P3_reg3_reg[4]/NET0131  ;
  assign n909 = ~\P3_reg3_reg[5]/NET0131  & n908 ;
  assign n910 = ~\P3_reg3_reg[6]/NET0131  & n909 ;
  assign n911 = ~\P3_reg3_reg[7]/NET0131  & n910 ;
  assign n912 = ~\P3_reg3_reg[8]/NET0131  & n911 ;
  assign n913 = ~\P3_reg3_reg[9]/NET0131  & n912 ;
  assign n914 = ~\P3_reg3_reg[10]/NET0131  & n913 ;
  assign n915 = ~\P3_reg3_reg[11]/NET0131  & ~\P3_reg3_reg[12]/NET0131  ;
  assign n916 = n914 & n915 ;
  assign n917 = ~\P3_reg3_reg[13]/NET0131  & ~\P3_reg3_reg[14]/NET0131  ;
  assign n918 = ~\P3_reg3_reg[15]/NET0131  & ~\P3_reg3_reg[16]/NET0131  ;
  assign n919 = n917 & n918 ;
  assign n920 = n916 & n919 ;
  assign n921 = ~\P3_reg3_reg[17]/NET0131  & ~\P3_reg3_reg[18]/NET0131  ;
  assign n922 = n920 & n921 ;
  assign n923 = ~\P3_reg3_reg[19]/NET0131  & n922 ;
  assign n924 = ~\P3_reg3_reg[20]/NET0131  & n923 ;
  assign n1228 = ~\P3_reg3_reg[21]/NET0131  & ~\P3_reg3_reg[22]/NET0131  ;
  assign n1229 = ~\P3_reg3_reg[23]/NET0131  & ~\P3_reg3_reg[24]/NET0131  ;
  assign n1230 = n1228 & n1229 ;
  assign n1231 = n924 & n1230 ;
  assign n1322 = ~\P3_reg3_reg[25]/NET0131  & ~\P3_reg3_reg[26]/NET0131  ;
  assign n1323 = ~\P3_reg3_reg[27]/NET0131  & ~\P3_reg3_reg[28]/NET0131  ;
  assign n1324 = n1322 & n1323 ;
  assign n1325 = n1231 & n1324 ;
  assign n1326 = n907 & n1325 ;
  assign n901 = ~n894 & n900 ;
  assign n1333 = \P3_reg2_reg[31]/NET0131  & n901 ;
  assign n903 = n894 & ~n900 ;
  assign n1331 = \P3_reg1_reg[31]/NET0131  & n903 ;
  assign n905 = ~n894 & ~n900 ;
  assign n1332 = \P3_reg0_reg[31]/NET0131  & n905 ;
  assign n1334 = ~n1331 & ~n1332 ;
  assign n1335 = ~n1333 & n1334 ;
  assign n1336 = ~n1326 & n1335 ;
  assign n767 = ~n724 & ~n733 ;
  assign n768 = \P1_addr_reg[19]/NET0131  & \P2_addr_reg[19]/NET0131  ;
  assign n769 = ~\P2_rd_reg/NET0131  & ~\P3_addr_reg[19]/NET0131  ;
  assign n770 = n768 & n769 ;
  assign n771 = ~\P1_addr_reg[19]/NET0131  & ~\P2_addr_reg[19]/NET0131  ;
  assign n772 = ~\P1_rd_reg/NET0131  & \P3_addr_reg[19]/NET0131  ;
  assign n773 = n771 & n772 ;
  assign n774 = ~n770 & ~n773 ;
  assign n1337 = \si[31]_pad  & n774 ;
  assign n813 = ~\P1_datao_reg[14]/NET0131  & \P2_datao_reg[14]/NET0131  ;
  assign n814 = \P1_datao_reg[13]/NET0131  & ~\P2_datao_reg[13]/NET0131  ;
  assign n815 = \P1_datao_reg[14]/NET0131  & ~\P2_datao_reg[14]/NET0131  ;
  assign n816 = ~n814 & ~n815 ;
  assign n817 = ~n813 & ~n816 ;
  assign n818 = ~\P1_datao_reg[12]/NET0131  & \P2_datao_reg[12]/NET0131  ;
  assign n819 = \P1_datao_reg[12]/NET0131  & ~\P2_datao_reg[12]/NET0131  ;
  assign n820 = \P1_datao_reg[11]/NET0131  & ~\P2_datao_reg[11]/NET0131  ;
  assign n821 = ~n819 & ~n820 ;
  assign n822 = ~n818 & ~n821 ;
  assign n823 = ~\P1_datao_reg[13]/NET0131  & \P2_datao_reg[13]/NET0131  ;
  assign n824 = ~n813 & ~n823 ;
  assign n825 = n822 & n824 ;
  assign n826 = ~n817 & ~n825 ;
  assign n827 = ~\P1_datao_reg[10]/NET0131  & \P2_datao_reg[10]/NET0131  ;
  assign n828 = \P1_datao_reg[10]/NET0131  & ~\P2_datao_reg[10]/NET0131  ;
  assign n829 = \P1_datao_reg[9]/NET0131  & ~\P2_datao_reg[9]/NET0131  ;
  assign n830 = ~n828 & ~n829 ;
  assign n831 = ~n827 & ~n830 ;
  assign n832 = ~\P1_datao_reg[7]/NET0131  & \P2_datao_reg[7]/NET0131  ;
  assign n833 = \P1_datao_reg[2]/NET0131  & ~\P2_datao_reg[2]/NET0131  ;
  assign n834 = \P1_datao_reg[1]/NET0131  & ~\P2_datao_reg[1]/NET0131  ;
  assign n835 = ~\P1_datao_reg[1]/NET0131  & \P2_datao_reg[1]/NET0131  ;
  assign n836 = ~\P1_datao_reg[0]/NET0131  & \P2_datao_reg[0]/NET0131  ;
  assign n837 = ~n835 & ~n836 ;
  assign n838 = ~n834 & ~n837 ;
  assign n839 = ~n833 & n838 ;
  assign n840 = ~\P1_datao_reg[3]/NET0131  & \P2_datao_reg[3]/NET0131  ;
  assign n841 = ~\P1_datao_reg[2]/NET0131  & \P2_datao_reg[2]/NET0131  ;
  assign n842 = ~n840 & ~n841 ;
  assign n843 = ~n839 & n842 ;
  assign n844 = \P1_datao_reg[3]/NET0131  & ~\P2_datao_reg[3]/NET0131  ;
  assign n845 = \P1_datao_reg[4]/NET0131  & ~\P2_datao_reg[4]/NET0131  ;
  assign n846 = ~n844 & ~n845 ;
  assign n847 = ~n843 & n846 ;
  assign n848 = ~\P1_datao_reg[6]/NET0131  & \P2_datao_reg[6]/NET0131  ;
  assign n849 = ~\P1_datao_reg[5]/NET0131  & \P2_datao_reg[5]/NET0131  ;
  assign n850 = ~\P1_datao_reg[4]/NET0131  & \P2_datao_reg[4]/NET0131  ;
  assign n851 = ~n849 & ~n850 ;
  assign n852 = ~n848 & n851 ;
  assign n853 = ~n847 & n852 ;
  assign n854 = \P1_datao_reg[6]/NET0131  & ~\P2_datao_reg[6]/NET0131  ;
  assign n855 = \P1_datao_reg[5]/NET0131  & ~\P2_datao_reg[5]/NET0131  ;
  assign n856 = ~n848 & n855 ;
  assign n857 = ~n854 & ~n856 ;
  assign n858 = ~n853 & n857 ;
  assign n859 = ~n832 & ~n858 ;
  assign n860 = \P1_datao_reg[8]/NET0131  & ~\P2_datao_reg[8]/NET0131  ;
  assign n861 = \P1_datao_reg[7]/NET0131  & ~\P2_datao_reg[7]/NET0131  ;
  assign n862 = ~n860 & ~n861 ;
  assign n863 = ~n859 & n862 ;
  assign n864 = ~\P1_datao_reg[8]/NET0131  & \P2_datao_reg[8]/NET0131  ;
  assign n865 = ~\P1_datao_reg[9]/NET0131  & \P2_datao_reg[9]/NET0131  ;
  assign n866 = ~n827 & ~n865 ;
  assign n867 = ~n864 & n866 ;
  assign n868 = ~n863 & n867 ;
  assign n869 = ~n831 & ~n868 ;
  assign n870 = ~\P1_datao_reg[11]/NET0131  & \P2_datao_reg[11]/NET0131  ;
  assign n871 = ~n818 & ~n870 ;
  assign n872 = n824 & n871 ;
  assign n873 = ~n869 & n872 ;
  assign n874 = n826 & ~n873 ;
  assign n779 = ~\P1_datao_reg[22]/NET0131  & \P2_datao_reg[22]/NET0131  ;
  assign n784 = ~\P1_datao_reg[21]/NET0131  & \P2_datao_reg[21]/NET0131  ;
  assign n785 = ~n779 & ~n784 ;
  assign n786 = ~\P1_datao_reg[20]/NET0131  & \P2_datao_reg[20]/NET0131  ;
  assign n793 = ~\P1_datao_reg[19]/NET0131  & \P2_datao_reg[19]/NET0131  ;
  assign n794 = ~n786 & ~n793 ;
  assign n795 = n785 & n794 ;
  assign n797 = ~\P1_datao_reg[17]/NET0131  & \P2_datao_reg[17]/NET0131  ;
  assign n798 = ~\P1_datao_reg[18]/NET0131  & \P2_datao_reg[18]/NET0131  ;
  assign n799 = ~n797 & ~n798 ;
  assign n805 = ~\P1_datao_reg[16]/NET0131  & \P2_datao_reg[16]/NET0131  ;
  assign n875 = ~\P1_datao_reg[15]/NET0131  & \P2_datao_reg[15]/NET0131  ;
  assign n876 = ~n805 & ~n875 ;
  assign n877 = n799 & n876 ;
  assign n878 = n795 & n877 ;
  assign n879 = ~n874 & n878 ;
  assign n1276 = ~\P1_datao_reg[30]/NET0131  & \P2_datao_reg[30]/NET0131  ;
  assign n1283 = ~\P1_datao_reg[29]/NET0131  & \P2_datao_reg[29]/NET0131  ;
  assign n1338 = ~n1276 & ~n1283 ;
  assign n1284 = ~\P1_datao_reg[28]/NET0131  & \P2_datao_reg[28]/NET0131  ;
  assign n1286 = ~\P1_datao_reg[27]/NET0131  & \P2_datao_reg[27]/NET0131  ;
  assign n1343 = ~n1284 & ~n1286 ;
  assign n1344 = n1338 & n1343 ;
  assign n776 = ~\P1_datao_reg[23]/NET0131  & \P2_datao_reg[23]/NET0131  ;
  assign n1208 = ~\P1_datao_reg[24]/NET0131  & \P2_datao_reg[24]/NET0131  ;
  assign n1244 = ~n776 & ~n1208 ;
  assign n1239 = ~\P1_datao_reg[25]/NET0131  & \P2_datao_reg[25]/NET0131  ;
  assign n1287 = ~\P1_datao_reg[26]/NET0131  & \P2_datao_reg[26]/NET0131  ;
  assign n1347 = ~n1239 & ~n1287 ;
  assign n1350 = n1244 & n1347 ;
  assign n1354 = n1344 & n1350 ;
  assign n1355 = n879 & n1354 ;
  assign n1240 = \P1_datao_reg[25]/NET0131  & ~\P2_datao_reg[25]/NET0131  ;
  assign n1304 = \P1_datao_reg[26]/NET0131  & ~\P2_datao_reg[26]/NET0131  ;
  assign n1345 = ~n1240 & ~n1304 ;
  assign n1346 = ~n1287 & ~n1345 ;
  assign n777 = \P1_datao_reg[23]/NET0131  & ~\P2_datao_reg[23]/NET0131  ;
  assign n1209 = \P1_datao_reg[24]/NET0131  & ~\P2_datao_reg[24]/NET0131  ;
  assign n1242 = ~n777 & ~n1209 ;
  assign n1243 = ~n1208 & ~n1242 ;
  assign n1348 = n1243 & n1347 ;
  assign n1349 = ~n1346 & ~n1348 ;
  assign n780 = \P1_datao_reg[22]/NET0131  & ~\P2_datao_reg[22]/NET0131  ;
  assign n781 = \P1_datao_reg[21]/NET0131  & ~\P2_datao_reg[21]/NET0131  ;
  assign n782 = ~n780 & ~n781 ;
  assign n783 = ~n779 & ~n782 ;
  assign n787 = \P1_datao_reg[20]/NET0131  & ~\P2_datao_reg[20]/NET0131  ;
  assign n788 = \P1_datao_reg[19]/NET0131  & ~\P2_datao_reg[19]/NET0131  ;
  assign n789 = ~n787 & ~n788 ;
  assign n790 = ~n786 & ~n789 ;
  assign n791 = n785 & n790 ;
  assign n792 = ~n783 & ~n791 ;
  assign n796 = \P1_datao_reg[18]/NET0131  & ~\P2_datao_reg[18]/NET0131  ;
  assign n800 = ~n796 & ~n799 ;
  assign n801 = \P1_datao_reg[17]/NET0131  & ~\P2_datao_reg[17]/NET0131  ;
  assign n802 = ~n796 & ~n801 ;
  assign n803 = ~n798 & ~n802 ;
  assign n804 = \P1_datao_reg[16]/NET0131  & ~\P2_datao_reg[16]/NET0131  ;
  assign n806 = \P1_datao_reg[15]/NET0131  & ~\P2_datao_reg[15]/NET0131  ;
  assign n807 = ~n805 & n806 ;
  assign n808 = ~n804 & ~n807 ;
  assign n809 = ~n803 & n808 ;
  assign n810 = ~n800 & ~n809 ;
  assign n811 = n795 & n810 ;
  assign n812 = n792 & ~n811 ;
  assign n1351 = ~n812 & n1350 ;
  assign n1352 = n1349 & ~n1351 ;
  assign n1353 = n1344 & ~n1352 ;
  assign n1277 = \P1_datao_reg[30]/NET0131  & ~\P2_datao_reg[30]/NET0131  ;
  assign n1279 = \P1_datao_reg[29]/NET0131  & ~\P2_datao_reg[29]/NET0131  ;
  assign n1303 = \P1_datao_reg[28]/NET0131  & ~\P2_datao_reg[28]/NET0131  ;
  assign n1305 = \P1_datao_reg[27]/NET0131  & ~\P2_datao_reg[27]/NET0131  ;
  assign n1339 = ~n1303 & ~n1305 ;
  assign n1340 = ~n1284 & ~n1339 ;
  assign n1341 = ~n1279 & ~n1340 ;
  assign n1342 = n1338 & ~n1341 ;
  assign n1356 = ~n1277 & ~n1342 ;
  assign n1357 = ~n1353 & n1356 ;
  assign n1358 = ~n1355 & n1357 ;
  assign n1359 = \P1_datao_reg[31]/NET0131  & ~n1358 ;
  assign n1360 = ~\P1_datao_reg[31]/NET0131  & n1358 ;
  assign n1361 = ~n1359 & ~n1360 ;
  assign n1363 = ~\P2_datao_reg[31]/NET0131  & n1361 ;
  assign n1362 = \P2_datao_reg[31]/NET0131  & ~n1361 ;
  assign n1364 = ~n774 & ~n1362 ;
  assign n1365 = ~n1363 & n1364 ;
  assign n1366 = ~n1337 & ~n1365 ;
  assign n1367 = ~n767 & ~n1366 ;
  assign n1479 = ~n1336 & ~n1367 ;
  assign n1275 = \si[30]_pad  & n774 ;
  assign n1278 = ~n1276 & ~n1277 ;
  assign n946 = ~n814 & ~n819 ;
  assign n947 = ~n823 & ~n946 ;
  assign n948 = ~n820 & ~n828 ;
  assign n949 = ~n870 & ~n948 ;
  assign n950 = ~n818 & ~n823 ;
  assign n951 = n949 & n950 ;
  assign n952 = ~n947 & ~n951 ;
  assign n953 = ~n829 & ~n860 ;
  assign n954 = ~n865 & ~n953 ;
  assign n955 = ~n838 & ~n841 ;
  assign n956 = ~n833 & ~n844 ;
  assign n957 = ~n955 & n956 ;
  assign n958 = ~n840 & ~n957 ;
  assign n959 = n851 & n958 ;
  assign n960 = n845 & ~n849 ;
  assign n961 = ~n855 & ~n960 ;
  assign n962 = ~n959 & n961 ;
  assign n963 = ~n848 & ~n962 ;
  assign n964 = ~n854 & ~n861 ;
  assign n965 = ~n963 & n964 ;
  assign n966 = ~n832 & ~n864 ;
  assign n967 = ~n865 & n966 ;
  assign n968 = ~n965 & n967 ;
  assign n969 = ~n954 & ~n968 ;
  assign n970 = ~n827 & ~n870 ;
  assign n971 = n950 & n970 ;
  assign n972 = ~n969 & n971 ;
  assign n973 = n952 & ~n972 ;
  assign n974 = ~n797 & ~n805 ;
  assign n975 = ~n813 & ~n875 ;
  assign n976 = n974 & n975 ;
  assign n977 = ~n973 & n976 ;
  assign n939 = ~n784 & ~n786 ;
  assign n944 = ~n793 & ~n798 ;
  assign n945 = n939 & n944 ;
  assign n1211 = ~n776 & ~n779 ;
  assign n1280 = ~n1208 & ~n1239 ;
  assign n1281 = n1211 & n1280 ;
  assign n1282 = n945 & n1281 ;
  assign n1285 = ~n1283 & ~n1284 ;
  assign n1288 = ~n1286 & ~n1287 ;
  assign n1289 = n1285 & n1288 ;
  assign n1290 = n1282 & n1289 ;
  assign n1291 = n977 & n1290 ;
  assign n1292 = ~n1209 & ~n1240 ;
  assign n1293 = ~n1239 & ~n1292 ;
  assign n1294 = ~n777 & ~n780 ;
  assign n1295 = ~n776 & n1280 ;
  assign n1296 = ~n1294 & n1295 ;
  assign n1297 = ~n1293 & ~n1296 ;
  assign n937 = ~n781 & ~n787 ;
  assign n938 = ~n784 & ~n937 ;
  assign n940 = ~n788 & ~n796 ;
  assign n941 = ~n793 & ~n940 ;
  assign n942 = n939 & n941 ;
  assign n943 = ~n938 & ~n942 ;
  assign n978 = ~n806 & ~n815 ;
  assign n979 = ~n875 & ~n978 ;
  assign n980 = ~n804 & ~n979 ;
  assign n981 = n974 & ~n980 ;
  assign n982 = ~n801 & ~n981 ;
  assign n1298 = n945 & ~n982 ;
  assign n1299 = n943 & ~n1298 ;
  assign n1300 = n1281 & ~n1299 ;
  assign n1301 = n1297 & ~n1300 ;
  assign n1302 = n1289 & ~n1301 ;
  assign n1306 = ~n1304 & ~n1305 ;
  assign n1307 = ~n1286 & ~n1306 ;
  assign n1308 = ~n1303 & ~n1307 ;
  assign n1309 = n1285 & ~n1308 ;
  assign n1310 = ~n1279 & ~n1309 ;
  assign n1311 = ~n1302 & n1310 ;
  assign n1312 = ~n1291 & n1311 ;
  assign n1314 = n1278 & ~n1312 ;
  assign n1313 = ~n1278 & n1312 ;
  assign n1315 = ~n774 & ~n1313 ;
  assign n1316 = ~n1314 & n1315 ;
  assign n1317 = ~n1275 & ~n1316 ;
  assign n1318 = ~n767 & ~n1317 ;
  assign n1321 = \P3_reg2_reg[30]/NET0131  & n901 ;
  assign n1319 = \P3_reg1_reg[30]/NET0131  & n903 ;
  assign n1320 = \P3_reg0_reg[30]/NET0131  & n905 ;
  assign n1327 = ~n1319 & ~n1320 ;
  assign n1328 = ~n1321 & n1327 ;
  assign n1329 = ~n1326 & n1328 ;
  assign n1330 = ~n1318 & ~n1329 ;
  assign n1368 = n1336 & n1367 ;
  assign n1369 = ~n1330 & ~n1368 ;
  assign n1480 = n1318 & n1329 ;
  assign n1370 = \si[29]_pad  & n774 ;
  assign n1371 = ~n1279 & ~n1283 ;
  assign n1004 = n794 & n803 ;
  assign n1005 = ~n790 & ~n1004 ;
  assign n1006 = ~n806 & ~n817 ;
  assign n1007 = n876 & ~n1006 ;
  assign n1008 = ~n804 & ~n1007 ;
  assign n1009 = n831 & n871 ;
  assign n1010 = ~n822 & ~n1009 ;
  assign n1011 = n858 & ~n861 ;
  assign n1012 = n966 & ~n1011 ;
  assign n1013 = ~n860 & ~n1012 ;
  assign n1014 = n866 & n871 ;
  assign n1015 = ~n1013 & n1014 ;
  assign n1016 = n1010 & ~n1015 ;
  assign n1017 = n824 & n876 ;
  assign n1018 = ~n1016 & n1017 ;
  assign n1019 = n1008 & ~n1018 ;
  assign n1020 = n794 & n799 ;
  assign n1021 = ~n1019 & n1020 ;
  assign n1022 = n1005 & ~n1021 ;
  assign n1247 = n785 & n1244 ;
  assign n1375 = n1343 & n1347 ;
  assign n1376 = n1247 & n1375 ;
  assign n1377 = ~n1022 & n1376 ;
  assign n1245 = n783 & n1244 ;
  assign n1246 = ~n1243 & ~n1245 ;
  assign n1372 = ~n1246 & n1347 ;
  assign n1373 = ~n1346 & ~n1372 ;
  assign n1374 = n1343 & ~n1373 ;
  assign n1378 = ~n1340 & ~n1374 ;
  assign n1379 = ~n1377 & n1378 ;
  assign n1381 = n1371 & ~n1379 ;
  assign n1380 = ~n1371 & n1379 ;
  assign n1382 = ~n774 & ~n1380 ;
  assign n1383 = ~n1381 & n1382 ;
  assign n1384 = ~n1370 & ~n1383 ;
  assign n1385 = ~n767 & ~n1384 ;
  assign n1388 = \P3_reg2_reg[29]/NET0131  & n901 ;
  assign n1386 = \P3_reg1_reg[29]/NET0131  & n903 ;
  assign n1387 = \P3_reg0_reg[29]/NET0131  & n905 ;
  assign n1389 = ~n1386 & ~n1387 ;
  assign n1390 = ~n1388 & n1389 ;
  assign n1391 = ~n1326 & n1390 ;
  assign n1392 = ~n1385 & ~n1391 ;
  assign n1394 = \si[28]_pad  & n774 ;
  assign n1395 = ~n1284 & ~n1303 ;
  assign n1041 = n968 & n970 ;
  assign n1042 = n954 & n970 ;
  assign n1043 = ~n949 & ~n1042 ;
  assign n1044 = ~n1041 & n1043 ;
  assign n1045 = n950 & n975 ;
  assign n1046 = ~n1044 & n1045 ;
  assign n1047 = n947 & n975 ;
  assign n1048 = ~n979 & ~n1047 ;
  assign n1049 = ~n1046 & n1048 ;
  assign n1050 = n944 & n974 ;
  assign n1051 = ~n1049 & n1050 ;
  assign n1052 = ~n801 & ~n804 ;
  assign n1053 = ~n797 & n944 ;
  assign n1054 = ~n1052 & n1053 ;
  assign n1055 = ~n941 & ~n1054 ;
  assign n1056 = ~n1051 & n1055 ;
  assign n1212 = n939 & n1211 ;
  assign n1213 = ~n1056 & n1212 ;
  assign n1396 = n1280 & n1288 ;
  assign n1397 = n1213 & n1396 ;
  assign n1214 = ~n780 & ~n938 ;
  assign n1215 = n1211 & ~n1214 ;
  assign n1216 = ~n777 & ~n1215 ;
  assign n1398 = ~n1216 & n1280 ;
  assign n1399 = ~n1293 & ~n1398 ;
  assign n1400 = n1288 & ~n1399 ;
  assign n1401 = ~n1307 & ~n1400 ;
  assign n1402 = ~n1397 & n1401 ;
  assign n1404 = n1395 & ~n1402 ;
  assign n1403 = ~n1395 & n1402 ;
  assign n1405 = ~n774 & ~n1403 ;
  assign n1406 = ~n1404 & n1405 ;
  assign n1407 = ~n1394 & ~n1406 ;
  assign n1408 = ~n767 & ~n1407 ;
  assign n1266 = ~\P3_reg3_reg[25]/NET0131  & n1231 ;
  assign n1412 = ~\P3_reg3_reg[26]/NET0131  & n1266 ;
  assign n1413 = ~\P3_reg3_reg[27]/NET0131  & n1412 ;
  assign n1414 = \P3_reg3_reg[28]/NET0131  & ~n1413 ;
  assign n1415 = ~n1325 & ~n1414 ;
  assign n1416 = n907 & ~n1415 ;
  assign n1411 = \P3_reg0_reg[28]/NET0131  & n905 ;
  assign n1409 = \P3_reg1_reg[28]/NET0131  & n903 ;
  assign n1410 = \P3_reg2_reg[28]/NET0131  & n901 ;
  assign n1417 = ~n1409 & ~n1410 ;
  assign n1418 = ~n1411 & n1417 ;
  assign n1419 = ~n1416 & n1418 ;
  assign n1420 = ~n1408 & ~n1419 ;
  assign n1493 = n1385 & n1391 ;
  assign n1993 = n1420 & ~n1493 ;
  assign n1994 = ~n1392 & ~n1993 ;
  assign n2006 = ~n1480 & ~n1994 ;
  assign n2007 = n1369 & ~n2006 ;
  assign n2008 = ~n1479 & ~n2007 ;
  assign n1207 = \si[24]_pad  & n774 ;
  assign n1210 = ~n1208 & ~n1209 ;
  assign n1217 = ~n1213 & n1216 ;
  assign n1219 = n1210 & ~n1217 ;
  assign n1218 = ~n1210 & n1217 ;
  assign n1220 = ~n774 & ~n1218 ;
  assign n1221 = ~n1219 & n1220 ;
  assign n1222 = ~n1207 & ~n1221 ;
  assign n1223 = ~n767 & ~n1222 ;
  assign n925 = ~\P3_reg3_reg[21]/NET0131  & n924 ;
  assign n926 = ~\P3_reg3_reg[22]/NET0131  & n925 ;
  assign n927 = ~\P3_reg3_reg[23]/NET0131  & n926 ;
  assign n1227 = \P3_reg3_reg[24]/NET0131  & ~n927 ;
  assign n1232 = ~n1227 & ~n1231 ;
  assign n1233 = n907 & ~n1232 ;
  assign n1226 = \P3_reg0_reg[24]/NET0131  & n905 ;
  assign n1224 = \P3_reg1_reg[24]/NET0131  & n903 ;
  assign n1225 = \P3_reg2_reg[24]/NET0131  & n901 ;
  assign n1234 = ~n1224 & ~n1225 ;
  assign n1235 = ~n1226 & n1234 ;
  assign n1236 = ~n1233 & n1235 ;
  assign n1237 = ~n1223 & ~n1236 ;
  assign n1238 = ~\si[25]_pad  & n774 ;
  assign n1241 = ~n1239 & ~n1240 ;
  assign n1251 = n1017 & n1020 ;
  assign n1252 = n1015 & n1251 ;
  assign n1248 = ~n1010 & n1017 ;
  assign n1249 = n1008 & ~n1248 ;
  assign n1250 = n1020 & ~n1249 ;
  assign n1253 = n1005 & ~n1250 ;
  assign n1254 = ~n1252 & n1253 ;
  assign n1255 = n1247 & ~n1254 ;
  assign n1256 = n1246 & ~n1255 ;
  assign n1258 = n1241 & n1256 ;
  assign n1257 = ~n1241 & ~n1256 ;
  assign n1259 = ~n774 & ~n1257 ;
  assign n1260 = ~n1258 & n1259 ;
  assign n1261 = ~n1238 & ~n1260 ;
  assign n1262 = ~n767 & n1261 ;
  assign n1267 = \P3_reg3_reg[25]/NET0131  & ~n1231 ;
  assign n1268 = ~n1266 & ~n1267 ;
  assign n1269 = n907 & ~n1268 ;
  assign n1265 = \P3_reg1_reg[25]/NET0131  & n903 ;
  assign n1263 = \P3_reg0_reg[25]/NET0131  & n905 ;
  assign n1264 = \P3_reg2_reg[25]/NET0131  & n901 ;
  assign n1270 = ~n1263 & ~n1264 ;
  assign n1271 = ~n1265 & n1270 ;
  assign n1272 = ~n1269 & n1271 ;
  assign n1273 = ~n1262 & ~n1272 ;
  assign n1274 = ~n1237 & ~n1273 ;
  assign n1449 = ~\si[26]_pad  & n774 ;
  assign n1450 = ~n1287 & ~n1304 ;
  assign n1456 = n976 & n1282 ;
  assign n1457 = n972 & n1456 ;
  assign n1451 = ~n952 & n976 ;
  assign n1452 = n982 & ~n1451 ;
  assign n1453 = n945 & ~n1452 ;
  assign n1454 = n943 & ~n1453 ;
  assign n1455 = n1281 & ~n1454 ;
  assign n1458 = n1297 & ~n1455 ;
  assign n1459 = ~n1457 & n1458 ;
  assign n1461 = n1450 & n1459 ;
  assign n1460 = ~n1450 & ~n1459 ;
  assign n1462 = ~n774 & ~n1460 ;
  assign n1463 = ~n1461 & n1462 ;
  assign n1464 = ~n1449 & ~n1463 ;
  assign n1465 = ~n767 & n1464 ;
  assign n1469 = \P3_reg3_reg[26]/NET0131  & ~n1266 ;
  assign n1470 = ~n1412 & ~n1469 ;
  assign n1471 = n907 & ~n1470 ;
  assign n1468 = \P3_reg0_reg[26]/NET0131  & n905 ;
  assign n1466 = \P3_reg1_reg[26]/NET0131  & n903 ;
  assign n1467 = \P3_reg2_reg[26]/NET0131  & n901 ;
  assign n1472 = ~n1466 & ~n1467 ;
  assign n1473 = ~n1468 & n1472 ;
  assign n1474 = ~n1471 & n1473 ;
  assign n1483 = n1465 & n1474 ;
  assign n1421 = ~\si[27]_pad  & n774 ;
  assign n1422 = ~n1286 & ~n1305 ;
  assign n1423 = n873 & n878 ;
  assign n1424 = ~n826 & n877 ;
  assign n1425 = ~n810 & ~n1424 ;
  assign n1426 = n795 & ~n1425 ;
  assign n1427 = n792 & ~n1426 ;
  assign n1428 = ~n1423 & n1427 ;
  assign n1429 = n1350 & ~n1428 ;
  assign n1430 = n1349 & ~n1429 ;
  assign n1432 = n1422 & n1430 ;
  assign n1431 = ~n1422 & ~n1430 ;
  assign n1433 = ~n774 & ~n1431 ;
  assign n1434 = ~n1432 & n1433 ;
  assign n1435 = ~n1421 & ~n1434 ;
  assign n1436 = ~n767 & n1435 ;
  assign n1440 = \P3_reg3_reg[27]/NET0131  & ~n1412 ;
  assign n1441 = ~n1413 & ~n1440 ;
  assign n1442 = n907 & ~n1441 ;
  assign n1439 = \P3_reg0_reg[27]/NET0131  & n905 ;
  assign n1437 = \P3_reg1_reg[27]/NET0131  & n903 ;
  assign n1438 = \P3_reg2_reg[27]/NET0131  & n901 ;
  assign n1443 = ~n1437 & ~n1438 ;
  assign n1444 = ~n1439 & n1443 ;
  assign n1445 = ~n1442 & n1444 ;
  assign n1484 = n1436 & n1445 ;
  assign n1485 = ~n1483 & ~n1484 ;
  assign n1487 = n1262 & n1272 ;
  assign n1949 = n1485 & ~n1487 ;
  assign n1950 = ~n1274 & n1949 ;
  assign n1446 = ~n1436 & ~n1445 ;
  assign n1475 = ~n1465 & ~n1474 ;
  assign n1948 = n1475 & ~n1484 ;
  assign n1951 = ~n1446 & ~n1948 ;
  assign n1952 = ~n1950 & n1951 ;
  assign n1488 = n1223 & n1236 ;
  assign n1954 = ~n1488 & n1949 ;
  assign n775 = \si[23]_pad  & n774 ;
  assign n778 = ~n776 & ~n777 ;
  assign n880 = n812 & ~n879 ;
  assign n882 = n778 & ~n880 ;
  assign n881 = ~n778 & n880 ;
  assign n883 = ~n774 & ~n881 ;
  assign n884 = ~n882 & n883 ;
  assign n885 = ~n775 & ~n884 ;
  assign n886 = ~n767 & ~n885 ;
  assign n928 = \P3_reg3_reg[23]/NET0131  & ~n926 ;
  assign n929 = ~n927 & ~n928 ;
  assign n930 = n907 & ~n929 ;
  assign n906 = \P3_reg0_reg[23]/NET0131  & n905 ;
  assign n902 = \P3_reg2_reg[23]/NET0131  & n901 ;
  assign n904 = \P3_reg1_reg[23]/NET0131  & n903 ;
  assign n931 = ~n902 & ~n904 ;
  assign n932 = ~n906 & n931 ;
  assign n933 = ~n930 & n932 ;
  assign n934 = n886 & n933 ;
  assign n935 = \si[22]_pad  & n774 ;
  assign n936 = ~n779 & ~n780 ;
  assign n983 = ~n977 & n982 ;
  assign n984 = n945 & ~n983 ;
  assign n985 = n943 & ~n984 ;
  assign n987 = n936 & ~n985 ;
  assign n986 = ~n936 & n985 ;
  assign n988 = ~n774 & ~n986 ;
  assign n989 = ~n987 & n988 ;
  assign n990 = ~n935 & ~n989 ;
  assign n991 = ~n767 & ~n990 ;
  assign n995 = \P3_reg3_reg[22]/NET0131  & ~n925 ;
  assign n996 = ~n926 & ~n995 ;
  assign n997 = n907 & ~n996 ;
  assign n994 = \P3_reg1_reg[22]/NET0131  & n903 ;
  assign n992 = \P3_reg2_reg[22]/NET0131  & n901 ;
  assign n993 = \P3_reg0_reg[22]/NET0131  & n905 ;
  assign n998 = ~n992 & ~n993 ;
  assign n999 = ~n994 & n998 ;
  assign n1000 = ~n997 & n999 ;
  assign n1001 = n991 & n1000 ;
  assign n1002 = ~n934 & ~n1001 ;
  assign n1003 = \si[21]_pad  & n774 ;
  assign n1023 = ~n781 & ~n784 ;
  assign n1025 = ~n1022 & n1023 ;
  assign n1024 = n1022 & ~n1023 ;
  assign n1026 = ~n774 & ~n1024 ;
  assign n1027 = ~n1025 & n1026 ;
  assign n1028 = ~n1003 & ~n1027 ;
  assign n1029 = ~n767 & ~n1028 ;
  assign n1033 = \P3_reg3_reg[21]/NET0131  & ~n924 ;
  assign n1034 = ~n925 & ~n1033 ;
  assign n1035 = n907 & ~n1034 ;
  assign n1032 = \P3_reg1_reg[21]/NET0131  & n903 ;
  assign n1030 = \P3_reg2_reg[21]/NET0131  & n901 ;
  assign n1031 = \P3_reg0_reg[21]/NET0131  & n905 ;
  assign n1036 = ~n1030 & ~n1031 ;
  assign n1037 = ~n1032 & n1036 ;
  assign n1038 = ~n1035 & n1037 ;
  assign n1039 = ~n1029 & ~n1038 ;
  assign n1040 = \si[20]_pad  & n774 ;
  assign n1057 = ~n786 & ~n787 ;
  assign n1059 = ~n1056 & n1057 ;
  assign n1058 = n1056 & ~n1057 ;
  assign n1060 = ~n774 & ~n1058 ;
  assign n1061 = ~n1059 & n1060 ;
  assign n1062 = ~n1040 & ~n1061 ;
  assign n1063 = ~n767 & ~n1062 ;
  assign n1067 = \P3_reg3_reg[20]/NET0131  & ~n923 ;
  assign n1068 = ~n924 & ~n1067 ;
  assign n1069 = n907 & ~n1068 ;
  assign n1066 = \P3_reg2_reg[20]/NET0131  & n901 ;
  assign n1064 = \P3_reg0_reg[20]/NET0131  & n905 ;
  assign n1065 = \P3_reg1_reg[20]/NET0131  & n903 ;
  assign n1070 = ~n1064 & ~n1065 ;
  assign n1071 = ~n1066 & n1070 ;
  assign n1072 = ~n1069 & n1071 ;
  assign n1073 = ~n1063 & ~n1072 ;
  assign n1074 = ~n1039 & ~n1073 ;
  assign n1075 = n1029 & n1038 ;
  assign n1076 = ~n1074 & ~n1075 ;
  assign n1077 = n1002 & n1076 ;
  assign n1078 = ~n991 & ~n1000 ;
  assign n1079 = ~n886 & ~n933 ;
  assign n1080 = ~n1078 & ~n1079 ;
  assign n1081 = ~n934 & ~n1080 ;
  assign n1082 = ~n1077 & ~n1081 ;
  assign n1083 = n1063 & n1072 ;
  assign n1084 = ~n1075 & ~n1083 ;
  assign n1085 = n1002 & n1084 ;
  assign n1087 = \P3_reg2_reg[19]/NET0131  & n901 ;
  assign n1088 = \P3_reg0_reg[19]/NET0131  & n905 ;
  assign n1093 = ~n1087 & ~n1088 ;
  assign n1089 = \P3_reg3_reg[19]/NET0131  & ~n922 ;
  assign n1090 = ~n923 & ~n1089 ;
  assign n1091 = n907 & ~n1090 ;
  assign n1092 = \P3_reg1_reg[19]/NET0131  & n903 ;
  assign n1094 = ~n1091 & ~n1092 ;
  assign n1095 = n1093 & n1094 ;
  assign n1096 = \si[19]_pad  & n774 ;
  assign n1097 = ~n788 & ~n793 ;
  assign n1098 = ~n874 & n877 ;
  assign n1099 = ~n810 & ~n1098 ;
  assign n1101 = n1097 & ~n1099 ;
  assign n1100 = ~n1097 & n1099 ;
  assign n1102 = ~n774 & ~n1100 ;
  assign n1103 = ~n1101 & n1102 ;
  assign n1104 = ~n1096 & ~n1103 ;
  assign n1105 = ~n767 & ~n1104 ;
  assign n1106 = ~\P3_IR_reg[19]/NET0131  & ~n662 ;
  assign n1107 = \P3_IR_reg[19]/NET0131  & n662 ;
  assign n1108 = ~n1106 & ~n1107 ;
  assign n1109 = n767 & n1108 ;
  assign n1110 = ~n1105 & ~n1109 ;
  assign n1111 = n1095 & ~n1110 ;
  assign n1112 = \P3_reg2_reg[18]/NET0131  & n901 ;
  assign n1113 = \P3_reg0_reg[18]/NET0131  & n905 ;
  assign n1119 = ~n1112 & ~n1113 ;
  assign n1114 = ~\P3_reg3_reg[17]/NET0131  & n920 ;
  assign n1115 = \P3_reg3_reg[18]/NET0131  & ~n1114 ;
  assign n1116 = ~n922 & ~n1115 ;
  assign n1117 = n907 & ~n1116 ;
  assign n1118 = \P3_reg1_reg[18]/NET0131  & n903 ;
  assign n1120 = ~n1117 & ~n1118 ;
  assign n1121 = n1119 & n1120 ;
  assign n1122 = \si[18]_pad  & n774 ;
  assign n1123 = ~n796 & ~n798 ;
  assign n1125 = ~n983 & n1123 ;
  assign n1124 = n983 & ~n1123 ;
  assign n1126 = ~n774 & ~n1124 ;
  assign n1127 = ~n1125 & n1126 ;
  assign n1128 = ~n1122 & ~n1127 ;
  assign n1129 = ~n767 & ~n1128 ;
  assign n1130 = ~\P3_IR_reg[17]/NET0131  & n680 ;
  assign n1131 = \P3_IR_reg[31]/NET0131  & ~n1130 ;
  assign n1132 = ~n677 & ~n1131 ;
  assign n1133 = \P3_IR_reg[18]/NET0131  & ~n1132 ;
  assign n1134 = ~\P3_IR_reg[18]/NET0131  & n1132 ;
  assign n1135 = ~n1133 & ~n1134 ;
  assign n1136 = n767 & n1135 ;
  assign n1137 = ~n1129 & ~n1136 ;
  assign n1138 = n1121 & ~n1137 ;
  assign n1139 = ~n1111 & ~n1138 ;
  assign n1140 = \P3_reg1_reg[17]/NET0131  & n903 ;
  assign n1141 = ~\P3_reg3_reg[1]/NET0131  & ~\P3_reg3_reg[2]/NET0131  ;
  assign n1142 = \P3_reg3_reg[3]/NET0131  & ~n1141 ;
  assign n1143 = n920 & ~n1142 ;
  assign n1144 = \P3_reg3_reg[17]/NET0131  & ~n1143 ;
  assign n1145 = n1114 & ~n1142 ;
  assign n1146 = ~n1144 & ~n1145 ;
  assign n1147 = n907 & ~n1146 ;
  assign n1150 = ~n1140 & ~n1147 ;
  assign n1148 = \P3_reg0_reg[17]/NET0131  & n905 ;
  assign n1149 = \P3_reg2_reg[17]/NET0131  & n901 ;
  assign n1151 = ~n1148 & ~n1149 ;
  assign n1152 = n1150 & n1151 ;
  assign n1153 = \si[17]_pad  & n774 ;
  assign n1154 = ~n797 & ~n801 ;
  assign n1156 = ~n1019 & n1154 ;
  assign n1155 = n1019 & ~n1154 ;
  assign n1157 = ~n774 & ~n1155 ;
  assign n1158 = ~n1156 & n1157 ;
  assign n1159 = ~n1153 & ~n1158 ;
  assign n1160 = ~n767 & ~n1159 ;
  assign n1161 = \P3_IR_reg[31]/NET0131  & ~n695 ;
  assign n1162 = \P3_IR_reg[17]/NET0131  & ~n1161 ;
  assign n1163 = ~\P3_IR_reg[17]/NET0131  & n1161 ;
  assign n1164 = ~n1162 & ~n1163 ;
  assign n1165 = n767 & ~n1164 ;
  assign n1166 = ~n1160 & ~n1165 ;
  assign n1170 = n1152 & ~n1166 ;
  assign n1167 = ~n1152 & n1166 ;
  assign n1171 = \si[16]_pad  & n774 ;
  assign n1172 = ~n804 & ~n805 ;
  assign n1174 = ~n1049 & n1172 ;
  assign n1173 = n1049 & ~n1172 ;
  assign n1175 = ~n774 & ~n1173 ;
  assign n1176 = ~n1174 & n1175 ;
  assign n1177 = ~n1171 & ~n1176 ;
  assign n1178 = ~n767 & ~n1177 ;
  assign n1179 = \P3_IR_reg[31]/NET0131  & ~n679 ;
  assign n1180 = ~n677 & ~n1179 ;
  assign n1181 = \P3_IR_reg[16]/NET0131  & ~n1180 ;
  assign n1182 = ~\P3_IR_reg[16]/NET0131  & n1180 ;
  assign n1183 = ~n1181 & ~n1182 ;
  assign n1184 = n767 & n1183 ;
  assign n1185 = ~n1178 & ~n1184 ;
  assign n1189 = ~\P3_reg3_reg[13]/NET0131  & n916 ;
  assign n1190 = ~\P3_reg3_reg[14]/NET0131  & n1189 ;
  assign n1191 = ~\P3_reg3_reg[15]/NET0131  & n1190 ;
  assign n1192 = \P3_reg3_reg[16]/NET0131  & ~n1191 ;
  assign n1193 = ~n920 & ~n1192 ;
  assign n1194 = n907 & ~n1193 ;
  assign n1188 = \P3_reg1_reg[16]/NET0131  & n903 ;
  assign n1186 = \P3_reg2_reg[16]/NET0131  & n901 ;
  assign n1187 = \P3_reg0_reg[16]/NET0131  & n905 ;
  assign n1195 = ~n1186 & ~n1187 ;
  assign n1196 = ~n1188 & n1195 ;
  assign n1197 = ~n1194 & n1196 ;
  assign n1497 = n1185 & ~n1197 ;
  assign n1955 = ~n1167 & ~n1497 ;
  assign n1956 = ~n1170 & ~n1955 ;
  assign n1957 = n1139 & n1956 ;
  assign n1202 = ~n1095 & n1110 ;
  assign n1168 = ~n1121 & n1137 ;
  assign n1958 = ~n1111 & n1168 ;
  assign n1959 = ~n1202 & ~n1958 ;
  assign n1960 = ~n1957 & n1959 ;
  assign n1961 = n1085 & ~n1960 ;
  assign n1962 = n1082 & ~n1961 ;
  assign n1198 = ~n1185 & n1197 ;
  assign n1199 = ~n1170 & ~n1198 ;
  assign n1963 = n1139 & n1199 ;
  assign n1964 = n1085 & n1963 ;
  assign n1498 = \P3_IR_reg[15]/NET0131  & ~\P3_IR_reg[31]/NET0131  ;
  assign n1499 = \P3_IR_reg[15]/NET0131  & ~n657 ;
  assign n1500 = \P3_IR_reg[31]/NET0131  & ~n658 ;
  assign n1501 = ~n1499 & n1500 ;
  assign n1502 = ~n1498 & ~n1501 ;
  assign n1503 = n767 & ~n1502 ;
  assign n1504 = \si[15]_pad  & n774 ;
  assign n1505 = ~n806 & ~n875 ;
  assign n1507 = ~n874 & n1505 ;
  assign n1506 = n874 & ~n1505 ;
  assign n1508 = ~n774 & ~n1506 ;
  assign n1509 = ~n1507 & n1508 ;
  assign n1510 = ~n1504 & ~n1509 ;
  assign n1511 = ~n767 & ~n1510 ;
  assign n1512 = ~n1503 & ~n1511 ;
  assign n1513 = \P3_reg3_reg[15]/NET0131  & ~n1190 ;
  assign n1514 = ~n1191 & ~n1513 ;
  assign n1515 = n907 & ~n1514 ;
  assign n1516 = \P3_reg0_reg[15]/NET0131  & n905 ;
  assign n1519 = ~n1515 & ~n1516 ;
  assign n1517 = \P3_reg2_reg[15]/NET0131  & n901 ;
  assign n1518 = \P3_reg1_reg[15]/NET0131  & n903 ;
  assign n1520 = ~n1517 & ~n1518 ;
  assign n1521 = n1519 & n1520 ;
  assign n1522 = ~n1512 & n1521 ;
  assign n1523 = \P3_reg2_reg[14]/NET0131  & n901 ;
  assign n1524 = \P3_reg3_reg[14]/NET0131  & ~n1189 ;
  assign n1525 = ~n1190 & ~n1524 ;
  assign n1526 = n907 & ~n1525 ;
  assign n1529 = ~n1523 & ~n1526 ;
  assign n1527 = \P3_reg1_reg[14]/NET0131  & n903 ;
  assign n1528 = \P3_reg0_reg[14]/NET0131  & n905 ;
  assign n1530 = ~n1527 & ~n1528 ;
  assign n1531 = n1529 & n1530 ;
  assign n1532 = \si[14]_pad  & n774 ;
  assign n1533 = ~n813 & ~n815 ;
  assign n1535 = ~n973 & n1533 ;
  assign n1534 = n973 & ~n1533 ;
  assign n1536 = ~n774 & ~n1534 ;
  assign n1537 = ~n1535 & n1536 ;
  assign n1538 = ~n1532 & ~n1537 ;
  assign n1539 = ~n767 & ~n1538 ;
  assign n1540 = ~\P3_IR_reg[14]/NET0131  & ~n677 ;
  assign n1541 = \P3_IR_reg[14]/NET0131  & n677 ;
  assign n1542 = ~n1540 & ~n1541 ;
  assign n1543 = n767 & n1542 ;
  assign n1544 = ~n1539 & ~n1543 ;
  assign n1545 = n1531 & ~n1544 ;
  assign n1546 = ~n1522 & ~n1545 ;
  assign n1547 = \si[13]_pad  & n774 ;
  assign n1548 = ~n814 & ~n823 ;
  assign n1550 = ~n1016 & n1548 ;
  assign n1549 = n1016 & ~n1548 ;
  assign n1551 = ~n774 & ~n1549 ;
  assign n1552 = ~n1550 & n1551 ;
  assign n1553 = ~n1547 & ~n1552 ;
  assign n1554 = ~n767 & ~n1553 ;
  assign n1555 = \P3_IR_reg[31]/NET0131  & ~n694 ;
  assign n1556 = \P3_IR_reg[13]/NET0131  & n1555 ;
  assign n1557 = ~\P3_IR_reg[13]/NET0131  & ~n1555 ;
  assign n1558 = ~n1556 & ~n1557 ;
  assign n1559 = n767 & n1558 ;
  assign n1560 = ~n1554 & ~n1559 ;
  assign n1561 = \P3_reg2_reg[13]/NET0131  & n901 ;
  assign n1562 = \P3_reg0_reg[13]/NET0131  & n905 ;
  assign n1567 = ~n1561 & ~n1562 ;
  assign n1563 = \P3_reg3_reg[13]/NET0131  & ~n916 ;
  assign n1564 = ~n1189 & ~n1563 ;
  assign n1565 = n907 & ~n1564 ;
  assign n1566 = \P3_reg1_reg[13]/NET0131  & n903 ;
  assign n1568 = ~n1565 & ~n1566 ;
  assign n1569 = n1567 & n1568 ;
  assign n1570 = n1560 & ~n1569 ;
  assign n1571 = \P3_IR_reg[31]/NET0131  & ~n675 ;
  assign n1572 = ~\P3_IR_reg[12]/NET0131  & ~n1571 ;
  assign n1573 = \P3_IR_reg[12]/NET0131  & n1571 ;
  assign n1574 = ~n1572 & ~n1573 ;
  assign n1575 = n767 & ~n1574 ;
  assign n1576 = \si[12]_pad  & n774 ;
  assign n1577 = ~n818 & ~n819 ;
  assign n1579 = ~n1044 & n1577 ;
  assign n1578 = n1044 & ~n1577 ;
  assign n1580 = ~n774 & ~n1578 ;
  assign n1581 = ~n1579 & n1580 ;
  assign n1582 = ~n1576 & ~n1581 ;
  assign n1583 = ~n767 & n1582 ;
  assign n1584 = ~n1575 & ~n1583 ;
  assign n1585 = \P3_reg2_reg[12]/NET0131  & n901 ;
  assign n1586 = \P3_reg0_reg[12]/NET0131  & n905 ;
  assign n1592 = ~n1585 & ~n1586 ;
  assign n1587 = ~\P3_reg3_reg[11]/NET0131  & n914 ;
  assign n1588 = \P3_reg3_reg[12]/NET0131  & ~n1587 ;
  assign n1589 = ~n916 & ~n1588 ;
  assign n1590 = n907 & ~n1589 ;
  assign n1591 = \P3_reg1_reg[12]/NET0131  & n903 ;
  assign n1593 = ~n1590 & ~n1591 ;
  assign n1594 = n1592 & n1593 ;
  assign n1595 = ~n1584 & ~n1594 ;
  assign n1596 = ~n1570 & ~n1595 ;
  assign n1597 = ~n1560 & n1569 ;
  assign n1598 = ~n1596 & ~n1597 ;
  assign n1599 = n1546 & n1598 ;
  assign n1600 = n1512 & ~n1521 ;
  assign n1601 = ~n1531 & n1544 ;
  assign n1602 = ~n1600 & ~n1601 ;
  assign n1603 = ~n1522 & ~n1602 ;
  assign n1604 = ~n1599 & ~n1603 ;
  assign n1713 = n1584 & n1594 ;
  assign n1714 = ~n1597 & ~n1713 ;
  assign n1980 = n1546 & n1714 ;
  assign n1629 = \P3_reg0_reg[10]/NET0131  & n905 ;
  assign n1630 = \P3_reg3_reg[10]/NET0131  & ~n913 ;
  assign n1631 = ~n914 & ~n1630 ;
  assign n1632 = n907 & ~n1631 ;
  assign n1635 = ~n1629 & ~n1632 ;
  assign n1633 = \P3_reg1_reg[10]/NET0131  & n903 ;
  assign n1634 = \P3_reg2_reg[10]/NET0131  & n901 ;
  assign n1636 = ~n1633 & ~n1634 ;
  assign n1637 = n1635 & n1636 ;
  assign n1638 = \si[10]_pad  & n774 ;
  assign n1639 = ~n827 & ~n828 ;
  assign n1641 = ~n969 & n1639 ;
  assign n1640 = n969 & ~n1639 ;
  assign n1642 = ~n774 & ~n1640 ;
  assign n1643 = ~n1641 & n1642 ;
  assign n1644 = ~n1638 & ~n1643 ;
  assign n1645 = ~n767 & ~n1644 ;
  assign n1646 = \P3_IR_reg[31]/NET0131  & ~n674 ;
  assign n1647 = \P3_IR_reg[10]/NET0131  & n1646 ;
  assign n1648 = ~\P3_IR_reg[10]/NET0131  & ~n1646 ;
  assign n1649 = ~n1647 & ~n1648 ;
  assign n1650 = n767 & n1649 ;
  assign n1651 = ~n1645 & ~n1650 ;
  assign n1652 = n1637 & ~n1651 ;
  assign n1605 = \P3_reg2_reg[11]/NET0131  & n901 ;
  assign n1606 = \P3_reg0_reg[11]/NET0131  & n905 ;
  assign n1611 = ~n1605 & ~n1606 ;
  assign n1607 = \P3_reg3_reg[11]/NET0131  & ~n914 ;
  assign n1608 = ~n1587 & ~n1607 ;
  assign n1609 = n907 & ~n1608 ;
  assign n1610 = \P3_reg1_reg[11]/NET0131  & n903 ;
  assign n1612 = ~n1609 & ~n1610 ;
  assign n1613 = n1611 & n1612 ;
  assign n1614 = \si[11]_pad  & n774 ;
  assign n1615 = ~n820 & ~n870 ;
  assign n1617 = ~n869 & n1615 ;
  assign n1616 = n869 & ~n1615 ;
  assign n1618 = ~n774 & ~n1616 ;
  assign n1619 = ~n1617 & n1618 ;
  assign n1620 = ~n1614 & ~n1619 ;
  assign n1621 = ~n767 & ~n1620 ;
  assign n1622 = \P3_IR_reg[31]/NET0131  & ~n653 ;
  assign n1623 = \P3_IR_reg[11]/NET0131  & n1622 ;
  assign n1624 = ~\P3_IR_reg[11]/NET0131  & ~n1622 ;
  assign n1625 = ~n1623 & ~n1624 ;
  assign n1626 = n767 & n1625 ;
  assign n1627 = ~n1621 & ~n1626 ;
  assign n1653 = n1613 & ~n1627 ;
  assign n1654 = ~n1652 & ~n1653 ;
  assign n1655 = \P3_reg2_reg[9]/NET0131  & n901 ;
  assign n1656 = \P3_reg3_reg[9]/NET0131  & ~n912 ;
  assign n1657 = ~n913 & ~n1656 ;
  assign n1658 = n907 & ~n1657 ;
  assign n1661 = ~n1655 & ~n1658 ;
  assign n1659 = \P3_reg0_reg[9]/NET0131  & n905 ;
  assign n1660 = \P3_reg1_reg[9]/NET0131  & n903 ;
  assign n1662 = ~n1659 & ~n1660 ;
  assign n1663 = n1661 & n1662 ;
  assign n1664 = \si[9]_pad  & n774 ;
  assign n1665 = ~n829 & ~n865 ;
  assign n1667 = ~n1013 & n1665 ;
  assign n1666 = n1013 & ~n1665 ;
  assign n1668 = ~n774 & ~n1666 ;
  assign n1669 = ~n1667 & n1668 ;
  assign n1670 = ~n1664 & ~n1669 ;
  assign n1671 = ~n767 & ~n1670 ;
  assign n1672 = \P3_IR_reg[31]/NET0131  & ~n691 ;
  assign n1673 = \P3_IR_reg[9]/NET0131  & n1672 ;
  assign n1674 = ~\P3_IR_reg[9]/NET0131  & ~n1672 ;
  assign n1675 = ~n1673 & ~n1674 ;
  assign n1676 = n767 & n1675 ;
  assign n1677 = ~n1671 & ~n1676 ;
  assign n1678 = n1663 & ~n1677 ;
  assign n1707 = ~n1663 & n1677 ;
  assign n1679 = \P3_reg1_reg[8]/NET0131  & n903 ;
  assign n1680 = \P3_reg3_reg[8]/NET0131  & ~n911 ;
  assign n1681 = ~n912 & ~n1680 ;
  assign n1682 = n907 & ~n1681 ;
  assign n1685 = ~n1679 & ~n1682 ;
  assign n1683 = \P3_reg2_reg[8]/NET0131  & n901 ;
  assign n1684 = \P3_reg0_reg[8]/NET0131  & n905 ;
  assign n1686 = ~n1683 & ~n1684 ;
  assign n1687 = n1685 & n1686 ;
  assign n1688 = \si[8]_pad  & n774 ;
  assign n1689 = ~n832 & ~n965 ;
  assign n1690 = ~n860 & ~n864 ;
  assign n1692 = n1689 & n1690 ;
  assign n1691 = ~n1689 & ~n1690 ;
  assign n1693 = ~n774 & ~n1691 ;
  assign n1694 = ~n1692 & n1693 ;
  assign n1695 = ~n1688 & ~n1694 ;
  assign n1696 = ~n767 & ~n1695 ;
  assign n1697 = \P3_IR_reg[31]/NET0131  & ~n648 ;
  assign n1698 = \P3_IR_reg[31]/NET0131  & ~n650 ;
  assign n1699 = ~n1697 & ~n1698 ;
  assign n1700 = \P3_IR_reg[8]/NET0131  & ~n1699 ;
  assign n1701 = ~\P3_IR_reg[8]/NET0131  & n1699 ;
  assign n1702 = ~n1700 & ~n1701 ;
  assign n1703 = n767 & n1702 ;
  assign n1704 = ~n1696 & ~n1703 ;
  assign n1923 = ~n1687 & n1704 ;
  assign n1924 = ~n1707 & ~n1923 ;
  assign n1981 = ~n1678 & ~n1924 ;
  assign n1982 = n1654 & n1981 ;
  assign n1628 = ~n1613 & n1627 ;
  assign n1708 = ~n1637 & n1651 ;
  assign n1922 = ~n1628 & ~n1708 ;
  assign n1983 = ~n1653 & ~n1922 ;
  assign n1984 = ~n1982 & ~n1983 ;
  assign n1721 = \P3_reg2_reg[7]/NET0131  & n901 ;
  assign n1722 = \P3_reg0_reg[7]/NET0131  & n905 ;
  assign n1727 = ~n1721 & ~n1722 ;
  assign n1723 = \P3_reg3_reg[7]/NET0131  & ~n910 ;
  assign n1724 = ~n911 & ~n1723 ;
  assign n1725 = n907 & ~n1724 ;
  assign n1726 = \P3_reg1_reg[7]/NET0131  & n903 ;
  assign n1728 = ~n1725 & ~n1726 ;
  assign n1729 = n1727 & n1728 ;
  assign n1730 = \si[7]_pad  & n774 ;
  assign n1731 = ~n832 & ~n861 ;
  assign n1733 = ~n858 & n1731 ;
  assign n1732 = n858 & ~n1731 ;
  assign n1734 = ~n774 & ~n1732 ;
  assign n1735 = ~n1733 & n1734 ;
  assign n1736 = ~n1730 & ~n1735 ;
  assign n1737 = ~n767 & ~n1736 ;
  assign n1738 = \P3_IR_reg[31]/NET0131  & \P3_IR_reg[6]/NET0131  ;
  assign n1739 = ~n1697 & ~n1738 ;
  assign n1740 = \P3_IR_reg[7]/NET0131  & ~n1739 ;
  assign n1741 = ~\P3_IR_reg[7]/NET0131  & n1739 ;
  assign n1742 = ~n1740 & ~n1741 ;
  assign n1743 = n767 & n1742 ;
  assign n1744 = ~n1737 & ~n1743 ;
  assign n1746 = n1729 & ~n1744 ;
  assign n1747 = \P3_reg2_reg[6]/NET0131  & n901 ;
  assign n1748 = \P3_reg0_reg[6]/NET0131  & n905 ;
  assign n1753 = ~n1747 & ~n1748 ;
  assign n1749 = \P3_reg3_reg[6]/NET0131  & ~n909 ;
  assign n1750 = ~n910 & ~n1749 ;
  assign n1751 = n907 & ~n1750 ;
  assign n1752 = \P3_reg1_reg[6]/NET0131  & n903 ;
  assign n1754 = ~n1751 & ~n1752 ;
  assign n1755 = n1753 & n1754 ;
  assign n1756 = \si[6]_pad  & n774 ;
  assign n1757 = ~n848 & ~n854 ;
  assign n1759 = ~n962 & n1757 ;
  assign n1758 = n962 & ~n1757 ;
  assign n1760 = ~n774 & ~n1758 ;
  assign n1761 = ~n1759 & n1760 ;
  assign n1762 = ~n1756 & ~n1761 ;
  assign n1763 = ~n767 & ~n1762 ;
  assign n1764 = \P3_IR_reg[6]/NET0131  & ~n1697 ;
  assign n1765 = ~\P3_IR_reg[6]/NET0131  & n1697 ;
  assign n1766 = ~n1764 & ~n1765 ;
  assign n1767 = n767 & ~n1766 ;
  assign n1768 = ~n1763 & ~n1767 ;
  assign n1769 = n1755 & ~n1768 ;
  assign n1770 = ~n1746 & ~n1769 ;
  assign n1798 = \P3_reg2_reg[4]/NET0131  & n901 ;
  assign n1799 = \P3_reg0_reg[4]/NET0131  & n905 ;
  assign n1804 = ~n1798 & ~n1799 ;
  assign n1800 = \P3_reg3_reg[3]/NET0131  & \P3_reg3_reg[4]/NET0131  ;
  assign n1801 = ~n908 & ~n1800 ;
  assign n1802 = n907 & ~n1801 ;
  assign n1803 = \P3_reg1_reg[4]/NET0131  & n903 ;
  assign n1805 = ~n1802 & ~n1803 ;
  assign n1806 = n1804 & n1805 ;
  assign n1807 = \si[4]_pad  & n774 ;
  assign n1808 = ~n845 & ~n850 ;
  assign n1810 = n958 & n1808 ;
  assign n1809 = ~n958 & ~n1808 ;
  assign n1811 = ~n774 & ~n1809 ;
  assign n1812 = ~n1810 & n1811 ;
  assign n1813 = ~n1807 & ~n1812 ;
  assign n1814 = ~n767 & ~n1813 ;
  assign n1815 = \P3_IR_reg[31]/NET0131  & ~n646 ;
  assign n1816 = \P3_IR_reg[4]/NET0131  & ~n1815 ;
  assign n1817 = ~\P3_IR_reg[4]/NET0131  & n1815 ;
  assign n1818 = ~n1816 & ~n1817 ;
  assign n1819 = n767 & ~n1818 ;
  assign n1820 = ~n1814 & ~n1819 ;
  assign n1821 = n1806 & ~n1820 ;
  assign n1771 = \P3_reg2_reg[5]/NET0131  & n901 ;
  assign n1772 = \P3_reg0_reg[5]/NET0131  & n905 ;
  assign n1777 = ~n1771 & ~n1772 ;
  assign n1773 = \P3_reg3_reg[5]/NET0131  & ~n908 ;
  assign n1774 = ~n909 & ~n1773 ;
  assign n1775 = n907 & ~n1774 ;
  assign n1776 = \P3_reg1_reg[5]/NET0131  & n903 ;
  assign n1778 = ~n1775 & ~n1776 ;
  assign n1779 = n1777 & n1778 ;
  assign n1780 = \si[5]_pad  & n774 ;
  assign n1781 = ~n847 & ~n850 ;
  assign n1782 = ~n849 & ~n855 ;
  assign n1784 = n1781 & n1782 ;
  assign n1783 = ~n1781 & ~n1782 ;
  assign n1785 = ~n774 & ~n1783 ;
  assign n1786 = ~n1784 & n1785 ;
  assign n1787 = ~n1780 & ~n1786 ;
  assign n1788 = ~n767 & ~n1787 ;
  assign n1789 = \P3_IR_reg[31]/NET0131  & ~n647 ;
  assign n1790 = ~\P3_IR_reg[5]/NET0131  & n1789 ;
  assign n1791 = \P3_IR_reg[5]/NET0131  & ~n1789 ;
  assign n1792 = ~n1790 & ~n1791 ;
  assign n1793 = n767 & ~n1792 ;
  assign n1794 = ~n1788 & ~n1793 ;
  assign n1822 = n1779 & ~n1794 ;
  assign n1823 = ~n1821 & ~n1822 ;
  assign n1824 = \P3_reg2_reg[2]/NET0131  & n901 ;
  assign n1825 = \P3_reg0_reg[2]/NET0131  & n905 ;
  assign n1828 = ~n1824 & ~n1825 ;
  assign n1826 = \P3_reg1_reg[2]/NET0131  & n903 ;
  assign n1827 = \P3_reg3_reg[2]/NET0131  & n907 ;
  assign n1829 = ~n1826 & ~n1827 ;
  assign n1830 = n1828 & n1829 ;
  assign n1831 = \si[2]_pad  & n774 ;
  assign n1832 = ~n833 & ~n841 ;
  assign n1834 = ~n838 & n1832 ;
  assign n1833 = n838 & ~n1832 ;
  assign n1835 = ~n774 & ~n1833 ;
  assign n1836 = ~n1834 & n1835 ;
  assign n1837 = ~n1831 & ~n1836 ;
  assign n1838 = ~n767 & ~n1837 ;
  assign n1839 = \P3_IR_reg[31]/NET0131  & ~n644 ;
  assign n1840 = ~\P3_IR_reg[2]/NET0131  & ~n1839 ;
  assign n1841 = \P3_IR_reg[2]/NET0131  & n1839 ;
  assign n1842 = ~n1840 & ~n1841 ;
  assign n1843 = n767 & n1842 ;
  assign n1844 = ~n1838 & ~n1843 ;
  assign n1845 = n1830 & ~n1844 ;
  assign n1846 = \P3_reg1_reg[3]/NET0131  & n903 ;
  assign n1847 = \P3_reg2_reg[3]/NET0131  & n901 ;
  assign n1850 = ~n1846 & ~n1847 ;
  assign n1848 = \P3_reg0_reg[3]/NET0131  & n905 ;
  assign n1849 = ~\P3_reg3_reg[3]/NET0131  & n907 ;
  assign n1851 = ~n1848 & ~n1849 ;
  assign n1852 = n1850 & n1851 ;
  assign n1853 = \P3_IR_reg[2]/NET0131  & \P3_IR_reg[31]/NET0131  ;
  assign n1854 = ~n1839 & ~n1853 ;
  assign n1855 = \P3_IR_reg[3]/NET0131  & ~n1854 ;
  assign n1856 = ~\P3_IR_reg[3]/NET0131  & n1854 ;
  assign n1857 = ~n1855 & ~n1856 ;
  assign n1858 = n767 & n1857 ;
  assign n1859 = n843 & ~n844 ;
  assign n1860 = ~n840 & ~n844 ;
  assign n1861 = ~n833 & ~n1860 ;
  assign n1862 = ~n955 & n1861 ;
  assign n1863 = ~n1859 & ~n1862 ;
  assign n1864 = ~n774 & ~n1863 ;
  assign n1865 = ~\si[3]_pad  & n774 ;
  assign n1866 = ~n1864 & ~n1865 ;
  assign n1867 = ~n767 & n1866 ;
  assign n1868 = ~n1858 & ~n1867 ;
  assign n1869 = n1852 & ~n1868 ;
  assign n1870 = ~n1845 & ~n1869 ;
  assign n1871 = \P3_reg1_reg[1]/NET0131  & n903 ;
  assign n1872 = \P3_reg3_reg[1]/NET0131  & n907 ;
  assign n1875 = ~n1871 & ~n1872 ;
  assign n1873 = \P3_reg2_reg[1]/NET0131  & n901 ;
  assign n1874 = \P3_reg0_reg[1]/NET0131  & n905 ;
  assign n1876 = ~n1873 & ~n1874 ;
  assign n1877 = n1875 & n1876 ;
  assign n1878 = \P3_IR_reg[1]/NET0131  & ~\P3_IR_reg[31]/NET0131  ;
  assign n1879 = \P3_IR_reg[0]/NET0131  & \P3_IR_reg[1]/NET0131  ;
  assign n1880 = n1839 & ~n1879 ;
  assign n1881 = ~n1878 & ~n1880 ;
  assign n1882 = n767 & ~n1881 ;
  assign n1883 = \si[1]_pad  & n774 ;
  assign n1884 = ~n834 & ~n835 ;
  assign n1886 = ~n836 & n1884 ;
  assign n1885 = n836 & ~n1884 ;
  assign n1887 = ~n774 & ~n1885 ;
  assign n1888 = ~n1886 & n1887 ;
  assign n1889 = ~n1883 & ~n1888 ;
  assign n1890 = ~n767 & ~n1889 ;
  assign n1891 = ~n1882 & ~n1890 ;
  assign n1910 = ~n1877 & n1891 ;
  assign n1892 = n1877 & ~n1891 ;
  assign n1893 = \P3_reg3_reg[0]/NET0131  & n907 ;
  assign n1894 = \P3_reg2_reg[0]/NET0131  & n901 ;
  assign n1897 = ~n1893 & ~n1894 ;
  assign n1895 = \P3_reg0_reg[0]/NET0131  & n905 ;
  assign n1896 = \P3_reg1_reg[0]/NET0131  & n903 ;
  assign n1898 = ~n1895 & ~n1896 ;
  assign n1899 = n1897 & n1898 ;
  assign n1900 = \si[0]_pad  & n774 ;
  assign n1901 = \P1_datao_reg[0]/NET0131  & ~\P2_datao_reg[0]/NET0131  ;
  assign n1902 = ~n836 & ~n1901 ;
  assign n1903 = ~n774 & ~n1902 ;
  assign n1904 = ~n1900 & ~n1903 ;
  assign n1905 = ~n767 & n1904 ;
  assign n1906 = ~\P3_IR_reg[0]/NET0131  & n767 ;
  assign n1907 = ~n1905 & ~n1906 ;
  assign n1965 = n1899 & n1907 ;
  assign n1966 = ~n1892 & ~n1965 ;
  assign n1967 = ~n1910 & ~n1966 ;
  assign n1968 = n1870 & ~n1967 ;
  assign n1911 = ~n1830 & n1844 ;
  assign n1915 = ~n1852 & n1868 ;
  assign n1969 = ~n1911 & ~n1915 ;
  assign n1970 = ~n1869 & ~n1969 ;
  assign n1971 = ~n1968 & ~n1970 ;
  assign n1972 = n1823 & ~n1971 ;
  assign n1795 = ~n1779 & n1794 ;
  assign n1916 = ~n1806 & n1820 ;
  assign n1973 = ~n1795 & ~n1916 ;
  assign n1974 = ~n1822 & ~n1973 ;
  assign n1975 = ~n1972 & ~n1974 ;
  assign n1976 = n1770 & ~n1975 ;
  assign n1745 = ~n1729 & n1744 ;
  assign n1796 = ~n1755 & n1768 ;
  assign n1977 = ~n1745 & ~n1796 ;
  assign n1978 = ~n1746 & ~n1977 ;
  assign n1979 = ~n1976 & ~n1978 ;
  assign n1705 = n1687 & ~n1704 ;
  assign n1706 = ~n1678 & ~n1705 ;
  assign n2009 = n1654 & n1706 ;
  assign n2010 = ~n1979 & n2009 ;
  assign n2011 = n1984 & ~n2010 ;
  assign n2012 = n1980 & ~n2011 ;
  assign n2013 = n1604 & ~n2012 ;
  assign n2014 = n1964 & ~n2013 ;
  assign n2015 = n1962 & ~n2014 ;
  assign n2016 = n1954 & ~n2015 ;
  assign n2017 = n1952 & ~n2016 ;
  assign n1481 = ~n1479 & ~n1480 ;
  assign n1494 = n1408 & n1419 ;
  assign n1495 = ~n1493 & ~n1494 ;
  assign n2018 = n1481 & n1495 ;
  assign n2019 = ~n2017 & n2018 ;
  assign n2020 = ~n2008 & ~n2019 ;
  assign n1943 = \P3_B_reg/NET0131  & n670 ;
  assign n2022 = n708 & ~n1943 ;
  assign n2023 = n2020 & n2022 ;
  assign n2021 = ~n708 & ~n2020 ;
  assign n2024 = ~n687 & ~n701 ;
  assign n2025 = ~n2021 & n2024 ;
  assign n2026 = ~n2023 & n2025 ;
  assign n1709 = ~n1707 & ~n1708 ;
  assign n1710 = ~n1706 & n1709 ;
  assign n1711 = n1654 & ~n1710 ;
  assign n1712 = ~n1628 & ~n1711 ;
  assign n1715 = ~n1570 & ~n1601 ;
  assign n1716 = ~n1714 & n1715 ;
  assign n1717 = n1546 & ~n1716 ;
  assign n1718 = ~n1600 & ~n1717 ;
  assign n1719 = ~n1712 & ~n1718 ;
  assign n1720 = n1604 & ~n1719 ;
  assign n1985 = n1980 & ~n1984 ;
  assign n1986 = n1604 & ~n1985 ;
  assign n1987 = n1979 & n1986 ;
  assign n1988 = ~n1720 & ~n1987 ;
  assign n1989 = n1964 & n1988 ;
  assign n1990 = n1962 & ~n1989 ;
  assign n1944 = ~n1329 & ~n1336 ;
  assign n1945 = n1318 & ~n1944 ;
  assign n1946 = ~n1479 & ~n1945 ;
  assign n1947 = n1495 & n1946 ;
  assign n1991 = n1947 & n1954 ;
  assign n1992 = ~n1990 & n1991 ;
  assign n1995 = n1946 & ~n1994 ;
  assign n1953 = n1947 & ~n1952 ;
  assign n1996 = ~n1330 & ~n1336 ;
  assign n1997 = n1367 & ~n1996 ;
  assign n1998 = ~n1953 & ~n1997 ;
  assign n1999 = ~n1995 & n1998 ;
  assign n2000 = ~n1992 & n1999 ;
  assign n2002 = n708 & ~n2000 ;
  assign n2001 = ~n708 & n2000 ;
  assign n2003 = ~n1943 & ~n2001 ;
  assign n2004 = ~n2002 & n2003 ;
  assign n2005 = n711 & ~n2004 ;
  assign n1393 = n1369 & ~n1392 ;
  assign n1447 = ~n1420 & ~n1446 ;
  assign n1448 = n1393 & n1447 ;
  assign n1476 = n1274 & ~n1475 ;
  assign n1477 = n1448 & n1476 ;
  assign n1797 = ~n1795 & ~n1796 ;
  assign n1908 = ~n1899 & ~n1907 ;
  assign n1909 = ~n1892 & n1908 ;
  assign n1912 = ~n1910 & ~n1911 ;
  assign n1913 = ~n1909 & n1912 ;
  assign n1914 = n1870 & ~n1913 ;
  assign n1917 = ~n1915 & ~n1916 ;
  assign n1918 = ~n1914 & n1917 ;
  assign n1919 = n1823 & ~n1918 ;
  assign n1920 = n1797 & ~n1919 ;
  assign n1921 = n1770 & ~n1920 ;
  assign n1925 = ~n1745 & n1924 ;
  assign n1926 = n1922 & n1925 ;
  assign n1927 = n1596 & n1926 ;
  assign n1928 = n1602 & n1927 ;
  assign n1929 = ~n1921 & n1928 ;
  assign n1930 = ~n1720 & ~n1929 ;
  assign n1203 = n1074 & ~n1202 ;
  assign n1204 = n1080 & n1203 ;
  assign n1169 = ~n1167 & ~n1168 ;
  assign n1931 = n1169 & ~n1497 ;
  assign n1932 = n1204 & n1931 ;
  assign n1933 = ~n1930 & n1932 ;
  assign n1934 = n1477 & n1933 ;
  assign n1086 = n1082 & ~n1085 ;
  assign n1200 = n1169 & ~n1199 ;
  assign n1201 = n1139 & ~n1200 ;
  assign n1205 = ~n1201 & n1204 ;
  assign n1206 = ~n1086 & ~n1205 ;
  assign n1478 = ~n1206 & n1477 ;
  assign n1486 = ~n1273 & ~n1475 ;
  assign n1489 = ~n1487 & ~n1488 ;
  assign n1490 = n1486 & ~n1489 ;
  assign n1491 = n1485 & ~n1490 ;
  assign n1492 = n1448 & ~n1491 ;
  assign n1482 = ~n1368 & ~n1481 ;
  assign n1496 = n1393 & ~n1495 ;
  assign n1935 = ~n1482 & ~n1496 ;
  assign n1936 = ~n1492 & n1935 ;
  assign n1937 = ~n1478 & n1936 ;
  assign n1938 = ~n1934 & n1937 ;
  assign n1940 = ~n708 & n1938 ;
  assign n766 = ~n670 & n735 ;
  assign n1939 = n708 & ~n1938 ;
  assign n1941 = n766 & ~n1939 ;
  assign n1942 = ~n1940 & n1941 ;
  assign n2132 = ~\P3_B_reg/NET0131  & ~n1938 ;
  assign n2133 = n712 & n735 ;
  assign n2134 = ~n2132 & n2133 ;
  assign n2091 = ~n1392 & ~n1493 ;
  assign n2069 = ~n1223 & n1236 ;
  assign n2070 = n1223 & ~n1236 ;
  assign n2071 = ~n2069 & ~n2070 ;
  assign n2122 = n1481 & ~n2071 ;
  assign n2123 = n2091 & n2122 ;
  assign n2030 = ~n1408 & n1419 ;
  assign n2031 = n1408 & ~n1419 ;
  assign n2032 = ~n2030 & ~n2031 ;
  assign n2036 = ~n1522 & ~n1600 ;
  assign n2051 = ~n1637 & ~n1651 ;
  assign n2052 = n1637 & n1651 ;
  assign n2053 = ~n2051 & ~n2052 ;
  assign n2048 = ~n1613 & ~n1627 ;
  assign n2049 = n1613 & n1627 ;
  assign n2050 = ~n2048 & ~n2049 ;
  assign n2054 = ~n1892 & ~n1910 ;
  assign n2055 = ~n1965 & n2054 ;
  assign n2096 = n1823 & ~n1908 ;
  assign n2033 = n1729 & n1744 ;
  assign n2034 = ~n1729 & ~n1744 ;
  assign n2035 = ~n2033 & ~n2034 ;
  assign n2097 = n1973 & ~n2035 ;
  assign n2100 = n2096 & n2097 ;
  assign n2101 = n2055 & n2100 ;
  assign n2104 = ~n2050 & n2101 ;
  assign n2105 = ~n2053 & n2104 ;
  assign n2108 = n2036 & n2105 ;
  assign n2040 = ~n1465 & n1474 ;
  assign n2041 = n1465 & ~n1474 ;
  assign n2042 = ~n2040 & ~n2041 ;
  assign n2046 = ~n1545 & ~n1601 ;
  assign n2109 = ~n2042 & n2046 ;
  assign n2110 = n2108 & n2109 ;
  assign n2056 = ~n1262 & n1272 ;
  assign n2057 = n1262 & ~n1272 ;
  assign n2058 = ~n2056 & ~n2057 ;
  assign n2082 = n1560 & n1569 ;
  assign n2083 = ~n1560 & ~n1569 ;
  assign n2084 = ~n2082 & ~n2083 ;
  assign n2075 = ~n1584 & n1594 ;
  assign n2076 = n1584 & ~n1594 ;
  assign n2077 = ~n2075 & ~n2076 ;
  assign n2065 = n1663 & n1677 ;
  assign n2066 = ~n1663 & ~n1677 ;
  assign n2067 = ~n2065 & ~n2066 ;
  assign n2062 = ~n1687 & ~n1704 ;
  assign n2063 = n1687 & n1704 ;
  assign n2064 = ~n2062 & ~n2063 ;
  assign n2068 = ~n1769 & ~n1796 ;
  assign n2037 = n1852 & n1868 ;
  assign n2038 = ~n1852 & ~n1868 ;
  assign n2039 = ~n2037 & ~n2038 ;
  assign n2047 = ~n1845 & ~n1911 ;
  assign n2098 = ~n2039 & n2047 ;
  assign n2099 = n2068 & n2098 ;
  assign n2102 = ~n2064 & n2099 ;
  assign n2103 = ~n2067 & n2102 ;
  assign n2106 = ~n2077 & n2103 ;
  assign n2107 = ~n2084 & n2106 ;
  assign n2111 = ~n2058 & n2107 ;
  assign n2114 = n2110 & n2111 ;
  assign n2072 = n1121 & n1137 ;
  assign n2073 = ~n1121 & ~n1137 ;
  assign n2074 = ~n2072 & ~n2073 ;
  assign n2079 = n1436 & ~n1445 ;
  assign n2080 = ~n1436 & n1445 ;
  assign n2081 = ~n2079 & ~n2080 ;
  assign n2115 = ~n2074 & ~n2081 ;
  assign n2118 = n2114 & n2115 ;
  assign n2043 = ~n991 & n1000 ;
  assign n2044 = n991 & ~n1000 ;
  assign n2045 = ~n2043 & ~n2044 ;
  assign n2088 = ~n886 & n933 ;
  assign n2089 = n886 & ~n933 ;
  assign n2090 = ~n2088 & ~n2089 ;
  assign n2059 = ~n1185 & ~n1197 ;
  assign n2060 = n1185 & n1197 ;
  assign n2061 = ~n2059 & ~n2060 ;
  assign n2078 = ~n1167 & ~n1170 ;
  assign n2112 = ~n2061 & n2078 ;
  assign n2113 = ~n2090 & n2112 ;
  assign n2119 = ~n2045 & n2113 ;
  assign n2120 = n2118 & n2119 ;
  assign n2093 = ~n1063 & n1072 ;
  assign n2094 = n1063 & ~n1072 ;
  assign n2095 = ~n2093 & ~n2094 ;
  assign n2085 = ~n1029 & n1038 ;
  assign n2086 = n1029 & ~n1038 ;
  assign n2087 = ~n2085 & ~n2086 ;
  assign n2092 = ~n1111 & ~n1202 ;
  assign n2116 = ~n2087 & n2092 ;
  assign n2117 = ~n2095 & n2116 ;
  assign n2121 = n1369 & n2117 ;
  assign n2124 = n2120 & n2121 ;
  assign n2125 = ~n2032 & n2124 ;
  assign n2126 = n2123 & n2125 ;
  assign n2128 = n2022 & n2126 ;
  assign n2127 = ~n708 & ~n2126 ;
  assign n2129 = ~n687 & n701 ;
  assign n2130 = ~n2127 & n2129 ;
  assign n2131 = ~n2128 & n2130 ;
  assign n2027 = \P3_B_reg/NET0131  & ~n711 ;
  assign n2028 = n736 & n2027 ;
  assign n2029 = n737 & ~n1938 ;
  assign n2135 = ~n2028 & ~n2029 ;
  assign n2136 = ~n2131 & n2135 ;
  assign n2137 = ~n2134 & n2136 ;
  assign n2138 = ~n1942 & n2137 ;
  assign n2139 = ~n2005 & n2138 ;
  assign n2140 = ~n2026 & n2139 ;
  assign n2141 = n765 & ~n2140 ;
  assign n2142 = ~n764 & ~n2141 ;
  assign n2143 = \P1_state_reg[0]/NET0131  & ~n670 ;
  assign n2144 = \P3_reg0_reg[29]/NET0131  & ~n2143 ;
  assign n2145 = ~n670 & n757 ;
  assign n2146 = \P3_reg0_reg[29]/NET0131  & n2145 ;
  assign n2147 = ~n670 & ~n757 ;
  assign n2148 = n745 & n752 ;
  assign n2151 = ~\P3_B_reg/NET0131  & n755 ;
  assign n2152 = n2148 & n2151 ;
  assign n2153 = ~\P3_d_reg[0]/NET0131  & ~n2152 ;
  assign n2154 = n752 & ~n2153 ;
  assign n2149 = \P3_B_reg/NET0131  & ~n755 ;
  assign n2150 = n2148 & n2149 ;
  assign n2155 = ~n752 & n755 ;
  assign n2156 = ~n2150 & ~n2155 ;
  assign n2157 = ~n2154 & n2156 ;
  assign n2158 = \P3_d_reg[1]/NET0131  & n752 ;
  assign n2159 = ~n745 & ~n752 ;
  assign n2160 = ~n2158 & ~n2159 ;
  assign n2161 = ~n2150 & n2160 ;
  assign n2162 = ~n2152 & n2161 ;
  assign n2163 = n2157 & n2162 ;
  assign n2164 = \P3_reg0_reg[29]/NET0131  & ~n2163 ;
  assign n2165 = ~n1705 & ~n1746 ;
  assign n2166 = ~n1821 & ~n1917 ;
  assign n2167 = n1912 & ~n1966 ;
  assign n2168 = ~n1821 & n1870 ;
  assign n2169 = ~n2167 & n2168 ;
  assign n2170 = ~n2166 & ~n2169 ;
  assign n2171 = ~n1769 & ~n1822 ;
  assign n2172 = ~n2170 & n2171 ;
  assign n2173 = n2165 & n2172 ;
  assign n2174 = ~n1769 & ~n1797 ;
  assign n2175 = n2165 & n2174 ;
  assign n2176 = ~n1745 & ~n1923 ;
  assign n2177 = ~n1705 & ~n2176 ;
  assign n2178 = ~n2175 & ~n2177 ;
  assign n2179 = ~n2173 & n2178 ;
  assign n2180 = ~n1653 & ~n1713 ;
  assign n2181 = ~n1652 & ~n1678 ;
  assign n2182 = n2180 & n2181 ;
  assign n2183 = ~n2179 & n2182 ;
  assign n2184 = ~n1652 & ~n1709 ;
  assign n2185 = n2180 & n2184 ;
  assign n2186 = n1628 & ~n1713 ;
  assign n2187 = ~n1595 & ~n2186 ;
  assign n2188 = ~n2185 & n2187 ;
  assign n2189 = ~n2183 & n2188 ;
  assign n2190 = ~n1198 & ~n1522 ;
  assign n2191 = ~n1545 & ~n1597 ;
  assign n2192 = n2190 & n2191 ;
  assign n2193 = ~n2189 & n2192 ;
  assign n2194 = ~n1545 & ~n1715 ;
  assign n2195 = n2190 & n2194 ;
  assign n2196 = ~n1198 & n1600 ;
  assign n2197 = ~n1497 & ~n2196 ;
  assign n2198 = ~n2195 & n2197 ;
  assign n2199 = ~n2193 & n2198 ;
  assign n2200 = ~n1083 & ~n1111 ;
  assign n2201 = ~n1138 & ~n1170 ;
  assign n2202 = n2200 & n2201 ;
  assign n2203 = ~n2199 & n2202 ;
  assign n2204 = ~n1138 & ~n1169 ;
  assign n2205 = n2200 & n2204 ;
  assign n2206 = ~n1083 & n1202 ;
  assign n2207 = ~n1073 & ~n2206 ;
  assign n2208 = ~n2205 & n2207 ;
  assign n2209 = ~n2203 & n2208 ;
  assign n2210 = ~n1494 & n1949 ;
  assign n2211 = ~n934 & ~n1488 ;
  assign n2212 = ~n1001 & ~n1075 ;
  assign n2213 = n2211 & n2212 ;
  assign n2214 = n2210 & n2213 ;
  assign n2215 = ~n2209 & n2214 ;
  assign n2216 = ~n1001 & n1039 ;
  assign n2217 = ~n1078 & ~n2216 ;
  assign n2218 = n2211 & ~n2217 ;
  assign n2219 = n1079 & ~n1488 ;
  assign n2220 = ~n1237 & ~n2219 ;
  assign n2221 = ~n2218 & n2220 ;
  assign n2222 = n2210 & ~n2221 ;
  assign n2223 = n1485 & ~n1486 ;
  assign n2224 = n1447 & ~n2223 ;
  assign n2225 = ~n1494 & ~n2224 ;
  assign n2226 = ~n2222 & ~n2225 ;
  assign n2227 = ~n2215 & n2226 ;
  assign n2228 = n2091 & ~n2227 ;
  assign n2229 = ~n2091 & n2227 ;
  assign n2230 = ~n2228 & ~n2229 ;
  assign n2231 = n2163 & n2230 ;
  assign n2232 = ~n2164 & ~n2231 ;
  assign n2233 = ~n735 & ~n736 ;
  assign n2234 = ~n688 & ~n2233 ;
  assign n2235 = ~n2232 & n2234 ;
  assign n2236 = ~n2157 & ~n2162 ;
  assign n2237 = \P3_reg0_reg[29]/NET0131  & ~n2236 ;
  assign n2238 = n724 & n733 ;
  assign n2239 = ~n767 & ~n2238 ;
  assign n2240 = ~n1419 & n2239 ;
  assign n2243 = ~n1336 & ~n1899 ;
  assign n2244 = ~n1877 & n2243 ;
  assign n2245 = ~n1830 & n2244 ;
  assign n2246 = ~n1852 & n2245 ;
  assign n2247 = ~n1779 & ~n1806 ;
  assign n2248 = n2246 & n2247 ;
  assign n2249 = ~n1687 & ~n1729 ;
  assign n2250 = ~n1755 & n2249 ;
  assign n2251 = n2248 & n2250 ;
  assign n2252 = ~n1637 & ~n1663 ;
  assign n2253 = n2251 & n2252 ;
  assign n2254 = ~n1594 & ~n1613 ;
  assign n2255 = n2253 & n2254 ;
  assign n2256 = ~n1521 & ~n1531 ;
  assign n2257 = ~n1152 & ~n1569 ;
  assign n2258 = ~n1197 & n2257 ;
  assign n2259 = n2256 & n2258 ;
  assign n2260 = n2255 & n2259 ;
  assign n2261 = ~n1095 & ~n1121 ;
  assign n2262 = ~n1038 & n2261 ;
  assign n2263 = ~n1072 & n2262 ;
  assign n2264 = n2260 & n2263 ;
  assign n2265 = ~n1000 & ~n1272 ;
  assign n2266 = ~n933 & n2265 ;
  assign n2267 = ~n1236 & n2266 ;
  assign n2268 = n2264 & n2267 ;
  assign n2269 = ~n1445 & ~n1474 ;
  assign n2270 = ~n1419 & n2269 ;
  assign n2271 = ~n1391 & n2270 ;
  assign n2272 = n2268 & n2271 ;
  assign n2274 = n1329 & ~n2272 ;
  assign n2241 = \P3_B_reg/NET0131  & n724 ;
  assign n2242 = ~n2239 & ~n2241 ;
  assign n2273 = ~n1329 & n2272 ;
  assign n2275 = n2242 & ~n2273 ;
  assign n2276 = ~n2274 & n2275 ;
  assign n2277 = ~n2240 & ~n2276 ;
  assign n2278 = n2236 & ~n2277 ;
  assign n2279 = ~n2237 & ~n2278 ;
  assign n2280 = n737 & ~n2279 ;
  assign n2281 = ~n701 & n708 ;
  assign n2282 = ~n670 & ~n687 ;
  assign n2283 = n2281 & n2282 ;
  assign n2284 = ~n710 & ~n2283 ;
  assign n2285 = ~n2281 & n2282 ;
  assign n2286 = ~n2163 & n2285 ;
  assign n2287 = n2284 & ~n2286 ;
  assign n2288 = \P3_reg0_reg[29]/NET0131  & ~n2287 ;
  assign n2289 = n2163 & n2285 ;
  assign n2290 = n1385 & n2289 ;
  assign n2397 = ~n2288 & ~n2290 ;
  assign n2398 = ~n2280 & n2397 ;
  assign n2399 = ~n2235 & n2398 ;
  assign n2291 = ~n1512 & ~n1521 ;
  assign n2292 = ~n2059 & ~n2291 ;
  assign n2293 = n1512 & n1521 ;
  assign n2294 = n1531 & n1544 ;
  assign n2295 = ~n1531 & ~n1544 ;
  assign n2296 = ~n2083 & ~n2295 ;
  assign n2297 = ~n2294 & ~n2296 ;
  assign n2298 = ~n2293 & n2297 ;
  assign n2299 = n2292 & ~n2298 ;
  assign n2300 = ~n2060 & ~n2299 ;
  assign n2305 = ~n1830 & ~n1844 ;
  assign n2306 = ~n1877 & ~n1891 ;
  assign n2307 = n1877 & n1891 ;
  assign n2308 = ~n1899 & n1907 ;
  assign n2309 = ~n2307 & n2308 ;
  assign n2310 = ~n2306 & ~n2309 ;
  assign n2311 = ~n2305 & n2310 ;
  assign n2312 = n1806 & n1820 ;
  assign n2313 = n1830 & n1844 ;
  assign n2314 = ~n2037 & ~n2313 ;
  assign n2315 = ~n2312 & n2314 ;
  assign n2316 = ~n2311 & n2315 ;
  assign n2317 = ~n1806 & ~n1820 ;
  assign n2318 = ~n2038 & ~n2317 ;
  assign n2319 = ~n2312 & ~n2318 ;
  assign n2320 = ~n2316 & ~n2319 ;
  assign n2301 = ~n2033 & ~n2063 ;
  assign n2302 = n1755 & n1768 ;
  assign n2303 = n1779 & n1794 ;
  assign n2304 = ~n2302 & ~n2303 ;
  assign n2321 = n2301 & n2304 ;
  assign n2322 = ~n2320 & n2321 ;
  assign n2323 = ~n1755 & ~n1768 ;
  assign n2324 = ~n1779 & ~n1794 ;
  assign n2325 = ~n2302 & n2324 ;
  assign n2326 = ~n2323 & ~n2325 ;
  assign n2327 = n2301 & ~n2326 ;
  assign n2328 = n2034 & ~n2063 ;
  assign n2329 = ~n2062 & ~n2328 ;
  assign n2330 = ~n2327 & n2329 ;
  assign n2331 = ~n2322 & n2330 ;
  assign n2332 = ~n2049 & ~n2075 ;
  assign n2333 = ~n2052 & ~n2065 ;
  assign n2334 = n2332 & n2333 ;
  assign n2335 = ~n2331 & n2334 ;
  assign n2336 = ~n2052 & n2066 ;
  assign n2337 = ~n2051 & ~n2336 ;
  assign n2338 = n2332 & ~n2337 ;
  assign n2339 = n2048 & ~n2075 ;
  assign n2340 = ~n2076 & ~n2339 ;
  assign n2341 = ~n2338 & n2340 ;
  assign n2342 = ~n2335 & n2341 ;
  assign n2343 = ~n2293 & ~n2294 ;
  assign n2344 = ~n2082 & n2343 ;
  assign n2345 = ~n2060 & n2344 ;
  assign n2346 = ~n2342 & n2345 ;
  assign n2347 = ~n2300 & ~n2346 ;
  assign n2348 = n1152 & n1166 ;
  assign n2349 = n1095 & n1110 ;
  assign n2350 = ~n2093 & ~n2349 ;
  assign n2351 = ~n2072 & n2350 ;
  assign n2352 = ~n2348 & n2351 ;
  assign n2353 = ~n2347 & n2352 ;
  assign n2354 = ~n1152 & ~n1166 ;
  assign n2355 = ~n2072 & n2354 ;
  assign n2356 = ~n2073 & ~n2355 ;
  assign n2357 = n2350 & ~n2356 ;
  assign n2358 = ~n1095 & ~n1110 ;
  assign n2359 = ~n2093 & n2358 ;
  assign n2360 = ~n2094 & ~n2359 ;
  assign n2361 = ~n2357 & n2360 ;
  assign n2362 = ~n2353 & n2361 ;
  assign n2363 = ~n2040 & ~n2056 ;
  assign n2364 = ~n2080 & n2363 ;
  assign n2365 = ~n2030 & n2364 ;
  assign n2366 = ~n2043 & ~n2088 ;
  assign n2367 = ~n2069 & n2366 ;
  assign n2368 = ~n2085 & n2367 ;
  assign n2369 = n2365 & n2368 ;
  assign n2370 = ~n2362 & n2369 ;
  assign n2371 = ~n2044 & ~n2086 ;
  assign n2372 = n2367 & ~n2371 ;
  assign n2373 = ~n2069 & n2089 ;
  assign n2374 = ~n2070 & ~n2373 ;
  assign n2375 = ~n2372 & n2374 ;
  assign n2376 = n2365 & ~n2375 ;
  assign n2377 = ~n2041 & ~n2057 ;
  assign n2378 = ~n2040 & ~n2377 ;
  assign n2379 = ~n2079 & ~n2378 ;
  assign n2380 = ~n2080 & ~n2379 ;
  assign n2381 = ~n2031 & ~n2380 ;
  assign n2382 = ~n2030 & ~n2381 ;
  assign n2383 = ~n2376 & ~n2382 ;
  assign n2384 = ~n2370 & n2383 ;
  assign n2385 = ~n2091 & n2384 ;
  assign n2386 = n2091 & ~n2384 ;
  assign n2387 = ~n2385 & ~n2386 ;
  assign n2388 = n2163 & ~n2387 ;
  assign n2389 = ~n2164 & ~n2388 ;
  assign n2390 = n670 & ~n2024 ;
  assign n2391 = ~n713 & ~n2390 ;
  assign n2392 = ~n2389 & n2391 ;
  assign n2393 = n712 & n2129 ;
  assign n2394 = n2236 & ~n2387 ;
  assign n2395 = ~n2237 & ~n2394 ;
  assign n2396 = n2393 & ~n2395 ;
  assign n2400 = ~n2392 & ~n2396 ;
  assign n2401 = n2399 & n2400 ;
  assign n2402 = n2147 & ~n2401 ;
  assign n2403 = ~n2146 & ~n2402 ;
  assign n2404 = \P1_state_reg[0]/NET0131  & ~n2403 ;
  assign n2405 = ~n2144 & ~n2404 ;
  assign n2406 = \P3_reg2_reg[28]/NET0131  & ~n2143 ;
  assign n2407 = \P3_reg2_reg[28]/NET0131  & n2145 ;
  assign n2408 = ~n2157 & n2162 ;
  assign n2409 = \P3_reg2_reg[28]/NET0131  & ~n2408 ;
  assign n2410 = n1963 & n2012 ;
  assign n2411 = ~n1604 & n1963 ;
  assign n2412 = n1960 & ~n2411 ;
  assign n2413 = ~n2410 & n2412 ;
  assign n2414 = n1085 & n1954 ;
  assign n2415 = ~n2413 & n2414 ;
  assign n2416 = ~n1082 & n1954 ;
  assign n2417 = n1952 & ~n2416 ;
  assign n2418 = ~n2415 & n2417 ;
  assign n2419 = n2032 & ~n2418 ;
  assign n2420 = ~n2032 & n2418 ;
  assign n2421 = ~n2419 & ~n2420 ;
  assign n2422 = n2408 & ~n2421 ;
  assign n2423 = ~n2409 & ~n2422 ;
  assign n2424 = ~n708 & n2129 ;
  assign n2425 = n670 & n2424 ;
  assign n2426 = ~n2423 & n2425 ;
  assign n2431 = ~n1445 & n2239 ;
  assign n2432 = n2268 & n2270 ;
  assign n2433 = n1391 & ~n2432 ;
  assign n2434 = ~n2239 & ~n2272 ;
  assign n2435 = ~n2433 & n2434 ;
  assign n2436 = ~n2431 & ~n2435 ;
  assign n2437 = n2408 & ~n2436 ;
  assign n2438 = ~n2409 & ~n2437 ;
  assign n2439 = n737 & ~n2438 ;
  assign n2427 = n2157 & ~n2162 ;
  assign n2441 = n2285 & n2427 ;
  assign n2442 = n1408 & n2441 ;
  assign n2428 = n2285 & ~n2427 ;
  assign n2429 = ~n710 & ~n2428 ;
  assign n2430 = \P3_reg2_reg[28]/NET0131  & ~n2429 ;
  assign n2440 = ~n1415 & n2283 ;
  assign n2520 = ~n2430 & ~n2440 ;
  assign n2521 = ~n2442 & n2520 ;
  assign n2522 = ~n2439 & n2521 ;
  assign n2523 = ~n2426 & n2522 ;
  assign n2443 = \P3_reg2_reg[28]/NET0131  & ~n2427 ;
  assign n2444 = ~n2049 & ~n2052 ;
  assign n2445 = n2062 & ~n2065 ;
  assign n2446 = ~n2066 & ~n2445 ;
  assign n2447 = n2444 & ~n2446 ;
  assign n2448 = ~n2049 & n2051 ;
  assign n2449 = ~n2048 & ~n2448 ;
  assign n2450 = ~n2447 & n2449 ;
  assign n2451 = ~n2310 & n2314 ;
  assign n2452 = ~n2037 & n2305 ;
  assign n2453 = ~n2038 & ~n2452 ;
  assign n2454 = ~n2451 & n2453 ;
  assign n2455 = ~n2303 & ~n2312 ;
  assign n2456 = ~n2454 & n2455 ;
  assign n2457 = ~n2317 & ~n2324 ;
  assign n2458 = ~n2303 & ~n2457 ;
  assign n2459 = ~n2456 & ~n2458 ;
  assign n2460 = ~n2033 & ~n2302 ;
  assign n2461 = ~n2459 & n2460 ;
  assign n2462 = ~n2033 & n2323 ;
  assign n2463 = ~n2034 & ~n2462 ;
  assign n2464 = ~n2461 & n2463 ;
  assign n2465 = ~n2063 & ~n2065 ;
  assign n2466 = ~n2464 & n2465 ;
  assign n2467 = n2444 & n2466 ;
  assign n2468 = n2450 & ~n2467 ;
  assign n2469 = ~n2060 & ~n2348 ;
  assign n2470 = ~n2072 & n2469 ;
  assign n2471 = ~n2349 & n2470 ;
  assign n2472 = ~n2075 & ~n2082 ;
  assign n2473 = n2343 & n2472 ;
  assign n2474 = n2471 & n2473 ;
  assign n2475 = ~n2468 & n2474 ;
  assign n2476 = ~n2076 & ~n2083 ;
  assign n2477 = n2344 & ~n2476 ;
  assign n2478 = ~n2291 & ~n2295 ;
  assign n2479 = ~n2293 & ~n2478 ;
  assign n2480 = ~n2477 & ~n2479 ;
  assign n2481 = n2471 & ~n2480 ;
  assign n2482 = ~n2073 & ~n2358 ;
  assign n2483 = n2059 & ~n2348 ;
  assign n2484 = ~n2354 & ~n2483 ;
  assign n2485 = ~n2072 & ~n2484 ;
  assign n2486 = n2482 & ~n2485 ;
  assign n2487 = ~n2349 & ~n2486 ;
  assign n2488 = ~n2481 & ~n2487 ;
  assign n2489 = ~n2475 & n2488 ;
  assign n2490 = ~n2069 & n2364 ;
  assign n2491 = ~n2085 & ~n2093 ;
  assign n2492 = n2366 & n2491 ;
  assign n2493 = n2490 & n2492 ;
  assign n2494 = ~n2489 & n2493 ;
  assign n2496 = ~n2085 & n2094 ;
  assign n2497 = ~n2086 & ~n2496 ;
  assign n2498 = n2366 & ~n2497 ;
  assign n2499 = n2044 & ~n2088 ;
  assign n2500 = ~n2089 & ~n2499 ;
  assign n2501 = ~n2498 & n2500 ;
  assign n2502 = n2490 & ~n2501 ;
  assign n2503 = ~n2057 & ~n2070 ;
  assign n2504 = n2364 & ~n2503 ;
  assign n2495 = n2041 & ~n2080 ;
  assign n2505 = ~n2079 & ~n2495 ;
  assign n2506 = ~n2504 & n2505 ;
  assign n2507 = ~n2502 & n2506 ;
  assign n2508 = ~n2494 & n2507 ;
  assign n2509 = n2032 & n2508 ;
  assign n2510 = ~n2032 & ~n2508 ;
  assign n2511 = ~n2509 & ~n2510 ;
  assign n2512 = n2427 & ~n2511 ;
  assign n2513 = ~n2443 & ~n2512 ;
  assign n2514 = n714 & ~n2513 ;
  assign n2515 = ~n2421 & n2427 ;
  assign n2516 = ~n2443 & ~n2515 ;
  assign n2517 = n736 & n2024 ;
  assign n2518 = ~n766 & ~n2517 ;
  assign n2519 = ~n2516 & ~n2518 ;
  assign n2524 = ~n2514 & ~n2519 ;
  assign n2525 = n2523 & n2524 ;
  assign n2526 = n2147 & ~n2525 ;
  assign n2527 = ~n2407 & ~n2526 ;
  assign n2528 = \P1_state_reg[0]/NET0131  & ~n2527 ;
  assign n2529 = ~n2406 & ~n2528 ;
  assign n2530 = ~n1441 & n2145 ;
  assign n2531 = ~n1441 & ~n2163 ;
  assign n2532 = n2304 & ~n2320 ;
  assign n2533 = n2326 & ~n2532 ;
  assign n2534 = n2301 & n2333 ;
  assign n2535 = ~n2533 & n2534 ;
  assign n2536 = ~n2329 & n2333 ;
  assign n2537 = n2337 & ~n2536 ;
  assign n2538 = ~n2535 & n2537 ;
  assign n2539 = ~n2082 & ~n2294 ;
  assign n2540 = n2332 & n2539 ;
  assign n2541 = ~n2538 & n2540 ;
  assign n2542 = ~n2340 & n2539 ;
  assign n2543 = ~n2297 & ~n2542 ;
  assign n2544 = ~n2541 & n2543 ;
  assign n2545 = ~n2293 & n2470 ;
  assign n2546 = ~n2544 & n2545 ;
  assign n2547 = ~n2292 & n2470 ;
  assign n2548 = n2356 & ~n2547 ;
  assign n2549 = ~n2546 & n2548 ;
  assign n2550 = ~n2085 & n2350 ;
  assign n2551 = ~n2043 & n2550 ;
  assign n2552 = ~n2088 & n2363 ;
  assign n2553 = ~n2069 & n2552 ;
  assign n2554 = n2551 & n2553 ;
  assign n2555 = ~n2549 & n2554 ;
  assign n2556 = ~n2085 & ~n2360 ;
  assign n2557 = n2371 & ~n2556 ;
  assign n2558 = ~n2043 & ~n2557 ;
  assign n2559 = n2553 & n2558 ;
  assign n2560 = n2363 & ~n2374 ;
  assign n2561 = ~n2378 & ~n2560 ;
  assign n2562 = ~n2559 & n2561 ;
  assign n2563 = ~n2555 & n2562 ;
  assign n2564 = n2081 & n2563 ;
  assign n2565 = ~n2081 & ~n2563 ;
  assign n2566 = ~n2564 & ~n2565 ;
  assign n2567 = n2163 & ~n2566 ;
  assign n2568 = ~n2531 & ~n2567 ;
  assign n2569 = n2393 & ~n2568 ;
  assign n2570 = n2268 & n2269 ;
  assign n2571 = n1419 & ~n2570 ;
  assign n2572 = ~n2239 & ~n2432 ;
  assign n2573 = ~n2571 & n2572 ;
  assign n2574 = ~n1474 & n2239 ;
  assign n2575 = ~n2573 & ~n2574 ;
  assign n2576 = n2163 & ~n2575 ;
  assign n2577 = ~n2531 & ~n2576 ;
  assign n2578 = n737 & ~n2577 ;
  assign n2579 = ~n2236 & ~n2281 ;
  assign n2580 = n2282 & ~n2579 ;
  assign n2581 = n1436 & n2580 ;
  assign n2582 = ~n2236 & n2285 ;
  assign n2583 = ~n710 & ~n2582 ;
  assign n2584 = ~n1441 & ~n2583 ;
  assign n2624 = ~n2581 & ~n2584 ;
  assign n2625 = ~n2578 & n2624 ;
  assign n2626 = ~n2569 & n2625 ;
  assign n2585 = ~n1441 & ~n2236 ;
  assign n2586 = ~n1483 & ~n1487 ;
  assign n2587 = n2211 & n2586 ;
  assign n2588 = ~n2172 & ~n2174 ;
  assign n2589 = n2165 & n2181 ;
  assign n2590 = ~n2588 & n2589 ;
  assign n2591 = n2177 & n2181 ;
  assign n2592 = ~n2184 & ~n2591 ;
  assign n2593 = ~n2590 & n2592 ;
  assign n2594 = n2180 & n2191 ;
  assign n2595 = ~n2593 & n2594 ;
  assign n2596 = ~n2187 & n2191 ;
  assign n2597 = ~n2194 & ~n2596 ;
  assign n2598 = ~n2595 & n2597 ;
  assign n2599 = n2190 & n2201 ;
  assign n2600 = ~n2598 & n2599 ;
  assign n2601 = ~n2197 & n2201 ;
  assign n2602 = ~n2204 & ~n2601 ;
  assign n2603 = ~n2600 & n2602 ;
  assign n2604 = n2200 & n2212 ;
  assign n2605 = ~n2603 & n2604 ;
  assign n2606 = n2587 & n2605 ;
  assign n2610 = ~n2220 & n2586 ;
  assign n2607 = ~n2207 & n2212 ;
  assign n2608 = n2217 & ~n2607 ;
  assign n2609 = n2587 & ~n2608 ;
  assign n2611 = ~n1483 & ~n1486 ;
  assign n2612 = ~n2609 & ~n2611 ;
  assign n2613 = ~n2610 & n2612 ;
  assign n2614 = ~n2606 & n2613 ;
  assign n2615 = n2081 & ~n2614 ;
  assign n2616 = ~n2081 & n2614 ;
  assign n2617 = ~n2615 & ~n2616 ;
  assign n2618 = n2236 & ~n2617 ;
  assign n2619 = ~n2585 & ~n2618 ;
  assign n2620 = n2234 & ~n2619 ;
  assign n2621 = n2236 & ~n2566 ;
  assign n2622 = ~n2585 & ~n2621 ;
  assign n2623 = n2391 & ~n2622 ;
  assign n2627 = ~n2620 & ~n2623 ;
  assign n2628 = n2626 & n2627 ;
  assign n2629 = n2147 & ~n2628 ;
  assign n2630 = ~n2530 & ~n2629 ;
  assign n2631 = \P1_state_reg[0]/NET0131  & ~n2630 ;
  assign n2632 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[27]/NET0131  ;
  assign n2633 = n765 & ~n1441 ;
  assign n2634 = ~n2632 & ~n2633 ;
  assign n2635 = ~n2631 & n2634 ;
  assign n2636 = ~n1415 & n2145 ;
  assign n2637 = ~n1415 & ~n2163 ;
  assign n2638 = n2163 & ~n2511 ;
  assign n2639 = ~n2637 & ~n2638 ;
  assign n2640 = n2393 & ~n2639 ;
  assign n2642 = n2163 & ~n2436 ;
  assign n2643 = ~n2637 & ~n2642 ;
  assign n2644 = n737 & ~n2643 ;
  assign n2641 = n1408 & n2580 ;
  assign n2645 = ~n1415 & ~n2583 ;
  assign n2653 = ~n2641 & ~n2645 ;
  assign n2654 = ~n2644 & n2653 ;
  assign n2655 = ~n2640 & n2654 ;
  assign n2646 = ~n1415 & ~n2236 ;
  assign n2647 = n2236 & ~n2421 ;
  assign n2648 = ~n2646 & ~n2647 ;
  assign n2649 = n2234 & ~n2648 ;
  assign n2650 = n2236 & ~n2511 ;
  assign n2651 = ~n2646 & ~n2650 ;
  assign n2652 = n2391 & ~n2651 ;
  assign n2656 = ~n2649 & ~n2652 ;
  assign n2657 = n2655 & n2656 ;
  assign n2658 = n2147 & ~n2657 ;
  assign n2659 = ~n2636 & ~n2658 ;
  assign n2660 = \P1_state_reg[0]/NET0131  & ~n2659 ;
  assign n2661 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[28]/NET0131  ;
  assign n2662 = n765 & ~n1415 ;
  assign n2663 = ~n2661 & ~n2662 ;
  assign n2664 = ~n2660 & n2663 ;
  assign n2665 = ~\P1_IR_reg[0]/NET0131  & ~\P1_IR_reg[1]/NET0131  ;
  assign n2666 = ~\P1_IR_reg[2]/NET0131  & n2665 ;
  assign n2667 = ~\P1_IR_reg[3]/NET0131  & n2666 ;
  assign n2668 = ~\P1_IR_reg[4]/NET0131  & ~\P1_IR_reg[5]/NET0131  ;
  assign n2669 = ~\P1_IR_reg[6]/NET0131  & n2668 ;
  assign n2670 = n2667 & n2669 ;
  assign n2671 = ~\P1_IR_reg[7]/NET0131  & ~\P1_IR_reg[8]/NET0131  ;
  assign n2672 = n2670 & n2671 ;
  assign n2673 = ~\P1_IR_reg[10]/NET0131  & ~\P1_IR_reg[9]/NET0131  ;
  assign n2674 = n2672 & n2673 ;
  assign n2675 = ~\P1_IR_reg[11]/NET0131  & ~\P1_IR_reg[12]/NET0131  ;
  assign n2676 = ~\P1_IR_reg[13]/NET0131  & n2675 ;
  assign n2677 = n2674 & n2676 ;
  assign n2678 = ~\P1_IR_reg[16]/NET0131  & ~\P1_IR_reg[17]/NET0131  ;
  assign n2679 = ~\P1_IR_reg[14]/NET0131  & ~\P1_IR_reg[15]/NET0131  ;
  assign n2680 = n2678 & n2679 ;
  assign n2681 = ~\P1_IR_reg[18]/NET0131  & ~\P1_IR_reg[19]/NET0131  ;
  assign n2682 = n2680 & n2681 ;
  assign n2683 = n2677 & n2682 ;
  assign n2684 = \P1_IR_reg[31]/NET0131  & ~n2683 ;
  assign n2685 = ~\P1_IR_reg[20]/NET0131  & ~\P1_IR_reg[21]/NET0131  ;
  assign n2703 = ~\P1_IR_reg[22]/NET0131  & ~\P1_IR_reg[23]/NET0131  ;
  assign n2704 = n2685 & n2703 ;
  assign n2705 = ~\P1_IR_reg[24]/NET0131  & ~\P1_IR_reg[25]/NET0131  ;
  assign n2706 = n2704 & n2705 ;
  assign n2707 = ~\P1_IR_reg[26]/NET0131  & n2706 ;
  assign n2708 = ~\P1_IR_reg[27]/NET0131  & n2707 ;
  assign n2709 = \P1_IR_reg[31]/NET0131  & ~n2708 ;
  assign n2710 = ~n2684 & ~n2709 ;
  assign n2711 = \P1_IR_reg[28]/NET0131  & ~n2710 ;
  assign n2712 = ~\P1_IR_reg[28]/NET0131  & n2710 ;
  assign n2713 = ~n2711 & ~n2712 ;
  assign n2714 = ~\P1_IR_reg[14]/NET0131  & n2676 ;
  assign n2715 = n2674 & n2714 ;
  assign n2716 = ~\P1_IR_reg[15]/NET0131  & ~\P1_IR_reg[18]/NET0131  ;
  assign n2717 = n2678 & n2716 ;
  assign n2718 = n2715 & n2717 ;
  assign n2719 = \P1_IR_reg[31]/NET0131  & ~n2718 ;
  assign n2720 = ~\P1_IR_reg[19]/NET0131  & n2707 ;
  assign n2721 = \P1_IR_reg[31]/NET0131  & ~n2720 ;
  assign n2722 = ~n2719 & ~n2721 ;
  assign n2723 = \P1_IR_reg[27]/NET0131  & ~n2722 ;
  assign n2724 = ~\P1_IR_reg[27]/NET0131  & n2722 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = ~n2713 & ~n2725 ;
  assign n2727 = \P2_datao_reg[22]/NET0131  & n774 ;
  assign n2728 = ~\P2_datao_reg[21]/NET0131  & ~\si[21]_pad  ;
  assign n2729 = \P2_datao_reg[21]/NET0131  & \si[21]_pad  ;
  assign n2730 = \P2_datao_reg[20]/NET0131  & \si[20]_pad  ;
  assign n2731 = ~n2729 & ~n2730 ;
  assign n2732 = ~n2728 & ~n2731 ;
  assign n2733 = ~\P2_datao_reg[19]/NET0131  & ~\si[19]_pad  ;
  assign n2734 = \P2_datao_reg[19]/NET0131  & \si[19]_pad  ;
  assign n2735 = \P2_datao_reg[18]/NET0131  & \si[18]_pad  ;
  assign n2736 = ~n2734 & ~n2735 ;
  assign n2737 = ~n2733 & ~n2736 ;
  assign n2738 = ~\P2_datao_reg[20]/NET0131  & ~\si[20]_pad  ;
  assign n2739 = ~n2728 & ~n2738 ;
  assign n2740 = n2737 & n2739 ;
  assign n2741 = ~n2732 & ~n2740 ;
  assign n2742 = ~\P2_datao_reg[18]/NET0131  & ~\si[18]_pad  ;
  assign n2743 = ~n2733 & ~n2742 ;
  assign n2744 = n2739 & n2743 ;
  assign n2745 = \P2_datao_reg[17]/NET0131  & \si[17]_pad  ;
  assign n2746 = ~\P2_datao_reg[17]/NET0131  & ~\si[17]_pad  ;
  assign n2747 = ~\P2_datao_reg[16]/NET0131  & ~\si[16]_pad  ;
  assign n2748 = ~n2746 & ~n2747 ;
  assign n2749 = \P2_datao_reg[16]/NET0131  & \si[16]_pad  ;
  assign n2750 = ~\P2_datao_reg[15]/NET0131  & ~\si[15]_pad  ;
  assign n2751 = \P2_datao_reg[15]/NET0131  & \si[15]_pad  ;
  assign n2752 = \P2_datao_reg[14]/NET0131  & \si[14]_pad  ;
  assign n2753 = ~n2751 & ~n2752 ;
  assign n2754 = ~n2750 & ~n2753 ;
  assign n2755 = ~n2749 & ~n2754 ;
  assign n2756 = n2748 & ~n2755 ;
  assign n2757 = ~n2745 & ~n2756 ;
  assign n2771 = \P2_datao_reg[5]/NET0131  & \si[5]_pad  ;
  assign n2772 = \P2_datao_reg[4]/NET0131  & \si[4]_pad  ;
  assign n2773 = \P2_datao_reg[3]/NET0131  & \si[3]_pad  ;
  assign n2774 = ~\P2_datao_reg[2]/NET0131  & ~\si[2]_pad  ;
  assign n2775 = \P2_datao_reg[2]/NET0131  & \si[2]_pad  ;
  assign n2776 = ~\P2_datao_reg[1]/NET0131  & ~\si[1]_pad  ;
  assign n2777 = \P2_datao_reg[1]/NET0131  & \si[1]_pad  ;
  assign n2778 = \P2_datao_reg[0]/NET0131  & \si[0]_pad  ;
  assign n2779 = ~n2777 & ~n2778 ;
  assign n2780 = ~n2776 & ~n2779 ;
  assign n2781 = ~n2775 & ~n2780 ;
  assign n2782 = ~n2774 & ~n2781 ;
  assign n2783 = ~n2773 & ~n2782 ;
  assign n2784 = ~\P2_datao_reg[3]/NET0131  & ~\si[3]_pad  ;
  assign n2785 = ~\P2_datao_reg[4]/NET0131  & ~\si[4]_pad  ;
  assign n2786 = ~n2784 & ~n2785 ;
  assign n2787 = ~n2783 & n2786 ;
  assign n2788 = ~n2772 & ~n2787 ;
  assign n2789 = ~n2771 & n2788 ;
  assign n2758 = ~\P2_datao_reg[9]/NET0131  & ~\si[9]_pad  ;
  assign n2763 = ~\P2_datao_reg[8]/NET0131  & ~\si[8]_pad  ;
  assign n2764 = ~\P2_datao_reg[7]/NET0131  & ~\si[7]_pad  ;
  assign n2765 = ~n2763 & ~n2764 ;
  assign n2766 = ~n2758 & n2765 ;
  assign n2790 = ~\P2_datao_reg[6]/NET0131  & ~\si[6]_pad  ;
  assign n2791 = ~\P2_datao_reg[5]/NET0131  & ~\si[5]_pad  ;
  assign n2792 = ~n2790 & ~n2791 ;
  assign n2793 = n2766 & n2792 ;
  assign n2794 = ~n2789 & n2793 ;
  assign n2759 = \P2_datao_reg[9]/NET0131  & \si[9]_pad  ;
  assign n2760 = \P2_datao_reg[8]/NET0131  & \si[8]_pad  ;
  assign n2761 = ~n2759 & ~n2760 ;
  assign n2762 = ~n2758 & ~n2761 ;
  assign n2767 = \P2_datao_reg[7]/NET0131  & \si[7]_pad  ;
  assign n2768 = \P2_datao_reg[6]/NET0131  & \si[6]_pad  ;
  assign n2769 = ~n2767 & ~n2768 ;
  assign n2770 = n2766 & ~n2769 ;
  assign n2795 = ~n2762 & ~n2770 ;
  assign n2796 = ~n2794 & n2795 ;
  assign n2797 = ~\P2_datao_reg[10]/NET0131  & ~\si[10]_pad  ;
  assign n2798 = ~\P2_datao_reg[13]/NET0131  & ~\si[13]_pad  ;
  assign n2799 = ~\P2_datao_reg[12]/NET0131  & ~\si[12]_pad  ;
  assign n2800 = ~\P2_datao_reg[11]/NET0131  & ~\si[11]_pad  ;
  assign n2801 = ~n2799 & ~n2800 ;
  assign n2802 = ~n2798 & n2801 ;
  assign n2803 = ~n2797 & n2802 ;
  assign n2804 = ~n2796 & n2803 ;
  assign n2805 = \P2_datao_reg[13]/NET0131  & \si[13]_pad  ;
  assign n2806 = \P2_datao_reg[12]/NET0131  & \si[12]_pad  ;
  assign n2807 = ~n2805 & ~n2806 ;
  assign n2808 = ~n2798 & ~n2807 ;
  assign n2809 = \P2_datao_reg[11]/NET0131  & \si[11]_pad  ;
  assign n2810 = \P2_datao_reg[10]/NET0131  & \si[10]_pad  ;
  assign n2811 = ~n2809 & ~n2810 ;
  assign n2812 = n2802 & ~n2811 ;
  assign n2813 = ~n2808 & ~n2812 ;
  assign n2814 = ~n2804 & n2813 ;
  assign n2815 = ~\P2_datao_reg[14]/NET0131  & ~\si[14]_pad  ;
  assign n2816 = ~n2750 & ~n2815 ;
  assign n2817 = n2748 & n2816 ;
  assign n2818 = ~n2814 & n2817 ;
  assign n2819 = n2757 & ~n2818 ;
  assign n2820 = n2744 & ~n2819 ;
  assign n2821 = n2741 & ~n2820 ;
  assign n2822 = \P2_datao_reg[22]/NET0131  & \si[22]_pad  ;
  assign n2823 = ~\P2_datao_reg[22]/NET0131  & ~\si[22]_pad  ;
  assign n2824 = ~n2822 & ~n2823 ;
  assign n2826 = n2821 & ~n2824 ;
  assign n2825 = ~n2821 & n2824 ;
  assign n2827 = ~n774 & ~n2825 ;
  assign n2828 = ~n2826 & n2827 ;
  assign n2829 = ~n2727 & ~n2828 ;
  assign n2830 = ~n2726 & ~n2829 ;
  assign n2831 = n2683 & n2706 ;
  assign n2832 = \P1_IR_reg[31]/NET0131  & ~n2831 ;
  assign n2833 = ~\P1_IR_reg[27]/NET0131  & ~\P1_IR_reg[28]/NET0131  ;
  assign n2834 = ~\P1_IR_reg[26]/NET0131  & n2833 ;
  assign n2835 = ~\P1_IR_reg[29]/NET0131  & n2834 ;
  assign n2836 = \P1_IR_reg[31]/NET0131  & ~n2835 ;
  assign n2837 = ~n2832 & ~n2836 ;
  assign n2838 = \P1_IR_reg[30]/NET0131  & ~n2837 ;
  assign n2839 = ~\P1_IR_reg[30]/NET0131  & n2837 ;
  assign n2840 = ~n2838 & ~n2839 ;
  assign n2693 = ~\P1_IR_reg[13]/NET0131  & ~\P1_IR_reg[20]/NET0131  ;
  assign n2694 = n2682 & n2693 ;
  assign n2695 = \P1_IR_reg[31]/NET0131  & ~n2694 ;
  assign n2691 = n2674 & n2675 ;
  assign n2841 = ~\P1_IR_reg[21]/NET0131  & ~\P1_IR_reg[24]/NET0131  ;
  assign n2842 = n2703 & n2841 ;
  assign n2843 = n2691 & n2842 ;
  assign n2844 = ~\P1_IR_reg[25]/NET0131  & n2834 ;
  assign n2845 = n2843 & n2844 ;
  assign n2846 = \P1_IR_reg[31]/NET0131  & ~n2845 ;
  assign n2847 = ~n2695 & ~n2846 ;
  assign n2848 = \P1_IR_reg[29]/NET0131  & ~n2847 ;
  assign n2849 = ~\P1_IR_reg[29]/NET0131  & n2847 ;
  assign n2850 = ~n2848 & ~n2849 ;
  assign n2857 = n2840 & n2850 ;
  assign n2858 = \P1_reg3_reg[19]/NET0131  & \P1_reg3_reg[20]/NET0131  ;
  assign n2859 = \P1_reg3_reg[3]/NET0131  & \P1_reg3_reg[4]/NET0131  ;
  assign n2860 = \P1_reg3_reg[5]/NET0131  & n2859 ;
  assign n2861 = \P1_reg3_reg[6]/NET0131  & n2860 ;
  assign n2862 = \P1_reg3_reg[7]/NET0131  & n2861 ;
  assign n2863 = \P1_reg3_reg[8]/NET0131  & n2862 ;
  assign n2864 = \P1_reg3_reg[9]/NET0131  & n2863 ;
  assign n2865 = \P1_reg3_reg[10]/NET0131  & n2864 ;
  assign n2866 = \P1_reg3_reg[11]/NET0131  & n2865 ;
  assign n2867 = \P1_reg3_reg[12]/NET0131  & n2866 ;
  assign n2868 = \P1_reg3_reg[13]/NET0131  & \P1_reg3_reg[14]/NET0131  ;
  assign n2869 = n2867 & n2868 ;
  assign n2870 = \P1_reg3_reg[15]/NET0131  & n2869 ;
  assign n2871 = \P1_reg3_reg[16]/NET0131  & n2870 ;
  assign n2872 = \P1_reg3_reg[17]/NET0131  & n2871 ;
  assign n2873 = \P1_reg3_reg[18]/NET0131  & n2872 ;
  assign n2874 = n2858 & n2873 ;
  assign n2875 = \P1_reg3_reg[21]/NET0131  & n2874 ;
  assign n2876 = ~\P1_reg3_reg[22]/NET0131  & ~n2875 ;
  assign n2878 = \P1_reg3_reg[18]/NET0131  & \P1_reg3_reg[21]/NET0131  ;
  assign n2879 = \P1_reg3_reg[22]/NET0131  & n2878 ;
  assign n2877 = \P1_reg3_reg[16]/NET0131  & \P1_reg3_reg[17]/NET0131  ;
  assign n2880 = n2858 & n2877 ;
  assign n2881 = n2879 & n2880 ;
  assign n2882 = n2870 & n2881 ;
  assign n2883 = ~n2876 & ~n2882 ;
  assign n2884 = n2857 & n2883 ;
  assign n2855 = ~n2840 & ~n2850 ;
  assign n2856 = \P1_reg0_reg[22]/NET0131  & n2855 ;
  assign n2851 = n2840 & ~n2850 ;
  assign n2852 = \P1_reg2_reg[22]/NET0131  & n2851 ;
  assign n2853 = ~n2840 & n2850 ;
  assign n2854 = \P1_reg1_reg[22]/NET0131  & n2853 ;
  assign n2885 = ~n2852 & ~n2854 ;
  assign n2886 = ~n2856 & n2885 ;
  assign n2887 = ~n2884 & n2886 ;
  assign n3957 = n2830 & n2887 ;
  assign n3259 = \P2_datao_reg[23]/NET0131  & n774 ;
  assign n3260 = ~n2728 & ~n2823 ;
  assign n3146 = ~n2730 & ~n2734 ;
  assign n3147 = ~n2738 & ~n3146 ;
  assign n3261 = ~n2729 & ~n3147 ;
  assign n3262 = n3260 & ~n3261 ;
  assign n3263 = ~n2822 & ~n3262 ;
  assign n2908 = ~n2768 & ~n2771 ;
  assign n2909 = ~n2790 & ~n2908 ;
  assign n2910 = ~n2783 & ~n2784 ;
  assign n2911 = ~n2772 & ~n2910 ;
  assign n2912 = ~n2785 & n2792 ;
  assign n2913 = ~n2911 & n2912 ;
  assign n2914 = ~n2909 & ~n2913 ;
  assign n2904 = ~n2758 & ~n2797 ;
  assign n2915 = n2765 & n2904 ;
  assign n2916 = ~n2914 & n2915 ;
  assign n2902 = ~n2759 & ~n2810 ;
  assign n2903 = ~n2797 & ~n2902 ;
  assign n2905 = ~n2763 & n2904 ;
  assign n2906 = ~n2760 & ~n2767 ;
  assign n2907 = n2905 & ~n2906 ;
  assign n2917 = ~n2903 & ~n2907 ;
  assign n2918 = ~n2916 & n2917 ;
  assign n2919 = n2802 & ~n2815 ;
  assign n2920 = ~n2918 & n2919 ;
  assign n2896 = ~n2752 & ~n2805 ;
  assign n2897 = ~n2815 & ~n2896 ;
  assign n2898 = ~n2798 & ~n2815 ;
  assign n2899 = ~n2799 & n2898 ;
  assign n2900 = ~n2806 & ~n2809 ;
  assign n2901 = n2899 & ~n2900 ;
  assign n2921 = ~n2897 & ~n2901 ;
  assign n2922 = ~n2920 & n2921 ;
  assign n2923 = ~n2742 & ~n2746 ;
  assign n2924 = ~n2747 & ~n2750 ;
  assign n2925 = n2923 & n2924 ;
  assign n2926 = ~n2922 & n2925 ;
  assign n2927 = ~n2735 & ~n2923 ;
  assign n2928 = ~n2735 & ~n2745 ;
  assign n2929 = ~n2742 & ~n2928 ;
  assign n2930 = ~n2747 & n2751 ;
  assign n2931 = ~n2749 & ~n2930 ;
  assign n2932 = ~n2929 & n2931 ;
  assign n2933 = ~n2927 & ~n2932 ;
  assign n2934 = ~n2926 & ~n2933 ;
  assign n3143 = ~n2733 & ~n2738 ;
  assign n3264 = n3143 & n3260 ;
  assign n3265 = ~n2934 & n3264 ;
  assign n3266 = n3263 & ~n3265 ;
  assign n2974 = \P2_datao_reg[23]/NET0131  & \si[23]_pad  ;
  assign n2975 = ~\P2_datao_reg[23]/NET0131  & ~\si[23]_pad  ;
  assign n3267 = ~n2974 & ~n2975 ;
  assign n3269 = n3266 & ~n3267 ;
  assign n3268 = ~n3266 & n3267 ;
  assign n3270 = ~n774 & ~n3268 ;
  assign n3271 = ~n3269 & n3270 ;
  assign n3272 = ~n3259 & ~n3271 ;
  assign n3273 = ~n2726 & ~n3272 ;
  assign n3274 = \P1_reg0_reg[23]/NET0131  & n2855 ;
  assign n3275 = \P1_reg1_reg[23]/NET0131  & n2853 ;
  assign n3281 = ~n3274 & ~n3275 ;
  assign n3276 = \P1_reg2_reg[23]/NET0131  & n2851 ;
  assign n3277 = \P1_reg3_reg[23]/NET0131  & n2882 ;
  assign n3278 = ~\P1_reg3_reg[23]/NET0131  & ~n2882 ;
  assign n3279 = ~n3277 & ~n3278 ;
  assign n3280 = n2857 & n3279 ;
  assign n3282 = ~n3276 & ~n3280 ;
  assign n3283 = n3281 & n3282 ;
  assign n3958 = n3273 & n3283 ;
  assign n3959 = ~n3957 & ~n3958 ;
  assign n3287 = \P2_datao_reg[21]/NET0131  & n774 ;
  assign n3050 = n2765 & n2792 ;
  assign n3051 = ~n2788 & n3050 ;
  assign n3052 = ~n2767 & ~n2909 ;
  assign n3053 = n2765 & ~n3052 ;
  assign n3054 = ~n2760 & ~n3053 ;
  assign n3055 = ~n3051 & n3054 ;
  assign n3056 = n2801 & n2904 ;
  assign n3057 = ~n3055 & n3056 ;
  assign n3058 = ~n2809 & ~n2903 ;
  assign n3059 = n2801 & ~n3058 ;
  assign n3060 = ~n2806 & ~n3059 ;
  assign n3061 = ~n3057 & n3060 ;
  assign n3062 = n2898 & n2924 ;
  assign n3063 = ~n3061 & n3062 ;
  assign n3048 = ~n2751 & ~n2897 ;
  assign n3049 = n2924 & ~n3048 ;
  assign n3064 = ~n2749 & ~n3049 ;
  assign n3065 = ~n3063 & n3064 ;
  assign n3144 = n2923 & n3143 ;
  assign n3145 = ~n3065 & n3144 ;
  assign n3148 = n2929 & n3143 ;
  assign n3149 = ~n3147 & ~n3148 ;
  assign n3150 = ~n3145 & n3149 ;
  assign n3288 = ~n2728 & ~n2729 ;
  assign n3290 = n3150 & ~n3288 ;
  assign n3289 = ~n3150 & n3288 ;
  assign n3291 = ~n774 & ~n3289 ;
  assign n3292 = ~n3290 & n3291 ;
  assign n3293 = ~n3287 & ~n3292 ;
  assign n3294 = ~n2726 & ~n3293 ;
  assign n3298 = ~\P1_reg3_reg[21]/NET0131  & ~n2874 ;
  assign n3299 = ~n2875 & ~n3298 ;
  assign n3300 = n2857 & n3299 ;
  assign n3297 = \P1_reg2_reg[21]/NET0131  & n2851 ;
  assign n3295 = \P1_reg1_reg[21]/NET0131  & n2853 ;
  assign n3296 = \P1_reg0_reg[21]/NET0131  & n2855 ;
  assign n3301 = ~n3295 & ~n3296 ;
  assign n3302 = ~n3297 & n3301 ;
  assign n3303 = ~n3300 & n3302 ;
  assign n3960 = n3294 & n3303 ;
  assign n3944 = ~n3294 & ~n3303 ;
  assign n3581 = \P2_datao_reg[20]/NET0131  & n774 ;
  assign n2984 = n2910 & n2912 ;
  assign n2983 = n2772 & n2792 ;
  assign n2985 = ~n2909 & ~n2983 ;
  assign n2986 = ~n2984 & n2985 ;
  assign n2987 = ~n2764 & ~n2986 ;
  assign n2988 = ~n2767 & ~n2987 ;
  assign n2989 = ~n2800 & n2905 ;
  assign n2990 = ~n2988 & n2989 ;
  assign n2991 = ~n2762 & ~n2810 ;
  assign n2992 = ~n2797 & ~n2800 ;
  assign n2993 = ~n2991 & n2992 ;
  assign n2994 = ~n2809 & ~n2993 ;
  assign n2995 = ~n2990 & n2994 ;
  assign n2996 = ~n2750 & n2899 ;
  assign n2997 = ~n2995 & n2996 ;
  assign n2998 = n2808 & n2816 ;
  assign n2999 = ~n2754 & ~n2998 ;
  assign n3000 = ~n2997 & n2999 ;
  assign n3001 = n2743 & n2748 ;
  assign n3002 = ~n3000 & n3001 ;
  assign n3003 = ~n2745 & ~n2749 ;
  assign n3004 = n2743 & ~n2746 ;
  assign n3005 = ~n3003 & n3004 ;
  assign n3006 = ~n2737 & ~n3005 ;
  assign n3007 = ~n3002 & n3006 ;
  assign n3582 = ~n2730 & ~n2738 ;
  assign n3584 = n3007 & ~n3582 ;
  assign n3583 = ~n3007 & n3582 ;
  assign n3585 = ~n774 & ~n3583 ;
  assign n3586 = ~n3584 & n3585 ;
  assign n3587 = ~n3581 & ~n3586 ;
  assign n3588 = ~n2726 & ~n3587 ;
  assign n2943 = \P1_reg3_reg[19]/NET0131  & n2873 ;
  assign n3592 = ~\P1_reg3_reg[20]/NET0131  & ~n2943 ;
  assign n3593 = ~n2874 & ~n3592 ;
  assign n3594 = n2857 & n3593 ;
  assign n3591 = \P1_reg1_reg[20]/NET0131  & n2853 ;
  assign n3589 = \P1_reg2_reg[20]/NET0131  & n2851 ;
  assign n3590 = \P1_reg0_reg[20]/NET0131  & n2855 ;
  assign n3595 = ~n3589 & ~n3590 ;
  assign n3596 = ~n3591 & n3595 ;
  assign n3597 = ~n3594 & n3596 ;
  assign n3945 = ~n3588 & ~n3597 ;
  assign n4022 = ~n3944 & ~n3945 ;
  assign n4023 = ~n3960 & ~n4022 ;
  assign n4024 = n3959 & n4023 ;
  assign n3941 = ~n3273 & ~n3283 ;
  assign n3942 = ~n2830 & ~n2887 ;
  assign n3943 = ~n3941 & ~n3942 ;
  assign n4025 = ~n3943 & ~n3958 ;
  assign n4026 = ~n4024 & ~n4025 ;
  assign n3961 = n3588 & n3597 ;
  assign n3962 = ~n3960 & ~n3961 ;
  assign n4027 = n3959 & n3962 ;
  assign n2891 = ~\P1_IR_reg[19]/NET0131  & ~n2719 ;
  assign n2892 = \P1_IR_reg[19]/NET0131  & n2719 ;
  assign n2893 = ~n2891 & ~n2892 ;
  assign n2894 = n2726 & ~n2893 ;
  assign n2895 = \P2_datao_reg[19]/NET0131  & n774 ;
  assign n2935 = ~n2733 & ~n2734 ;
  assign n2937 = ~n2934 & n2935 ;
  assign n2936 = n2934 & ~n2935 ;
  assign n2938 = ~n774 & ~n2936 ;
  assign n2939 = ~n2937 & n2938 ;
  assign n2940 = ~n2895 & ~n2939 ;
  assign n2941 = ~n2726 & n2940 ;
  assign n2942 = ~n2894 & ~n2941 ;
  assign n2944 = ~\P1_reg3_reg[19]/NET0131  & ~n2873 ;
  assign n2945 = ~n2943 & ~n2944 ;
  assign n2946 = n2857 & n2945 ;
  assign n2949 = \P1_reg2_reg[19]/NET0131  & n2851 ;
  assign n2947 = \P1_reg0_reg[19]/NET0131  & n2855 ;
  assign n2948 = \P1_reg1_reg[19]/NET0131  & n2853 ;
  assign n2950 = ~n2947 & ~n2948 ;
  assign n2951 = ~n2949 & n2950 ;
  assign n2952 = ~n2946 & n2951 ;
  assign n3967 = n2942 & n2952 ;
  assign n3085 = \P1_IR_reg[31]/NET0131  & ~n2677 ;
  assign n3086 = \P1_IR_reg[31]/NET0131  & ~n2680 ;
  assign n3087 = ~n3085 & ~n3086 ;
  assign n3088 = \P1_IR_reg[18]/NET0131  & ~n3087 ;
  assign n3089 = ~\P1_IR_reg[18]/NET0131  & n3087 ;
  assign n3090 = ~n3088 & ~n3089 ;
  assign n3091 = n2726 & ~n3090 ;
  assign n3092 = \P2_datao_reg[18]/NET0131  & n774 ;
  assign n3093 = ~n2735 & ~n2742 ;
  assign n3095 = ~n2819 & n3093 ;
  assign n3094 = n2819 & ~n3093 ;
  assign n3096 = ~n774 & ~n3094 ;
  assign n3097 = ~n3095 & n3096 ;
  assign n3098 = ~n3092 & ~n3097 ;
  assign n3099 = ~n2726 & n3098 ;
  assign n3100 = ~n3091 & ~n3099 ;
  assign n3101 = ~\P1_reg3_reg[18]/NET0131  & ~n2872 ;
  assign n3102 = ~n2873 & ~n3101 ;
  assign n3103 = n2857 & n3102 ;
  assign n3106 = \P1_reg2_reg[18]/NET0131  & n2851 ;
  assign n3104 = \P1_reg1_reg[18]/NET0131  & n2853 ;
  assign n3105 = \P1_reg0_reg[18]/NET0131  & n2855 ;
  assign n3107 = ~n3104 & ~n3105 ;
  assign n3108 = ~n3106 & n3107 ;
  assign n3109 = ~n3103 & n3108 ;
  assign n3968 = n3100 & n3109 ;
  assign n3969 = ~n3967 & ~n3968 ;
  assign n2692 = \P1_IR_reg[31]/NET0131  & ~n2691 ;
  assign n3038 = ~\P1_IR_reg[13]/NET0131  & n2679 ;
  assign n3039 = ~\P1_IR_reg[16]/NET0131  & n3038 ;
  assign n3040 = \P1_IR_reg[31]/NET0131  & ~n3039 ;
  assign n3041 = ~n2692 & ~n3040 ;
  assign n3042 = \P1_IR_reg[17]/NET0131  & ~n3041 ;
  assign n3043 = ~\P1_IR_reg[17]/NET0131  & n3041 ;
  assign n3044 = ~n3042 & ~n3043 ;
  assign n3045 = n2726 & ~n3044 ;
  assign n3046 = \P2_datao_reg[17]/NET0131  & n774 ;
  assign n3047 = ~n2745 & ~n2746 ;
  assign n3067 = n3047 & ~n3065 ;
  assign n3066 = ~n3047 & n3065 ;
  assign n3068 = ~n774 & ~n3066 ;
  assign n3069 = ~n3067 & n3068 ;
  assign n3070 = ~n3046 & ~n3069 ;
  assign n3071 = ~n2726 & n3070 ;
  assign n3072 = ~n3045 & ~n3071 ;
  assign n3073 = \P1_reg1_reg[17]/NET0131  & n2853 ;
  assign n3074 = \P1_reg0_reg[17]/NET0131  & n2855 ;
  assign n3079 = ~n3073 & ~n3074 ;
  assign n3075 = \P1_reg2_reg[17]/NET0131  & n2851 ;
  assign n3076 = ~\P1_reg3_reg[17]/NET0131  & ~n2871 ;
  assign n3077 = ~n2872 & ~n3076 ;
  assign n3078 = n2857 & n3077 ;
  assign n3080 = ~n3075 & ~n3078 ;
  assign n3081 = n3079 & n3080 ;
  assign n3970 = n3072 & n3081 ;
  assign n3180 = \P1_IR_reg[31]/NET0131  & ~n3038 ;
  assign n3181 = ~n2692 & ~n3180 ;
  assign n3182 = \P1_IR_reg[16]/NET0131  & ~n3181 ;
  assign n3183 = ~\P1_IR_reg[16]/NET0131  & n3181 ;
  assign n3184 = ~n3182 & ~n3183 ;
  assign n3185 = n2726 & ~n3184 ;
  assign n3186 = \P2_datao_reg[16]/NET0131  & n774 ;
  assign n3187 = ~n2747 & ~n2749 ;
  assign n3189 = ~n3000 & n3187 ;
  assign n3188 = n3000 & ~n3187 ;
  assign n3190 = ~n774 & ~n3188 ;
  assign n3191 = ~n3189 & n3190 ;
  assign n3192 = ~n3186 & ~n3191 ;
  assign n3193 = ~n2726 & n3192 ;
  assign n3194 = ~n3185 & ~n3193 ;
  assign n3195 = \P1_reg2_reg[16]/NET0131  & n2851 ;
  assign n3196 = \P1_reg0_reg[16]/NET0131  & n2855 ;
  assign n3201 = ~n3195 & ~n3196 ;
  assign n3197 = \P1_reg1_reg[16]/NET0131  & n2853 ;
  assign n3198 = ~\P1_reg3_reg[16]/NET0131  & ~n2870 ;
  assign n3199 = ~n2871 & ~n3198 ;
  assign n3200 = n2857 & n3199 ;
  assign n3202 = ~n3197 & ~n3200 ;
  assign n3203 = n3201 & n3202 ;
  assign n3950 = ~n3194 & ~n3203 ;
  assign n3951 = ~n3072 & ~n3081 ;
  assign n4028 = ~n3950 & ~n3951 ;
  assign n4029 = ~n3970 & ~n4028 ;
  assign n4030 = n3969 & n4029 ;
  assign n3946 = ~n2942 & ~n2952 ;
  assign n3952 = ~n3100 & ~n3109 ;
  assign n4031 = n3952 & ~n3967 ;
  assign n4032 = ~n3946 & ~n4031 ;
  assign n4033 = ~n4030 & n4032 ;
  assign n3971 = n3194 & n3203 ;
  assign n3972 = ~n3970 & ~n3971 ;
  assign n4034 = n3969 & n3972 ;
  assign n3207 = \P1_IR_reg[14]/NET0131  & ~n3085 ;
  assign n3208 = ~\P1_IR_reg[14]/NET0131  & n3085 ;
  assign n3209 = ~n3207 & ~n3208 ;
  assign n3210 = n2726 & n3209 ;
  assign n3211 = \P2_datao_reg[14]/NET0131  & n774 ;
  assign n3212 = ~n2752 & ~n2815 ;
  assign n3214 = ~n2814 & n3212 ;
  assign n3213 = n2814 & ~n3212 ;
  assign n3215 = ~n774 & ~n3213 ;
  assign n3216 = ~n3214 & n3215 ;
  assign n3217 = ~n3211 & ~n3216 ;
  assign n3218 = ~n2726 & n3217 ;
  assign n3219 = ~n3210 & ~n3218 ;
  assign n3220 = \P1_reg0_reg[14]/NET0131  & n2855 ;
  assign n3221 = \P1_reg3_reg[13]/NET0131  & n2867 ;
  assign n3222 = ~\P1_reg3_reg[14]/NET0131  & ~n3221 ;
  assign n3223 = ~n2869 & ~n3222 ;
  assign n3224 = n2857 & n3223 ;
  assign n3227 = ~n3220 & ~n3224 ;
  assign n3225 = \P1_reg2_reg[14]/NET0131  & n2851 ;
  assign n3226 = \P1_reg1_reg[14]/NET0131  & n2853 ;
  assign n3228 = ~n3225 & ~n3226 ;
  assign n3229 = n3227 & n3228 ;
  assign n3873 = n3219 & n3229 ;
  assign n3601 = \P1_IR_reg[31]/NET0131  & ~n2715 ;
  assign n3602 = \P1_IR_reg[15]/NET0131  & n3601 ;
  assign n3603 = ~\P1_IR_reg[15]/NET0131  & ~n3601 ;
  assign n3604 = ~n3602 & ~n3603 ;
  assign n3605 = n2726 & ~n3604 ;
  assign n3606 = \P2_datao_reg[15]/NET0131  & n774 ;
  assign n3607 = ~n2750 & ~n2751 ;
  assign n3609 = ~n2922 & n3607 ;
  assign n3608 = n2922 & ~n3607 ;
  assign n3610 = ~n774 & ~n3608 ;
  assign n3611 = ~n3609 & n3610 ;
  assign n3612 = ~n3606 & ~n3611 ;
  assign n3613 = ~n2726 & n3612 ;
  assign n3614 = ~n3605 & ~n3613 ;
  assign n3615 = \P1_reg2_reg[15]/NET0131  & n2851 ;
  assign n3616 = \P1_reg1_reg[15]/NET0131  & n2853 ;
  assign n3621 = ~n3615 & ~n3616 ;
  assign n3617 = ~\P1_reg3_reg[15]/NET0131  & ~n2869 ;
  assign n3618 = ~n2870 & ~n3617 ;
  assign n3619 = n2857 & n3618 ;
  assign n3620 = \P1_reg0_reg[15]/NET0131  & n2855 ;
  assign n3622 = ~n3619 & ~n3620 ;
  assign n3623 = n3621 & n3622 ;
  assign n3874 = n3614 & n3623 ;
  assign n3875 = ~n3873 & ~n3874 ;
  assign n3333 = ~\P1_IR_reg[13]/NET0131  & ~n2692 ;
  assign n3334 = \P1_IR_reg[13]/NET0131  & n2692 ;
  assign n3335 = ~n3333 & ~n3334 ;
  assign n3336 = n2726 & ~n3335 ;
  assign n3337 = \P2_datao_reg[13]/NET0131  & n774 ;
  assign n3338 = ~n2798 & ~n2805 ;
  assign n3340 = ~n3061 & n3338 ;
  assign n3339 = n3061 & ~n3338 ;
  assign n3341 = ~n774 & ~n3339 ;
  assign n3342 = ~n3340 & n3341 ;
  assign n3343 = ~n3337 & ~n3342 ;
  assign n3344 = ~n2726 & n3343 ;
  assign n3345 = ~n3336 & ~n3344 ;
  assign n3346 = \P1_reg2_reg[13]/NET0131  & n2851 ;
  assign n3347 = \P1_reg0_reg[13]/NET0131  & n2855 ;
  assign n3352 = ~n3346 & ~n3347 ;
  assign n3348 = ~\P1_reg3_reg[13]/NET0131  & ~n2867 ;
  assign n3349 = ~n3221 & ~n3348 ;
  assign n3350 = n2857 & n3349 ;
  assign n3351 = \P1_reg1_reg[13]/NET0131  & n2853 ;
  assign n3353 = ~n3350 & ~n3351 ;
  assign n3354 = n3352 & n3353 ;
  assign n3876 = ~n3345 & ~n3354 ;
  assign n3877 = n3345 & n3354 ;
  assign n3233 = \P1_IR_reg[31]/NET0131  & ~n2674 ;
  assign n3627 = \P1_IR_reg[11]/NET0131  & \P1_IR_reg[31]/NET0131  ;
  assign n3628 = ~n3233 & ~n3627 ;
  assign n3629 = \P1_IR_reg[12]/NET0131  & ~n3628 ;
  assign n3630 = ~\P1_IR_reg[12]/NET0131  & n3628 ;
  assign n3631 = ~n3629 & ~n3630 ;
  assign n3632 = n2726 & ~n3631 ;
  assign n3633 = \P2_datao_reg[12]/NET0131  & n774 ;
  assign n3634 = ~n2799 & ~n2806 ;
  assign n3636 = ~n2995 & n3634 ;
  assign n3635 = n2995 & ~n3634 ;
  assign n3637 = ~n774 & ~n3635 ;
  assign n3638 = ~n3636 & n3637 ;
  assign n3639 = ~n3633 & ~n3638 ;
  assign n3640 = ~n2726 & n3639 ;
  assign n3641 = ~n3632 & ~n3640 ;
  assign n3642 = \P1_reg2_reg[12]/NET0131  & n2851 ;
  assign n3643 = \P1_reg1_reg[12]/NET0131  & n2853 ;
  assign n3648 = ~n3642 & ~n3643 ;
  assign n3644 = ~\P1_reg3_reg[12]/NET0131  & ~n2866 ;
  assign n3645 = ~n2867 & ~n3644 ;
  assign n3646 = n2857 & n3645 ;
  assign n3647 = \P1_reg0_reg[12]/NET0131  & n2855 ;
  assign n3649 = ~n3646 & ~n3647 ;
  assign n3650 = n3648 & n3649 ;
  assign n3878 = ~n3641 & ~n3650 ;
  assign n3879 = ~n3877 & n3878 ;
  assign n3880 = ~n3876 & ~n3879 ;
  assign n3881 = n3875 & ~n3880 ;
  assign n3882 = ~n3614 & ~n3623 ;
  assign n3883 = ~n3219 & ~n3229 ;
  assign n3884 = ~n3874 & n3883 ;
  assign n3885 = ~n3882 & ~n3884 ;
  assign n3886 = ~n3881 & n3885 ;
  assign n3900 = n3641 & n3650 ;
  assign n3901 = ~n3877 & ~n3900 ;
  assign n4035 = n3875 & n3901 ;
  assign n3234 = \P1_IR_reg[11]/NET0131  & ~n3233 ;
  assign n3235 = ~\P1_IR_reg[11]/NET0131  & n3233 ;
  assign n3236 = ~n3234 & ~n3235 ;
  assign n3237 = n2726 & n3236 ;
  assign n3238 = \P2_datao_reg[11]/NET0131  & n774 ;
  assign n3239 = ~n2800 & ~n2809 ;
  assign n3241 = ~n2918 & n3239 ;
  assign n3240 = n2918 & ~n3239 ;
  assign n3242 = ~n774 & ~n3240 ;
  assign n3243 = ~n3241 & n3242 ;
  assign n3244 = ~n3238 & ~n3243 ;
  assign n3245 = ~n2726 & n3244 ;
  assign n3246 = ~n3237 & ~n3245 ;
  assign n3247 = \P1_reg2_reg[11]/NET0131  & n2851 ;
  assign n3248 = \P1_reg1_reg[11]/NET0131  & n2853 ;
  assign n3253 = ~n3247 & ~n3248 ;
  assign n3249 = ~\P1_reg3_reg[11]/NET0131  & ~n2865 ;
  assign n3250 = ~n2866 & ~n3249 ;
  assign n3251 = n2857 & n3250 ;
  assign n3252 = \P1_reg0_reg[11]/NET0131  & n2855 ;
  assign n3254 = ~n3251 & ~n3252 ;
  assign n3255 = n3253 & n3254 ;
  assign n3888 = n3246 & n3255 ;
  assign n3307 = \P1_IR_reg[31]/NET0131  & ~n2672 ;
  assign n3654 = \P1_IR_reg[31]/NET0131  & \P1_IR_reg[9]/NET0131  ;
  assign n3655 = ~n3307 & ~n3654 ;
  assign n3656 = \P1_IR_reg[10]/NET0131  & ~n3655 ;
  assign n3657 = ~\P1_IR_reg[10]/NET0131  & n3655 ;
  assign n3658 = ~n3656 & ~n3657 ;
  assign n3659 = n2726 & ~n3658 ;
  assign n3660 = \P2_datao_reg[10]/NET0131  & n774 ;
  assign n3661 = ~n2797 & ~n2810 ;
  assign n3663 = ~n2796 & n3661 ;
  assign n3662 = n2796 & ~n3661 ;
  assign n3664 = ~n774 & ~n3662 ;
  assign n3665 = ~n3663 & n3664 ;
  assign n3666 = ~n3660 & ~n3665 ;
  assign n3667 = ~n2726 & n3666 ;
  assign n3668 = ~n3659 & ~n3667 ;
  assign n3669 = \P1_reg1_reg[10]/NET0131  & n2853 ;
  assign n3670 = \P1_reg2_reg[10]/NET0131  & n2851 ;
  assign n3675 = ~n3669 & ~n3670 ;
  assign n3671 = ~\P1_reg3_reg[10]/NET0131  & ~n2864 ;
  assign n3672 = ~n2865 & ~n3671 ;
  assign n3673 = n2857 & n3672 ;
  assign n3674 = \P1_reg0_reg[10]/NET0131  & n2855 ;
  assign n3676 = ~n3673 & ~n3674 ;
  assign n3677 = n3675 & n3676 ;
  assign n3889 = n3668 & n3677 ;
  assign n3890 = ~n3888 & ~n3889 ;
  assign n3308 = \P1_IR_reg[9]/NET0131  & ~n3307 ;
  assign n3309 = ~\P1_IR_reg[9]/NET0131  & n3307 ;
  assign n3310 = ~n3308 & ~n3309 ;
  assign n3311 = n2726 & n3310 ;
  assign n3312 = \P2_datao_reg[9]/NET0131  & n774 ;
  assign n3313 = ~n2758 & ~n2759 ;
  assign n3315 = ~n3055 & n3313 ;
  assign n3314 = n3055 & ~n3313 ;
  assign n3316 = ~n774 & ~n3314 ;
  assign n3317 = ~n3315 & n3316 ;
  assign n3318 = ~n3312 & ~n3317 ;
  assign n3319 = ~n2726 & n3318 ;
  assign n3320 = ~n3311 & ~n3319 ;
  assign n3321 = \P1_reg2_reg[9]/NET0131  & n2851 ;
  assign n3322 = \P1_reg1_reg[9]/NET0131  & n2853 ;
  assign n3327 = ~n3321 & ~n3322 ;
  assign n3323 = ~\P1_reg3_reg[9]/NET0131  & ~n2863 ;
  assign n3324 = ~n2864 & ~n3323 ;
  assign n3325 = n2857 & n3324 ;
  assign n3326 = \P1_reg0_reg[9]/NET0131  & n2855 ;
  assign n3328 = ~n3325 & ~n3326 ;
  assign n3329 = n3327 & n3328 ;
  assign n3891 = n3320 & n3329 ;
  assign n3894 = ~n3320 & ~n3329 ;
  assign n3555 = \P1_IR_reg[31]/NET0131  & ~n2670 ;
  assign n3799 = \P1_IR_reg[31]/NET0131  & \P1_IR_reg[7]/NET0131  ;
  assign n3800 = ~n3555 & ~n3799 ;
  assign n3801 = \P1_IR_reg[8]/NET0131  & ~n3800 ;
  assign n3802 = ~\P1_IR_reg[8]/NET0131  & n3800 ;
  assign n3803 = ~n3801 & ~n3802 ;
  assign n3804 = n2726 & ~n3803 ;
  assign n3805 = \P2_datao_reg[8]/NET0131  & n774 ;
  assign n3806 = ~n2760 & ~n2763 ;
  assign n3808 = ~n2988 & n3806 ;
  assign n3807 = n2988 & ~n3806 ;
  assign n3809 = ~n774 & ~n3807 ;
  assign n3810 = ~n3808 & n3809 ;
  assign n3811 = ~n3805 & ~n3810 ;
  assign n3812 = ~n2726 & n3811 ;
  assign n3813 = ~n3804 & ~n3812 ;
  assign n3814 = \P1_reg1_reg[8]/NET0131  & n2853 ;
  assign n3815 = \P1_reg2_reg[8]/NET0131  & n2851 ;
  assign n3820 = ~n3814 & ~n3815 ;
  assign n3816 = \P1_reg0_reg[8]/NET0131  & n2855 ;
  assign n3817 = ~\P1_reg3_reg[8]/NET0131  & ~n2862 ;
  assign n3818 = ~n2863 & ~n3817 ;
  assign n3819 = n2857 & n3818 ;
  assign n3821 = ~n3816 & ~n3819 ;
  assign n3822 = n3820 & n3821 ;
  assign n3932 = ~n3813 & ~n3822 ;
  assign n3933 = ~n3894 & ~n3932 ;
  assign n4036 = ~n3891 & ~n3933 ;
  assign n4037 = n3890 & n4036 ;
  assign n3887 = ~n3246 & ~n3255 ;
  assign n3895 = ~n3668 & ~n3677 ;
  assign n4038 = ~n3888 & n3895 ;
  assign n4039 = ~n3887 & ~n4038 ;
  assign n4040 = ~n4037 & n4039 ;
  assign n3358 = \P1_reg0_reg[2]/NET0131  & n2855 ;
  assign n3359 = \P1_reg3_reg[2]/NET0131  & n2857 ;
  assign n3362 = ~n3358 & ~n3359 ;
  assign n3360 = \P1_reg2_reg[2]/NET0131  & n2851 ;
  assign n3361 = \P1_reg1_reg[2]/NET0131  & n2853 ;
  assign n3363 = ~n3360 & ~n3361 ;
  assign n3364 = n3362 & n3363 ;
  assign n3365 = \P2_datao_reg[2]/NET0131  & n774 ;
  assign n3366 = ~n2774 & ~n2775 ;
  assign n3368 = n2780 & n3366 ;
  assign n3367 = ~n2780 & ~n3366 ;
  assign n3369 = ~n774 & ~n3367 ;
  assign n3370 = ~n3368 & n3369 ;
  assign n3371 = ~n3365 & ~n3370 ;
  assign n3372 = ~n2726 & ~n3371 ;
  assign n3373 = \P1_IR_reg[31]/NET0131  & ~n2665 ;
  assign n3374 = \P1_IR_reg[2]/NET0131  & ~n3373 ;
  assign n3375 = ~\P1_IR_reg[2]/NET0131  & n3373 ;
  assign n3376 = ~n3374 & ~n3375 ;
  assign n3377 = n2726 & ~n3376 ;
  assign n3378 = ~n3372 & ~n3377 ;
  assign n3379 = n3364 & ~n3378 ;
  assign n3750 = \P1_reg2_reg[3]/NET0131  & n2851 ;
  assign n3751 = \P1_reg1_reg[3]/NET0131  & n2853 ;
  assign n3754 = ~n3750 & ~n3751 ;
  assign n3752 = ~\P1_reg3_reg[3]/NET0131  & n2857 ;
  assign n3753 = \P1_reg0_reg[3]/NET0131  & n2855 ;
  assign n3755 = ~n3752 & ~n3753 ;
  assign n3756 = n3754 & n3755 ;
  assign n3757 = \P2_datao_reg[3]/NET0131  & n774 ;
  assign n3758 = ~n2773 & ~n2784 ;
  assign n3760 = n2782 & n3758 ;
  assign n3759 = ~n2782 & ~n3758 ;
  assign n3761 = ~n774 & ~n3759 ;
  assign n3762 = ~n3760 & n3761 ;
  assign n3763 = ~n3757 & ~n3762 ;
  assign n3764 = ~n2726 & ~n3763 ;
  assign n3765 = \P1_IR_reg[31]/NET0131  & ~n2666 ;
  assign n3766 = \P1_IR_reg[3]/NET0131  & ~n3765 ;
  assign n3767 = ~\P1_IR_reg[3]/NET0131  & n3765 ;
  assign n3768 = ~n3766 & ~n3767 ;
  assign n3769 = n2726 & ~n3768 ;
  assign n3770 = ~n3764 & ~n3769 ;
  assign n3771 = n3756 & ~n3770 ;
  assign n3922 = ~n3379 & ~n3771 ;
  assign n3698 = \P1_reg1_reg[1]/NET0131  & n2853 ;
  assign n3699 = \P1_reg3_reg[1]/NET0131  & n2857 ;
  assign n3702 = ~n3698 & ~n3699 ;
  assign n3700 = \P1_reg2_reg[1]/NET0131  & n2851 ;
  assign n3701 = \P1_reg0_reg[1]/NET0131  & n2855 ;
  assign n3703 = ~n3700 & ~n3701 ;
  assign n3704 = n3702 & n3703 ;
  assign n3705 = \P1_IR_reg[1]/NET0131  & ~\P1_IR_reg[31]/NET0131  ;
  assign n3706 = \P1_IR_reg[0]/NET0131  & \P1_IR_reg[1]/NET0131  ;
  assign n3707 = n3373 & ~n3706 ;
  assign n3708 = ~n3705 & ~n3707 ;
  assign n3709 = n2726 & ~n3708 ;
  assign n3710 = ~\P2_datao_reg[1]/NET0131  & n774 ;
  assign n3711 = ~n2776 & ~n2777 ;
  assign n3713 = ~n2778 & n3711 ;
  assign n3712 = n2778 & ~n3711 ;
  assign n3714 = ~n774 & ~n3712 ;
  assign n3715 = ~n3713 & n3714 ;
  assign n3716 = ~n3710 & ~n3715 ;
  assign n3717 = ~n2726 & n3716 ;
  assign n3718 = ~n3709 & ~n3717 ;
  assign n3720 = n3704 & ~n3718 ;
  assign n3681 = \P1_reg3_reg[0]/NET0131  & n2857 ;
  assign n3682 = \P1_reg0_reg[0]/NET0131  & n2855 ;
  assign n3685 = ~n3681 & ~n3682 ;
  assign n3683 = \P1_reg2_reg[0]/NET0131  & n2851 ;
  assign n3684 = \P1_reg1_reg[0]/NET0131  & n2853 ;
  assign n3686 = ~n3683 & ~n3684 ;
  assign n3687 = n3685 & n3686 ;
  assign n3688 = \si[0]_pad  & ~n774 ;
  assign n3689 = ~\P2_datao_reg[0]/NET0131  & ~n3688 ;
  assign n3690 = ~n774 & n2778 ;
  assign n3691 = ~n3689 & ~n3690 ;
  assign n3692 = ~n2726 & n3691 ;
  assign n3693 = \P1_IR_reg[0]/NET0131  & n2726 ;
  assign n3694 = ~n3692 & ~n3693 ;
  assign n3695 = n3687 & ~n3694 ;
  assign n3719 = ~n3704 & n3718 ;
  assign n4041 = n3695 & ~n3719 ;
  assign n4042 = ~n3720 & ~n4041 ;
  assign n4043 = n3922 & n4042 ;
  assign n3380 = ~n3364 & n3378 ;
  assign n3772 = ~n3756 & n3770 ;
  assign n3924 = ~n3380 & ~n3772 ;
  assign n4044 = ~n3771 & ~n3924 ;
  assign n4045 = ~n4043 & ~n4044 ;
  assign n3556 = \P1_IR_reg[7]/NET0131  & ~n3555 ;
  assign n3557 = ~\P1_IR_reg[7]/NET0131  & n3555 ;
  assign n3558 = ~n3556 & ~n3557 ;
  assign n3559 = n2726 & n3558 ;
  assign n3560 = \P2_datao_reg[7]/NET0131  & n774 ;
  assign n3561 = ~n2764 & ~n2767 ;
  assign n3563 = ~n2914 & n3561 ;
  assign n3562 = n2914 & ~n3561 ;
  assign n3564 = ~n774 & ~n3562 ;
  assign n3565 = ~n3563 & n3564 ;
  assign n3566 = ~n3560 & ~n3565 ;
  assign n3567 = ~n2726 & n3566 ;
  assign n3568 = ~n3559 & ~n3567 ;
  assign n3569 = \P1_reg2_reg[7]/NET0131  & n2851 ;
  assign n3570 = \P1_reg1_reg[7]/NET0131  & n2853 ;
  assign n3575 = ~n3569 & ~n3570 ;
  assign n3571 = \P1_reg0_reg[7]/NET0131  & n2855 ;
  assign n3572 = ~\P1_reg3_reg[7]/NET0131  & ~n2861 ;
  assign n3573 = ~n2862 & ~n3572 ;
  assign n3574 = n2857 & n3573 ;
  assign n3576 = ~n3571 & ~n3574 ;
  assign n3577 = n3575 & n3576 ;
  assign n3909 = n3568 & n3577 ;
  assign n3722 = ~\P2_datao_reg[6]/NET0131  & n774 ;
  assign n3723 = ~n2768 & ~n2790 ;
  assign n3724 = ~n2789 & ~n2791 ;
  assign n3726 = n3723 & ~n3724 ;
  assign n3725 = ~n3723 & n3724 ;
  assign n3727 = ~n774 & ~n3725 ;
  assign n3728 = ~n3726 & n3727 ;
  assign n3729 = ~n3722 & ~n3728 ;
  assign n3730 = ~n2726 & ~n3729 ;
  assign n3121 = \P1_IR_reg[31]/NET0131  & ~n2667 ;
  assign n3731 = \P1_IR_reg[31]/NET0131  & ~n2668 ;
  assign n3732 = ~n3121 & ~n3731 ;
  assign n3733 = \P1_IR_reg[6]/NET0131  & ~n3732 ;
  assign n3734 = ~\P1_IR_reg[6]/NET0131  & n3732 ;
  assign n3735 = ~n3733 & ~n3734 ;
  assign n3736 = n2726 & ~n3735 ;
  assign n3737 = ~n3730 & ~n3736 ;
  assign n3738 = ~\P1_reg3_reg[6]/NET0131  & ~n2860 ;
  assign n3739 = ~n2861 & ~n3738 ;
  assign n3740 = n2857 & n3739 ;
  assign n3741 = \P1_reg2_reg[6]/NET0131  & n2851 ;
  assign n3744 = ~n3740 & ~n3741 ;
  assign n3742 = \P1_reg0_reg[6]/NET0131  & n2855 ;
  assign n3743 = \P1_reg1_reg[6]/NET0131  & n2853 ;
  assign n3745 = ~n3742 & ~n3743 ;
  assign n3746 = n3744 & n3745 ;
  assign n3910 = n3737 & n3746 ;
  assign n3911 = ~n3909 & ~n3910 ;
  assign n3774 = ~\P2_datao_reg[4]/NET0131  & n774 ;
  assign n3775 = ~n2772 & ~n2785 ;
  assign n3777 = ~n2910 & n3775 ;
  assign n3776 = n2910 & ~n3775 ;
  assign n3778 = ~n774 & ~n3776 ;
  assign n3779 = ~n3777 & n3778 ;
  assign n3780 = ~n3774 & ~n3779 ;
  assign n3781 = ~n2726 & n3780 ;
  assign n3782 = ~\P1_IR_reg[4]/NET0131  & ~n3121 ;
  assign n3122 = \P1_IR_reg[31]/NET0131  & \P1_IR_reg[4]/NET0131  ;
  assign n3783 = ~n2667 & n3122 ;
  assign n3784 = ~n3782 & ~n3783 ;
  assign n3785 = n2726 & n3784 ;
  assign n3786 = ~n3781 & ~n3785 ;
  assign n3787 = \P1_reg2_reg[4]/NET0131  & n2851 ;
  assign n3788 = \P1_reg0_reg[4]/NET0131  & n2855 ;
  assign n3793 = ~n3787 & ~n3788 ;
  assign n3789 = \P1_reg1_reg[4]/NET0131  & n2853 ;
  assign n3790 = ~\P1_reg3_reg[3]/NET0131  & ~\P1_reg3_reg[4]/NET0131  ;
  assign n3791 = ~n2859 & ~n3790 ;
  assign n3792 = n2857 & n3791 ;
  assign n3794 = ~n3789 & ~n3792 ;
  assign n3795 = n3793 & n3794 ;
  assign n3796 = ~n3786 & n3795 ;
  assign n3113 = \P2_datao_reg[5]/NET0131  & n774 ;
  assign n3114 = ~n2771 & ~n2791 ;
  assign n3116 = ~n2788 & n3114 ;
  assign n3115 = n2788 & ~n3114 ;
  assign n3117 = ~n774 & ~n3115 ;
  assign n3118 = ~n3116 & n3117 ;
  assign n3119 = ~n3113 & ~n3118 ;
  assign n3120 = ~n2726 & ~n3119 ;
  assign n3123 = ~n3121 & ~n3122 ;
  assign n3124 = \P1_IR_reg[5]/NET0131  & ~n3123 ;
  assign n3125 = ~\P1_IR_reg[5]/NET0131  & n3123 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = n2726 & n3126 ;
  assign n3128 = ~n3120 & ~n3127 ;
  assign n3129 = \P1_reg2_reg[5]/NET0131  & n2851 ;
  assign n3130 = \P1_reg1_reg[5]/NET0131  & n2853 ;
  assign n3135 = ~n3129 & ~n3130 ;
  assign n3131 = \P1_reg0_reg[5]/NET0131  & n2855 ;
  assign n3132 = ~\P1_reg3_reg[5]/NET0131  & ~n2859 ;
  assign n3133 = ~n2860 & ~n3132 ;
  assign n3134 = n2857 & n3133 ;
  assign n3136 = ~n3131 & ~n3134 ;
  assign n3137 = n3135 & n3136 ;
  assign n3912 = ~n3128 & n3137 ;
  assign n3913 = ~n3796 & ~n3912 ;
  assign n4046 = n3911 & n3913 ;
  assign n4047 = ~n4045 & n4046 ;
  assign n3797 = n3786 & ~n3795 ;
  assign n3914 = n3128 & ~n3137 ;
  assign n3920 = ~n3797 & ~n3914 ;
  assign n4048 = ~n3912 & ~n3920 ;
  assign n4049 = n3911 & n4048 ;
  assign n3908 = ~n3568 & ~n3577 ;
  assign n3915 = ~n3737 & ~n3746 ;
  assign n3921 = ~n3908 & ~n3915 ;
  assign n4050 = ~n3909 & ~n3921 ;
  assign n4051 = ~n4049 & ~n4050 ;
  assign n4052 = ~n4047 & n4051 ;
  assign n3892 = n3813 & n3822 ;
  assign n3893 = ~n3891 & ~n3892 ;
  assign n4053 = n3890 & n3893 ;
  assign n4054 = ~n4052 & n4053 ;
  assign n4055 = n4040 & ~n4054 ;
  assign n4056 = n4035 & ~n4055 ;
  assign n4057 = n3886 & ~n4056 ;
  assign n4058 = n4034 & ~n4057 ;
  assign n4059 = n4033 & ~n4058 ;
  assign n4060 = n4027 & ~n4059 ;
  assign n4061 = n4026 & ~n4060 ;
  assign n3441 = ~\P2_datao_reg[30]/NET0131  & ~\si[30]_pad  ;
  assign n2960 = ~\P2_datao_reg[27]/NET0131  & ~\si[27]_pad  ;
  assign n2957 = ~\P2_datao_reg[28]/NET0131  & ~\si[28]_pad  ;
  assign n3383 = ~\P2_datao_reg[29]/NET0131  & ~\si[29]_pad  ;
  assign n3442 = ~n2957 & ~n3383 ;
  assign n3443 = ~n2960 & n3442 ;
  assign n3444 = ~n3441 & n3443 ;
  assign n2965 = ~\P2_datao_reg[26]/NET0131  & ~\si[26]_pad  ;
  assign n2967 = ~\P2_datao_reg[25]/NET0131  & ~\si[25]_pad  ;
  assign n2972 = ~\P2_datao_reg[24]/NET0131  & ~\si[24]_pad  ;
  assign n2973 = ~n2967 & ~n2972 ;
  assign n3418 = n2973 & ~n2975 ;
  assign n3419 = ~n2965 & n3418 ;
  assign n3445 = n3264 & n3419 ;
  assign n3446 = n3444 & n3445 ;
  assign n3447 = n2926 & n3446 ;
  assign n2961 = \P2_datao_reg[26]/NET0131  & \si[26]_pad  ;
  assign n2968 = \P2_datao_reg[25]/NET0131  & \si[25]_pad  ;
  assign n3387 = ~n2961 & ~n2968 ;
  assign n3388 = ~n2965 & ~n3387 ;
  assign n2969 = \P2_datao_reg[24]/NET0131  & \si[24]_pad  ;
  assign n3154 = ~n2969 & ~n2974 ;
  assign n3155 = ~n2972 & ~n3154 ;
  assign n3389 = ~n2965 & ~n2967 ;
  assign n3416 = n3155 & n3389 ;
  assign n3417 = ~n3388 & ~n3416 ;
  assign n3451 = n2933 & n3264 ;
  assign n3452 = n3263 & ~n3451 ;
  assign n3453 = n3419 & ~n3452 ;
  assign n3454 = n3417 & ~n3453 ;
  assign n3455 = n3444 & ~n3454 ;
  assign n3384 = \P2_datao_reg[29]/NET0131  & \si[29]_pad  ;
  assign n2958 = \P2_datao_reg[28]/NET0131  & \si[28]_pad  ;
  assign n2962 = \P2_datao_reg[27]/NET0131  & \si[27]_pad  ;
  assign n3386 = ~n2958 & ~n2962 ;
  assign n3448 = ~n3386 & n3442 ;
  assign n3449 = ~n3384 & ~n3448 ;
  assign n3450 = ~n3441 & ~n3449 ;
  assign n3456 = \P2_datao_reg[30]/NET0131  & \si[30]_pad  ;
  assign n3457 = ~n3450 & ~n3456 ;
  assign n3458 = ~n3455 & n3457 ;
  assign n3459 = ~n3447 & n3458 ;
  assign n3460 = ~\si[31]_pad  & ~n3459 ;
  assign n3461 = \si[31]_pad  & n3459 ;
  assign n3462 = ~n3460 & ~n3461 ;
  assign n3463 = ~n774 & ~n3462 ;
  assign n3464 = \P2_datao_reg[31]/NET0131  & n3463 ;
  assign n3465 = ~\P2_datao_reg[31]/NET0131  & ~n3463 ;
  assign n3466 = ~n3464 & ~n3465 ;
  assign n3467 = ~n2726 & n3466 ;
  assign n3023 = \P1_reg3_reg[23]/NET0131  & \P1_reg3_reg[24]/NET0131  ;
  assign n3024 = \P1_reg3_reg[25]/NET0131  & \P1_reg3_reg[26]/NET0131  ;
  assign n3025 = \P1_reg3_reg[27]/NET0131  & n3024 ;
  assign n3026 = n3023 & n3025 ;
  assign n3027 = n2882 & n3026 ;
  assign n3028 = \P1_reg3_reg[28]/NET0131  & n3027 ;
  assign n3405 = n2857 & n3028 ;
  assign n3468 = \P1_reg2_reg[31]/NET0131  & n2851 ;
  assign n3471 = ~n3405 & ~n3468 ;
  assign n3469 = \P1_reg0_reg[31]/NET0131  & n2855 ;
  assign n3470 = \P1_reg1_reg[31]/NET0131  & n2853 ;
  assign n3472 = ~n3469 & ~n3470 ;
  assign n3473 = n3471 & n3472 ;
  assign n3552 = ~n3467 & ~n3473 ;
  assign n3475 = \P2_datao_reg[30]/NET0131  & n774 ;
  assign n3476 = ~n3441 & ~n3456 ;
  assign n3487 = ~n2965 & n3443 ;
  assign n3484 = ~n2823 & n3418 ;
  assign n3489 = n2744 & n3484 ;
  assign n3490 = n3487 & n3489 ;
  assign n3491 = n2818 & n3490 ;
  assign n2970 = ~n2968 & ~n2969 ;
  assign n2971 = ~n2967 & ~n2970 ;
  assign n3479 = ~n2822 & ~n2974 ;
  assign n3480 = n3418 & ~n3479 ;
  assign n3481 = ~n2971 & ~n3480 ;
  assign n3482 = n2744 & ~n2757 ;
  assign n3483 = n2741 & ~n3482 ;
  assign n3485 = ~n3483 & n3484 ;
  assign n3486 = n3481 & ~n3485 ;
  assign n3488 = ~n3486 & n3487 ;
  assign n2963 = ~n2961 & ~n2962 ;
  assign n2964 = ~n2960 & ~n2963 ;
  assign n3477 = ~n2958 & ~n2964 ;
  assign n3478 = n3442 & ~n3477 ;
  assign n3492 = ~n3384 & ~n3478 ;
  assign n3493 = ~n3488 & n3492 ;
  assign n3494 = ~n3491 & n3493 ;
  assign n3496 = n3476 & ~n3494 ;
  assign n3495 = ~n3476 & n3494 ;
  assign n3497 = ~n774 & ~n3495 ;
  assign n3498 = ~n3496 & n3497 ;
  assign n3499 = ~n3475 & ~n3498 ;
  assign n3500 = ~n2726 & ~n3499 ;
  assign n3501 = \P1_reg2_reg[30]/NET0131  & n2851 ;
  assign n3504 = ~n3405 & ~n3501 ;
  assign n3502 = \P1_reg0_reg[30]/NET0131  & n2855 ;
  assign n3503 = \P1_reg1_reg[30]/NET0131  & n2853 ;
  assign n3505 = ~n3502 & ~n3503 ;
  assign n3506 = n3504 & n3505 ;
  assign n3553 = n3500 & n3506 ;
  assign n3554 = ~n3552 & ~n3553 ;
  assign n3382 = \P2_datao_reg[29]/NET0131  & n774 ;
  assign n3385 = ~n3383 & ~n3384 ;
  assign n2976 = ~n2823 & ~n2975 ;
  assign n3151 = ~n2972 & n2976 ;
  assign n3152 = ~n2728 & n3151 ;
  assign n3153 = ~n3150 & n3152 ;
  assign n2966 = ~n2960 & ~n2965 ;
  assign n3393 = n2966 & ~n2967 ;
  assign n3394 = n3153 & n3393 ;
  assign n3156 = ~n2729 & ~n2822 ;
  assign n3157 = n3151 & ~n3156 ;
  assign n3158 = ~n3155 & ~n3157 ;
  assign n3390 = ~n3158 & n3389 ;
  assign n3391 = ~n3388 & ~n3390 ;
  assign n3392 = ~n2960 & ~n3391 ;
  assign n3395 = n3386 & ~n3392 ;
  assign n3396 = ~n3394 & n3395 ;
  assign n3397 = ~n2957 & ~n3396 ;
  assign n3399 = n3385 & n3397 ;
  assign n3398 = ~n3385 & ~n3397 ;
  assign n3400 = ~n774 & ~n3398 ;
  assign n3401 = ~n3399 & n3400 ;
  assign n3402 = ~n3382 & ~n3401 ;
  assign n3403 = ~n2726 & ~n3402 ;
  assign n3404 = \P1_reg1_reg[29]/NET0131  & n2853 ;
  assign n3408 = ~n3404 & ~n3405 ;
  assign n3406 = \P1_reg0_reg[29]/NET0131  & n2855 ;
  assign n3407 = \P1_reg2_reg[29]/NET0131  & n2851 ;
  assign n3409 = ~n3406 & ~n3407 ;
  assign n3410 = n3408 & n3409 ;
  assign n3411 = n3403 & n3410 ;
  assign n2956 = \P2_datao_reg[28]/NET0131  & n774 ;
  assign n2959 = ~n2957 & ~n2958 ;
  assign n3008 = n2739 & n2976 ;
  assign n3009 = ~n3007 & n3008 ;
  assign n3010 = n2966 & n2973 ;
  assign n3011 = n3009 & n3010 ;
  assign n2977 = ~n2732 & ~n2822 ;
  assign n2978 = n2976 & ~n2977 ;
  assign n2979 = ~n2974 & ~n2978 ;
  assign n2980 = n2973 & ~n2979 ;
  assign n2981 = ~n2971 & ~n2980 ;
  assign n2982 = n2966 & ~n2981 ;
  assign n3012 = ~n2964 & ~n2982 ;
  assign n3013 = ~n3011 & n3012 ;
  assign n3015 = n2959 & ~n3013 ;
  assign n3014 = ~n2959 & n3013 ;
  assign n3016 = ~n774 & ~n3014 ;
  assign n3017 = ~n3015 & n3016 ;
  assign n3018 = ~n2956 & ~n3017 ;
  assign n3019 = ~n2726 & ~n3018 ;
  assign n3029 = ~\P1_reg3_reg[28]/NET0131  & ~n3027 ;
  assign n3030 = ~n3028 & ~n3029 ;
  assign n3031 = n2857 & n3030 ;
  assign n3022 = \P1_reg0_reg[28]/NET0131  & n2855 ;
  assign n3020 = \P1_reg2_reg[28]/NET0131  & n2851 ;
  assign n3021 = \P1_reg1_reg[28]/NET0131  & n2853 ;
  assign n3032 = ~n3020 & ~n3021 ;
  assign n3033 = ~n3022 & n3032 ;
  assign n3034 = ~n3031 & n3033 ;
  assign n4001 = n3019 & n3034 ;
  assign n4002 = ~n3411 & ~n4001 ;
  assign n4016 = n3554 & n4002 ;
  assign n3414 = \P2_datao_reg[27]/NET0131  & n774 ;
  assign n3415 = ~n2960 & ~n2962 ;
  assign n3420 = ~n3266 & n3419 ;
  assign n3421 = n3417 & ~n3420 ;
  assign n3423 = n3415 & ~n3421 ;
  assign n3422 = ~n3415 & n3421 ;
  assign n3424 = ~n774 & ~n3422 ;
  assign n3425 = ~n3423 & n3424 ;
  assign n3426 = ~n3414 & ~n3425 ;
  assign n3427 = ~n2726 & ~n3426 ;
  assign n3169 = n2882 & n3023 ;
  assign n3171 = \P1_reg3_reg[25]/NET0131  & n3169 ;
  assign n3431 = \P1_reg3_reg[26]/NET0131  & n3171 ;
  assign n3432 = ~\P1_reg3_reg[27]/NET0131  & ~n3431 ;
  assign n3433 = ~n3027 & ~n3432 ;
  assign n3434 = n2857 & n3433 ;
  assign n3430 = \P1_reg1_reg[27]/NET0131  & n2853 ;
  assign n3428 = \P1_reg0_reg[27]/NET0131  & n2855 ;
  assign n3429 = \P1_reg2_reg[27]/NET0131  & n2851 ;
  assign n3435 = ~n3428 & ~n3429 ;
  assign n3436 = ~n3430 & n3435 ;
  assign n3437 = ~n3434 & n3436 ;
  assign n3986 = n3427 & n3437 ;
  assign n3509 = \P2_datao_reg[26]/NET0131  & n774 ;
  assign n3510 = ~n2961 & ~n2965 ;
  assign n3511 = ~n2821 & n3484 ;
  assign n3512 = n3481 & ~n3511 ;
  assign n3514 = n3510 & ~n3512 ;
  assign n3513 = ~n3510 & n3512 ;
  assign n3515 = ~n774 & ~n3513 ;
  assign n3516 = ~n3514 & n3515 ;
  assign n3517 = ~n3509 & ~n3516 ;
  assign n3518 = ~n2726 & ~n3517 ;
  assign n3522 = ~\P1_reg3_reg[26]/NET0131  & ~n3171 ;
  assign n3523 = ~n3431 & ~n3522 ;
  assign n3524 = n2857 & n3523 ;
  assign n3521 = \P1_reg0_reg[26]/NET0131  & n2855 ;
  assign n3519 = \P1_reg2_reg[26]/NET0131  & n2851 ;
  assign n3520 = \P1_reg1_reg[26]/NET0131  & n2853 ;
  assign n3525 = ~n3519 & ~n3520 ;
  assign n3526 = ~n3521 & n3525 ;
  assign n3527 = ~n3524 & n3526 ;
  assign n3987 = n3518 & n3527 ;
  assign n3988 = ~n3986 & ~n3987 ;
  assign n3141 = \P2_datao_reg[25]/NET0131  & n774 ;
  assign n3142 = ~n2967 & ~n2968 ;
  assign n3159 = ~n3153 & n3158 ;
  assign n3161 = n3142 & ~n3159 ;
  assign n3160 = ~n3142 & n3159 ;
  assign n3162 = ~n774 & ~n3160 ;
  assign n3163 = ~n3161 & n3162 ;
  assign n3164 = ~n3141 & ~n3163 ;
  assign n3165 = ~n2726 & ~n3164 ;
  assign n3170 = ~\P1_reg3_reg[25]/NET0131  & ~n3169 ;
  assign n3172 = ~n3170 & ~n3171 ;
  assign n3173 = n2857 & n3172 ;
  assign n3168 = \P1_reg1_reg[25]/NET0131  & n2853 ;
  assign n3166 = \P1_reg0_reg[25]/NET0131  & n2855 ;
  assign n3167 = \P1_reg2_reg[25]/NET0131  & n2851 ;
  assign n3174 = ~n3166 & ~n3167 ;
  assign n3175 = ~n3168 & n3174 ;
  assign n3176 = ~n3173 & n3175 ;
  assign n3989 = n3165 & n3176 ;
  assign n3531 = \P2_datao_reg[24]/NET0131  & n774 ;
  assign n3532 = ~n2969 & ~n2972 ;
  assign n3533 = n2979 & ~n3009 ;
  assign n3535 = n3532 & ~n3533 ;
  assign n3534 = ~n3532 & n3533 ;
  assign n3536 = ~n774 & ~n3534 ;
  assign n3537 = ~n3535 & n3536 ;
  assign n3538 = ~n3531 & ~n3537 ;
  assign n3539 = ~n2726 & ~n3538 ;
  assign n3543 = ~\P1_reg3_reg[24]/NET0131  & ~n3277 ;
  assign n3544 = ~n3169 & ~n3543 ;
  assign n3545 = n2857 & n3544 ;
  assign n3542 = \P1_reg2_reg[24]/NET0131  & n2851 ;
  assign n3540 = \P1_reg1_reg[24]/NET0131  & n2853 ;
  assign n3541 = \P1_reg0_reg[24]/NET0131  & n2855 ;
  assign n3546 = ~n3540 & ~n3541 ;
  assign n3547 = ~n3542 & n3546 ;
  assign n3548 = ~n3545 & n3547 ;
  assign n3990 = n3539 & n3548 ;
  assign n3991 = ~n3989 & ~n3990 ;
  assign n4062 = n3988 & n3991 ;
  assign n4063 = n4016 & n4062 ;
  assign n4064 = ~n4061 & n4063 ;
  assign n3978 = ~n3518 & ~n3527 ;
  assign n3979 = ~n3427 & ~n3437 ;
  assign n3980 = ~n3978 & ~n3979 ;
  assign n3981 = ~n3165 & ~n3176 ;
  assign n3982 = ~n3539 & ~n3548 ;
  assign n3983 = ~n3981 & ~n3982 ;
  assign n4017 = ~n3983 & ~n3989 ;
  assign n4018 = ~n3987 & n4017 ;
  assign n4019 = n3980 & ~n4018 ;
  assign n4020 = ~n3986 & ~n4019 ;
  assign n4021 = n4016 & n4020 ;
  assign n3474 = n3467 & n3473 ;
  assign n3507 = ~n3500 & ~n3506 ;
  assign n3412 = ~n3403 & ~n3410 ;
  assign n3997 = ~n3019 & ~n3034 ;
  assign n3998 = ~n3412 & ~n3997 ;
  assign n4013 = ~n3411 & ~n3998 ;
  assign n4014 = ~n3507 & ~n4013 ;
  assign n4015 = n3554 & ~n4014 ;
  assign n4065 = ~n3474 & ~n4015 ;
  assign n4066 = ~n4021 & n4065 ;
  assign n4067 = ~n4064 & n4066 ;
  assign n4068 = ~\P1_B_reg/NET0131  & n4067 ;
  assign n2700 = ~\P1_IR_reg[20]/NET0131  & ~n2684 ;
  assign n2701 = \P1_IR_reg[20]/NET0131  & n2684 ;
  assign n2702 = ~n2700 & ~n2701 ;
  assign n3861 = ~\P1_IR_reg[19]/NET0131  & ~\P1_IR_reg[22]/NET0131  ;
  assign n3862 = n2685 & n3861 ;
  assign n3863 = \P1_IR_reg[31]/NET0131  & ~n3862 ;
  assign n3864 = ~n2719 & ~n3863 ;
  assign n3865 = \P1_IR_reg[23]/NET0131  & ~n3864 ;
  assign n3866 = ~\P1_IR_reg[23]/NET0131  & n3864 ;
  assign n3867 = ~n3865 & ~n3866 ;
  assign n4069 = n2702 & n3867 ;
  assign n2686 = \P1_IR_reg[31]/NET0131  & ~n2685 ;
  assign n2687 = ~n2684 & ~n2686 ;
  assign n2688 = \P1_IR_reg[22]/NET0131  & ~n2687 ;
  assign n2689 = ~\P1_IR_reg[22]/NET0131  & n2687 ;
  assign n2690 = ~n2688 & ~n2689 ;
  assign n2696 = ~n2692 & ~n2695 ;
  assign n2697 = \P1_IR_reg[21]/NET0131  & ~n2696 ;
  assign n2698 = ~\P1_IR_reg[21]/NET0131  & n2696 ;
  assign n2699 = ~n2697 & ~n2698 ;
  assign n4070 = ~n2690 & ~n2699 ;
  assign n4071 = n4069 & n4070 ;
  assign n4072 = ~n4068 & n4071 ;
  assign n2888 = ~n2830 & n2887 ;
  assign n2889 = n2830 & ~n2887 ;
  assign n2890 = ~n2888 & ~n2889 ;
  assign n3624 = ~n3614 & n3623 ;
  assign n3625 = n3614 & ~n3623 ;
  assign n3626 = ~n3624 & ~n3625 ;
  assign n3082 = n3072 & ~n3081 ;
  assign n3083 = ~n3072 & n3081 ;
  assign n3084 = ~n3082 & ~n3083 ;
  assign n3138 = ~n3128 & ~n3137 ;
  assign n3139 = n3128 & n3137 ;
  assign n3140 = ~n3138 & ~n3139 ;
  assign n3330 = n3320 & ~n3329 ;
  assign n3331 = ~n3320 & n3329 ;
  assign n3332 = ~n3330 & ~n3331 ;
  assign n3826 = ~n3140 & ~n3332 ;
  assign n3381 = ~n3379 & ~n3380 ;
  assign n3578 = ~n3568 & n3577 ;
  assign n3579 = n3568 & ~n3577 ;
  assign n3580 = ~n3578 & ~n3579 ;
  assign n3827 = n3381 & ~n3580 ;
  assign n3833 = n3826 & n3827 ;
  assign n3256 = ~n3246 & n3255 ;
  assign n3257 = n3246 & ~n3255 ;
  assign n3258 = ~n3256 & ~n3257 ;
  assign n3355 = ~n3345 & n3354 ;
  assign n3356 = n3345 & ~n3354 ;
  assign n3357 = ~n3355 & ~n3356 ;
  assign n3834 = ~n3258 & ~n3357 ;
  assign n3835 = n3833 & n3834 ;
  assign n3839 = ~n3084 & n3835 ;
  assign n3840 = ~n3626 & n3839 ;
  assign n3844 = ~n2890 & n3840 ;
  assign n2953 = ~n2942 & n2952 ;
  assign n2954 = n2942 & ~n2952 ;
  assign n2955 = ~n2953 & ~n2954 ;
  assign n3598 = ~n3588 & n3597 ;
  assign n3599 = n3588 & ~n3597 ;
  assign n3600 = ~n3598 & ~n3599 ;
  assign n3845 = ~n2955 & ~n3600 ;
  assign n3846 = n3844 & n3845 ;
  assign n3177 = ~n3165 & n3176 ;
  assign n3178 = n3165 & ~n3176 ;
  assign n3179 = ~n3177 & ~n3178 ;
  assign n3110 = ~n3100 & n3109 ;
  assign n3111 = n3100 & ~n3109 ;
  assign n3112 = ~n3110 & ~n3111 ;
  assign n3823 = ~n3813 & n3822 ;
  assign n3824 = n3813 & ~n3822 ;
  assign n3825 = ~n3823 & ~n3824 ;
  assign n3773 = ~n3771 & ~n3772 ;
  assign n3798 = ~n3796 & ~n3797 ;
  assign n3830 = n3773 & n3798 ;
  assign n3831 = ~n3825 & n3830 ;
  assign n3678 = ~n3668 & n3677 ;
  assign n3679 = n3668 & ~n3677 ;
  assign n3680 = ~n3678 & ~n3679 ;
  assign n3696 = ~n3687 & n3694 ;
  assign n3697 = ~n3695 & ~n3696 ;
  assign n3828 = ~n3680 & n3697 ;
  assign n3721 = ~n3719 & ~n3720 ;
  assign n3747 = ~n3737 & n3746 ;
  assign n3748 = n3737 & ~n3746 ;
  assign n3749 = ~n3747 & ~n3748 ;
  assign n3829 = n3721 & ~n3749 ;
  assign n3832 = n3828 & n3829 ;
  assign n3836 = n3831 & n3832 ;
  assign n3230 = ~n3219 & n3229 ;
  assign n3231 = n3219 & ~n3229 ;
  assign n3232 = ~n3230 & ~n3231 ;
  assign n3651 = ~n3641 & n3650 ;
  assign n3652 = n3641 & ~n3650 ;
  assign n3653 = ~n3651 & ~n3652 ;
  assign n3837 = ~n3232 & ~n3653 ;
  assign n3838 = n3836 & n3837 ;
  assign n3841 = ~n3112 & n3838 ;
  assign n3204 = n3194 & ~n3203 ;
  assign n3205 = ~n3194 & n3203 ;
  assign n3206 = ~n3204 & ~n3205 ;
  assign n3304 = ~n3294 & n3303 ;
  assign n3305 = n3294 & ~n3303 ;
  assign n3306 = ~n3304 & ~n3305 ;
  assign n3842 = ~n3206 & ~n3306 ;
  assign n3843 = n3841 & n3842 ;
  assign n3847 = ~n3179 & n3843 ;
  assign n3850 = n3846 & n3847 ;
  assign n3528 = n3518 & ~n3527 ;
  assign n3529 = ~n3518 & n3527 ;
  assign n3530 = ~n3528 & ~n3529 ;
  assign n3549 = ~n3539 & n3548 ;
  assign n3550 = n3539 & ~n3548 ;
  assign n3551 = ~n3549 & ~n3550 ;
  assign n3851 = ~n3530 & ~n3551 ;
  assign n3852 = n3850 & n3851 ;
  assign n3035 = ~n3019 & n3034 ;
  assign n3036 = n3019 & ~n3034 ;
  assign n3037 = ~n3035 & ~n3036 ;
  assign n3284 = n3273 & ~n3283 ;
  assign n3285 = ~n3273 & n3283 ;
  assign n3286 = ~n3284 & ~n3285 ;
  assign n3508 = ~n3474 & ~n3507 ;
  assign n3848 = ~n3286 & n3508 ;
  assign n3849 = n3554 & n3848 ;
  assign n3853 = ~n3037 & n3849 ;
  assign n3413 = ~n3411 & ~n3412 ;
  assign n3438 = n3427 & ~n3437 ;
  assign n3439 = ~n3427 & n3437 ;
  assign n3440 = ~n3438 & ~n3439 ;
  assign n3854 = n3413 & ~n3440 ;
  assign n3855 = n3853 & n3854 ;
  assign n3856 = n3852 & n3855 ;
  assign n3858 = n2702 & n3856 ;
  assign n3857 = ~n2702 & ~n3856 ;
  assign n3859 = n2699 & ~n3857 ;
  assign n3860 = ~n3858 & n3859 ;
  assign n3868 = ~n2699 & n2702 ;
  assign n3869 = \P1_B_reg/NET0131  & n3867 ;
  assign n3870 = ~n3868 & n3869 ;
  assign n3871 = ~n3860 & ~n3870 ;
  assign n3872 = ~n2690 & ~n3871 ;
  assign n3896 = ~n3894 & ~n3895 ;
  assign n3897 = ~n3893 & n3896 ;
  assign n3898 = n3890 & ~n3897 ;
  assign n3899 = ~n3887 & ~n3898 ;
  assign n3902 = ~n3876 & ~n3883 ;
  assign n3903 = ~n3901 & n3902 ;
  assign n3904 = n3875 & ~n3903 ;
  assign n3905 = ~n3882 & ~n3904 ;
  assign n3906 = ~n3899 & ~n3905 ;
  assign n3907 = n3886 & ~n3906 ;
  assign n3916 = ~n3914 & ~n3915 ;
  assign n3917 = ~n3913 & n3916 ;
  assign n3918 = n3911 & ~n3917 ;
  assign n3919 = ~n3908 & ~n3918 ;
  assign n3923 = ~n3772 & ~n3922 ;
  assign n3925 = n3696 & ~n3720 ;
  assign n3926 = ~n3719 & n3924 ;
  assign n3927 = ~n3925 & n3926 ;
  assign n3928 = ~n3923 & ~n3927 ;
  assign n3929 = n3920 & n3921 ;
  assign n3930 = ~n3928 & n3929 ;
  assign n3931 = ~n3919 & ~n3930 ;
  assign n3935 = ~n3895 & n3933 ;
  assign n3936 = ~n3882 & n3935 ;
  assign n3934 = ~n3878 & ~n3887 ;
  assign n3937 = n3902 & n3934 ;
  assign n3938 = n3936 & n3937 ;
  assign n3939 = ~n3931 & n3938 ;
  assign n3940 = ~n3907 & ~n3939 ;
  assign n3947 = ~n3945 & ~n3946 ;
  assign n3948 = ~n3944 & n3947 ;
  assign n3949 = n3943 & n3948 ;
  assign n3953 = ~n3951 & ~n3952 ;
  assign n3954 = ~n3950 & n3953 ;
  assign n3955 = n3949 & n3954 ;
  assign n3956 = ~n3940 & n3955 ;
  assign n3963 = ~n3942 & ~n3944 ;
  assign n3964 = ~n3962 & n3963 ;
  assign n3965 = n3959 & ~n3964 ;
  assign n3966 = ~n3941 & ~n3965 ;
  assign n3973 = n3953 & ~n3972 ;
  assign n3974 = n3969 & ~n3973 ;
  assign n3975 = n3949 & ~n3974 ;
  assign n3976 = ~n3966 & ~n3975 ;
  assign n3977 = ~n3956 & n3976 ;
  assign n3984 = n3980 & n3983 ;
  assign n3985 = ~n3977 & n3984 ;
  assign n3992 = ~n3978 & ~n3981 ;
  assign n3993 = ~n3991 & n3992 ;
  assign n3994 = n3988 & ~n3993 ;
  assign n3995 = ~n3979 & ~n3994 ;
  assign n3996 = ~n3985 & ~n3995 ;
  assign n3999 = n3508 & n3998 ;
  assign n4000 = ~n3996 & n3999 ;
  assign n4003 = ~n3412 & ~n3507 ;
  assign n4004 = ~n4002 & n4003 ;
  assign n4005 = n3554 & ~n4004 ;
  assign n4006 = ~n3474 & ~n4005 ;
  assign n4007 = ~n4000 & ~n4006 ;
  assign n4008 = ~\P1_B_reg/NET0131  & n4007 ;
  assign n4009 = ~n2699 & ~n2702 ;
  assign n4010 = n3867 & n4009 ;
  assign n4011 = n2690 & n4010 ;
  assign n4012 = ~n4008 & n4011 ;
  assign n4122 = ~n3872 & ~n4012 ;
  assign n4125 = ~n4072 & n4122 ;
  assign n4074 = n2702 & ~n4007 ;
  assign n4073 = ~n2702 & n4007 ;
  assign n4075 = n2690 & ~n2699 ;
  assign n4076 = ~n3867 & n4075 ;
  assign n4077 = ~n4073 & n4076 ;
  assign n4078 = ~n4074 & n4077 ;
  assign n4080 = n4027 & n4034 ;
  assign n4081 = n4035 & ~n4040 ;
  assign n4082 = n3886 & ~n4081 ;
  assign n4083 = n4052 & n4082 ;
  assign n4084 = ~n3907 & ~n4083 ;
  assign n4085 = n4080 & n4084 ;
  assign n4086 = n4027 & ~n4033 ;
  assign n4087 = n4026 & ~n4086 ;
  assign n4088 = ~n4085 & n4087 ;
  assign n4089 = n4062 & ~n4088 ;
  assign n4090 = ~n4020 & ~n4089 ;
  assign n4091 = ~n3473 & ~n3506 ;
  assign n4092 = n3500 & ~n4091 ;
  assign n4093 = ~n3552 & ~n4092 ;
  assign n4094 = n4002 & n4093 ;
  assign n4095 = ~n4090 & n4094 ;
  assign n4096 = n4013 & n4093 ;
  assign n4097 = ~n3473 & ~n3507 ;
  assign n4098 = n3467 & ~n4097 ;
  assign n4099 = ~n4096 & ~n4098 ;
  assign n4100 = ~n4095 & n4099 ;
  assign n4102 = ~n2702 & ~n4100 ;
  assign n4101 = n2702 & n4100 ;
  assign n4079 = n2690 & n2699 ;
  assign n4103 = ~n3867 & n4079 ;
  assign n4104 = ~n4101 & n4103 ;
  assign n4105 = ~n4102 & n4104 ;
  assign n4126 = ~n4078 & ~n4105 ;
  assign n4127 = n4125 & n4126 ;
  assign n4117 = ~n2699 & n4007 ;
  assign n4116 = n2699 & ~n4100 ;
  assign n4118 = ~\P1_B_reg/NET0131  & ~n4116 ;
  assign n4119 = ~n4117 & n4118 ;
  assign n4120 = n2690 & n4069 ;
  assign n4121 = ~n4119 & n4120 ;
  assign n4114 = ~n2690 & n4009 ;
  assign n4115 = n4067 & n4114 ;
  assign n4106 = ~\P1_B_reg/NET0131  & ~n4100 ;
  assign n4107 = ~n2702 & n3867 ;
  assign n4108 = n4079 & n4107 ;
  assign n4109 = ~n4106 & n4108 ;
  assign n4110 = ~n2690 & ~n3867 ;
  assign n4111 = ~n2699 & n4110 ;
  assign n4112 = n2702 & n4111 ;
  assign n4113 = ~n4067 & n4112 ;
  assign n4123 = ~n4109 & ~n4113 ;
  assign n4124 = ~n4115 & n4123 ;
  assign n4128 = ~n4121 & n4124 ;
  assign n4129 = n4127 & n4128 ;
  assign n4130 = \P1_state_reg[0]/NET0131  & n3867 ;
  assign n4131 = ~n4129 & n4130 ;
  assign n4132 = \P1_B_reg/NET0131  & ~n4130 ;
  assign n4133 = ~n4131 & ~n4132 ;
  assign n4134 = \P3_reg2_reg[27]/NET0131  & n2145 ;
  assign n4135 = \P3_reg2_reg[27]/NET0131  & ~n2408 ;
  assign n4136 = n2408 & ~n2617 ;
  assign n4137 = ~n4135 & ~n4136 ;
  assign n4138 = n2425 & ~n4137 ;
  assign n4139 = n2408 & ~n2575 ;
  assign n4140 = ~n4135 & ~n4139 ;
  assign n4141 = n737 & ~n4140 ;
  assign n4144 = n1436 & n2441 ;
  assign n4142 = \P3_reg2_reg[27]/NET0131  & ~n2429 ;
  assign n4143 = ~n1441 & n2283 ;
  assign n4152 = ~n4142 & ~n4143 ;
  assign n4153 = ~n4144 & n4152 ;
  assign n4154 = ~n4141 & n4153 ;
  assign n4155 = ~n4138 & n4154 ;
  assign n4145 = \P3_reg2_reg[27]/NET0131  & ~n2427 ;
  assign n4146 = n2427 & ~n2566 ;
  assign n4147 = ~n4145 & ~n4146 ;
  assign n4148 = n714 & ~n4147 ;
  assign n4149 = n2427 & ~n2617 ;
  assign n4150 = ~n4145 & ~n4149 ;
  assign n4151 = ~n2518 & ~n4150 ;
  assign n4156 = ~n4148 & ~n4151 ;
  assign n4157 = n4155 & n4156 ;
  assign n4158 = n2147 & ~n4157 ;
  assign n4159 = ~n4134 & ~n4158 ;
  assign n4160 = \P1_state_reg[0]/NET0131  & ~n4159 ;
  assign n4161 = \P3_reg2_reg[27]/NET0131  & ~n2143 ;
  assign n4162 = ~n4160 & ~n4161 ;
  assign n4163 = ~\P2_IR_reg[0]/NET0131  & ~\P2_IR_reg[1]/NET0131  ;
  assign n4164 = ~\P2_IR_reg[2]/NET0131  & n4163 ;
  assign n4165 = ~\P2_IR_reg[3]/NET0131  & n4164 ;
  assign n4166 = ~\P2_IR_reg[4]/NET0131  & n4165 ;
  assign n4167 = ~\P2_IR_reg[5]/NET0131  & n4166 ;
  assign n4168 = ~\P2_IR_reg[6]/NET0131  & ~\P2_IR_reg[7]/NET0131  ;
  assign n4169 = ~\P2_IR_reg[8]/NET0131  & n4168 ;
  assign n4170 = n4167 & n4169 ;
  assign n4171 = ~\P2_IR_reg[10]/NET0131  & ~\P2_IR_reg[11]/NET0131  ;
  assign n4172 = ~\P2_IR_reg[12]/NET0131  & ~\P2_IR_reg[9]/NET0131  ;
  assign n4173 = n4171 & n4172 ;
  assign n4174 = n4170 & n4173 ;
  assign n4175 = ~\P2_IR_reg[16]/NET0131  & ~\P2_IR_reg[17]/NET0131  ;
  assign n4176 = ~\P2_IR_reg[18]/NET0131  & n4175 ;
  assign n4177 = ~\P2_IR_reg[19]/NET0131  & n4176 ;
  assign n4178 = ~\P2_IR_reg[13]/NET0131  & ~\P2_IR_reg[14]/NET0131  ;
  assign n4179 = ~\P2_IR_reg[15]/NET0131  & n4178 ;
  assign n4180 = ~\P2_IR_reg[20]/NET0131  & n4179 ;
  assign n4181 = n4177 & n4180 ;
  assign n4182 = n4174 & n4181 ;
  assign n4183 = \P2_IR_reg[31]/NET0131  & ~n4182 ;
  assign n4184 = ~\P2_IR_reg[21]/NET0131  & ~\P2_IR_reg[22]/NET0131  ;
  assign n4185 = ~\P2_IR_reg[23]/NET0131  & n4184 ;
  assign n4186 = \P2_IR_reg[31]/NET0131  & ~n4185 ;
  assign n4187 = ~n4183 & ~n4186 ;
  assign n4188 = \P2_IR_reg[24]/NET0131  & ~n4187 ;
  assign n4189 = ~\P2_IR_reg[24]/NET0131  & n4187 ;
  assign n4190 = ~n4188 & ~n4189 ;
  assign n4191 = \P2_B_reg/NET0131  & ~n4190 ;
  assign n4192 = ~\P2_IR_reg[24]/NET0131  & n4185 ;
  assign n4193 = n4182 & n4192 ;
  assign n4194 = \P2_IR_reg[31]/NET0131  & ~n4193 ;
  assign n4195 = \P2_IR_reg[25]/NET0131  & ~n4194 ;
  assign n4196 = ~\P2_IR_reg[25]/NET0131  & n4194 ;
  assign n4197 = ~n4195 & ~n4196 ;
  assign n4198 = n4191 & n4197 ;
  assign n4199 = ~\P2_d_reg[0]/NET0131  & ~n4198 ;
  assign n4200 = ~\P2_IR_reg[25]/NET0131  & n4192 ;
  assign n4201 = n4182 & n4200 ;
  assign n4202 = \P2_IR_reg[31]/NET0131  & ~n4201 ;
  assign n4203 = \P2_IR_reg[26]/NET0131  & ~n4202 ;
  assign n4204 = ~\P2_IR_reg[26]/NET0131  & n4202 ;
  assign n4205 = ~n4203 & ~n4204 ;
  assign n4206 = ~n4199 & ~n4205 ;
  assign n4208 = \P2_B_reg/NET0131  & ~n4205 ;
  assign n4207 = ~n4197 & ~n4205 ;
  assign n4209 = n4190 & ~n4207 ;
  assign n4210 = ~n4208 & n4209 ;
  assign n4211 = ~n4206 & ~n4210 ;
  assign n4212 = n4197 & n4205 ;
  assign n4213 = ~\P2_B_reg/NET0131  & n4190 ;
  assign n4214 = ~n4191 & ~n4213 ;
  assign n4215 = n4197 & ~n4214 ;
  assign n4216 = ~\P2_d_reg[1]/NET0131  & ~n4205 ;
  assign n4217 = ~n4215 & n4216 ;
  assign n4218 = ~n4212 & ~n4217 ;
  assign n4219 = n4211 & n4218 ;
  assign n4220 = \P2_reg2_reg[29]/NET0131  & ~n4219 ;
  assign n4221 = ~\P2_IR_reg[26]/NET0131  & n4201 ;
  assign n4222 = \P2_IR_reg[31]/NET0131  & ~n4221 ;
  assign n4223 = ~\P2_IR_reg[27]/NET0131  & ~n4222 ;
  assign n4224 = \P2_IR_reg[27]/NET0131  & n4222 ;
  assign n4225 = ~n4223 & ~n4224 ;
  assign n4226 = ~\P2_IR_reg[26]/NET0131  & ~\P2_IR_reg[27]/NET0131  ;
  assign n4227 = \P2_IR_reg[31]/NET0131  & ~n4226 ;
  assign n4228 = ~n4202 & ~n4227 ;
  assign n4229 = \P2_IR_reg[28]/NET0131  & ~n4228 ;
  assign n4230 = ~\P2_IR_reg[28]/NET0131  & n4228 ;
  assign n4231 = ~n4229 & ~n4230 ;
  assign n4232 = ~n4225 & ~n4231 ;
  assign n4233 = \P1_datao_reg[29]/NET0131  & ~n774 ;
  assign n4234 = \P1_datao_reg[29]/NET0131  & \si[29]_pad  ;
  assign n4235 = ~\P1_datao_reg[29]/NET0131  & ~\si[29]_pad  ;
  assign n4236 = ~n4234 & ~n4235 ;
  assign n4237 = ~\P1_datao_reg[28]/NET0131  & ~\si[28]_pad  ;
  assign n4238 = ~\P1_datao_reg[27]/NET0131  & ~\si[27]_pad  ;
  assign n4239 = ~\P1_datao_reg[26]/NET0131  & ~\si[26]_pad  ;
  assign n4240 = ~\P1_datao_reg[25]/NET0131  & ~\si[25]_pad  ;
  assign n4241 = ~n4239 & ~n4240 ;
  assign n4242 = ~n4238 & n4241 ;
  assign n4243 = ~\P1_datao_reg[12]/NET0131  & ~\si[12]_pad  ;
  assign n4244 = \P1_datao_reg[12]/NET0131  & \si[12]_pad  ;
  assign n4245 = \P1_datao_reg[11]/NET0131  & \si[11]_pad  ;
  assign n4246 = ~n4244 & ~n4245 ;
  assign n4247 = ~\P1_datao_reg[11]/NET0131  & ~\si[11]_pad  ;
  assign n4248 = ~\P1_datao_reg[10]/NET0131  & ~\si[10]_pad  ;
  assign n4249 = \P1_datao_reg[10]/NET0131  & \si[10]_pad  ;
  assign n4250 = \P1_datao_reg[9]/NET0131  & \si[9]_pad  ;
  assign n4251 = ~n4249 & ~n4250 ;
  assign n4252 = ~n4248 & ~n4251 ;
  assign n4253 = ~n4247 & n4252 ;
  assign n4254 = n4246 & ~n4253 ;
  assign n4255 = ~n4243 & ~n4254 ;
  assign n4256 = \P1_datao_reg[4]/NET0131  & \si[4]_pad  ;
  assign n4257 = \P1_datao_reg[3]/NET0131  & \si[3]_pad  ;
  assign n4258 = ~\P1_datao_reg[2]/NET0131  & ~\si[2]_pad  ;
  assign n4259 = \P1_datao_reg[2]/NET0131  & \si[2]_pad  ;
  assign n4260 = ~\P1_datao_reg[1]/NET0131  & ~\si[1]_pad  ;
  assign n4261 = \P1_datao_reg[1]/NET0131  & \si[1]_pad  ;
  assign n4262 = \P1_datao_reg[0]/NET0131  & \si[0]_pad  ;
  assign n4263 = ~n4261 & ~n4262 ;
  assign n4264 = ~n4260 & ~n4263 ;
  assign n4265 = ~n4259 & ~n4264 ;
  assign n4266 = ~n4258 & ~n4265 ;
  assign n4267 = ~n4257 & ~n4266 ;
  assign n4268 = ~\P1_datao_reg[3]/NET0131  & ~\si[3]_pad  ;
  assign n4269 = ~\P1_datao_reg[4]/NET0131  & ~\si[4]_pad  ;
  assign n4270 = ~n4268 & ~n4269 ;
  assign n4271 = ~n4267 & n4270 ;
  assign n4272 = ~n4256 & ~n4271 ;
  assign n4273 = ~\P1_datao_reg[6]/NET0131  & ~\si[6]_pad  ;
  assign n4274 = ~\P1_datao_reg[5]/NET0131  & ~\si[5]_pad  ;
  assign n4275 = ~n4273 & ~n4274 ;
  assign n4276 = ~\P1_datao_reg[7]/NET0131  & ~\si[7]_pad  ;
  assign n4277 = ~\P1_datao_reg[8]/NET0131  & ~\si[8]_pad  ;
  assign n4278 = ~n4276 & ~n4277 ;
  assign n4279 = n4275 & n4278 ;
  assign n4280 = ~n4272 & n4279 ;
  assign n4281 = \P1_datao_reg[8]/NET0131  & \si[8]_pad  ;
  assign n4282 = \P1_datao_reg[6]/NET0131  & \si[6]_pad  ;
  assign n4283 = \P1_datao_reg[5]/NET0131  & \si[5]_pad  ;
  assign n4284 = ~n4282 & ~n4283 ;
  assign n4285 = ~n4273 & ~n4284 ;
  assign n4286 = \P1_datao_reg[7]/NET0131  & \si[7]_pad  ;
  assign n4287 = ~n4285 & ~n4286 ;
  assign n4288 = n4278 & ~n4287 ;
  assign n4289 = ~n4281 & ~n4288 ;
  assign n4290 = ~n4280 & n4289 ;
  assign n4291 = ~\P1_datao_reg[9]/NET0131  & ~\si[9]_pad  ;
  assign n4292 = ~n4248 & ~n4291 ;
  assign n4293 = ~n4247 & n4292 ;
  assign n4294 = ~n4243 & n4293 ;
  assign n4295 = ~n4290 & n4294 ;
  assign n4296 = ~n4255 & ~n4295 ;
  assign n4297 = ~\P1_datao_reg[13]/NET0131  & ~\si[13]_pad  ;
  assign n4298 = ~\P1_datao_reg[16]/NET0131  & ~\si[16]_pad  ;
  assign n4299 = ~\P1_datao_reg[15]/NET0131  & ~\si[15]_pad  ;
  assign n4300 = ~\P1_datao_reg[14]/NET0131  & ~\si[14]_pad  ;
  assign n4301 = ~n4299 & ~n4300 ;
  assign n4302 = ~n4298 & n4301 ;
  assign n4303 = ~n4297 & n4302 ;
  assign n4304 = ~n4296 & n4303 ;
  assign n4305 = \P1_datao_reg[15]/NET0131  & \si[15]_pad  ;
  assign n4306 = \P1_datao_reg[16]/NET0131  & \si[16]_pad  ;
  assign n4307 = ~n4305 & ~n4306 ;
  assign n4308 = ~n4298 & ~n4307 ;
  assign n4309 = \P1_datao_reg[13]/NET0131  & \si[13]_pad  ;
  assign n4310 = \P1_datao_reg[14]/NET0131  & \si[14]_pad  ;
  assign n4311 = ~n4309 & ~n4310 ;
  assign n4312 = n4302 & ~n4311 ;
  assign n4313 = ~n4308 & ~n4312 ;
  assign n4314 = ~n4304 & n4313 ;
  assign n4315 = ~\P1_datao_reg[19]/NET0131  & ~\si[19]_pad  ;
  assign n4316 = ~\P1_datao_reg[20]/NET0131  & ~\si[20]_pad  ;
  assign n4317 = ~n4315 & ~n4316 ;
  assign n4318 = ~\P1_datao_reg[18]/NET0131  & ~\si[18]_pad  ;
  assign n4319 = ~\P1_datao_reg[17]/NET0131  & ~\si[17]_pad  ;
  assign n4320 = ~n4318 & ~n4319 ;
  assign n4321 = n4317 & n4320 ;
  assign n4322 = ~n4314 & n4321 ;
  assign n4323 = \P1_datao_reg[17]/NET0131  & \si[17]_pad  ;
  assign n4324 = \P1_datao_reg[18]/NET0131  & \si[18]_pad  ;
  assign n4325 = ~n4323 & ~n4324 ;
  assign n4326 = ~n4318 & ~n4325 ;
  assign n4327 = n4317 & n4326 ;
  assign n4328 = \P1_datao_reg[19]/NET0131  & \si[19]_pad  ;
  assign n4329 = \P1_datao_reg[20]/NET0131  & \si[20]_pad  ;
  assign n4330 = ~n4328 & ~n4329 ;
  assign n4331 = ~n4316 & ~n4330 ;
  assign n4332 = ~n4327 & ~n4331 ;
  assign n4333 = ~n4322 & n4332 ;
  assign n4334 = ~\P1_datao_reg[23]/NET0131  & ~\si[23]_pad  ;
  assign n4335 = ~\P1_datao_reg[24]/NET0131  & ~\si[24]_pad  ;
  assign n4336 = ~n4334 & ~n4335 ;
  assign n4337 = ~\P1_datao_reg[22]/NET0131  & ~\si[22]_pad  ;
  assign n4338 = ~\P1_datao_reg[21]/NET0131  & ~\si[21]_pad  ;
  assign n4339 = ~n4337 & ~n4338 ;
  assign n4340 = n4336 & n4339 ;
  assign n4341 = ~n4333 & n4340 ;
  assign n4342 = n4242 & n4341 ;
  assign n4343 = \P1_datao_reg[27]/NET0131  & \si[27]_pad  ;
  assign n4344 = \P1_datao_reg[28]/NET0131  & \si[28]_pad  ;
  assign n4345 = ~n4343 & ~n4344 ;
  assign n4346 = \P1_datao_reg[25]/NET0131  & \si[25]_pad  ;
  assign n4347 = \P1_datao_reg[26]/NET0131  & \si[26]_pad  ;
  assign n4348 = ~n4346 & ~n4347 ;
  assign n4349 = ~n4239 & ~n4348 ;
  assign n4350 = \P1_datao_reg[22]/NET0131  & \si[22]_pad  ;
  assign n4351 = \P1_datao_reg[21]/NET0131  & \si[21]_pad  ;
  assign n4352 = ~n4350 & ~n4351 ;
  assign n4353 = ~n4337 & ~n4352 ;
  assign n4354 = n4336 & n4353 ;
  assign n4355 = \P1_datao_reg[23]/NET0131  & \si[23]_pad  ;
  assign n4356 = \P1_datao_reg[24]/NET0131  & \si[24]_pad  ;
  assign n4357 = ~n4355 & ~n4356 ;
  assign n4358 = ~n4335 & ~n4357 ;
  assign n4359 = ~n4354 & ~n4358 ;
  assign n4360 = n4241 & ~n4359 ;
  assign n4361 = ~n4349 & ~n4360 ;
  assign n4362 = ~n4238 & ~n4361 ;
  assign n4363 = n4345 & ~n4362 ;
  assign n4364 = ~n4342 & n4363 ;
  assign n4365 = ~n4237 & ~n4364 ;
  assign n4367 = n4236 & n4365 ;
  assign n4366 = ~n4236 & ~n4365 ;
  assign n4368 = n774 & ~n4366 ;
  assign n4369 = ~n4367 & n4368 ;
  assign n4370 = ~n4233 & ~n4369 ;
  assign n4371 = ~n4232 & ~n4370 ;
  assign n4372 = ~\P2_IR_reg[28]/NET0131  & ~\P2_IR_reg[29]/NET0131  ;
  assign n4373 = n4226 & n4372 ;
  assign n4374 = \P2_IR_reg[31]/NET0131  & ~n4373 ;
  assign n4375 = ~n4202 & ~n4374 ;
  assign n4376 = \P2_IR_reg[30]/NET0131  & ~n4375 ;
  assign n4377 = ~\P2_IR_reg[30]/NET0131  & n4375 ;
  assign n4378 = ~n4376 & ~n4377 ;
  assign n4379 = ~\P2_IR_reg[25]/NET0131  & ~\P2_IR_reg[28]/NET0131  ;
  assign n4380 = n4226 & n4379 ;
  assign n4381 = \P2_IR_reg[31]/NET0131  & ~n4380 ;
  assign n4382 = ~n4194 & ~n4381 ;
  assign n4383 = \P2_IR_reg[29]/NET0131  & ~n4382 ;
  assign n4384 = ~\P2_IR_reg[29]/NET0131  & n4382 ;
  assign n4385 = ~n4383 & ~n4384 ;
  assign n4386 = n4378 & n4385 ;
  assign n4387 = \P2_reg3_reg[3]/NET0131  & \P2_reg3_reg[4]/NET0131  ;
  assign n4388 = \P2_reg3_reg[5]/NET0131  & n4387 ;
  assign n4389 = \P2_reg3_reg[6]/NET0131  & n4388 ;
  assign n4390 = \P2_reg3_reg[7]/NET0131  & n4389 ;
  assign n4391 = \P2_reg3_reg[8]/NET0131  & n4390 ;
  assign n4392 = \P2_reg3_reg[9]/NET0131  & n4391 ;
  assign n4393 = \P2_reg3_reg[10]/NET0131  & n4392 ;
  assign n4394 = \P2_reg3_reg[11]/NET0131  & n4393 ;
  assign n4395 = \P2_reg3_reg[12]/NET0131  & \P2_reg3_reg[13]/NET0131  ;
  assign n4396 = n4394 & n4395 ;
  assign n4397 = \P2_reg3_reg[14]/NET0131  & \P2_reg3_reg[15]/NET0131  ;
  assign n4398 = \P2_reg3_reg[16]/NET0131  & n4397 ;
  assign n4399 = n4396 & n4398 ;
  assign n4400 = \P2_reg3_reg[17]/NET0131  & \P2_reg3_reg[18]/NET0131  ;
  assign n4401 = \P2_reg3_reg[19]/NET0131  & n4400 ;
  assign n4402 = n4399 & n4401 ;
  assign n4403 = \P2_reg3_reg[20]/NET0131  & n4402 ;
  assign n4404 = \P2_reg3_reg[21]/NET0131  & \P2_reg3_reg[22]/NET0131  ;
  assign n4405 = \P2_reg3_reg[23]/NET0131  & \P2_reg3_reg[24]/NET0131  ;
  assign n4406 = n4404 & n4405 ;
  assign n4407 = n4403 & n4406 ;
  assign n4408 = \P2_reg3_reg[25]/NET0131  & \P2_reg3_reg[26]/NET0131  ;
  assign n4409 = \P2_reg3_reg[27]/NET0131  & \P2_reg3_reg[28]/NET0131  ;
  assign n4410 = n4408 & n4409 ;
  assign n4411 = n4407 & n4410 ;
  assign n4412 = n4386 & n4411 ;
  assign n4413 = n4378 & ~n4385 ;
  assign n4414 = \P2_reg2_reg[29]/NET0131  & n4413 ;
  assign n4419 = ~n4412 & ~n4414 ;
  assign n4415 = ~n4378 & n4385 ;
  assign n4416 = \P2_reg1_reg[29]/NET0131  & n4415 ;
  assign n4417 = ~n4378 & ~n4385 ;
  assign n4418 = \P2_reg0_reg[29]/NET0131  & n4417 ;
  assign n4420 = ~n4416 & ~n4418 ;
  assign n4421 = n4419 & n4420 ;
  assign n4422 = n4371 & n4421 ;
  assign n4423 = ~n4371 & ~n4421 ;
  assign n4424 = ~n4422 & ~n4423 ;
  assign n4718 = \P2_reg0_reg[19]/NET0131  & n4417 ;
  assign n4719 = \P2_reg3_reg[17]/NET0131  & n4399 ;
  assign n4720 = \P2_reg3_reg[18]/NET0131  & n4719 ;
  assign n4721 = ~\P2_reg3_reg[19]/NET0131  & ~n4720 ;
  assign n4722 = ~n4402 & ~n4721 ;
  assign n4723 = n4386 & n4722 ;
  assign n4726 = ~n4718 & ~n4723 ;
  assign n4724 = \P2_reg2_reg[19]/NET0131  & n4413 ;
  assign n4725 = \P2_reg1_reg[19]/NET0131  & n4415 ;
  assign n4727 = ~n4724 & ~n4725 ;
  assign n4728 = n4726 & n4727 ;
  assign n4729 = n4174 & n4179 ;
  assign n4730 = \P2_IR_reg[31]/NET0131  & ~n4729 ;
  assign n4731 = \P2_IR_reg[31]/NET0131  & ~n4176 ;
  assign n4732 = ~n4730 & ~n4731 ;
  assign n4733 = \P2_IR_reg[19]/NET0131  & ~n4732 ;
  assign n4734 = ~\P2_IR_reg[19]/NET0131  & n4732 ;
  assign n4735 = ~n4733 & ~n4734 ;
  assign n4736 = n4232 & ~n4735 ;
  assign n4737 = \P1_datao_reg[19]/NET0131  & ~n774 ;
  assign n4447 = ~n4243 & ~n4297 ;
  assign n4506 = ~n4247 & n4447 ;
  assign n4433 = n4270 & n4275 ;
  assign n4510 = n4266 & n4433 ;
  assign n4511 = ~n4256 & ~n4257 ;
  assign n4512 = ~n4269 & n4275 ;
  assign n4513 = ~n4511 & n4512 ;
  assign n4514 = ~n4285 & ~n4513 ;
  assign n4515 = ~n4510 & n4514 ;
  assign n4516 = n4278 & n4292 ;
  assign n4517 = ~n4515 & n4516 ;
  assign n4507 = ~n4281 & ~n4286 ;
  assign n4508 = ~n4277 & n4292 ;
  assign n4509 = ~n4507 & n4508 ;
  assign n4518 = ~n4252 & ~n4509 ;
  assign n4519 = ~n4517 & n4518 ;
  assign n4520 = n4506 & ~n4519 ;
  assign n4521 = ~n4246 & n4447 ;
  assign n4522 = n4311 & ~n4521 ;
  assign n4523 = ~n4520 & n4522 ;
  assign n4524 = n4302 & n4320 ;
  assign n4525 = ~n4523 & n4524 ;
  assign n4505 = n4308 & n4320 ;
  assign n4526 = ~n4326 & ~n4505 ;
  assign n4527 = ~n4525 & n4526 ;
  assign n4738 = ~n4315 & ~n4328 ;
  assign n4740 = n4527 & ~n4738 ;
  assign n4739 = ~n4527 & n4738 ;
  assign n4741 = n774 & ~n4739 ;
  assign n4742 = ~n4740 & n4741 ;
  assign n4743 = ~n4737 & ~n4742 ;
  assign n4744 = ~n4232 & n4743 ;
  assign n4745 = ~n4736 & ~n4744 ;
  assign n4746 = n4728 & ~n4745 ;
  assign n4747 = \P1_datao_reg[20]/NET0131  & ~n774 ;
  assign n4434 = ~n4267 & n4433 ;
  assign n4435 = n4256 & n4275 ;
  assign n4436 = n4287 & ~n4435 ;
  assign n4437 = ~n4434 & n4436 ;
  assign n4438 = n4278 & n4293 ;
  assign n4439 = ~n4437 & n4438 ;
  assign n4440 = ~n4247 & ~n4248 ;
  assign n4441 = ~n4250 & ~n4281 ;
  assign n4442 = ~n4291 & ~n4441 ;
  assign n4443 = ~n4249 & ~n4442 ;
  assign n4444 = n4440 & ~n4443 ;
  assign n4445 = ~n4245 & ~n4444 ;
  assign n4446 = ~n4439 & n4445 ;
  assign n4448 = n4301 & n4447 ;
  assign n4449 = ~n4446 & n4448 ;
  assign n4450 = ~n4244 & ~n4309 ;
  assign n4451 = ~n4297 & ~n4450 ;
  assign n4452 = n4301 & n4451 ;
  assign n4453 = ~n4305 & ~n4310 ;
  assign n4454 = ~n4299 & ~n4453 ;
  assign n4455 = ~n4452 & ~n4454 ;
  assign n4456 = ~n4449 & n4455 ;
  assign n4457 = ~n4315 & ~n4318 ;
  assign n4458 = ~n4298 & ~n4319 ;
  assign n4459 = n4457 & n4458 ;
  assign n4460 = ~n4456 & n4459 ;
  assign n4461 = ~n4306 & ~n4323 ;
  assign n4462 = ~n4319 & ~n4461 ;
  assign n4463 = n4457 & n4462 ;
  assign n4464 = ~n4324 & ~n4328 ;
  assign n4465 = ~n4315 & ~n4464 ;
  assign n4466 = ~n4463 & ~n4465 ;
  assign n4467 = ~n4460 & n4466 ;
  assign n4748 = ~n4316 & ~n4329 ;
  assign n4750 = n4467 & ~n4748 ;
  assign n4749 = ~n4467 & n4748 ;
  assign n4751 = n774 & ~n4749 ;
  assign n4752 = ~n4750 & n4751 ;
  assign n4753 = ~n4747 & ~n4752 ;
  assign n4754 = ~n4232 & ~n4753 ;
  assign n4755 = \P2_reg1_reg[20]/NET0131  & n4415 ;
  assign n4756 = ~\P2_reg3_reg[20]/NET0131  & ~n4402 ;
  assign n4757 = ~n4403 & ~n4756 ;
  assign n4758 = n4386 & n4757 ;
  assign n4761 = ~n4755 & ~n4758 ;
  assign n4759 = \P2_reg2_reg[20]/NET0131  & n4413 ;
  assign n4760 = \P2_reg0_reg[20]/NET0131  & n4417 ;
  assign n4762 = ~n4759 & ~n4760 ;
  assign n4763 = n4761 & n4762 ;
  assign n4764 = ~n4754 & n4763 ;
  assign n4765 = ~n4746 & ~n4764 ;
  assign n4766 = \P2_reg0_reg[17]/NET0131  & n4417 ;
  assign n4767 = \P2_reg1_reg[17]/NET0131  & n4415 ;
  assign n4772 = ~n4766 & ~n4767 ;
  assign n4768 = \P2_reg2_reg[17]/NET0131  & n4413 ;
  assign n4769 = ~\P2_reg3_reg[17]/NET0131  & ~n4399 ;
  assign n4770 = ~n4719 & ~n4769 ;
  assign n4771 = n4386 & n4770 ;
  assign n4773 = ~n4768 & ~n4771 ;
  assign n4774 = n4772 & n4773 ;
  assign n4775 = \P2_IR_reg[16]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n4776 = ~n4730 & ~n4775 ;
  assign n4777 = \P2_IR_reg[17]/NET0131  & ~n4776 ;
  assign n4778 = ~\P2_IR_reg[17]/NET0131  & n4776 ;
  assign n4779 = ~n4777 & ~n4778 ;
  assign n4780 = n4232 & ~n4779 ;
  assign n4781 = \P1_datao_reg[17]/NET0131  & ~n774 ;
  assign n4782 = ~n4319 & ~n4323 ;
  assign n4784 = ~n4314 & n4782 ;
  assign n4783 = n4314 & ~n4782 ;
  assign n4785 = n774 & ~n4783 ;
  assign n4786 = ~n4784 & n4785 ;
  assign n4787 = ~n4781 & ~n4786 ;
  assign n4788 = ~n4232 & n4787 ;
  assign n4789 = ~n4780 & ~n4788 ;
  assign n4790 = n4774 & ~n4789 ;
  assign n4791 = \P2_reg0_reg[18]/NET0131  & n4417 ;
  assign n4792 = ~\P2_reg3_reg[18]/NET0131  & ~n4719 ;
  assign n4793 = ~n4720 & ~n4792 ;
  assign n4794 = n4386 & n4793 ;
  assign n4797 = ~n4791 & ~n4794 ;
  assign n4795 = \P2_reg2_reg[18]/NET0131  & n4413 ;
  assign n4796 = \P2_reg1_reg[18]/NET0131  & n4415 ;
  assign n4798 = ~n4795 & ~n4796 ;
  assign n4799 = n4797 & n4798 ;
  assign n4800 = \P2_IR_reg[31]/NET0131  & ~n4175 ;
  assign n4801 = ~n4730 & ~n4800 ;
  assign n4802 = \P2_IR_reg[18]/NET0131  & ~n4801 ;
  assign n4803 = ~\P2_IR_reg[18]/NET0131  & n4801 ;
  assign n4804 = ~n4802 & ~n4803 ;
  assign n4805 = n4232 & ~n4804 ;
  assign n4806 = \P1_datao_reg[18]/NET0131  & ~n774 ;
  assign n4559 = ~n4256 & ~n4283 ;
  assign n4560 = ~n4271 & n4559 ;
  assign n4561 = n4279 & ~n4291 ;
  assign n4562 = ~n4560 & n4561 ;
  assign n4563 = ~n4282 & ~n4286 ;
  assign n4564 = n4278 & ~n4291 ;
  assign n4565 = ~n4563 & n4564 ;
  assign n4566 = ~n4442 & ~n4565 ;
  assign n4567 = ~n4562 & n4566 ;
  assign n4568 = n4440 & n4447 ;
  assign n4569 = ~n4567 & n4568 ;
  assign n4557 = ~n4245 & ~n4249 ;
  assign n4558 = n4506 & ~n4557 ;
  assign n4570 = ~n4451 & ~n4558 ;
  assign n4571 = ~n4569 & n4570 ;
  assign n4572 = n4302 & ~n4319 ;
  assign n4573 = ~n4571 & n4572 ;
  assign n4556 = n4454 & n4458 ;
  assign n4574 = ~n4462 & ~n4556 ;
  assign n4575 = ~n4573 & n4574 ;
  assign n4807 = ~n4318 & ~n4324 ;
  assign n4809 = n4575 & ~n4807 ;
  assign n4808 = ~n4575 & n4807 ;
  assign n4810 = n774 & ~n4808 ;
  assign n4811 = ~n4809 & n4810 ;
  assign n4812 = ~n4806 & ~n4811 ;
  assign n4813 = ~n4232 & n4812 ;
  assign n4814 = ~n4805 & ~n4813 ;
  assign n4815 = n4799 & ~n4814 ;
  assign n4816 = ~n4790 & ~n4815 ;
  assign n4817 = n4765 & n4816 ;
  assign n4818 = \P2_reg2_reg[14]/NET0131  & n4413 ;
  assign n4819 = \P2_reg3_reg[14]/NET0131  & n4396 ;
  assign n4820 = ~\P2_reg3_reg[14]/NET0131  & ~n4396 ;
  assign n4821 = ~n4819 & ~n4820 ;
  assign n4822 = n4386 & n4821 ;
  assign n4825 = ~n4818 & ~n4822 ;
  assign n4823 = \P2_reg1_reg[14]/NET0131  & n4415 ;
  assign n4824 = \P2_reg0_reg[14]/NET0131  & n4417 ;
  assign n4826 = ~n4823 & ~n4824 ;
  assign n4827 = n4825 & n4826 ;
  assign n4828 = \P2_IR_reg[31]/NET0131  & ~n4174 ;
  assign n4829 = \P2_IR_reg[13]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n4830 = ~n4828 & ~n4829 ;
  assign n4831 = \P2_IR_reg[14]/NET0131  & ~n4830 ;
  assign n4832 = ~\P2_IR_reg[14]/NET0131  & n4830 ;
  assign n4833 = ~n4831 & ~n4832 ;
  assign n4834 = n4232 & ~n4833 ;
  assign n4835 = \P1_datao_reg[14]/NET0131  & ~n774 ;
  assign n4836 = ~n4300 & ~n4310 ;
  assign n4838 = ~n4571 & n4836 ;
  assign n4837 = n4571 & ~n4836 ;
  assign n4839 = n774 & ~n4837 ;
  assign n4840 = ~n4838 & n4839 ;
  assign n4841 = ~n4835 & ~n4840 ;
  assign n4842 = ~n4232 & n4841 ;
  assign n4843 = ~n4834 & ~n4842 ;
  assign n4844 = n4827 & ~n4843 ;
  assign n4845 = \P2_reg2_reg[13]/NET0131  & n4413 ;
  assign n4846 = \P2_reg1_reg[13]/NET0131  & n4415 ;
  assign n4852 = ~n4845 & ~n4846 ;
  assign n4847 = \P2_reg3_reg[12]/NET0131  & n4394 ;
  assign n4848 = ~\P2_reg3_reg[13]/NET0131  & ~n4847 ;
  assign n4849 = ~n4396 & ~n4848 ;
  assign n4850 = n4386 & n4849 ;
  assign n4851 = \P2_reg0_reg[13]/NET0131  & n4417 ;
  assign n4853 = ~n4850 & ~n4851 ;
  assign n4854 = n4852 & n4853 ;
  assign n4855 = \P2_IR_reg[13]/NET0131  & ~n4828 ;
  assign n4856 = ~\P2_IR_reg[13]/NET0131  & n4828 ;
  assign n4857 = ~n4855 & ~n4856 ;
  assign n4858 = n4232 & n4857 ;
  assign n4859 = \P1_datao_reg[13]/NET0131  & ~n774 ;
  assign n4860 = ~n4297 & ~n4309 ;
  assign n4862 = ~n4296 & n4860 ;
  assign n4861 = n4296 & ~n4860 ;
  assign n4863 = n774 & ~n4861 ;
  assign n4864 = ~n4862 & n4863 ;
  assign n4865 = ~n4859 & ~n4864 ;
  assign n4866 = ~n4232 & n4865 ;
  assign n4867 = ~n4858 & ~n4866 ;
  assign n4868 = n4854 & ~n4867 ;
  assign n4869 = ~n4844 & ~n4868 ;
  assign n4870 = \P2_reg0_reg[16]/NET0131  & n4417 ;
  assign n4871 = \P2_reg2_reg[16]/NET0131  & n4413 ;
  assign n4877 = ~n4870 & ~n4871 ;
  assign n4872 = \P2_reg1_reg[16]/NET0131  & n4415 ;
  assign n4873 = \P2_reg3_reg[15]/NET0131  & n4819 ;
  assign n4874 = ~\P2_reg3_reg[16]/NET0131  & ~n4873 ;
  assign n4875 = ~n4399 & ~n4874 ;
  assign n4876 = n4386 & n4875 ;
  assign n4878 = ~n4872 & ~n4876 ;
  assign n4879 = n4877 & n4878 ;
  assign n4880 = \P2_IR_reg[16]/NET0131  & ~n4730 ;
  assign n4881 = ~\P2_IR_reg[16]/NET0131  & n4730 ;
  assign n4882 = ~n4880 & ~n4881 ;
  assign n4883 = n4232 & n4882 ;
  assign n4884 = \P1_datao_reg[16]/NET0131  & ~n774 ;
  assign n4885 = ~n4298 & ~n4306 ;
  assign n4887 = ~n4456 & n4885 ;
  assign n4886 = n4456 & ~n4885 ;
  assign n4888 = n774 & ~n4886 ;
  assign n4889 = ~n4887 & n4888 ;
  assign n4890 = ~n4884 & ~n4889 ;
  assign n4891 = ~n4232 & n4890 ;
  assign n4892 = ~n4883 & ~n4891 ;
  assign n4893 = n4879 & ~n4892 ;
  assign n4894 = \P2_reg1_reg[15]/NET0131  & n4415 ;
  assign n4895 = \P2_reg2_reg[15]/NET0131  & n4413 ;
  assign n4900 = ~n4894 & ~n4895 ;
  assign n4896 = \P2_reg0_reg[15]/NET0131  & n4417 ;
  assign n4897 = ~\P2_reg3_reg[15]/NET0131  & ~n4819 ;
  assign n4898 = ~n4873 & ~n4897 ;
  assign n4899 = n4386 & n4898 ;
  assign n4901 = ~n4896 & ~n4899 ;
  assign n4902 = n4900 & n4901 ;
  assign n4903 = \P2_IR_reg[31]/NET0131  & ~n4178 ;
  assign n4904 = ~n4828 & ~n4903 ;
  assign n4905 = \P2_IR_reg[15]/NET0131  & ~n4904 ;
  assign n4906 = ~\P2_IR_reg[15]/NET0131  & n4904 ;
  assign n4907 = ~n4905 & ~n4906 ;
  assign n4908 = n4232 & ~n4907 ;
  assign n4909 = \P1_datao_reg[15]/NET0131  & ~n774 ;
  assign n4910 = ~n4300 & ~n4523 ;
  assign n4911 = ~n4299 & ~n4305 ;
  assign n4913 = n4910 & n4911 ;
  assign n4912 = ~n4910 & ~n4911 ;
  assign n4914 = n774 & ~n4912 ;
  assign n4915 = ~n4913 & n4914 ;
  assign n4916 = ~n4909 & ~n4915 ;
  assign n4917 = ~n4232 & n4916 ;
  assign n4918 = ~n4908 & ~n4917 ;
  assign n4919 = n4902 & ~n4918 ;
  assign n4920 = ~n4893 & ~n4919 ;
  assign n4921 = n4869 & n4920 ;
  assign n4922 = n4817 & n4921 ;
  assign n4923 = \P2_reg0_reg[11]/NET0131  & n4417 ;
  assign n4924 = \P2_reg2_reg[11]/NET0131  & n4413 ;
  assign n4929 = ~n4923 & ~n4924 ;
  assign n4925 = ~\P2_reg3_reg[11]/NET0131  & ~n4393 ;
  assign n4926 = ~n4394 & ~n4925 ;
  assign n4927 = n4386 & n4926 ;
  assign n4928 = \P2_reg1_reg[11]/NET0131  & n4415 ;
  assign n4930 = ~n4927 & ~n4928 ;
  assign n4931 = n4929 & n4930 ;
  assign n4932 = ~\P2_IR_reg[9]/NET0131  & n4170 ;
  assign n4933 = \P2_IR_reg[31]/NET0131  & ~n4932 ;
  assign n4934 = \P2_IR_reg[10]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n4935 = ~n4933 & ~n4934 ;
  assign n4936 = \P2_IR_reg[11]/NET0131  & ~n4935 ;
  assign n4937 = ~\P2_IR_reg[11]/NET0131  & n4935 ;
  assign n4938 = ~n4936 & ~n4937 ;
  assign n4939 = n4232 & ~n4938 ;
  assign n4940 = \P1_datao_reg[11]/NET0131  & ~n774 ;
  assign n4941 = ~n4245 & ~n4247 ;
  assign n4943 = ~n4519 & n4941 ;
  assign n4942 = n4519 & ~n4941 ;
  assign n4944 = n774 & ~n4942 ;
  assign n4945 = ~n4943 & n4944 ;
  assign n4946 = ~n4940 & ~n4945 ;
  assign n4947 = ~n4232 & n4946 ;
  assign n4948 = ~n4939 & ~n4947 ;
  assign n4949 = n4931 & ~n4948 ;
  assign n4950 = \P2_reg0_reg[12]/NET0131  & n4417 ;
  assign n4951 = ~\P2_reg3_reg[12]/NET0131  & ~n4394 ;
  assign n4952 = ~n4847 & ~n4951 ;
  assign n4953 = n4386 & n4952 ;
  assign n4956 = ~n4950 & ~n4953 ;
  assign n4954 = \P2_reg2_reg[12]/NET0131  & n4413 ;
  assign n4955 = \P2_reg1_reg[12]/NET0131  & n4415 ;
  assign n4957 = ~n4954 & ~n4955 ;
  assign n4958 = n4956 & n4957 ;
  assign n4959 = \P2_IR_reg[31]/NET0131  & ~n4171 ;
  assign n4960 = ~n4933 & ~n4959 ;
  assign n4961 = \P2_IR_reg[12]/NET0131  & ~n4960 ;
  assign n4962 = ~\P2_IR_reg[12]/NET0131  & n4960 ;
  assign n4963 = ~n4961 & ~n4962 ;
  assign n4964 = n4232 & ~n4963 ;
  assign n4965 = \P1_datao_reg[12]/NET0131  & ~n774 ;
  assign n4966 = ~n4243 & ~n4244 ;
  assign n4968 = ~n4446 & n4966 ;
  assign n4967 = n4446 & ~n4966 ;
  assign n4969 = n774 & ~n4967 ;
  assign n4970 = ~n4968 & n4969 ;
  assign n4971 = ~n4965 & ~n4970 ;
  assign n4972 = ~n4232 & n4971 ;
  assign n4973 = ~n4964 & ~n4972 ;
  assign n4974 = n4958 & ~n4973 ;
  assign n4975 = ~n4949 & ~n4974 ;
  assign n4976 = \P2_reg1_reg[10]/NET0131  & n4415 ;
  assign n4977 = ~\P2_reg3_reg[10]/NET0131  & ~n4392 ;
  assign n4978 = ~n4393 & ~n4977 ;
  assign n4979 = n4386 & n4978 ;
  assign n4982 = ~n4976 & ~n4979 ;
  assign n4980 = \P2_reg0_reg[10]/NET0131  & n4417 ;
  assign n4981 = \P2_reg2_reg[10]/NET0131  & n4413 ;
  assign n4983 = ~n4980 & ~n4981 ;
  assign n4984 = n4982 & n4983 ;
  assign n4985 = \P1_datao_reg[10]/NET0131  & ~n774 ;
  assign n4986 = ~n4248 & ~n4249 ;
  assign n4988 = ~n4567 & n4986 ;
  assign n4987 = n4567 & ~n4986 ;
  assign n4989 = n774 & ~n4987 ;
  assign n4990 = ~n4988 & n4989 ;
  assign n4991 = ~n4985 & ~n4990 ;
  assign n4992 = ~n4232 & ~n4991 ;
  assign n4993 = \P2_IR_reg[10]/NET0131  & ~n4933 ;
  assign n4994 = ~\P2_IR_reg[10]/NET0131  & n4933 ;
  assign n4995 = ~n4993 & ~n4994 ;
  assign n4996 = n4232 & ~n4995 ;
  assign n4997 = ~n4992 & ~n4996 ;
  assign n4998 = ~n4984 & ~n4997 ;
  assign n4999 = n4984 & n4997 ;
  assign n5000 = \P2_reg0_reg[9]/NET0131  & n4417 ;
  assign n5001 = \P2_reg1_reg[9]/NET0131  & n4415 ;
  assign n5006 = ~n5000 & ~n5001 ;
  assign n5002 = ~\P2_reg3_reg[9]/NET0131  & ~n4391 ;
  assign n5003 = ~n4392 & ~n5002 ;
  assign n5004 = n4386 & n5003 ;
  assign n5005 = \P2_reg2_reg[9]/NET0131  & n4413 ;
  assign n5007 = ~n5004 & ~n5005 ;
  assign n5008 = n5006 & n5007 ;
  assign n5009 = \P2_IR_reg[31]/NET0131  & ~n4170 ;
  assign n5010 = \P2_IR_reg[9]/NET0131  & n5009 ;
  assign n5011 = ~\P2_IR_reg[9]/NET0131  & ~n5009 ;
  assign n5012 = ~n5010 & ~n5011 ;
  assign n5013 = n4232 & ~n5012 ;
  assign n5014 = \P1_datao_reg[9]/NET0131  & ~n774 ;
  assign n5015 = ~n4250 & ~n4291 ;
  assign n5017 = ~n4290 & n5015 ;
  assign n5016 = n4290 & ~n5015 ;
  assign n5018 = n774 & ~n5016 ;
  assign n5019 = ~n5017 & n5018 ;
  assign n5020 = ~n5014 & ~n5019 ;
  assign n5021 = ~n4232 & n5020 ;
  assign n5022 = ~n5013 & ~n5021 ;
  assign n5023 = ~n5008 & n5022 ;
  assign n5024 = ~n4999 & n5023 ;
  assign n5025 = ~n4998 & ~n5024 ;
  assign n5026 = n4975 & ~n5025 ;
  assign n5027 = ~n4958 & n4973 ;
  assign n5028 = ~n4931 & n4948 ;
  assign n5029 = ~n5027 & ~n5028 ;
  assign n5030 = ~n4974 & ~n5029 ;
  assign n5031 = ~n5026 & ~n5030 ;
  assign n5032 = ~\P2_reg3_reg[8]/NET0131  & ~n4390 ;
  assign n5033 = ~n4391 & ~n5032 ;
  assign n5034 = n4386 & n5033 ;
  assign n5035 = \P2_reg0_reg[8]/NET0131  & n4417 ;
  assign n5038 = ~n5034 & ~n5035 ;
  assign n5036 = \P2_reg2_reg[8]/NET0131  & n4413 ;
  assign n5037 = \P2_reg1_reg[8]/NET0131  & n4415 ;
  assign n5039 = ~n5036 & ~n5037 ;
  assign n5040 = n5038 & n5039 ;
  assign n5041 = \P1_datao_reg[8]/NET0131  & ~n774 ;
  assign n5042 = ~n4276 & ~n4437 ;
  assign n5043 = ~n4277 & ~n4281 ;
  assign n5045 = n5042 & n5043 ;
  assign n5044 = ~n5042 & ~n5043 ;
  assign n5046 = n774 & ~n5044 ;
  assign n5047 = ~n5045 & n5046 ;
  assign n5048 = ~n5041 & ~n5047 ;
  assign n5049 = ~n4232 & ~n5048 ;
  assign n5050 = ~\P2_IR_reg[6]/NET0131  & n4167 ;
  assign n5051 = \P2_IR_reg[31]/NET0131  & ~n5050 ;
  assign n5052 = \P2_IR_reg[31]/NET0131  & \P2_IR_reg[7]/NET0131  ;
  assign n5053 = ~n5051 & ~n5052 ;
  assign n5054 = \P2_IR_reg[8]/NET0131  & ~n5053 ;
  assign n5055 = ~\P2_IR_reg[8]/NET0131  & n5053 ;
  assign n5056 = ~n5054 & ~n5055 ;
  assign n5057 = n4232 & n5056 ;
  assign n5058 = ~n5049 & ~n5057 ;
  assign n5059 = n5040 & n5058 ;
  assign n5060 = \P2_reg2_reg[7]/NET0131  & n4413 ;
  assign n5061 = \P2_reg1_reg[7]/NET0131  & n4415 ;
  assign n5066 = ~n5060 & ~n5061 ;
  assign n5062 = ~\P2_reg3_reg[7]/NET0131  & ~n4389 ;
  assign n5063 = ~n4390 & ~n5062 ;
  assign n5064 = n4386 & n5063 ;
  assign n5065 = \P2_reg0_reg[7]/NET0131  & n4417 ;
  assign n5067 = ~n5064 & ~n5065 ;
  assign n5068 = n5066 & n5067 ;
  assign n5069 = \P1_datao_reg[7]/NET0131  & ~n774 ;
  assign n5070 = ~n4276 & ~n4286 ;
  assign n5072 = ~n4515 & n5070 ;
  assign n5071 = n4515 & ~n5070 ;
  assign n5073 = n774 & ~n5071 ;
  assign n5074 = ~n5072 & n5073 ;
  assign n5075 = ~n5069 & ~n5074 ;
  assign n5076 = ~n4232 & ~n5075 ;
  assign n5077 = ~\P2_IR_reg[7]/NET0131  & ~n5051 ;
  assign n5078 = ~n5050 & n5052 ;
  assign n5079 = ~n5077 & ~n5078 ;
  assign n5080 = n4232 & n5079 ;
  assign n5081 = ~n5076 & ~n5080 ;
  assign n5082 = n5068 & n5081 ;
  assign n5083 = ~n5059 & ~n5082 ;
  assign n5133 = \P2_reg1_reg[2]/NET0131  & n4415 ;
  assign n5134 = \P2_reg3_reg[2]/NET0131  & n4386 ;
  assign n5137 = ~n5133 & ~n5134 ;
  assign n5135 = \P2_reg0_reg[2]/NET0131  & n4417 ;
  assign n5136 = \P2_reg2_reg[2]/NET0131  & n4413 ;
  assign n5138 = ~n5135 & ~n5136 ;
  assign n5139 = n5137 & n5138 ;
  assign n5140 = \P1_datao_reg[2]/NET0131  & ~n774 ;
  assign n5141 = ~n4258 & ~n4259 ;
  assign n5143 = n4264 & n5141 ;
  assign n5142 = ~n4264 & ~n5141 ;
  assign n5144 = n774 & ~n5142 ;
  assign n5145 = ~n5143 & n5144 ;
  assign n5146 = ~n5140 & ~n5145 ;
  assign n5147 = ~n4232 & ~n5146 ;
  assign n5148 = \P2_IR_reg[31]/NET0131  & ~n4163 ;
  assign n5149 = \P2_IR_reg[2]/NET0131  & n5148 ;
  assign n5150 = ~\P2_IR_reg[2]/NET0131  & ~n5148 ;
  assign n5151 = ~n5149 & ~n5150 ;
  assign n5152 = n4232 & n5151 ;
  assign n5153 = ~n5147 & ~n5152 ;
  assign n5154 = ~n5139 & ~n5153 ;
  assign n5155 = \P2_reg0_reg[1]/NET0131  & n4417 ;
  assign n5156 = \P2_reg3_reg[1]/NET0131  & n4386 ;
  assign n5159 = ~n5155 & ~n5156 ;
  assign n5157 = \P2_reg1_reg[1]/NET0131  & n4415 ;
  assign n5158 = \P2_reg2_reg[1]/NET0131  & n4413 ;
  assign n5160 = ~n5157 & ~n5158 ;
  assign n5161 = n5159 & n5160 ;
  assign n5162 = \P2_IR_reg[0]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n5163 = \P2_IR_reg[1]/NET0131  & ~n5162 ;
  assign n5164 = ~\P2_IR_reg[1]/NET0131  & n5162 ;
  assign n5165 = ~n5163 & ~n5164 ;
  assign n5166 = n4232 & ~n5165 ;
  assign n5167 = ~\P1_datao_reg[1]/NET0131  & ~n774 ;
  assign n5168 = ~n4260 & ~n4261 ;
  assign n5170 = ~n4262 & n5168 ;
  assign n5169 = n4262 & ~n5168 ;
  assign n5171 = n774 & ~n5169 ;
  assign n5172 = ~n5170 & n5171 ;
  assign n5173 = ~n5167 & ~n5172 ;
  assign n5174 = ~n4232 & n5173 ;
  assign n5175 = ~n5166 & ~n5174 ;
  assign n5176 = ~n5161 & ~n5175 ;
  assign n5177 = n5161 & n5175 ;
  assign n5178 = \P2_reg3_reg[0]/NET0131  & n4386 ;
  assign n5179 = \P2_reg2_reg[0]/NET0131  & n4413 ;
  assign n5182 = ~n5178 & ~n5179 ;
  assign n5180 = \P2_reg0_reg[0]/NET0131  & n4417 ;
  assign n5181 = \P2_reg1_reg[0]/NET0131  & n4415 ;
  assign n5183 = ~n5180 & ~n5181 ;
  assign n5184 = n5182 & n5183 ;
  assign n5185 = ~\P1_datao_reg[0]/NET0131  & ~n1900 ;
  assign n5186 = n774 & n4262 ;
  assign n5187 = ~n5185 & ~n5186 ;
  assign n5188 = ~n4232 & n5187 ;
  assign n5189 = \P2_IR_reg[0]/NET0131  & n4232 ;
  assign n5190 = ~n5188 & ~n5189 ;
  assign n5191 = ~n5184 & ~n5190 ;
  assign n5192 = ~n5177 & n5191 ;
  assign n5193 = ~n5176 & ~n5192 ;
  assign n5194 = ~n5154 & n5193 ;
  assign n5195 = \P2_reg2_reg[4]/NET0131  & n4413 ;
  assign n5196 = \P2_reg1_reg[4]/NET0131  & n4415 ;
  assign n5201 = ~n5195 & ~n5196 ;
  assign n5197 = \P2_reg0_reg[4]/NET0131  & n4417 ;
  assign n5198 = ~\P2_reg3_reg[3]/NET0131  & ~\P2_reg3_reg[4]/NET0131  ;
  assign n5199 = ~n4387 & ~n5198 ;
  assign n5200 = n4386 & n5199 ;
  assign n5202 = ~n5197 & ~n5200 ;
  assign n5203 = n5201 & n5202 ;
  assign n5204 = \P2_IR_reg[31]/NET0131  & ~n4165 ;
  assign n5205 = \P2_IR_reg[4]/NET0131  & ~n5204 ;
  assign n5206 = ~\P2_IR_reg[4]/NET0131  & n5204 ;
  assign n5207 = ~n5205 & ~n5206 ;
  assign n5208 = n4232 & ~n5207 ;
  assign n5209 = ~\P1_datao_reg[4]/NET0131  & ~n774 ;
  assign n5210 = ~n4267 & ~n4268 ;
  assign n5211 = ~n4256 & ~n4269 ;
  assign n5213 = n5210 & ~n5211 ;
  assign n5212 = ~n5210 & n5211 ;
  assign n5214 = n774 & ~n5212 ;
  assign n5215 = ~n5213 & n5214 ;
  assign n5216 = ~n5209 & ~n5215 ;
  assign n5217 = ~n4232 & n5216 ;
  assign n5218 = ~n5208 & ~n5217 ;
  assign n5219 = n5203 & n5218 ;
  assign n5220 = \P2_reg0_reg[3]/NET0131  & n4417 ;
  assign n5221 = ~\P2_reg3_reg[3]/NET0131  & n4386 ;
  assign n5224 = ~n5220 & ~n5221 ;
  assign n5222 = \P2_reg1_reg[3]/NET0131  & n4415 ;
  assign n5223 = \P2_reg2_reg[3]/NET0131  & n4413 ;
  assign n5225 = ~n5222 & ~n5223 ;
  assign n5226 = n5224 & n5225 ;
  assign n5227 = \P1_datao_reg[3]/NET0131  & ~n774 ;
  assign n5228 = ~n4257 & ~n4268 ;
  assign n5230 = n4266 & n5228 ;
  assign n5229 = ~n4266 & ~n5228 ;
  assign n5231 = n774 & ~n5229 ;
  assign n5232 = ~n5230 & n5231 ;
  assign n5233 = ~n5227 & ~n5232 ;
  assign n5234 = ~n4232 & ~n5233 ;
  assign n5235 = \P2_IR_reg[31]/NET0131  & ~n4164 ;
  assign n5236 = \P2_IR_reg[3]/NET0131  & n5235 ;
  assign n5237 = ~\P2_IR_reg[3]/NET0131  & ~n5235 ;
  assign n5238 = ~n5236 & ~n5237 ;
  assign n5239 = n4232 & n5238 ;
  assign n5240 = ~n5234 & ~n5239 ;
  assign n5241 = n5226 & n5240 ;
  assign n5242 = n5139 & n5153 ;
  assign n5243 = ~n5241 & ~n5242 ;
  assign n5244 = ~n5219 & n5243 ;
  assign n5245 = ~n5194 & n5244 ;
  assign n5246 = ~n5203 & ~n5218 ;
  assign n5247 = ~n5226 & ~n5240 ;
  assign n5248 = ~n5246 & ~n5247 ;
  assign n5249 = ~n5219 & ~n5248 ;
  assign n5250 = ~n5245 & ~n5249 ;
  assign n5084 = \P2_reg2_reg[6]/NET0131  & n4413 ;
  assign n5085 = \P2_reg1_reg[6]/NET0131  & n4415 ;
  assign n5090 = ~n5084 & ~n5085 ;
  assign n5086 = \P2_reg0_reg[6]/NET0131  & n4417 ;
  assign n5087 = ~\P2_reg3_reg[6]/NET0131  & ~n4388 ;
  assign n5088 = ~n4389 & ~n5087 ;
  assign n5089 = n4386 & n5088 ;
  assign n5091 = ~n5086 & ~n5089 ;
  assign n5092 = n5090 & n5091 ;
  assign n5093 = \P2_IR_reg[31]/NET0131  & ~n4167 ;
  assign n5094 = \P2_IR_reg[6]/NET0131  & ~n5093 ;
  assign n5095 = ~\P2_IR_reg[6]/NET0131  & n5093 ;
  assign n5096 = ~n5094 & ~n5095 ;
  assign n5097 = n4232 & ~n5096 ;
  assign n5098 = ~\P1_datao_reg[6]/NET0131  & ~n774 ;
  assign n5099 = ~n4273 & ~n4282 ;
  assign n5100 = ~n4274 & ~n4560 ;
  assign n5102 = n5099 & ~n5100 ;
  assign n5101 = ~n5099 & n5100 ;
  assign n5103 = n774 & ~n5101 ;
  assign n5104 = ~n5102 & n5103 ;
  assign n5105 = ~n5098 & ~n5104 ;
  assign n5106 = ~n4232 & n5105 ;
  assign n5107 = ~n5097 & ~n5106 ;
  assign n5108 = n5092 & n5107 ;
  assign n5109 = ~\P2_reg3_reg[5]/NET0131  & ~n4387 ;
  assign n5110 = ~n4388 & ~n5109 ;
  assign n5111 = n4386 & n5110 ;
  assign n5112 = \P2_reg1_reg[5]/NET0131  & n4415 ;
  assign n5115 = ~n5111 & ~n5112 ;
  assign n5113 = \P2_reg2_reg[5]/NET0131  & n4413 ;
  assign n5114 = \P2_reg0_reg[5]/NET0131  & n4417 ;
  assign n5116 = ~n5113 & ~n5114 ;
  assign n5117 = n5115 & n5116 ;
  assign n5118 = \P2_IR_reg[31]/NET0131  & ~n4166 ;
  assign n5119 = ~\P2_IR_reg[5]/NET0131  & ~n5118 ;
  assign n5120 = \P2_IR_reg[5]/NET0131  & n5118 ;
  assign n5121 = ~n5119 & ~n5120 ;
  assign n5122 = n4232 & ~n5121 ;
  assign n5123 = \P1_datao_reg[5]/NET0131  & ~n774 ;
  assign n5124 = ~n4274 & ~n4283 ;
  assign n5126 = ~n4272 & n5124 ;
  assign n5125 = n4272 & ~n5124 ;
  assign n5127 = n774 & ~n5125 ;
  assign n5128 = ~n5126 & n5127 ;
  assign n5129 = ~n5123 & ~n5128 ;
  assign n5130 = ~n4232 & n5129 ;
  assign n5131 = ~n5122 & ~n5130 ;
  assign n5132 = n5117 & ~n5131 ;
  assign n5251 = ~n5108 & ~n5132 ;
  assign n5252 = ~n5250 & n5251 ;
  assign n5253 = n5083 & n5252 ;
  assign n5254 = ~n5092 & ~n5107 ;
  assign n5255 = ~n5117 & n5131 ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5257 = ~n5108 & ~n5256 ;
  assign n5258 = n5083 & n5257 ;
  assign n5259 = ~n5040 & ~n5058 ;
  assign n5260 = ~n5068 & ~n5081 ;
  assign n5261 = ~n5059 & n5260 ;
  assign n5262 = ~n5259 & ~n5261 ;
  assign n5263 = ~n5258 & n5262 ;
  assign n5264 = ~n5253 & n5263 ;
  assign n5265 = n5008 & ~n5022 ;
  assign n5266 = ~n4999 & ~n5265 ;
  assign n5267 = n4975 & n5266 ;
  assign n5268 = ~n5264 & n5267 ;
  assign n5269 = n5031 & ~n5268 ;
  assign n5270 = n4922 & ~n5269 ;
  assign n5271 = ~n4827 & n4843 ;
  assign n5272 = ~n4854 & n4867 ;
  assign n5273 = ~n5271 & ~n5272 ;
  assign n5274 = ~n4844 & ~n5273 ;
  assign n5275 = n4920 & n5274 ;
  assign n5276 = ~n4879 & n4892 ;
  assign n5277 = ~n4902 & n4918 ;
  assign n5278 = ~n5276 & ~n5277 ;
  assign n5279 = ~n4893 & ~n5278 ;
  assign n5280 = ~n5275 & ~n5279 ;
  assign n5281 = n4817 & ~n5280 ;
  assign n5282 = ~n4799 & n4814 ;
  assign n5283 = ~n4774 & n4789 ;
  assign n5284 = ~n5282 & ~n5283 ;
  assign n5285 = ~n4815 & ~n5284 ;
  assign n5286 = n4765 & n5285 ;
  assign n5287 = n4754 & ~n4763 ;
  assign n5288 = ~n4728 & n4745 ;
  assign n5289 = ~n4764 & n5288 ;
  assign n5290 = ~n5287 & ~n5289 ;
  assign n5291 = ~n5286 & n5290 ;
  assign n5292 = ~n5281 & n5291 ;
  assign n5293 = ~n5270 & n5292 ;
  assign n4503 = \P1_datao_reg[27]/NET0131  & ~n774 ;
  assign n4504 = ~n4238 & ~n4343 ;
  assign n4528 = n4317 & n4339 ;
  assign n4529 = ~n4527 & n4528 ;
  assign n4530 = n4331 & n4339 ;
  assign n4531 = ~n4353 & ~n4530 ;
  assign n4532 = ~n4529 & n4531 ;
  assign n4533 = n4241 & n4336 ;
  assign n4534 = ~n4532 & n4533 ;
  assign n4535 = n4241 & n4358 ;
  assign n4536 = ~n4349 & ~n4535 ;
  assign n4537 = ~n4534 & n4536 ;
  assign n4539 = n4504 & ~n4537 ;
  assign n4538 = ~n4504 & n4537 ;
  assign n4540 = n774 & ~n4538 ;
  assign n4541 = ~n4539 & n4540 ;
  assign n4542 = ~n4503 & ~n4541 ;
  assign n4543 = ~n4232 & ~n4542 ;
  assign n4491 = \P2_reg3_reg[25]/NET0131  & n4407 ;
  assign n4492 = \P2_reg3_reg[26]/NET0131  & n4491 ;
  assign n4493 = \P2_reg3_reg[27]/NET0131  & n4492 ;
  assign n4547 = ~\P2_reg3_reg[27]/NET0131  & ~n4492 ;
  assign n4548 = ~n4493 & ~n4547 ;
  assign n4549 = n4386 & n4548 ;
  assign n4546 = \P2_reg0_reg[27]/NET0131  & n4417 ;
  assign n4544 = \P2_reg2_reg[27]/NET0131  & n4413 ;
  assign n4545 = \P2_reg1_reg[27]/NET0131  & n4415 ;
  assign n4550 = ~n4544 & ~n4545 ;
  assign n4551 = ~n4546 & n4550 ;
  assign n4552 = ~n4549 & n4551 ;
  assign n4553 = ~n4543 & n4552 ;
  assign n4554 = \P1_datao_reg[26]/NET0131  & ~n774 ;
  assign n4555 = ~n4239 & ~n4347 ;
  assign n4468 = ~n4316 & ~n4338 ;
  assign n4576 = n4457 & n4468 ;
  assign n4577 = ~n4575 & n4576 ;
  assign n4474 = ~n4329 & ~n4351 ;
  assign n4475 = ~n4338 & ~n4474 ;
  assign n4578 = n4465 & n4468 ;
  assign n4579 = ~n4475 & ~n4578 ;
  assign n4580 = ~n4577 & n4579 ;
  assign n4469 = ~n4334 & ~n4337 ;
  assign n4581 = ~n4240 & ~n4335 ;
  assign n4582 = n4469 & n4581 ;
  assign n4583 = ~n4580 & n4582 ;
  assign n4428 = ~n4346 & ~n4356 ;
  assign n4429 = ~n4240 & ~n4428 ;
  assign n4472 = ~n4350 & ~n4355 ;
  assign n4473 = ~n4334 & ~n4472 ;
  assign n4584 = n4473 & n4581 ;
  assign n4585 = ~n4429 & ~n4584 ;
  assign n4586 = ~n4583 & n4585 ;
  assign n4588 = n4555 & ~n4586 ;
  assign n4587 = ~n4555 & n4586 ;
  assign n4589 = n774 & ~n4587 ;
  assign n4590 = ~n4588 & n4589 ;
  assign n4591 = ~n4554 & ~n4590 ;
  assign n4592 = ~n4232 & ~n4591 ;
  assign n4596 = ~\P2_reg3_reg[26]/NET0131  & ~n4491 ;
  assign n4597 = ~n4492 & ~n4596 ;
  assign n4598 = n4386 & n4597 ;
  assign n4595 = \P2_reg2_reg[26]/NET0131  & n4413 ;
  assign n4593 = \P2_reg1_reg[26]/NET0131  & n4415 ;
  assign n4594 = \P2_reg0_reg[26]/NET0131  & n4417 ;
  assign n4599 = ~n4593 & ~n4594 ;
  assign n4600 = ~n4595 & n4599 ;
  assign n4601 = ~n4598 & n4600 ;
  assign n4602 = ~n4592 & n4601 ;
  assign n4603 = ~n4553 & ~n4602 ;
  assign n4605 = \P1_datao_reg[25]/NET0131  & ~n774 ;
  assign n4606 = ~n4240 & ~n4346 ;
  assign n4607 = ~n4341 & n4359 ;
  assign n4609 = n4606 & ~n4607 ;
  assign n4608 = ~n4606 & n4607 ;
  assign n4610 = n774 & ~n4608 ;
  assign n4611 = ~n4609 & n4610 ;
  assign n4612 = ~n4605 & ~n4611 ;
  assign n4613 = ~n4232 & ~n4612 ;
  assign n4617 = ~\P2_reg3_reg[25]/NET0131  & ~n4407 ;
  assign n4618 = ~n4491 & ~n4617 ;
  assign n4619 = n4386 & n4618 ;
  assign n4616 = \P2_reg0_reg[25]/NET0131  & n4417 ;
  assign n4614 = \P2_reg2_reg[25]/NET0131  & n4413 ;
  assign n4615 = \P2_reg1_reg[25]/NET0131  & n4415 ;
  assign n4620 = ~n4614 & ~n4615 ;
  assign n4621 = ~n4616 & n4620 ;
  assign n4622 = ~n4619 & n4621 ;
  assign n4626 = ~n4613 & n4622 ;
  assign n4627 = n4603 & ~n4626 ;
  assign n4425 = \P1_datao_reg[28]/NET0131  & ~n774 ;
  assign n4426 = ~n4237 & ~n4344 ;
  assign n4427 = ~n4343 & ~n4347 ;
  assign n4430 = ~n4239 & n4429 ;
  assign n4431 = n4427 & ~n4430 ;
  assign n4432 = ~n4238 & ~n4431 ;
  assign n4470 = n4468 & n4469 ;
  assign n4471 = ~n4467 & n4470 ;
  assign n4476 = n4469 & n4475 ;
  assign n4477 = ~n4473 & ~n4476 ;
  assign n4478 = ~n4471 & n4477 ;
  assign n4479 = n4242 & ~n4335 ;
  assign n4480 = ~n4478 & n4479 ;
  assign n4481 = ~n4432 & ~n4480 ;
  assign n4483 = n4426 & ~n4481 ;
  assign n4482 = ~n4426 & n4481 ;
  assign n4484 = n774 & ~n4482 ;
  assign n4485 = ~n4483 & n4484 ;
  assign n4486 = ~n4425 & ~n4485 ;
  assign n4487 = ~n4232 & ~n4486 ;
  assign n4494 = ~\P2_reg3_reg[28]/NET0131  & ~n4493 ;
  assign n4495 = \P2_reg3_reg[28]/NET0131  & n4493 ;
  assign n4496 = ~n4494 & ~n4495 ;
  assign n4497 = n4386 & n4496 ;
  assign n4490 = \P2_reg0_reg[28]/NET0131  & n4417 ;
  assign n4488 = \P2_reg1_reg[28]/NET0131  & n4415 ;
  assign n4489 = \P2_reg2_reg[28]/NET0131  & n4413 ;
  assign n4498 = ~n4488 & ~n4489 ;
  assign n4499 = ~n4490 & n4498 ;
  assign n4500 = ~n4497 & n4499 ;
  assign n4502 = ~n4487 & n4500 ;
  assign n4628 = \P1_datao_reg[24]/NET0131  & ~n774 ;
  assign n4629 = ~n4335 & ~n4356 ;
  assign n4631 = n4478 & ~n4629 ;
  assign n4630 = ~n4478 & n4629 ;
  assign n4632 = n774 & ~n4630 ;
  assign n4633 = ~n4631 & n4632 ;
  assign n4634 = ~n4628 & ~n4633 ;
  assign n4635 = ~n4232 & ~n4634 ;
  assign n4639 = \P2_reg3_reg[21]/NET0131  & n4403 ;
  assign n4640 = \P2_reg3_reg[22]/NET0131  & n4639 ;
  assign n4641 = \P2_reg3_reg[23]/NET0131  & n4640 ;
  assign n4642 = ~\P2_reg3_reg[24]/NET0131  & ~n4641 ;
  assign n4643 = ~n4407 & ~n4642 ;
  assign n4644 = n4386 & n4643 ;
  assign n4638 = \P2_reg2_reg[24]/NET0131  & n4413 ;
  assign n4636 = \P2_reg0_reg[24]/NET0131  & n4417 ;
  assign n4637 = \P2_reg1_reg[24]/NET0131  & n4415 ;
  assign n4645 = ~n4636 & ~n4637 ;
  assign n4646 = ~n4638 & n4645 ;
  assign n4647 = ~n4644 & n4646 ;
  assign n4648 = ~n4635 & n4647 ;
  assign n4649 = \P1_datao_reg[23]/NET0131  & ~n774 ;
  assign n4650 = ~n4334 & ~n4355 ;
  assign n4652 = n4532 & ~n4650 ;
  assign n4651 = ~n4532 & n4650 ;
  assign n4653 = n774 & ~n4651 ;
  assign n4654 = ~n4652 & n4653 ;
  assign n4655 = ~n4649 & ~n4654 ;
  assign n4656 = ~n4232 & ~n4655 ;
  assign n4660 = ~\P2_reg3_reg[23]/NET0131  & ~n4640 ;
  assign n4661 = ~n4641 & ~n4660 ;
  assign n4662 = n4386 & n4661 ;
  assign n4659 = \P2_reg0_reg[23]/NET0131  & n4417 ;
  assign n4657 = \P2_reg2_reg[23]/NET0131  & n4413 ;
  assign n4658 = \P2_reg1_reg[23]/NET0131  & n4415 ;
  assign n4663 = ~n4657 & ~n4658 ;
  assign n4664 = ~n4659 & n4663 ;
  assign n4665 = ~n4662 & n4664 ;
  assign n4666 = ~n4656 & n4665 ;
  assign n4667 = ~n4648 & ~n4666 ;
  assign n4668 = \P1_datao_reg[22]/NET0131  & ~n774 ;
  assign n4669 = ~n4337 & ~n4350 ;
  assign n4671 = n4580 & ~n4669 ;
  assign n4670 = ~n4580 & n4669 ;
  assign n4672 = n774 & ~n4670 ;
  assign n4673 = ~n4671 & n4672 ;
  assign n4674 = ~n4668 & ~n4673 ;
  assign n4675 = ~n4232 & ~n4674 ;
  assign n4679 = ~\P2_reg3_reg[22]/NET0131  & ~n4639 ;
  assign n4680 = ~n4640 & ~n4679 ;
  assign n4681 = n4386 & n4680 ;
  assign n4678 = \P2_reg0_reg[22]/NET0131  & n4417 ;
  assign n4676 = \P2_reg1_reg[22]/NET0131  & n4415 ;
  assign n4677 = \P2_reg2_reg[22]/NET0131  & n4413 ;
  assign n4682 = ~n4676 & ~n4677 ;
  assign n4683 = ~n4678 & n4682 ;
  assign n4684 = ~n4681 & n4683 ;
  assign n4686 = ~n4675 & n4684 ;
  assign n4687 = \P1_datao_reg[21]/NET0131  & ~n774 ;
  assign n4688 = ~n4338 & ~n4351 ;
  assign n4690 = ~n4333 & n4688 ;
  assign n4689 = n4333 & ~n4688 ;
  assign n4691 = n774 & ~n4689 ;
  assign n4692 = ~n4690 & n4691 ;
  assign n4693 = ~n4687 & ~n4692 ;
  assign n4694 = ~n4232 & ~n4693 ;
  assign n4695 = \P2_reg2_reg[21]/NET0131  & n4413 ;
  assign n4696 = ~\P2_reg3_reg[21]/NET0131  & ~n4403 ;
  assign n4697 = ~n4639 & ~n4696 ;
  assign n4698 = n4386 & n4697 ;
  assign n4701 = ~n4695 & ~n4698 ;
  assign n4699 = \P2_reg1_reg[21]/NET0131  & n4415 ;
  assign n4700 = \P2_reg0_reg[21]/NET0131  & n4417 ;
  assign n4702 = ~n4699 & ~n4700 ;
  assign n4703 = n4701 & n4702 ;
  assign n5294 = ~n4694 & n4703 ;
  assign n5295 = ~n4686 & ~n5294 ;
  assign n5296 = n4667 & n5295 ;
  assign n5297 = ~n4502 & n5296 ;
  assign n5298 = n4627 & n5297 ;
  assign n5299 = ~n5293 & n5298 ;
  assign n4501 = n4487 & ~n4500 ;
  assign n4685 = n4675 & ~n4684 ;
  assign n4704 = n4694 & ~n4703 ;
  assign n4705 = ~n4686 & n4704 ;
  assign n4706 = ~n4685 & ~n4705 ;
  assign n4707 = n4667 & ~n4706 ;
  assign n4708 = n4635 & ~n4647 ;
  assign n4709 = n4656 & ~n4665 ;
  assign n4710 = ~n4648 & n4709 ;
  assign n4711 = ~n4708 & ~n4710 ;
  assign n4712 = ~n4707 & n4711 ;
  assign n4713 = n4627 & ~n4712 ;
  assign n4604 = n4592 & ~n4601 ;
  assign n4623 = n4613 & ~n4622 ;
  assign n4624 = ~n4604 & ~n4623 ;
  assign n4625 = n4603 & ~n4624 ;
  assign n4714 = n4543 & ~n4552 ;
  assign n4715 = ~n4625 & ~n4714 ;
  assign n4716 = ~n4713 & n4715 ;
  assign n4717 = ~n4502 & ~n4716 ;
  assign n5300 = ~n4501 & ~n4717 ;
  assign n5301 = ~n5299 & n5300 ;
  assign n5302 = n4424 & ~n5301 ;
  assign n5303 = ~n4424 & n5301 ;
  assign n5304 = ~n5302 & ~n5303 ;
  assign n5305 = n4219 & ~n5304 ;
  assign n5306 = ~n4220 & ~n5305 ;
  assign n5307 = \P2_IR_reg[21]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n5308 = ~n4183 & ~n5307 ;
  assign n5309 = \P2_IR_reg[22]/NET0131  & ~n5308 ;
  assign n5310 = ~\P2_IR_reg[22]/NET0131  & n5308 ;
  assign n5311 = ~n5309 & ~n5310 ;
  assign n5312 = \P2_IR_reg[31]/NET0131  & ~n4184 ;
  assign n5313 = ~n4183 & ~n5312 ;
  assign n5314 = \P2_IR_reg[23]/NET0131  & ~n5313 ;
  assign n5315 = ~\P2_IR_reg[23]/NET0131  & n5313 ;
  assign n5316 = ~n5314 & ~n5315 ;
  assign n5317 = n5311 & n5316 ;
  assign n5318 = \P2_IR_reg[31]/NET0131  & ~n4177 ;
  assign n5319 = ~n4730 & ~n5318 ;
  assign n5320 = \P2_IR_reg[20]/NET0131  & ~n5319 ;
  assign n5321 = ~\P2_IR_reg[20]/NET0131  & n5319 ;
  assign n5322 = ~n5320 & ~n5321 ;
  assign n5323 = n5316 & ~n5322 ;
  assign n5324 = \P2_IR_reg[21]/NET0131  & ~n4183 ;
  assign n5325 = ~\P2_IR_reg[21]/NET0131  & n4183 ;
  assign n5326 = ~n5324 & ~n5325 ;
  assign n5327 = n5311 & n5326 ;
  assign n5328 = ~n5323 & ~n5327 ;
  assign n5329 = ~n5317 & ~n5328 ;
  assign n5330 = ~n5306 & n5329 ;
  assign n5331 = n4231 & ~n4500 ;
  assign n5334 = \P2_reg0_reg[30]/NET0131  & n4417 ;
  assign n5337 = ~n4412 & ~n5334 ;
  assign n5335 = \P2_reg1_reg[30]/NET0131  & n4415 ;
  assign n5336 = \P2_reg2_reg[30]/NET0131  & n4413 ;
  assign n5338 = ~n5335 & ~n5336 ;
  assign n5339 = n5337 & n5338 ;
  assign n5340 = \P2_reg2_reg[31]/NET0131  & n4413 ;
  assign n5343 = ~n4412 & ~n5340 ;
  assign n5341 = \P2_reg1_reg[31]/NET0131  & n4415 ;
  assign n5342 = \P2_reg0_reg[31]/NET0131  & n4417 ;
  assign n5344 = ~n5341 & ~n5342 ;
  assign n5345 = n5343 & n5344 ;
  assign n5346 = ~n5184 & ~n5345 ;
  assign n5347 = ~n5161 & n5346 ;
  assign n5348 = ~n5139 & n5347 ;
  assign n5349 = ~n5226 & n5348 ;
  assign n5350 = ~n5117 & ~n5203 ;
  assign n5351 = n5349 & n5350 ;
  assign n5352 = ~n5092 & n5351 ;
  assign n5353 = ~n5068 & n5352 ;
  assign n5354 = ~n4931 & ~n4984 ;
  assign n5355 = ~n5008 & ~n5040 ;
  assign n5356 = n5354 & n5355 ;
  assign n5357 = n5353 & n5356 ;
  assign n5358 = ~n4827 & ~n4854 ;
  assign n5359 = ~n4902 & ~n4958 ;
  assign n5360 = n5358 & n5359 ;
  assign n5361 = n5357 & n5360 ;
  assign n5362 = ~n4774 & ~n4879 ;
  assign n5363 = ~n4799 & n5362 ;
  assign n5364 = n5361 & n5363 ;
  assign n5366 = ~n4684 & ~n4703 ;
  assign n5367 = ~n4665 & n5366 ;
  assign n5368 = ~n4647 & n5367 ;
  assign n5365 = ~n4728 & ~n4763 ;
  assign n5369 = ~n4622 & n5365 ;
  assign n5370 = n5368 & n5369 ;
  assign n5371 = n5364 & n5370 ;
  assign n5372 = ~n4500 & ~n4552 ;
  assign n5373 = ~n4421 & n5372 ;
  assign n5374 = ~n4601 & n5373 ;
  assign n5375 = n5371 & n5374 ;
  assign n5377 = n5339 & ~n5375 ;
  assign n5332 = ~\P2_B_reg/NET0131  & ~n4231 ;
  assign n5333 = ~n4232 & ~n5332 ;
  assign n5376 = ~n5339 & n5375 ;
  assign n5378 = ~n5333 & ~n5376 ;
  assign n5379 = ~n5377 & n5378 ;
  assign n5380 = ~n5331 & ~n5379 ;
  assign n5381 = n4219 & ~n5380 ;
  assign n5382 = ~n4220 & ~n5381 ;
  assign n5383 = n5323 & n5327 ;
  assign n5384 = ~n5382 & n5383 ;
  assign n5385 = n4728 & n4745 ;
  assign n5386 = n4754 & n4763 ;
  assign n5387 = ~n5385 & ~n5386 ;
  assign n5388 = n4774 & n4789 ;
  assign n5389 = n4799 & n4814 ;
  assign n5390 = ~n5388 & ~n5389 ;
  assign n5391 = n5387 & n5390 ;
  assign n5392 = n4854 & n4867 ;
  assign n5393 = n4827 & n4843 ;
  assign n5394 = n4902 & n4918 ;
  assign n5395 = n4879 & n4892 ;
  assign n5396 = ~n5394 & ~n5395 ;
  assign n5397 = ~n5393 & n5396 ;
  assign n5398 = ~n5392 & n5397 ;
  assign n5399 = n5391 & n5398 ;
  assign n5400 = n4958 & n4973 ;
  assign n5401 = ~n4958 & ~n4973 ;
  assign n5402 = ~n4931 & ~n4948 ;
  assign n5403 = ~n5401 & ~n5402 ;
  assign n5404 = n4931 & n4948 ;
  assign n5405 = n4984 & ~n4997 ;
  assign n5406 = ~n5008 & ~n5022 ;
  assign n5407 = ~n4984 & n4997 ;
  assign n5408 = ~n5406 & ~n5407 ;
  assign n5409 = ~n5405 & ~n5408 ;
  assign n5410 = ~n5404 & n5409 ;
  assign n5411 = n5403 & ~n5410 ;
  assign n5412 = ~n5400 & ~n5411 ;
  assign n5413 = n5203 & ~n5218 ;
  assign n5414 = ~n5226 & n5240 ;
  assign n5415 = ~n5203 & n5218 ;
  assign n5416 = ~n5414 & ~n5415 ;
  assign n5417 = ~n5413 & ~n5416 ;
  assign n5418 = n5161 & ~n5175 ;
  assign n5419 = n5184 & ~n5190 ;
  assign n5420 = ~n5418 & ~n5419 ;
  assign n5421 = ~n5161 & n5175 ;
  assign n5422 = ~n5139 & n5153 ;
  assign n5423 = ~n5421 & ~n5422 ;
  assign n5424 = ~n5420 & n5423 ;
  assign n5425 = n5226 & ~n5240 ;
  assign n5426 = n5139 & ~n5153 ;
  assign n5427 = ~n5425 & ~n5426 ;
  assign n5428 = ~n5413 & n5427 ;
  assign n5429 = ~n5424 & n5428 ;
  assign n5430 = ~n5417 & ~n5429 ;
  assign n5431 = n5068 & ~n5081 ;
  assign n5432 = n5040 & ~n5058 ;
  assign n5433 = ~n5431 & ~n5432 ;
  assign n5434 = n5092 & ~n5107 ;
  assign n5435 = n5117 & n5131 ;
  assign n5436 = ~n5434 & ~n5435 ;
  assign n5437 = n5433 & n5436 ;
  assign n5438 = ~n5430 & n5437 ;
  assign n5439 = ~n5117 & ~n5131 ;
  assign n5440 = ~n5092 & n5107 ;
  assign n5441 = ~n5439 & ~n5440 ;
  assign n5442 = ~n5434 & ~n5441 ;
  assign n5443 = n5433 & n5442 ;
  assign n5444 = ~n5040 & n5058 ;
  assign n5445 = ~n5068 & n5081 ;
  assign n5446 = ~n5444 & ~n5445 ;
  assign n5447 = ~n5432 & ~n5446 ;
  assign n5448 = ~n5443 & ~n5447 ;
  assign n5449 = ~n5438 & n5448 ;
  assign n5450 = ~n5404 & ~n5405 ;
  assign n5451 = n5008 & n5022 ;
  assign n5452 = ~n5400 & ~n5451 ;
  assign n5453 = n5450 & n5452 ;
  assign n5454 = ~n5449 & n5453 ;
  assign n5455 = ~n5412 & ~n5454 ;
  assign n5456 = n5399 & ~n5455 ;
  assign n5457 = ~n4879 & ~n4892 ;
  assign n5458 = ~n4902 & ~n4918 ;
  assign n5459 = ~n5457 & ~n5458 ;
  assign n5460 = ~n5395 & ~n5459 ;
  assign n5461 = ~n4827 & ~n4843 ;
  assign n5462 = ~n4854 & ~n4867 ;
  assign n5463 = ~n5461 & ~n5462 ;
  assign n5464 = n5397 & ~n5463 ;
  assign n5465 = ~n5460 & ~n5464 ;
  assign n5466 = n5391 & ~n5465 ;
  assign n5467 = ~n4799 & ~n4814 ;
  assign n5468 = ~n4774 & ~n4789 ;
  assign n5469 = ~n5467 & ~n5468 ;
  assign n5470 = ~n5389 & ~n5469 ;
  assign n5471 = n5387 & n5470 ;
  assign n5472 = ~n4754 & ~n4763 ;
  assign n5473 = ~n4728 & ~n4745 ;
  assign n5474 = ~n5472 & ~n5473 ;
  assign n5475 = ~n5386 & ~n5474 ;
  assign n5476 = ~n5471 & ~n5475 ;
  assign n5477 = ~n5466 & n5476 ;
  assign n5478 = ~n5456 & n5477 ;
  assign n5479 = n4675 & n4684 ;
  assign n5480 = n4694 & n4703 ;
  assign n5481 = ~n5479 & ~n5480 ;
  assign n5482 = n4656 & n4665 ;
  assign n5483 = n4635 & n4647 ;
  assign n5484 = ~n5482 & ~n5483 ;
  assign n5485 = n5481 & n5484 ;
  assign n5486 = n4613 & n4622 ;
  assign n5487 = n4592 & n4601 ;
  assign n5488 = ~n5486 & ~n5487 ;
  assign n5489 = n4543 & n4552 ;
  assign n5490 = n4487 & n4500 ;
  assign n5491 = ~n5489 & ~n5490 ;
  assign n5492 = n5488 & n5491 ;
  assign n5493 = n5485 & n5492 ;
  assign n5494 = ~n5478 & n5493 ;
  assign n5506 = ~n4592 & ~n4601 ;
  assign n5507 = ~n4613 & ~n4622 ;
  assign n5508 = ~n5506 & ~n5507 ;
  assign n5509 = ~n5487 & ~n5508 ;
  assign n5510 = n5491 & n5509 ;
  assign n5495 = ~n4675 & ~n4684 ;
  assign n5496 = ~n4694 & ~n4703 ;
  assign n5497 = ~n5495 & ~n5496 ;
  assign n5498 = ~n5479 & ~n5497 ;
  assign n5499 = n5484 & n5498 ;
  assign n5500 = ~n4635 & ~n4647 ;
  assign n5501 = ~n4656 & ~n4665 ;
  assign n5502 = ~n5500 & ~n5501 ;
  assign n5503 = ~n5483 & ~n5502 ;
  assign n5504 = ~n5499 & ~n5503 ;
  assign n5505 = n5492 & ~n5504 ;
  assign n5511 = ~n4487 & ~n4500 ;
  assign n5512 = ~n4543 & ~n4552 ;
  assign n5513 = ~n5490 & n5512 ;
  assign n5514 = ~n5511 & ~n5513 ;
  assign n5515 = ~n5505 & n5514 ;
  assign n5516 = ~n5510 & n5515 ;
  assign n5517 = ~n5494 & n5516 ;
  assign n5518 = ~n4424 & n5517 ;
  assign n5519 = n4424 & ~n5517 ;
  assign n5520 = ~n5518 & ~n5519 ;
  assign n5521 = n4219 & n5520 ;
  assign n5522 = ~n4220 & ~n5521 ;
  assign n5523 = n5311 & ~n5326 ;
  assign n5524 = n5316 & n5322 ;
  assign n5525 = ~n5523 & ~n5524 ;
  assign n5526 = ~n5317 & ~n5525 ;
  assign n5527 = ~n5522 & n5526 ;
  assign n5529 = n5175 & n5190 ;
  assign n5530 = n5153 & n5529 ;
  assign n5531 = n5240 & n5530 ;
  assign n5532 = n5218 & n5531 ;
  assign n5533 = n5107 & ~n5131 ;
  assign n5534 = n5532 & n5533 ;
  assign n5535 = n5058 & n5081 ;
  assign n5536 = n5534 & n5535 ;
  assign n5537 = n4997 & ~n5022 ;
  assign n5538 = n5536 & n5537 ;
  assign n5539 = ~n4948 & ~n4973 ;
  assign n5540 = n5538 & n5539 ;
  assign n5541 = ~n4843 & ~n4918 ;
  assign n5542 = ~n4867 & ~n4892 ;
  assign n5543 = n5541 & n5542 ;
  assign n5544 = n5540 & n5543 ;
  assign n5528 = ~n4745 & ~n4814 ;
  assign n5545 = ~n4754 & ~n4789 ;
  assign n5546 = n5528 & n5545 ;
  assign n5547 = n5544 & n5546 ;
  assign n5548 = ~n4635 & ~n4656 ;
  assign n5549 = ~n4675 & ~n4694 ;
  assign n5550 = n5548 & n5549 ;
  assign n5551 = ~n4613 & n5550 ;
  assign n5552 = ~n4592 & n5551 ;
  assign n5553 = n5547 & n5552 ;
  assign n5554 = ~n4543 & n5553 ;
  assign n5555 = ~n4487 & n5554 ;
  assign n5556 = n4371 & ~n5555 ;
  assign n5557 = ~n4371 & n5555 ;
  assign n5558 = ~n5556 & ~n5557 ;
  assign n5559 = n4219 & n5558 ;
  assign n5560 = ~n4220 & ~n5559 ;
  assign n5561 = ~n5322 & n5326 ;
  assign n5562 = ~n5311 & ~n5316 ;
  assign n5563 = n5561 & n5562 ;
  assign n5564 = ~n5560 & n5563 ;
  assign n5565 = ~n5326 & n5562 ;
  assign n5566 = n4371 & n5565 ;
  assign n5567 = n4219 & n5566 ;
  assign n5568 = n5317 & ~n5561 ;
  assign n5569 = ~n4219 & n5565 ;
  assign n5570 = ~n5568 & ~n5569 ;
  assign n5571 = \P2_reg2_reg[29]/NET0131  & ~n5570 ;
  assign n5572 = ~n5311 & n5326 ;
  assign n5573 = ~n5316 & n5322 ;
  assign n5574 = n5572 & n5573 ;
  assign n5575 = n4411 & n5574 ;
  assign n5576 = ~n5571 & ~n5575 ;
  assign n5577 = ~n5567 & n5576 ;
  assign n5578 = ~n5564 & n5577 ;
  assign n5579 = ~n5527 & n5578 ;
  assign n5580 = ~n5384 & n5579 ;
  assign n5581 = ~n5330 & n5580 ;
  assign n5582 = n4190 & n4207 ;
  assign n5583 = ~n5316 & ~n5582 ;
  assign n5584 = ~n5581 & n5583 ;
  assign n5585 = ~n5316 & n5582 ;
  assign n5586 = \P2_reg2_reg[29]/NET0131  & n5585 ;
  assign n5587 = ~n5584 & ~n5586 ;
  assign n5588 = \P1_state_reg[0]/NET0131  & ~n5587 ;
  assign n5589 = \P1_state_reg[0]/NET0131  & ~n5316 ;
  assign n5590 = \P2_reg2_reg[29]/NET0131  & ~n5589 ;
  assign n5591 = ~n5588 & ~n5590 ;
  assign n5594 = ~n1232 & n2145 ;
  assign n5595 = ~n1232 & ~n2236 ;
  assign n5627 = n1963 & ~n1986 ;
  assign n5628 = n1960 & ~n5627 ;
  assign n5629 = n1085 & ~n5628 ;
  assign n5625 = n1980 & n2010 ;
  assign n5626 = n1964 & n5625 ;
  assign n5630 = n1082 & ~n5626 ;
  assign n5631 = ~n5629 & n5630 ;
  assign n5632 = n2071 & ~n5631 ;
  assign n5633 = ~n2071 & n5631 ;
  assign n5634 = ~n5632 & ~n5633 ;
  assign n5635 = n2236 & ~n5634 ;
  assign n5636 = ~n5595 & ~n5635 ;
  assign n5637 = n2234 & ~n5636 ;
  assign n5610 = ~n1232 & ~n2163 ;
  assign n5614 = ~n933 & n2239 ;
  assign n5615 = ~n1000 & n2264 ;
  assign n5616 = ~n933 & n5615 ;
  assign n5617 = ~n1236 & n5616 ;
  assign n5618 = ~n1272 & ~n2239 ;
  assign n5619 = ~n5617 & ~n5618 ;
  assign n5620 = ~n2268 & ~n5619 ;
  assign n5621 = ~n5614 & ~n5620 ;
  assign n5622 = n2163 & ~n5621 ;
  assign n5623 = ~n5610 & ~n5622 ;
  assign n5624 = n737 & ~n5623 ;
  assign n5638 = ~n1232 & ~n2583 ;
  assign n5639 = n1223 & n2580 ;
  assign n5640 = ~n5638 & ~n5639 ;
  assign n5641 = ~n5624 & n5640 ;
  assign n5642 = ~n5637 & n5641 ;
  assign n5599 = n2467 & n2474 ;
  assign n5596 = ~n2450 & n2473 ;
  assign n5597 = n2480 & ~n5596 ;
  assign n5598 = n2471 & ~n5597 ;
  assign n5600 = ~n2487 & ~n5598 ;
  assign n5601 = ~n5599 & n5600 ;
  assign n5602 = n2492 & ~n5601 ;
  assign n5603 = n2501 & ~n5602 ;
  assign n5604 = n2071 & n5603 ;
  assign n5605 = ~n2071 & ~n5603 ;
  assign n5606 = ~n5604 & ~n5605 ;
  assign n5607 = n2236 & ~n5606 ;
  assign n5608 = ~n5595 & ~n5607 ;
  assign n5609 = n2391 & ~n5608 ;
  assign n5611 = n2163 & ~n5606 ;
  assign n5612 = ~n5610 & ~n5611 ;
  assign n5613 = n2393 & ~n5612 ;
  assign n5643 = ~n5609 & ~n5613 ;
  assign n5644 = n5642 & n5643 ;
  assign n5645 = n2147 & ~n5644 ;
  assign n5646 = ~n5594 & ~n5645 ;
  assign n5647 = \P1_state_reg[0]/NET0131  & ~n5646 ;
  assign n5592 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[24]/NET0131  ;
  assign n5593 = n765 & ~n1232 ;
  assign n5648 = ~n5592 & ~n5593 ;
  assign n5649 = ~n5647 & n5648 ;
  assign n5650 = \P3_reg2_reg[25]/NET0131  & ~n2143 ;
  assign n5651 = \P3_reg2_reg[25]/NET0131  & n2145 ;
  assign n5652 = \P3_reg2_reg[25]/NET0131  & ~n2408 ;
  assign n5653 = ~n2209 & n2213 ;
  assign n5654 = n2221 & ~n5653 ;
  assign n5655 = n2058 & ~n5654 ;
  assign n5656 = ~n2058 & n5654 ;
  assign n5657 = ~n5655 & ~n5656 ;
  assign n5658 = n2408 & ~n5657 ;
  assign n5659 = ~n5652 & ~n5658 ;
  assign n5660 = n2425 & ~n5659 ;
  assign n5675 = ~n1474 & n2268 ;
  assign n5674 = n1474 & ~n2268 ;
  assign n5676 = ~n2239 & ~n5674 ;
  assign n5677 = ~n5675 & n5676 ;
  assign n5678 = ~n1236 & n2239 ;
  assign n5679 = ~n5677 & ~n5678 ;
  assign n5680 = n2408 & ~n5679 ;
  assign n5681 = ~n5652 & ~n5680 ;
  assign n5682 = n737 & ~n5681 ;
  assign n5684 = n1262 & n2441 ;
  assign n5673 = \P3_reg2_reg[25]/NET0131  & ~n2429 ;
  assign n5683 = ~n1268 & n2283 ;
  assign n5685 = ~n5673 & ~n5683 ;
  assign n5686 = ~n5684 & n5685 ;
  assign n5687 = ~n5682 & n5686 ;
  assign n5688 = ~n5660 & n5687 ;
  assign n5661 = \P3_reg2_reg[25]/NET0131  & ~n2427 ;
  assign n5662 = n2427 & ~n5657 ;
  assign n5663 = ~n5661 & ~n5662 ;
  assign n5664 = ~n2518 & ~n5663 ;
  assign n5665 = ~n2362 & n2368 ;
  assign n5666 = n2375 & ~n5665 ;
  assign n5667 = n2058 & n5666 ;
  assign n5668 = ~n2058 & ~n5666 ;
  assign n5669 = ~n5667 & ~n5668 ;
  assign n5670 = n2427 & ~n5669 ;
  assign n5671 = ~n5661 & ~n5670 ;
  assign n5672 = n714 & ~n5671 ;
  assign n5689 = ~n5664 & ~n5672 ;
  assign n5690 = n5688 & n5689 ;
  assign n5691 = n2147 & ~n5690 ;
  assign n5692 = ~n5651 & ~n5691 ;
  assign n5693 = \P1_state_reg[0]/NET0131  & ~n5692 ;
  assign n5694 = ~n5650 & ~n5693 ;
  assign n5695 = \P3_reg2_reg[26]/NET0131  & ~n2143 ;
  assign n5696 = \P3_reg2_reg[26]/NET0131  & n2145 ;
  assign n5697 = \P3_reg2_reg[26]/NET0131  & ~n2427 ;
  assign n5698 = n1002 & n1489 ;
  assign n5699 = n1706 & n1770 ;
  assign n5700 = ~n1975 & n5699 ;
  assign n5701 = n1706 & n1978 ;
  assign n5702 = ~n1981 & ~n5701 ;
  assign n5703 = ~n5700 & n5702 ;
  assign n5704 = n1654 & n1714 ;
  assign n5705 = ~n5703 & n5704 ;
  assign n5706 = n1714 & n1983 ;
  assign n5707 = ~n1598 & ~n5706 ;
  assign n5708 = ~n5705 & n5707 ;
  assign n5709 = n1199 & n1546 ;
  assign n5710 = ~n5708 & n5709 ;
  assign n5711 = n1199 & n1603 ;
  assign n5712 = ~n1956 & ~n5711 ;
  assign n5713 = ~n5710 & n5712 ;
  assign n5714 = n1084 & n1139 ;
  assign n5715 = ~n5713 & n5714 ;
  assign n5716 = n5698 & n5715 ;
  assign n5717 = n1084 & ~n1959 ;
  assign n5718 = ~n1076 & ~n5717 ;
  assign n5719 = n5698 & ~n5718 ;
  assign n5720 = n1081 & ~n1488 ;
  assign n5721 = n1274 & ~n5720 ;
  assign n5722 = ~n1487 & ~n5721 ;
  assign n5723 = ~n5719 & ~n5722 ;
  assign n5724 = ~n5716 & n5723 ;
  assign n5725 = n2042 & ~n5724 ;
  assign n5726 = ~n2042 & n5724 ;
  assign n5727 = ~n5725 & ~n5726 ;
  assign n5728 = n2427 & ~n5727 ;
  assign n5729 = ~n5697 & ~n5728 ;
  assign n5730 = ~n2518 & ~n5729 ;
  assign n5761 = \P3_reg2_reg[26]/NET0131  & ~n2408 ;
  assign n5766 = ~n1272 & n2239 ;
  assign n5767 = n1445 & ~n5675 ;
  assign n5768 = ~n2239 & ~n2570 ;
  assign n5769 = ~n5767 & n5768 ;
  assign n5770 = ~n5766 & ~n5769 ;
  assign n5771 = n2408 & ~n5770 ;
  assign n5772 = ~n5761 & ~n5771 ;
  assign n5773 = n737 & ~n5772 ;
  assign n5765 = n1465 & n2441 ;
  assign n5774 = \P3_reg2_reg[26]/NET0131  & ~n2429 ;
  assign n5775 = ~n1470 & n2283 ;
  assign n5776 = ~n5774 & ~n5775 ;
  assign n5777 = ~n5765 & n5776 ;
  assign n5778 = ~n5773 & n5777 ;
  assign n5779 = ~n5730 & n5778 ;
  assign n5731 = ~n2482 & n2550 ;
  assign n5732 = n2497 & ~n5731 ;
  assign n5733 = n2367 & ~n5732 ;
  assign n5734 = ~n2069 & ~n2500 ;
  assign n5735 = n2503 & ~n5734 ;
  assign n5736 = ~n5733 & n5735 ;
  assign n5737 = ~n2056 & ~n5736 ;
  assign n5738 = n2446 & ~n2466 ;
  assign n5739 = n2444 & n2472 ;
  assign n5740 = ~n5738 & n5739 ;
  assign n5741 = n2343 & n2469 ;
  assign n5742 = n5740 & n5741 ;
  assign n5743 = ~n2075 & ~n2449 ;
  assign n5744 = n2476 & ~n5743 ;
  assign n5745 = ~n2082 & ~n5744 ;
  assign n5746 = n5741 & n5745 ;
  assign n5747 = n2469 & n2479 ;
  assign n5748 = n2484 & ~n5747 ;
  assign n5749 = ~n5746 & n5748 ;
  assign n5750 = ~n5742 & n5749 ;
  assign n5751 = ~n2056 & n2351 ;
  assign n5752 = n2368 & n5751 ;
  assign n5753 = ~n5750 & n5752 ;
  assign n5754 = ~n5737 & ~n5753 ;
  assign n5755 = n2042 & n5754 ;
  assign n5756 = ~n2042 & ~n5754 ;
  assign n5757 = ~n5755 & ~n5756 ;
  assign n5758 = n2427 & ~n5757 ;
  assign n5759 = ~n5697 & ~n5758 ;
  assign n5760 = n714 & ~n5759 ;
  assign n5762 = n2408 & ~n5727 ;
  assign n5763 = ~n5761 & ~n5762 ;
  assign n5764 = n2425 & ~n5763 ;
  assign n5780 = ~n5760 & ~n5764 ;
  assign n5781 = n5779 & n5780 ;
  assign n5782 = n2147 & ~n5781 ;
  assign n5783 = ~n5696 & ~n5782 ;
  assign n5784 = \P1_state_reg[0]/NET0131  & ~n5783 ;
  assign n5785 = ~n5695 & ~n5784 ;
  assign n5786 = \P1_state_reg[0]/NET0131  & n5316 ;
  assign n5787 = \P2_B_reg/NET0131  & ~n5786 ;
  assign n5861 = ~\P1_datao_reg[30]/NET0131  & ~\si[30]_pad  ;
  assign n5862 = ~n4235 & ~n4237 ;
  assign n5863 = ~n4238 & n5862 ;
  assign n5864 = ~n5861 & n5863 ;
  assign n5865 = ~n4537 & n5864 ;
  assign n5866 = ~n4345 & n5862 ;
  assign n5867 = ~n4234 & ~n5866 ;
  assign n5868 = ~n5861 & ~n5867 ;
  assign n5869 = \P1_datao_reg[30]/NET0131  & \si[30]_pad  ;
  assign n5870 = ~n5868 & ~n5869 ;
  assign n5871 = ~n5865 & n5870 ;
  assign n5872 = ~n1337 & n5871 ;
  assign n5873 = ~\si[31]_pad  & n774 ;
  assign n5874 = ~n5871 & ~n5873 ;
  assign n5875 = ~n5872 & ~n5874 ;
  assign n5876 = \P1_datao_reg[31]/NET0131  & ~n5875 ;
  assign n5877 = ~\P1_datao_reg[31]/NET0131  & n5875 ;
  assign n5878 = ~n5876 & ~n5877 ;
  assign n5879 = ~n4232 & ~n5878 ;
  assign n5947 = n5345 & n5879 ;
  assign n5880 = ~n5345 & ~n5879 ;
  assign n5881 = \P1_datao_reg[30]/NET0131  & ~n774 ;
  assign n5882 = ~n5861 & ~n5869 ;
  assign n5883 = ~n4239 & n5863 ;
  assign n5884 = ~n4586 & n5883 ;
  assign n5886 = ~n4427 & n5863 ;
  assign n5885 = ~n4235 & n4344 ;
  assign n5887 = ~n4234 & ~n5885 ;
  assign n5888 = ~n5886 & n5887 ;
  assign n5889 = ~n5884 & n5888 ;
  assign n5891 = n5882 & ~n5889 ;
  assign n5890 = ~n5882 & n5889 ;
  assign n5892 = n774 & ~n5890 ;
  assign n5893 = ~n5891 & n5892 ;
  assign n5894 = ~n5881 & ~n5893 ;
  assign n5895 = ~n4232 & ~n5894 ;
  assign n5953 = n5339 & n5895 ;
  assign n5954 = ~n5880 & ~n5953 ;
  assign n5904 = ~n5339 & ~n5895 ;
  assign n5955 = ~n4423 & ~n5904 ;
  assign n5956 = ~n4422 & ~n5490 ;
  assign n5788 = ~n5487 & ~n5489 ;
  assign n5789 = ~n5483 & ~n5486 ;
  assign n5790 = n5788 & n5789 ;
  assign n5791 = ~n5458 & ~n5461 ;
  assign n5792 = ~n5394 & ~n5791 ;
  assign n5793 = ~n5393 & ~n5394 ;
  assign n5794 = ~n5401 & ~n5462 ;
  assign n5795 = ~n5392 & ~n5794 ;
  assign n5796 = n5793 & n5795 ;
  assign n5797 = ~n5792 & ~n5796 ;
  assign n5798 = ~n5402 & ~n5407 ;
  assign n5799 = ~n5404 & ~n5798 ;
  assign n5800 = ~n5406 & ~n5444 ;
  assign n5801 = ~n5451 & ~n5800 ;
  assign n5802 = n5450 & n5801 ;
  assign n5803 = ~n5799 & ~n5802 ;
  assign n5804 = ~n5392 & ~n5400 ;
  assign n5805 = ~n5393 & n5804 ;
  assign n5806 = ~n5394 & n5805 ;
  assign n5807 = ~n5803 & n5806 ;
  assign n5808 = n5797 & ~n5807 ;
  assign n5809 = ~n5431 & ~n5434 ;
  assign n5810 = ~n5413 & ~n5435 ;
  assign n5811 = ~n5420 & ~n5421 ;
  assign n5812 = n5427 & ~n5811 ;
  assign n5813 = ~n5414 & ~n5422 ;
  assign n5814 = ~n5425 & ~n5813 ;
  assign n5815 = ~n5812 & ~n5814 ;
  assign n5816 = n5810 & ~n5815 ;
  assign n5817 = n5809 & n5816 ;
  assign n5818 = ~n5415 & ~n5439 ;
  assign n5819 = ~n5435 & ~n5818 ;
  assign n5820 = n5809 & n5819 ;
  assign n5821 = ~n5431 & n5440 ;
  assign n5822 = ~n5445 & ~n5821 ;
  assign n5823 = ~n5820 & n5822 ;
  assign n5824 = ~n5817 & n5823 ;
  assign n5825 = ~n5432 & ~n5451 ;
  assign n5826 = n5450 & n5825 ;
  assign n5827 = ~n5824 & n5826 ;
  assign n5828 = n5806 & n5827 ;
  assign n5829 = n5808 & ~n5828 ;
  assign n5830 = ~n5479 & ~n5482 ;
  assign n5831 = ~n5386 & ~n5480 ;
  assign n5832 = n5830 & n5831 ;
  assign n5833 = ~n5385 & ~n5389 ;
  assign n5834 = ~n5388 & ~n5395 ;
  assign n5835 = n5833 & n5834 ;
  assign n5836 = n5832 & n5835 ;
  assign n5837 = ~n5829 & n5836 ;
  assign n5838 = ~n5457 & ~n5468 ;
  assign n5839 = ~n5388 & ~n5838 ;
  assign n5840 = n5833 & n5839 ;
  assign n5841 = ~n5467 & ~n5473 ;
  assign n5842 = ~n5385 & ~n5841 ;
  assign n5843 = ~n5840 & ~n5842 ;
  assign n5844 = n5832 & ~n5843 ;
  assign n5845 = ~n5472 & ~n5496 ;
  assign n5846 = ~n5480 & ~n5845 ;
  assign n5847 = n5830 & n5846 ;
  assign n5848 = ~n5495 & ~n5501 ;
  assign n5849 = ~n5482 & ~n5848 ;
  assign n5850 = ~n5847 & ~n5849 ;
  assign n5851 = ~n5844 & n5850 ;
  assign n5852 = ~n5837 & n5851 ;
  assign n5853 = n5790 & ~n5852 ;
  assign n5854 = ~n5506 & ~n5512 ;
  assign n5855 = ~n5500 & ~n5507 ;
  assign n5856 = ~n5486 & ~n5855 ;
  assign n5857 = ~n5487 & n5856 ;
  assign n5858 = n5854 & ~n5857 ;
  assign n5859 = ~n5489 & ~n5858 ;
  assign n6054 = ~n5511 & ~n5859 ;
  assign n6055 = ~n5853 & n6054 ;
  assign n6056 = n5956 & ~n6055 ;
  assign n6057 = n5955 & ~n6056 ;
  assign n6058 = n5954 & ~n6057 ;
  assign n6059 = ~n5947 & ~n6058 ;
  assign n6063 = ~n5322 & ~n6059 ;
  assign n6060 = \P2_B_reg/NET0131  & n5316 ;
  assign n6061 = n5322 & ~n6060 ;
  assign n6062 = n6059 & n6061 ;
  assign n6064 = n5572 & ~n6062 ;
  assign n6065 = ~n6063 & n6064 ;
  assign n5860 = ~n5853 & ~n5859 ;
  assign n5896 = ~n5339 & ~n5345 ;
  assign n5897 = n5895 & ~n5896 ;
  assign n5898 = ~n4422 & ~n5880 ;
  assign n5899 = ~n5897 & n5898 ;
  assign n5900 = ~n5490 & n5899 ;
  assign n5901 = ~n5860 & n5900 ;
  assign n5902 = ~n4423 & ~n5511 ;
  assign n5903 = n5899 & ~n5902 ;
  assign n5905 = ~n5345 & ~n5904 ;
  assign n5906 = n5879 & ~n5905 ;
  assign n5907 = ~n5903 & ~n5906 ;
  assign n5908 = ~n5901 & n5907 ;
  assign n5968 = ~n5316 & ~n5322 ;
  assign n6051 = n5908 & ~n5968 ;
  assign n6050 = ~n5573 & ~n5908 ;
  assign n6052 = n5523 & ~n6050 ;
  assign n6053 = ~n6051 & n6052 ;
  assign n6047 = ~\P2_B_reg/NET0131  & n5908 ;
  assign n6048 = n5523 & n5524 ;
  assign n6049 = ~n6047 & n6048 ;
  assign n5909 = ~\P2_B_reg/NET0131  & ~n5908 ;
  assign n5910 = n5323 & n5523 ;
  assign n5911 = ~n5909 & n5910 ;
  assign n5912 = n5469 & ~n5834 ;
  assign n5913 = n5833 & ~n5912 ;
  assign n5914 = n5474 & ~n5913 ;
  assign n5915 = n5831 & ~n5914 ;
  assign n5916 = n5497 & ~n5915 ;
  assign n5917 = n5830 & ~n5916 ;
  assign n5918 = ~n5501 & ~n5917 ;
  assign n5919 = ~n5184 & n5190 ;
  assign n5920 = ~n5418 & n5919 ;
  assign n5921 = n5423 & ~n5920 ;
  assign n5922 = n5427 & ~n5921 ;
  assign n5923 = n5416 & ~n5922 ;
  assign n5924 = n5810 & ~n5923 ;
  assign n5925 = n5441 & ~n5924 ;
  assign n5926 = n5809 & ~n5925 ;
  assign n5927 = ~n5445 & n5798 ;
  assign n5928 = n5800 & n5927 ;
  assign n5929 = n5791 & n5794 ;
  assign n5930 = n5928 & n5929 ;
  assign n5931 = ~n5926 & n5930 ;
  assign n5935 = ~n5393 & ~n5463 ;
  assign n5936 = ~n5458 & ~n5805 ;
  assign n5937 = ~n5935 & n5936 ;
  assign n5932 = n5408 & ~n5825 ;
  assign n5933 = n5450 & ~n5932 ;
  assign n5934 = ~n5402 & ~n5933 ;
  assign n5938 = ~n5394 & ~n5934 ;
  assign n5939 = ~n5937 & n5938 ;
  assign n5940 = n5797 & ~n5939 ;
  assign n5941 = ~n5931 & ~n5940 ;
  assign n5942 = n5838 & n5841 ;
  assign n5943 = n5845 & n5942 ;
  assign n5944 = n5848 & n5943 ;
  assign n5945 = ~n5941 & n5944 ;
  assign n5946 = ~n5918 & ~n5945 ;
  assign n5948 = ~n5904 & ~n5947 ;
  assign n5949 = n5902 & n5948 ;
  assign n5950 = n5854 & n5855 ;
  assign n5951 = n5949 & n5950 ;
  assign n5952 = ~n5946 & n5951 ;
  assign n5957 = n5955 & ~n5956 ;
  assign n5958 = n5954 & ~n5957 ;
  assign n5959 = ~n5947 & ~n5958 ;
  assign n5960 = n5508 & ~n5789 ;
  assign n5961 = n5788 & ~n5960 ;
  assign n5962 = ~n5512 & ~n5961 ;
  assign n5963 = n5949 & n5962 ;
  assign n5964 = ~n5959 & ~n5963 ;
  assign n5965 = ~n5952 & n5964 ;
  assign n5966 = n5327 & n5573 ;
  assign n5967 = n5965 & ~n5966 ;
  assign n5969 = n5327 & n5968 ;
  assign n5970 = ~n5965 & ~n5969 ;
  assign n5971 = ~n5967 & ~n5970 ;
  assign n5982 = ~n4553 & ~n4714 ;
  assign n5990 = ~n4815 & ~n5282 ;
  assign n5979 = ~n4790 & ~n5283 ;
  assign n5986 = ~n4666 & ~n4709 ;
  assign n6018 = ~n5979 & ~n5986 ;
  assign n6019 = ~n5990 & n6018 ;
  assign n5993 = ~n5059 & ~n5259 ;
  assign n5994 = ~n5413 & ~n5415 ;
  assign n6005 = ~n5993 & n5994 ;
  assign n5995 = ~n5241 & ~n5247 ;
  assign n5996 = ~n4974 & ~n5027 ;
  assign n6006 = ~n5995 & ~n5996 ;
  assign n6007 = n6005 & n6006 ;
  assign n5980 = ~n5082 & ~n5260 ;
  assign n5981 = ~n5434 & ~n5440 ;
  assign n6003 = ~n5980 & n5981 ;
  assign n5991 = ~n4949 & ~n5028 ;
  assign n5992 = ~n5405 & ~n5407 ;
  assign n6004 = ~n5991 & n5992 ;
  assign n6008 = n6003 & n6004 ;
  assign n6014 = n6007 & n6008 ;
  assign n5978 = ~n4764 & ~n5287 ;
  assign n5987 = ~n4746 & ~n5288 ;
  assign n6015 = ~n5978 & ~n5987 ;
  assign n6016 = n6014 & n6015 ;
  assign n6000 = ~n4868 & ~n5272 ;
  assign n5997 = ~n4893 & ~n5276 ;
  assign n5999 = ~n4844 & ~n5271 ;
  assign n6011 = ~n5997 & ~n5999 ;
  assign n6012 = ~n6000 & n6011 ;
  assign n5974 = ~n5154 & ~n5242 ;
  assign n6001 = ~n5919 & ~n5974 ;
  assign n5975 = ~n5023 & ~n5265 ;
  assign n5976 = ~n5132 & ~n5255 ;
  assign n6002 = ~n5975 & ~n5976 ;
  assign n6009 = n6001 & n6002 ;
  assign n5972 = ~n5418 & ~n5421 ;
  assign n5973 = ~n5419 & n5972 ;
  assign n5988 = ~n4919 & ~n5277 ;
  assign n6010 = n5973 & ~n5988 ;
  assign n6013 = n6009 & n6010 ;
  assign n6017 = n6012 & n6013 ;
  assign n6020 = n6016 & n6017 ;
  assign n6023 = n6019 & n6020 ;
  assign n6024 = ~n5982 & n6023 ;
  assign n5977 = ~n4602 & ~n4604 ;
  assign n5989 = ~n4704 & ~n5294 ;
  assign n5983 = ~n4685 & ~n4686 ;
  assign n5984 = ~n4648 & ~n4708 ;
  assign n6021 = ~n5983 & ~n5984 ;
  assign n6022 = ~n5989 & n6021 ;
  assign n6025 = ~n5977 & n6022 ;
  assign n5985 = ~n4501 & ~n4502 ;
  assign n5998 = ~n4623 & ~n4626 ;
  assign n6026 = ~n5985 & ~n5998 ;
  assign n6027 = n6025 & n6026 ;
  assign n6028 = n6024 & n6027 ;
  assign n6029 = n4424 & n5948 ;
  assign n6030 = n5954 & n6029 ;
  assign n6031 = n6028 & n6030 ;
  assign n6039 = ~\P2_B_reg/NET0131  & n6031 ;
  assign n6036 = ~n5311 & ~n5326 ;
  assign n6040 = n5524 & n6036 ;
  assign n6041 = ~n6039 & n6040 ;
  assign n6037 = ~n5322 & n6036 ;
  assign n6038 = n6031 & n6037 ;
  assign n6032 = n5322 & n5565 ;
  assign n6033 = ~n6031 & n6032 ;
  assign n6034 = \P2_B_reg/NET0131  & ~n5311 ;
  assign n6035 = n5323 & n6034 ;
  assign n6066 = ~n6033 & ~n6035 ;
  assign n6067 = ~n6038 & n6066 ;
  assign n6068 = ~n6041 & n6067 ;
  assign n6069 = ~n5971 & n6068 ;
  assign n6042 = ~\P2_B_reg/NET0131  & n5965 ;
  assign n6043 = n5383 & ~n6042 ;
  assign n6044 = ~\P2_B_reg/NET0131  & ~n5965 ;
  assign n6045 = n5327 & n5524 ;
  assign n6046 = ~n6044 & n6045 ;
  assign n6070 = ~n6043 & ~n6046 ;
  assign n6071 = n6069 & n6070 ;
  assign n6072 = ~n5911 & n6071 ;
  assign n6073 = ~n6049 & n6072 ;
  assign n6074 = ~n6053 & n6073 ;
  assign n6075 = ~n6065 & n6074 ;
  assign n6076 = n5786 & ~n6075 ;
  assign n6077 = ~n5787 & ~n6076 ;
  assign n6078 = \P1_state_reg[0]/NET0131  & ~n3867 ;
  assign n6079 = \P1_reg2_reg[29]/NET0131  & ~n6078 ;
  assign n6088 = \P1_IR_reg[31]/NET0131  & ~n2704 ;
  assign n6089 = ~n2684 & ~n6088 ;
  assign n6090 = \P1_IR_reg[24]/NET0131  & ~n6089 ;
  assign n6091 = ~\P1_IR_reg[24]/NET0131  & n6089 ;
  assign n6092 = ~n6090 & ~n6091 ;
  assign n6080 = \P1_IR_reg[26]/NET0131  & ~n2832 ;
  assign n6081 = ~\P1_IR_reg[26]/NET0131  & n2832 ;
  assign n6082 = ~n6080 & ~n6081 ;
  assign n6083 = \P1_IR_reg[31]/NET0131  & ~n2843 ;
  assign n6084 = ~n2695 & ~n6083 ;
  assign n6085 = \P1_IR_reg[25]/NET0131  & ~n6084 ;
  assign n6086 = ~\P1_IR_reg[25]/NET0131  & n6084 ;
  assign n6087 = ~n6085 & ~n6086 ;
  assign n6093 = ~n6082 & n6087 ;
  assign n6094 = n6092 & n6093 ;
  assign n6095 = ~n3867 & n6094 ;
  assign n6096 = \P1_reg2_reg[29]/NET0131  & n6095 ;
  assign n6097 = ~n3867 & ~n6094 ;
  assign n6098 = ~n6082 & ~n6087 ;
  assign n6102 = ~\P1_B_reg/NET0131  & n6092 ;
  assign n6103 = n6098 & n6102 ;
  assign n6099 = \P1_B_reg/NET0131  & ~n6092 ;
  assign n6100 = n6098 & n6099 ;
  assign n6101 = n6082 & n6092 ;
  assign n6104 = \P1_d_reg[0]/NET0131  & ~n6082 ;
  assign n6105 = ~n6101 & ~n6104 ;
  assign n6106 = ~n6100 & n6105 ;
  assign n6107 = ~n6103 & n6106 ;
  assign n6108 = n6082 & n6087 ;
  assign n6109 = \P1_d_reg[1]/NET0131  & ~n6082 ;
  assign n6110 = ~n6108 & ~n6109 ;
  assign n6111 = ~n6100 & n6110 ;
  assign n6112 = ~n6103 & n6111 ;
  assign n6113 = n6107 & ~n6112 ;
  assign n6114 = \P1_reg2_reg[29]/NET0131  & ~n6113 ;
  assign n6115 = ~n2953 & ~n3598 ;
  assign n6116 = ~n3083 & ~n3110 ;
  assign n6117 = n6115 & n6116 ;
  assign n6118 = ~n3230 & ~n3355 ;
  assign n6119 = ~n3205 & ~n3624 ;
  assign n6120 = n6118 & n6119 ;
  assign n6121 = n6117 & n6120 ;
  assign n6122 = ~n3256 & ~n3651 ;
  assign n6123 = n3330 & ~n3678 ;
  assign n6124 = ~n3679 & ~n6123 ;
  assign n6125 = n6122 & ~n6124 ;
  assign n6126 = n3257 & ~n3651 ;
  assign n6127 = ~n3652 & ~n6126 ;
  assign n6128 = ~n6125 & n6127 ;
  assign n6129 = n3786 & n3795 ;
  assign n6130 = n3756 & n3770 ;
  assign n6131 = ~n6129 & ~n6130 ;
  assign n6132 = ~n3364 & ~n3378 ;
  assign n6133 = n3364 & n3378 ;
  assign n6134 = n3704 & n3718 ;
  assign n6135 = ~n3704 & ~n3718 ;
  assign n6136 = ~n3687 & ~n3694 ;
  assign n6137 = ~n6135 & ~n6136 ;
  assign n6138 = ~n6134 & ~n6137 ;
  assign n6139 = ~n6133 & n6138 ;
  assign n6140 = ~n6132 & ~n6139 ;
  assign n6141 = n6131 & ~n6140 ;
  assign n6142 = ~n3786 & ~n3795 ;
  assign n6143 = ~n3756 & ~n3770 ;
  assign n6144 = ~n6129 & n6143 ;
  assign n6145 = ~n6142 & ~n6144 ;
  assign n6146 = ~n6141 & n6145 ;
  assign n6147 = ~n3139 & ~n3747 ;
  assign n6148 = ~n3578 & ~n3823 ;
  assign n6149 = n6147 & n6148 ;
  assign n6150 = ~n6146 & n6149 ;
  assign n6151 = ~n3138 & ~n3748 ;
  assign n6152 = ~n3747 & ~n6151 ;
  assign n6153 = n6148 & n6152 ;
  assign n6154 = n3579 & ~n3823 ;
  assign n6155 = ~n3824 & ~n6154 ;
  assign n6156 = ~n6153 & n6155 ;
  assign n6157 = ~n6150 & n6156 ;
  assign n6158 = ~n3331 & ~n3678 ;
  assign n6159 = n6122 & n6158 ;
  assign n6160 = ~n6157 & n6159 ;
  assign n6161 = n6128 & ~n6160 ;
  assign n6162 = n6121 & ~n6161 ;
  assign n6163 = ~n3230 & n3356 ;
  assign n6164 = ~n3231 & ~n6163 ;
  assign n6165 = n6119 & ~n6164 ;
  assign n6166 = ~n3204 & ~n3625 ;
  assign n6167 = ~n3205 & ~n6166 ;
  assign n6168 = ~n6165 & ~n6167 ;
  assign n6169 = n6117 & ~n6168 ;
  assign n6170 = ~n3082 & ~n3111 ;
  assign n6171 = ~n3110 & ~n6170 ;
  assign n6172 = n6115 & n6171 ;
  assign n6173 = n2954 & ~n3598 ;
  assign n6174 = ~n3599 & ~n6173 ;
  assign n6175 = ~n6172 & n6174 ;
  assign n6176 = ~n6169 & n6175 ;
  assign n6177 = ~n6162 & n6176 ;
  assign n6178 = ~n3177 & ~n3529 ;
  assign n6179 = ~n3035 & ~n3439 ;
  assign n6180 = n6178 & n6179 ;
  assign n6181 = ~n2888 & ~n3285 ;
  assign n6182 = ~n3549 & n6181 ;
  assign n6183 = ~n3304 & n6182 ;
  assign n6184 = n6180 & n6183 ;
  assign n6185 = ~n6177 & n6184 ;
  assign n6192 = ~n3178 & ~n3528 ;
  assign n6193 = ~n3529 & ~n6192 ;
  assign n6194 = ~n3438 & ~n6193 ;
  assign n6195 = n6179 & ~n6194 ;
  assign n6186 = ~n2889 & ~n3305 ;
  assign n6187 = n6182 & ~n6186 ;
  assign n6188 = n3284 & ~n3549 ;
  assign n6189 = ~n3550 & ~n6188 ;
  assign n6190 = ~n6187 & n6189 ;
  assign n6191 = n6180 & ~n6190 ;
  assign n6196 = ~n3036 & ~n6191 ;
  assign n6197 = ~n6195 & n6196 ;
  assign n6198 = ~n6185 & n6197 ;
  assign n6199 = ~n3413 & n6198 ;
  assign n6200 = n3413 & ~n6198 ;
  assign n6201 = ~n6199 & ~n6200 ;
  assign n6202 = n6113 & ~n6201 ;
  assign n6203 = ~n6114 & ~n6202 ;
  assign n6204 = n2690 & n3867 ;
  assign n6205 = ~n4069 & ~n4079 ;
  assign n6206 = ~n4110 & n6205 ;
  assign n6207 = ~n6204 & n6206 ;
  assign n6208 = ~n6203 & n6207 ;
  assign n6209 = ~n3889 & ~n3891 ;
  assign n6210 = ~n3888 & ~n3900 ;
  assign n6211 = n6209 & n6210 ;
  assign n6212 = ~n3771 & ~n3796 ;
  assign n6213 = ~n3379 & n4042 ;
  assign n6214 = ~n3380 & ~n6213 ;
  assign n6215 = n6212 & ~n6214 ;
  assign n6216 = ~n3772 & ~n3797 ;
  assign n6217 = ~n3796 & ~n6216 ;
  assign n6218 = ~n6215 & ~n6217 ;
  assign n6219 = ~n3892 & ~n3909 ;
  assign n6220 = ~n3910 & ~n3912 ;
  assign n6221 = n6219 & n6220 ;
  assign n6222 = ~n6218 & n6221 ;
  assign n6223 = n6211 & n6222 ;
  assign n6224 = ~n3910 & ~n3916 ;
  assign n6225 = n6219 & n6224 ;
  assign n6226 = ~n3892 & n3908 ;
  assign n6227 = ~n3932 & ~n6226 ;
  assign n6228 = ~n6225 & n6227 ;
  assign n6229 = n6211 & ~n6228 ;
  assign n6230 = ~n3889 & ~n3896 ;
  assign n6231 = n6210 & n6230 ;
  assign n6232 = ~n3900 & ~n3934 ;
  assign n6233 = ~n6231 & ~n6232 ;
  assign n6234 = ~n6229 & n6233 ;
  assign n6235 = ~n6223 & n6234 ;
  assign n6236 = ~n3961 & ~n3967 ;
  assign n6237 = ~n3968 & ~n3970 ;
  assign n6238 = n6236 & n6237 ;
  assign n6239 = ~n3874 & ~n3971 ;
  assign n6240 = ~n3873 & ~n3877 ;
  assign n6241 = n6239 & n6240 ;
  assign n6242 = n6238 & n6241 ;
  assign n6243 = ~n6235 & n6242 ;
  assign n6244 = ~n3873 & ~n3902 ;
  assign n6245 = n6239 & n6244 ;
  assign n6246 = n3882 & ~n3971 ;
  assign n6247 = ~n3950 & ~n6246 ;
  assign n6248 = ~n6245 & n6247 ;
  assign n6249 = n6238 & ~n6248 ;
  assign n6250 = ~n3953 & ~n3968 ;
  assign n6251 = n6236 & n6250 ;
  assign n6252 = ~n3947 & ~n3961 ;
  assign n6253 = ~n6251 & ~n6252 ;
  assign n6254 = ~n6249 & n6253 ;
  assign n6255 = ~n6243 & n6254 ;
  assign n6256 = ~n3957 & ~n3960 ;
  assign n6257 = ~n3958 & ~n3990 ;
  assign n6258 = n6256 & n6257 ;
  assign n6259 = ~n3987 & ~n3989 ;
  assign n6260 = ~n3986 & ~n4001 ;
  assign n6261 = n6259 & n6260 ;
  assign n6262 = n6258 & n6261 ;
  assign n6263 = ~n6255 & n6262 ;
  assign n6264 = ~n3957 & ~n3963 ;
  assign n6265 = n6257 & n6264 ;
  assign n6266 = n3941 & ~n3990 ;
  assign n6267 = ~n3982 & ~n6266 ;
  assign n6268 = ~n6265 & n6267 ;
  assign n6269 = n6261 & ~n6268 ;
  assign n6270 = ~n3987 & ~n3992 ;
  assign n6271 = n6260 & n6270 ;
  assign n6272 = n3979 & ~n4001 ;
  assign n6273 = ~n3997 & ~n6272 ;
  assign n6274 = ~n6271 & n6273 ;
  assign n6275 = ~n6269 & n6274 ;
  assign n6276 = ~n6263 & n6275 ;
  assign n6277 = n3413 & ~n6276 ;
  assign n6278 = ~n3413 & n6276 ;
  assign n6279 = ~n6277 & ~n6278 ;
  assign n6280 = n6113 & n6279 ;
  assign n6281 = ~n6114 & ~n6280 ;
  assign n6282 = ~n6204 & ~n6205 ;
  assign n6283 = ~n6281 & n6282 ;
  assign n6284 = n2713 & ~n3034 ;
  assign n6285 = ~n3473 & ~n3687 ;
  assign n6286 = ~n3704 & n6285 ;
  assign n6287 = ~n3364 & n6286 ;
  assign n6288 = ~n3756 & n6287 ;
  assign n6289 = ~n3137 & ~n3795 ;
  assign n6290 = n6288 & n6289 ;
  assign n6291 = ~n3746 & n6290 ;
  assign n6292 = ~n3577 & ~n3822 ;
  assign n6293 = n6291 & n6292 ;
  assign n6294 = ~n3255 & ~n3650 ;
  assign n6295 = ~n3354 & ~n3677 ;
  assign n6296 = n6294 & n6295 ;
  assign n6297 = ~n3203 & ~n3229 ;
  assign n6298 = ~n3329 & ~n3623 ;
  assign n6299 = n6297 & n6298 ;
  assign n6300 = n6296 & n6299 ;
  assign n6301 = n6293 & n6300 ;
  assign n6302 = ~n3081 & ~n3109 ;
  assign n6303 = n6301 & n6302 ;
  assign n6305 = ~n3303 & ~n3597 ;
  assign n6306 = ~n2887 & ~n2952 ;
  assign n6307 = n6305 & n6306 ;
  assign n6308 = ~n3283 & n6307 ;
  assign n6309 = ~n3548 & n6308 ;
  assign n6304 = ~n3176 & ~n3527 ;
  assign n6310 = ~n3437 & n6304 ;
  assign n6311 = n6309 & n6310 ;
  assign n6312 = n6303 & n6311 ;
  assign n6313 = ~n3034 & n6312 ;
  assign n6314 = ~n3410 & n6313 ;
  assign n6315 = n3506 & ~n6314 ;
  assign n6316 = ~n3410 & ~n3506 ;
  assign n6317 = n6313 & n6316 ;
  assign n6318 = \P1_B_reg/NET0131  & n2725 ;
  assign n6319 = ~n2713 & ~n6318 ;
  assign n6320 = ~n6317 & n6319 ;
  assign n6321 = ~n6315 & n6320 ;
  assign n6322 = ~n6284 & ~n6321 ;
  assign n6323 = n6113 & ~n6322 ;
  assign n6324 = ~n6114 & ~n6323 ;
  assign n6325 = n4011 & ~n6324 ;
  assign n6328 = n3694 & n3718 ;
  assign n6329 = n3378 & n6328 ;
  assign n6330 = n3770 & n6329 ;
  assign n6331 = n3786 & n6330 ;
  assign n6332 = n3128 & n6331 ;
  assign n6333 = ~n3737 & n6332 ;
  assign n6334 = ~n3568 & n6333 ;
  assign n6335 = ~n3813 & n6334 ;
  assign n6336 = ~n3320 & n6335 ;
  assign n6337 = ~n3246 & ~n3668 ;
  assign n6338 = n6336 & n6337 ;
  assign n6339 = ~n3219 & ~n3345 ;
  assign n6340 = ~n3641 & n6339 ;
  assign n6341 = n6338 & n6340 ;
  assign n6342 = ~n3072 & ~n3614 ;
  assign n6343 = ~n3100 & n6342 ;
  assign n6344 = ~n3194 & n6343 ;
  assign n6345 = n6341 & n6344 ;
  assign n6346 = ~n2830 & ~n3294 ;
  assign n6347 = ~n2942 & ~n3588 ;
  assign n6348 = ~n3273 & n6347 ;
  assign n6349 = n6346 & n6348 ;
  assign n6350 = n6345 & n6349 ;
  assign n6326 = ~n3165 & ~n3518 ;
  assign n6327 = ~n3427 & n6326 ;
  assign n6351 = ~n3019 & ~n3539 ;
  assign n6352 = n6327 & n6351 ;
  assign n6353 = n6350 & n6352 ;
  assign n6354 = ~n3403 & n6353 ;
  assign n6355 = n3403 & ~n6353 ;
  assign n6356 = ~n6354 & ~n6355 ;
  assign n6357 = n6113 & n6356 ;
  assign n6358 = ~n6114 & ~n6357 ;
  assign n6359 = ~n3867 & n4114 ;
  assign n6360 = ~n6358 & n6359 ;
  assign n6363 = n3403 & n6113 ;
  assign n6364 = ~n6114 & ~n6363 ;
  assign n6365 = n2699 & n4110 ;
  assign n6366 = ~n6364 & n6365 ;
  assign n6361 = ~n4009 & n6204 ;
  assign n6362 = \P1_reg2_reg[29]/NET0131  & n6361 ;
  assign n6367 = n3028 & n4112 ;
  assign n6368 = ~n6362 & ~n6367 ;
  assign n6369 = ~n6366 & n6368 ;
  assign n6370 = ~n6360 & n6369 ;
  assign n6371 = ~n6325 & n6370 ;
  assign n6372 = ~n6283 & n6371 ;
  assign n6373 = ~n6208 & n6372 ;
  assign n6374 = n6097 & ~n6373 ;
  assign n6375 = ~n6096 & ~n6374 ;
  assign n6376 = \P1_state_reg[0]/NET0131  & ~n6375 ;
  assign n6377 = ~n6079 & ~n6376 ;
  assign n6378 = \P2_reg1_reg[29]/NET0131  & ~n5589 ;
  assign n6379 = \P2_reg1_reg[29]/NET0131  & n5585 ;
  assign n6380 = ~n4211 & ~n4218 ;
  assign n6381 = \P2_reg1_reg[29]/NET0131  & ~n6380 ;
  assign n6382 = ~n5304 & n6380 ;
  assign n6383 = ~n6381 & ~n6382 ;
  assign n6384 = n5329 & ~n6383 ;
  assign n6385 = ~n5380 & n6380 ;
  assign n6386 = ~n6381 & ~n6385 ;
  assign n6387 = n5383 & ~n6386 ;
  assign n6388 = n5520 & n5526 ;
  assign n6389 = n5558 & n5563 ;
  assign n6390 = ~n5566 & ~n6389 ;
  assign n6391 = ~n6388 & n6390 ;
  assign n6392 = n6380 & ~n6391 ;
  assign n6393 = n5526 & ~n6380 ;
  assign n6394 = ~n5568 & ~n5574 ;
  assign n6395 = ~n5563 & ~n5565 ;
  assign n6396 = ~n6380 & ~n6395 ;
  assign n6397 = n6394 & ~n6396 ;
  assign n6398 = ~n6393 & n6397 ;
  assign n6399 = \P2_reg1_reg[29]/NET0131  & ~n6398 ;
  assign n6400 = ~n6392 & ~n6399 ;
  assign n6401 = ~n6387 & n6400 ;
  assign n6402 = ~n6384 & n6401 ;
  assign n6403 = n5583 & ~n6402 ;
  assign n6404 = ~n6379 & ~n6403 ;
  assign n6405 = \P1_state_reg[0]/NET0131  & ~n6404 ;
  assign n6406 = ~n6378 & ~n6405 ;
  assign n6407 = \P1_reg0_reg[29]/NET0131  & ~n6078 ;
  assign n6408 = \P1_reg0_reg[29]/NET0131  & n6095 ;
  assign n6409 = n6107 & n6112 ;
  assign n6410 = \P1_reg0_reg[29]/NET0131  & ~n6409 ;
  assign n6411 = ~n6201 & n6409 ;
  assign n6412 = ~n6410 & ~n6411 ;
  assign n6413 = n6207 & ~n6412 ;
  assign n6414 = n6279 & n6409 ;
  assign n6415 = ~n6410 & ~n6414 ;
  assign n6416 = n6282 & ~n6415 ;
  assign n6417 = n4011 & ~n6322 ;
  assign n6418 = n3403 & n6365 ;
  assign n6419 = n6356 & n6359 ;
  assign n6420 = ~n6418 & ~n6419 ;
  assign n6421 = ~n6417 & n6420 ;
  assign n6422 = n6409 & ~n6421 ;
  assign n6423 = n6365 & ~n6409 ;
  assign n6424 = ~n4112 & ~n6361 ;
  assign n6425 = ~n6423 & n6424 ;
  assign n6426 = ~n4110 & ~n6204 ;
  assign n6427 = n4009 & ~n6426 ;
  assign n6428 = ~n6409 & n6427 ;
  assign n6429 = n6425 & ~n6428 ;
  assign n6430 = \P1_reg0_reg[29]/NET0131  & ~n6429 ;
  assign n6431 = ~n6422 & ~n6430 ;
  assign n6432 = ~n6416 & n6431 ;
  assign n6433 = ~n6413 & n6432 ;
  assign n6434 = n6097 & ~n6433 ;
  assign n6435 = ~n6408 & ~n6434 ;
  assign n6436 = \P1_state_reg[0]/NET0131  & ~n6435 ;
  assign n6437 = ~n6407 & ~n6436 ;
  assign n6438 = \P3_reg1_reg[29]/NET0131  & ~n2143 ;
  assign n6439 = \P3_reg1_reg[29]/NET0131  & n2145 ;
  assign n6440 = \P3_reg1_reg[29]/NET0131  & ~n2408 ;
  assign n6441 = n2230 & n2408 ;
  assign n6442 = ~n6440 & ~n6441 ;
  assign n6443 = ~n2518 & ~n6442 ;
  assign n6444 = \P3_reg1_reg[29]/NET0131  & ~n2427 ;
  assign n6445 = ~n2277 & n2427 ;
  assign n6446 = ~n6444 & ~n6445 ;
  assign n6447 = n737 & ~n6446 ;
  assign n6448 = n2285 & ~n2408 ;
  assign n6449 = n2284 & ~n6448 ;
  assign n6450 = \P3_reg1_reg[29]/NET0131  & ~n6449 ;
  assign n6451 = n2285 & n2408 ;
  assign n6452 = n1385 & n6451 ;
  assign n6459 = ~n6450 & ~n6452 ;
  assign n6460 = ~n6447 & n6459 ;
  assign n6461 = ~n6443 & n6460 ;
  assign n6453 = ~n2387 & n2408 ;
  assign n6454 = ~n6440 & ~n6453 ;
  assign n6455 = n714 & ~n6454 ;
  assign n6456 = n2230 & n2427 ;
  assign n6457 = ~n6444 & ~n6456 ;
  assign n6458 = n2425 & ~n6457 ;
  assign n6462 = ~n6455 & ~n6458 ;
  assign n6463 = n6461 & n6462 ;
  assign n6464 = n2147 & ~n6463 ;
  assign n6465 = ~n6439 & ~n6464 ;
  assign n6466 = \P1_state_reg[0]/NET0131  & ~n6465 ;
  assign n6467 = ~n6438 & ~n6466 ;
  assign n6468 = \P3_reg2_reg[24]/NET0131  & ~n2143 ;
  assign n6469 = \P3_reg2_reg[24]/NET0131  & n2145 ;
  assign n6470 = \P3_reg2_reg[24]/NET0131  & ~n2427 ;
  assign n6471 = n2427 & ~n5606 ;
  assign n6472 = ~n6470 & ~n6471 ;
  assign n6473 = n714 & ~n6472 ;
  assign n6474 = \P3_reg2_reg[24]/NET0131  & ~n2408 ;
  assign n6475 = n2408 & ~n5634 ;
  assign n6476 = ~n6474 & ~n6475 ;
  assign n6477 = n2425 & ~n6476 ;
  assign n6480 = n1223 & n2441 ;
  assign n6478 = \P3_reg2_reg[24]/NET0131  & ~n2429 ;
  assign n6479 = ~n1232 & n2283 ;
  assign n6487 = ~n6478 & ~n6479 ;
  assign n6488 = ~n6480 & n6487 ;
  assign n6489 = ~n6477 & n6488 ;
  assign n6481 = n2427 & ~n5634 ;
  assign n6482 = ~n6470 & ~n6481 ;
  assign n6483 = ~n2518 & ~n6482 ;
  assign n6484 = n2408 & ~n5621 ;
  assign n6485 = ~n6474 & ~n6484 ;
  assign n6486 = n737 & ~n6485 ;
  assign n6490 = ~n6483 & ~n6486 ;
  assign n6491 = n6489 & n6490 ;
  assign n6492 = ~n6473 & n6491 ;
  assign n6493 = n2147 & ~n6492 ;
  assign n6494 = ~n6469 & ~n6493 ;
  assign n6495 = \P1_state_reg[0]/NET0131  & ~n6494 ;
  assign n6496 = ~n6468 & ~n6495 ;
  assign n6497 = \P3_reg2_reg[29]/NET0131  & ~n2143 ;
  assign n6498 = \P3_reg2_reg[29]/NET0131  & n2145 ;
  assign n6499 = \P3_reg2_reg[29]/NET0131  & ~n2427 ;
  assign n6500 = ~n6456 & ~n6499 ;
  assign n6501 = ~n2518 & ~n6500 ;
  assign n6502 = \P3_reg2_reg[29]/NET0131  & ~n2408 ;
  assign n6508 = ~n2277 & n2408 ;
  assign n6509 = ~n6502 & ~n6508 ;
  assign n6510 = n737 & ~n6509 ;
  assign n6511 = n1385 & n2441 ;
  assign n6512 = \P3_reg2_reg[29]/NET0131  & ~n2429 ;
  assign n6513 = n1325 & n2283 ;
  assign n6514 = ~n6512 & ~n6513 ;
  assign n6515 = ~n6511 & n6514 ;
  assign n6516 = ~n6510 & n6515 ;
  assign n6517 = ~n6501 & n6516 ;
  assign n6503 = ~n6441 & ~n6502 ;
  assign n6504 = n2425 & ~n6503 ;
  assign n6505 = ~n2387 & n2427 ;
  assign n6506 = ~n6499 & ~n6505 ;
  assign n6507 = n714 & ~n6506 ;
  assign n6518 = ~n6504 & ~n6507 ;
  assign n6519 = n6517 & n6518 ;
  assign n6520 = n2147 & ~n6519 ;
  assign n6521 = ~n6498 & ~n6520 ;
  assign n6522 = \P1_state_reg[0]/NET0131  & ~n6521 ;
  assign n6523 = ~n6497 & ~n6522 ;
  assign n6526 = ~n1090 & n2145 ;
  assign n6528 = ~n1090 & ~n2163 ;
  assign n6529 = n2092 & ~n2549 ;
  assign n6530 = ~n2092 & n2549 ;
  assign n6531 = ~n6529 & ~n6530 ;
  assign n6532 = n2163 & ~n6531 ;
  assign n6533 = ~n6528 & ~n6532 ;
  assign n6534 = n2393 & ~n6533 ;
  assign n6535 = ~n1090 & ~n2236 ;
  assign n6550 = n2092 & ~n2603 ;
  assign n6551 = ~n2092 & n2603 ;
  assign n6552 = ~n6550 & ~n6551 ;
  assign n6553 = n2236 & n6552 ;
  assign n6554 = ~n6535 & ~n6553 ;
  assign n6555 = n2234 & ~n6554 ;
  assign n6527 = ~n1110 & n2580 ;
  assign n6556 = ~n1090 & ~n2583 ;
  assign n6557 = ~n6527 & ~n6556 ;
  assign n6558 = ~n6555 & n6557 ;
  assign n6559 = ~n6534 & n6558 ;
  assign n6536 = n2236 & ~n6531 ;
  assign n6537 = ~n6535 & ~n6536 ;
  assign n6538 = n2391 & ~n6537 ;
  assign n6539 = ~n1121 & n2260 ;
  assign n6540 = ~n1095 & n6539 ;
  assign n6542 = n1072 & ~n6540 ;
  assign n6541 = ~n1072 & n6540 ;
  assign n6543 = ~n2239 & ~n6541 ;
  assign n6544 = ~n6542 & n6543 ;
  assign n6545 = ~n1121 & n2239 ;
  assign n6546 = ~n6544 & ~n6545 ;
  assign n6547 = n2163 & ~n6546 ;
  assign n6548 = ~n6528 & ~n6547 ;
  assign n6549 = n737 & ~n6548 ;
  assign n6560 = ~n6538 & ~n6549 ;
  assign n6561 = n6559 & n6560 ;
  assign n6562 = n2147 & ~n6561 ;
  assign n6563 = ~n6526 & ~n6562 ;
  assign n6564 = \P1_state_reg[0]/NET0131  & ~n6563 ;
  assign n6524 = n765 & ~n1090 ;
  assign n6525 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[19]/NET0131  ;
  assign n6565 = ~n6524 & ~n6525 ;
  assign n6566 = ~n6564 & n6565 ;
  assign n6567 = n3433 & n6095 ;
  assign n6568 = ~n6107 & ~n6112 ;
  assign n6569 = n3433 & ~n6568 ;
  assign n6570 = n6212 & n6220 ;
  assign n6571 = ~n6214 & n6570 ;
  assign n6572 = n6217 & n6220 ;
  assign n6573 = ~n6224 & ~n6572 ;
  assign n6574 = ~n6571 & n6573 ;
  assign n6575 = n6209 & n6219 ;
  assign n6576 = ~n6574 & n6575 ;
  assign n6577 = n6209 & ~n6227 ;
  assign n6578 = ~n6230 & ~n6577 ;
  assign n6579 = ~n6576 & n6578 ;
  assign n6580 = n6210 & n6240 ;
  assign n6581 = ~n6579 & n6580 ;
  assign n6582 = n6232 & n6240 ;
  assign n6583 = ~n6244 & ~n6582 ;
  assign n6584 = ~n6581 & n6583 ;
  assign n6585 = n6237 & n6239 ;
  assign n6586 = ~n6584 & n6585 ;
  assign n6587 = n6237 & ~n6247 ;
  assign n6588 = ~n6250 & ~n6587 ;
  assign n6589 = ~n6586 & n6588 ;
  assign n6590 = n6236 & n6256 ;
  assign n6591 = n6257 & n6259 ;
  assign n6592 = n6590 & n6591 ;
  assign n6593 = ~n6589 & n6592 ;
  assign n6595 = n6252 & n6256 ;
  assign n6596 = ~n6264 & ~n6595 ;
  assign n6597 = n6591 & ~n6596 ;
  assign n6594 = n6259 & ~n6267 ;
  assign n6598 = ~n6270 & ~n6594 ;
  assign n6599 = ~n6597 & n6598 ;
  assign n6600 = ~n6593 & n6599 ;
  assign n6601 = n3440 & ~n6600 ;
  assign n6602 = ~n3440 & n6600 ;
  assign n6603 = ~n6601 & ~n6602 ;
  assign n6604 = n6568 & ~n6603 ;
  assign n6605 = ~n6569 & ~n6604 ;
  assign n6606 = n6282 & ~n6605 ;
  assign n6607 = n6116 & n6119 ;
  assign n6608 = n6131 & n6147 ;
  assign n6609 = ~n6140 & n6608 ;
  assign n6610 = ~n6145 & n6147 ;
  assign n6611 = ~n6152 & ~n6610 ;
  assign n6612 = ~n6609 & n6611 ;
  assign n6613 = n6148 & n6158 ;
  assign n6614 = ~n6612 & n6613 ;
  assign n6615 = ~n6155 & n6158 ;
  assign n6616 = n6124 & ~n6615 ;
  assign n6617 = ~n6614 & n6616 ;
  assign n6618 = n6118 & n6122 ;
  assign n6619 = ~n6617 & n6618 ;
  assign n6620 = n6607 & n6619 ;
  assign n6621 = n6118 & ~n6127 ;
  assign n6622 = n6164 & ~n6621 ;
  assign n6623 = n6607 & ~n6622 ;
  assign n6624 = n6116 & n6167 ;
  assign n6625 = ~n6171 & ~n6624 ;
  assign n6626 = ~n6623 & n6625 ;
  assign n6627 = ~n6620 & n6626 ;
  assign n6628 = ~n3549 & n6178 ;
  assign n6629 = ~n3285 & n6628 ;
  assign n6630 = ~n2888 & ~n3304 ;
  assign n6631 = n6115 & n6630 ;
  assign n6632 = n6629 & n6631 ;
  assign n6633 = ~n6627 & n6632 ;
  assign n6634 = ~n3304 & ~n6174 ;
  assign n6635 = n6186 & ~n6634 ;
  assign n6636 = ~n2888 & ~n6635 ;
  assign n6637 = n6629 & n6636 ;
  assign n6638 = n6178 & ~n6189 ;
  assign n6639 = ~n6193 & ~n6638 ;
  assign n6640 = ~n6637 & n6639 ;
  assign n6641 = ~n6633 & n6640 ;
  assign n6642 = n3440 & n6641 ;
  assign n6643 = ~n3440 & ~n6641 ;
  assign n6644 = ~n6642 & ~n6643 ;
  assign n6645 = n6568 & ~n6644 ;
  assign n6646 = ~n6569 & ~n6645 ;
  assign n6647 = n6207 & ~n6646 ;
  assign n6651 = ~n3539 & n6350 ;
  assign n6652 = n6326 & n6651 ;
  assign n6653 = n3427 & ~n6652 ;
  assign n6654 = n6327 & n6651 ;
  assign n6655 = n6359 & ~n6654 ;
  assign n6656 = ~n6653 & n6655 ;
  assign n6657 = n3034 & ~n6312 ;
  assign n6658 = ~n6313 & ~n6657 ;
  assign n6659 = ~n2713 & ~n6658 ;
  assign n6660 = n2713 & n3527 ;
  assign n6661 = n4011 & ~n6660 ;
  assign n6662 = ~n6659 & n6661 ;
  assign n6663 = ~n6656 & ~n6662 ;
  assign n6664 = n6568 & ~n6663 ;
  assign n6648 = n6365 & n6568 ;
  assign n6649 = ~n4112 & ~n6648 ;
  assign n6650 = n3427 & ~n6649 ;
  assign n6665 = n6365 & ~n6568 ;
  assign n6666 = ~n6361 & ~n6665 ;
  assign n6667 = n6427 & ~n6568 ;
  assign n6668 = n6666 & ~n6667 ;
  assign n6669 = n3433 & ~n6668 ;
  assign n6670 = ~n6650 & ~n6669 ;
  assign n6671 = ~n6664 & n6670 ;
  assign n6672 = ~n6647 & n6671 ;
  assign n6673 = ~n6606 & n6672 ;
  assign n6674 = n6097 & ~n6673 ;
  assign n6675 = ~n6567 & ~n6674 ;
  assign n6676 = \P1_state_reg[0]/NET0131  & ~n6675 ;
  assign n6677 = \P1_reg3_reg[27]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6678 = n3433 & n4130 ;
  assign n6679 = ~n6677 & ~n6678 ;
  assign n6680 = ~n6676 & n6679 ;
  assign n6681 = \P1_reg1_reg[29]/NET0131  & ~n6078 ;
  assign n6682 = \P1_reg1_reg[29]/NET0131  & n6095 ;
  assign n6683 = ~n6107 & n6112 ;
  assign n6684 = \P1_reg1_reg[29]/NET0131  & ~n6683 ;
  assign n6685 = ~n6201 & n6683 ;
  assign n6686 = ~n6684 & ~n6685 ;
  assign n6687 = n6207 & ~n6686 ;
  assign n6688 = n6279 & n6683 ;
  assign n6689 = ~n6684 & ~n6688 ;
  assign n6690 = n6282 & ~n6689 ;
  assign n6691 = ~n6421 & n6683 ;
  assign n6692 = n4011 & ~n6683 ;
  assign n6693 = ~n3868 & n4110 ;
  assign n6694 = ~n6683 & n6693 ;
  assign n6695 = n6424 & ~n6694 ;
  assign n6696 = ~n6692 & n6695 ;
  assign n6697 = \P1_reg1_reg[29]/NET0131  & ~n6696 ;
  assign n6698 = ~n6691 & ~n6697 ;
  assign n6699 = ~n6690 & n6698 ;
  assign n6700 = ~n6687 & n6699 ;
  assign n6701 = n6097 & ~n6700 ;
  assign n6702 = ~n6682 & ~n6701 ;
  assign n6703 = \P1_state_reg[0]/NET0131  & ~n6702 ;
  assign n6704 = ~n6681 & ~n6703 ;
  assign n6705 = \P2_reg0_reg[29]/NET0131  & ~n5589 ;
  assign n6706 = n4211 & ~n4218 ;
  assign n6707 = \P2_reg0_reg[29]/NET0131  & ~n6706 ;
  assign n6708 = ~n5304 & n6706 ;
  assign n6709 = ~n6707 & ~n6708 ;
  assign n6710 = n5329 & ~n6709 ;
  assign n6711 = ~n5380 & n6706 ;
  assign n6712 = ~n6707 & ~n6711 ;
  assign n6713 = n5383 & ~n6712 ;
  assign n6714 = ~n6391 & n6706 ;
  assign n6715 = n5526 & ~n6706 ;
  assign n6716 = ~n6395 & ~n6706 ;
  assign n6717 = n6394 & ~n6716 ;
  assign n6718 = ~n6715 & n6717 ;
  assign n6719 = \P2_reg0_reg[29]/NET0131  & ~n6718 ;
  assign n6720 = ~n6714 & ~n6719 ;
  assign n6721 = ~n6713 & n6720 ;
  assign n6722 = ~n6710 & n6721 ;
  assign n6723 = n5583 & ~n6722 ;
  assign n6724 = \P2_reg0_reg[29]/NET0131  & n5585 ;
  assign n6725 = ~n6723 & ~n6724 ;
  assign n6726 = \P1_state_reg[0]/NET0131  & ~n6725 ;
  assign n6727 = ~n6705 & ~n6726 ;
  assign n6728 = \P2_reg2_reg[28]/NET0131  & ~n5589 ;
  assign n6729 = \P2_reg2_reg[28]/NET0131  & n5585 ;
  assign n6730 = \P2_reg2_reg[28]/NET0131  & ~n4219 ;
  assign n6731 = ~n5082 & ~n5108 ;
  assign n6732 = ~n5193 & n5243 ;
  assign n6733 = ~n5154 & ~n5247 ;
  assign n6734 = ~n5241 & ~n6733 ;
  assign n6735 = ~n6732 & ~n6734 ;
  assign n6736 = ~n5132 & ~n5219 ;
  assign n6737 = ~n6735 & n6736 ;
  assign n6738 = ~n5246 & ~n5255 ;
  assign n6739 = ~n5132 & ~n6738 ;
  assign n6740 = ~n6737 & ~n6739 ;
  assign n6741 = n6731 & ~n6740 ;
  assign n6742 = ~n5082 & n5254 ;
  assign n6743 = ~n5260 & ~n6742 ;
  assign n6744 = ~n6741 & n6743 ;
  assign n6745 = ~n5059 & ~n5265 ;
  assign n6746 = ~n4949 & ~n4999 ;
  assign n6747 = n6745 & n6746 ;
  assign n6748 = ~n6744 & n6747 ;
  assign n6749 = n5259 & ~n5265 ;
  assign n6750 = ~n5023 & ~n6749 ;
  assign n6751 = n6746 & ~n6750 ;
  assign n6752 = ~n4949 & n4998 ;
  assign n6753 = ~n5028 & ~n6752 ;
  assign n6754 = ~n6751 & n6753 ;
  assign n6755 = ~n6748 & n6754 ;
  assign n6756 = ~n4868 & ~n4974 ;
  assign n6757 = ~n4844 & ~n4919 ;
  assign n6758 = n6756 & n6757 ;
  assign n6759 = ~n4746 & ~n4815 ;
  assign n6760 = ~n4790 & ~n4893 ;
  assign n6761 = n6759 & n6760 ;
  assign n6762 = n6758 & n6761 ;
  assign n6763 = ~n6755 & n6762 ;
  assign n6764 = ~n5027 & ~n5272 ;
  assign n6765 = ~n4868 & ~n6764 ;
  assign n6766 = n6757 & n6765 ;
  assign n6767 = ~n5271 & ~n5277 ;
  assign n6768 = ~n4919 & ~n6767 ;
  assign n6769 = ~n6766 & ~n6768 ;
  assign n6770 = n6761 & ~n6769 ;
  assign n6771 = ~n5276 & ~n5283 ;
  assign n6772 = ~n4790 & ~n6771 ;
  assign n6773 = n6759 & n6772 ;
  assign n6774 = ~n4746 & n5282 ;
  assign n6775 = ~n5288 & ~n6774 ;
  assign n6776 = ~n6773 & n6775 ;
  assign n6777 = ~n6770 & n6776 ;
  assign n6778 = ~n6763 & n6777 ;
  assign n6779 = ~n4764 & ~n5294 ;
  assign n6780 = ~n4666 & ~n4686 ;
  assign n6781 = n6779 & n6780 ;
  assign n6782 = ~n4648 & n6781 ;
  assign n6783 = n4627 & n6782 ;
  assign n6784 = ~n6778 & n6783 ;
  assign n6785 = ~n4623 & ~n4708 ;
  assign n6786 = ~n4685 & ~n4709 ;
  assign n6787 = n5287 & ~n5294 ;
  assign n6788 = ~n4704 & ~n6787 ;
  assign n6789 = ~n4686 & ~n6788 ;
  assign n6790 = n6786 & ~n6789 ;
  assign n6791 = ~n4666 & ~n6790 ;
  assign n6792 = ~n4648 & n6791 ;
  assign n6793 = n6785 & ~n6792 ;
  assign n6794 = n4627 & ~n6793 ;
  assign n6795 = ~n4553 & n4604 ;
  assign n6796 = ~n4714 & ~n6795 ;
  assign n6797 = ~n6794 & n6796 ;
  assign n6798 = ~n6784 & n6797 ;
  assign n6799 = n5985 & n6798 ;
  assign n6800 = ~n5985 & ~n6798 ;
  assign n6801 = ~n6799 & ~n6800 ;
  assign n6802 = n4219 & ~n6801 ;
  assign n6803 = ~n6730 & ~n6802 ;
  assign n6804 = n5329 & ~n6803 ;
  assign n6805 = n5803 & ~n5827 ;
  assign n6806 = n5806 & n5835 ;
  assign n6807 = ~n6805 & n6806 ;
  assign n6808 = ~n5797 & n5835 ;
  assign n6809 = n5843 & ~n6808 ;
  assign n6810 = ~n6807 & n6809 ;
  assign n6811 = n5790 & n5832 ;
  assign n6812 = ~n6810 & n6811 ;
  assign n6813 = n5790 & ~n5850 ;
  assign n6814 = ~n5859 & ~n6813 ;
  assign n6815 = ~n6812 & n6814 ;
  assign n6816 = n5985 & ~n6815 ;
  assign n6817 = ~n5985 & n6815 ;
  assign n6818 = ~n6816 & ~n6817 ;
  assign n6819 = n4219 & ~n6818 ;
  assign n6820 = ~n6730 & ~n6819 ;
  assign n6821 = n5526 & ~n6820 ;
  assign n6822 = n4231 & ~n4552 ;
  assign n6823 = ~n4601 & n5372 ;
  assign n6824 = n5371 & n6823 ;
  assign n6825 = n4421 & ~n6824 ;
  assign n6826 = ~n4231 & ~n5375 ;
  assign n6827 = ~n6825 & n6826 ;
  assign n6828 = ~n6822 & ~n6827 ;
  assign n6829 = n5383 & ~n6828 ;
  assign n6830 = n4487 & n5565 ;
  assign n6831 = n4487 & ~n5554 ;
  assign n6832 = ~n5555 & ~n6831 ;
  assign n6833 = n5563 & n6832 ;
  assign n6834 = ~n6830 & ~n6833 ;
  assign n6835 = ~n6829 & n6834 ;
  assign n6836 = n4219 & ~n6835 ;
  assign n6837 = n4496 & n5574 ;
  assign n6838 = ~n4219 & ~n6395 ;
  assign n6839 = ~n5568 & ~n6838 ;
  assign n6840 = ~n4219 & n5383 ;
  assign n6841 = n6839 & ~n6840 ;
  assign n6842 = \P2_reg2_reg[28]/NET0131  & ~n6841 ;
  assign n6843 = ~n6837 & ~n6842 ;
  assign n6844 = ~n6836 & n6843 ;
  assign n6845 = ~n6821 & n6844 ;
  assign n6846 = ~n6804 & n6845 ;
  assign n6847 = n5583 & ~n6846 ;
  assign n6848 = ~n6729 & ~n6847 ;
  assign n6849 = \P1_state_reg[0]/NET0131  & ~n6848 ;
  assign n6850 = ~n6728 & ~n6849 ;
  assign n6851 = \P3_reg0_reg[27]/NET0131  & ~n2163 ;
  assign n6852 = n2163 & ~n2617 ;
  assign n6853 = ~n6851 & ~n6852 ;
  assign n6854 = n2234 & ~n6853 ;
  assign n6855 = \P3_reg0_reg[27]/NET0131  & ~n2236 ;
  assign n6856 = n2236 & ~n2575 ;
  assign n6857 = ~n6855 & ~n6856 ;
  assign n6858 = n737 & ~n6857 ;
  assign n6859 = n1436 & n2289 ;
  assign n6860 = \P3_reg0_reg[27]/NET0131  & ~n2287 ;
  assign n6865 = ~n6859 & ~n6860 ;
  assign n6866 = ~n6858 & n6865 ;
  assign n6867 = ~n6854 & n6866 ;
  assign n6861 = ~n2621 & ~n6855 ;
  assign n6862 = n2393 & ~n6861 ;
  assign n6863 = ~n2567 & ~n6851 ;
  assign n6864 = n2391 & ~n6863 ;
  assign n6868 = ~n6862 & ~n6864 ;
  assign n6869 = n6867 & n6868 ;
  assign n6870 = n2147 & ~n6869 ;
  assign n6871 = \P3_reg0_reg[27]/NET0131  & n2145 ;
  assign n6872 = ~n6870 & ~n6871 ;
  assign n6873 = \P1_state_reg[0]/NET0131  & ~n6872 ;
  assign n6874 = \P3_reg0_reg[27]/NET0131  & ~n2143 ;
  assign n6875 = ~n6873 & ~n6874 ;
  assign n6876 = \P3_reg0_reg[28]/NET0131  & ~n2143 ;
  assign n6877 = \P3_reg0_reg[28]/NET0131  & n2145 ;
  assign n6878 = \P3_reg0_reg[28]/NET0131  & ~n2236 ;
  assign n6879 = ~n2650 & ~n6878 ;
  assign n6880 = n2393 & ~n6879 ;
  assign n6882 = n2236 & ~n2436 ;
  assign n6883 = ~n6878 & ~n6882 ;
  assign n6884 = n737 & ~n6883 ;
  assign n6881 = \P3_reg0_reg[28]/NET0131  & ~n2287 ;
  assign n6885 = n1408 & n2289 ;
  assign n6892 = ~n6881 & ~n6885 ;
  assign n6893 = ~n6884 & n6892 ;
  assign n6894 = ~n6880 & n6893 ;
  assign n6886 = \P3_reg0_reg[28]/NET0131  & ~n2163 ;
  assign n6887 = ~n2638 & ~n6886 ;
  assign n6888 = n2391 & ~n6887 ;
  assign n6889 = n2163 & ~n2421 ;
  assign n6890 = ~n6886 & ~n6889 ;
  assign n6891 = n2234 & ~n6890 ;
  assign n6895 = ~n6888 & ~n6891 ;
  assign n6896 = n6894 & n6895 ;
  assign n6897 = n2147 & ~n6896 ;
  assign n6898 = ~n6877 & ~n6897 ;
  assign n6899 = \P1_state_reg[0]/NET0131  & ~n6898 ;
  assign n6900 = ~n6876 & ~n6899 ;
  assign n6901 = \P3_reg1_reg[28]/NET0131  & ~n2143 ;
  assign n6902 = \P3_reg1_reg[28]/NET0131  & n2145 ;
  assign n6903 = \P3_reg1_reg[28]/NET0131  & ~n2427 ;
  assign n6904 = ~n2515 & ~n6903 ;
  assign n6905 = n2425 & ~n6904 ;
  assign n6907 = n2427 & ~n2436 ;
  assign n6908 = ~n6903 & ~n6907 ;
  assign n6909 = n737 & ~n6908 ;
  assign n6906 = n1408 & n6451 ;
  assign n6910 = \P3_reg1_reg[28]/NET0131  & ~n6449 ;
  assign n6917 = ~n6906 & ~n6910 ;
  assign n6918 = ~n6909 & n6917 ;
  assign n6919 = ~n6905 & n6918 ;
  assign n6911 = \P3_reg1_reg[28]/NET0131  & ~n2408 ;
  assign n6912 = ~n2422 & ~n6911 ;
  assign n6913 = ~n2518 & ~n6912 ;
  assign n6914 = n2408 & ~n2511 ;
  assign n6915 = ~n6911 & ~n6914 ;
  assign n6916 = n714 & ~n6915 ;
  assign n6920 = ~n6913 & ~n6916 ;
  assign n6921 = n6919 & n6920 ;
  assign n6922 = n2147 & ~n6921 ;
  assign n6923 = ~n6902 & ~n6922 ;
  assign n6924 = \P1_state_reg[0]/NET0131  & ~n6923 ;
  assign n6925 = ~n6901 & ~n6924 ;
  assign n6926 = \P3_reg1_reg[27]/NET0131  & ~n2408 ;
  assign n6927 = ~n4136 & ~n6926 ;
  assign n6928 = ~n2518 & ~n6927 ;
  assign n6929 = \P3_reg1_reg[27]/NET0131  & ~n2427 ;
  assign n6930 = n2427 & ~n2575 ;
  assign n6931 = ~n6929 & ~n6930 ;
  assign n6932 = n737 & ~n6931 ;
  assign n6933 = \P3_reg1_reg[27]/NET0131  & ~n6449 ;
  assign n6934 = n1436 & n6451 ;
  assign n6940 = ~n6933 & ~n6934 ;
  assign n6941 = ~n6932 & n6940 ;
  assign n6942 = ~n6928 & n6941 ;
  assign n6935 = ~n4149 & ~n6929 ;
  assign n6936 = n2425 & ~n6935 ;
  assign n6937 = n2408 & ~n2566 ;
  assign n6938 = ~n6926 & ~n6937 ;
  assign n6939 = n714 & ~n6938 ;
  assign n6943 = ~n6936 & ~n6939 ;
  assign n6944 = n6942 & n6943 ;
  assign n6945 = n2147 & ~n6944 ;
  assign n6946 = \P3_reg1_reg[27]/NET0131  & n2145 ;
  assign n6947 = ~n6945 & ~n6946 ;
  assign n6948 = \P1_state_reg[0]/NET0131  & ~n6947 ;
  assign n6949 = \P3_reg1_reg[27]/NET0131  & ~n2143 ;
  assign n6950 = ~n6948 & ~n6949 ;
  assign n6953 = n3544 & n6095 ;
  assign n6954 = n3544 & ~n6568 ;
  assign n6968 = ~n3304 & n3599 ;
  assign n6969 = ~n3305 & ~n6968 ;
  assign n6970 = n6181 & ~n6969 ;
  assign n6971 = n2889 & ~n3285 ;
  assign n6972 = ~n3284 & ~n6971 ;
  assign n6973 = ~n6970 & n6972 ;
  assign n6974 = ~n3304 & ~n3598 ;
  assign n6975 = n6181 & n6974 ;
  assign n6983 = ~n3578 & ~n3747 ;
  assign n6984 = ~n6130 & ~n6133 ;
  assign n6985 = n6138 & n6984 ;
  assign n6986 = ~n6132 & ~n6143 ;
  assign n6987 = ~n6130 & ~n6986 ;
  assign n6988 = ~n6985 & ~n6987 ;
  assign n6989 = ~n3139 & ~n6129 ;
  assign n6990 = ~n6988 & n6989 ;
  assign n6991 = n6983 & n6990 ;
  assign n6992 = ~n3139 & n6142 ;
  assign n6993 = ~n3138 & ~n6992 ;
  assign n6994 = n6983 & ~n6993 ;
  assign n6995 = ~n3579 & ~n3748 ;
  assign n6996 = ~n3578 & ~n6995 ;
  assign n6997 = ~n6994 & ~n6996 ;
  assign n6998 = ~n6991 & n6997 ;
  assign n6999 = ~n3256 & ~n3678 ;
  assign n7000 = ~n3331 & ~n3823 ;
  assign n7001 = n6999 & n7000 ;
  assign n7002 = ~n6998 & n7001 ;
  assign n6976 = ~n2953 & ~n3110 ;
  assign n7003 = ~n3083 & ~n3205 ;
  assign n7004 = n6976 & n7003 ;
  assign n7005 = ~n3230 & ~n3624 ;
  assign n7006 = ~n3355 & ~n3651 ;
  assign n7007 = n7005 & n7006 ;
  assign n7008 = n7004 & n7007 ;
  assign n7009 = n7002 & n7008 ;
  assign n6977 = ~n3083 & n3204 ;
  assign n6978 = ~n3082 & ~n6977 ;
  assign n6979 = n6976 & ~n6978 ;
  assign n6980 = ~n2953 & n3111 ;
  assign n6981 = ~n2954 & ~n6980 ;
  assign n6982 = ~n6979 & n6981 ;
  assign n7010 = ~n3356 & ~n3652 ;
  assign n7011 = ~n3355 & ~n7010 ;
  assign n7012 = n7005 & n7011 ;
  assign n7013 = ~n3231 & ~n3625 ;
  assign n7014 = ~n3624 & ~n7013 ;
  assign n7015 = ~n7012 & ~n7014 ;
  assign n7016 = ~n3331 & n3824 ;
  assign n7017 = ~n3330 & ~n7016 ;
  assign n7018 = n6999 & ~n7017 ;
  assign n7019 = ~n3256 & n3679 ;
  assign n7020 = ~n3257 & ~n7019 ;
  assign n7021 = ~n7018 & n7020 ;
  assign n7022 = n7007 & ~n7021 ;
  assign n7023 = n7015 & ~n7022 ;
  assign n7024 = n7004 & ~n7023 ;
  assign n7025 = n6982 & ~n7024 ;
  assign n7026 = ~n7009 & n7025 ;
  assign n7027 = n6975 & ~n7026 ;
  assign n7028 = n6973 & ~n7027 ;
  assign n7029 = n3551 & n7028 ;
  assign n7030 = ~n3551 & ~n7028 ;
  assign n7031 = ~n7029 & ~n7030 ;
  assign n7032 = n6568 & ~n7031 ;
  assign n7033 = ~n6954 & ~n7032 ;
  assign n7034 = n6207 & ~n7033 ;
  assign n6958 = n4035 & n4054 ;
  assign n6959 = n4080 & n6958 ;
  assign n6955 = n4034 & ~n4082 ;
  assign n6956 = n4033 & ~n6955 ;
  assign n6957 = n4027 & ~n6956 ;
  assign n6960 = n4026 & ~n6957 ;
  assign n6961 = ~n6959 & n6960 ;
  assign n6962 = n3551 & ~n6961 ;
  assign n6963 = ~n3551 & n6961 ;
  assign n6964 = ~n6962 & ~n6963 ;
  assign n6965 = n6568 & ~n6964 ;
  assign n6966 = ~n6954 & ~n6965 ;
  assign n6967 = n6282 & ~n6966 ;
  assign n7038 = n6303 & n6309 ;
  assign n7039 = ~n3176 & n7038 ;
  assign n7040 = n3176 & ~n7038 ;
  assign n7041 = ~n7039 & ~n7040 ;
  assign n7042 = ~n2713 & ~n7041 ;
  assign n7043 = n2713 & n3283 ;
  assign n7044 = ~n7042 & ~n7043 ;
  assign n7045 = n6568 & n7044 ;
  assign n7046 = ~n6954 & ~n7045 ;
  assign n7047 = n4011 & ~n7046 ;
  assign n7048 = n3539 & ~n6350 ;
  assign n7049 = ~n6651 & ~n7048 ;
  assign n7050 = n6359 & n7049 ;
  assign n7051 = n6568 & n7050 ;
  assign n7035 = n6359 & ~n6568 ;
  assign n7036 = n6666 & ~n7035 ;
  assign n7037 = n3544 & ~n7036 ;
  assign n7052 = n3539 & ~n6649 ;
  assign n7053 = ~n7037 & ~n7052 ;
  assign n7054 = ~n7051 & n7053 ;
  assign n7055 = ~n7047 & n7054 ;
  assign n7056 = ~n6967 & n7055 ;
  assign n7057 = ~n7034 & n7056 ;
  assign n7058 = n6097 & ~n7057 ;
  assign n7059 = ~n6953 & ~n7058 ;
  assign n7060 = \P1_state_reg[0]/NET0131  & ~n7059 ;
  assign n6951 = \P1_reg3_reg[24]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6952 = n3544 & n4130 ;
  assign n7061 = ~n6951 & ~n6952 ;
  assign n7062 = ~n7060 & n7061 ;
  assign n7065 = n3172 & n6095 ;
  assign n7066 = n3172 & ~n6568 ;
  assign n7083 = n6121 & n6160 ;
  assign n7084 = n6120 & ~n6128 ;
  assign n7085 = n6168 & ~n7084 ;
  assign n7086 = n6117 & ~n7085 ;
  assign n7087 = n6175 & ~n7086 ;
  assign n7088 = ~n7083 & n7087 ;
  assign n7089 = n6183 & ~n7088 ;
  assign n7090 = n6190 & ~n7089 ;
  assign n7091 = n3179 & n7090 ;
  assign n7092 = ~n3179 & ~n7090 ;
  assign n7093 = ~n7091 & ~n7092 ;
  assign n7094 = n6568 & ~n7093 ;
  assign n7095 = ~n7066 & ~n7094 ;
  assign n7096 = n6207 & ~n7095 ;
  assign n7067 = ~n6222 & n6228 ;
  assign n7068 = n6211 & ~n7067 ;
  assign n7069 = n6242 & n7068 ;
  assign n7070 = ~n6233 & n6241 ;
  assign n7071 = n6248 & ~n7070 ;
  assign n7072 = n6238 & ~n7071 ;
  assign n7073 = n6253 & ~n7072 ;
  assign n7074 = ~n7069 & n7073 ;
  assign n7075 = n6258 & ~n7074 ;
  assign n7076 = n6268 & ~n7075 ;
  assign n7077 = n3179 & ~n7076 ;
  assign n7078 = ~n3179 & n7076 ;
  assign n7079 = ~n7077 & ~n7078 ;
  assign n7080 = n6568 & ~n7079 ;
  assign n7081 = ~n7066 & ~n7080 ;
  assign n7082 = n6282 & ~n7081 ;
  assign n7098 = n3527 & ~n7039 ;
  assign n7099 = n6304 & n7038 ;
  assign n7100 = ~n7098 & ~n7099 ;
  assign n7101 = ~n2713 & ~n7100 ;
  assign n7102 = n2713 & n3548 ;
  assign n7103 = ~n7101 & ~n7102 ;
  assign n7104 = n6568 & n7103 ;
  assign n7105 = ~n7066 & ~n7104 ;
  assign n7106 = n4011 & ~n7105 ;
  assign n7107 = n3165 & ~n6651 ;
  assign n7108 = ~n3165 & n6651 ;
  assign n7109 = ~n7107 & ~n7108 ;
  assign n7110 = n6568 & n7109 ;
  assign n7111 = ~n7066 & ~n7110 ;
  assign n7112 = n6359 & ~n7111 ;
  assign n7097 = n3172 & ~n6666 ;
  assign n7113 = n3165 & ~n6649 ;
  assign n7114 = ~n7097 & ~n7113 ;
  assign n7115 = ~n7112 & n7114 ;
  assign n7116 = ~n7106 & n7115 ;
  assign n7117 = ~n7082 & n7116 ;
  assign n7118 = ~n7096 & n7117 ;
  assign n7119 = n6097 & ~n7118 ;
  assign n7120 = ~n7065 & ~n7119 ;
  assign n7121 = \P1_state_reg[0]/NET0131  & ~n7120 ;
  assign n7063 = \P1_reg3_reg[25]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7064 = n3172 & n4130 ;
  assign n7122 = ~n7063 & ~n7064 ;
  assign n7123 = ~n7121 & n7122 ;
  assign n7124 = n3523 & n6095 ;
  assign n7125 = n3523 & ~n6568 ;
  assign n7126 = n3913 & ~n4045 ;
  assign n7127 = ~n4048 & ~n7126 ;
  assign n7128 = n3893 & n3911 ;
  assign n7129 = ~n7127 & n7128 ;
  assign n7130 = n3893 & n4050 ;
  assign n7131 = ~n4036 & ~n7130 ;
  assign n7132 = ~n7129 & n7131 ;
  assign n7133 = n3890 & n3901 ;
  assign n7134 = ~n7132 & n7133 ;
  assign n7135 = n3901 & ~n4039 ;
  assign n7136 = n3880 & ~n7135 ;
  assign n7137 = ~n7134 & n7136 ;
  assign n7138 = n3875 & n3972 ;
  assign n7139 = ~n7137 & n7138 ;
  assign n7140 = ~n3885 & n3972 ;
  assign n7141 = ~n4029 & ~n7140 ;
  assign n7142 = ~n7139 & n7141 ;
  assign n7143 = n3959 & n3991 ;
  assign n7144 = n3962 & n3969 ;
  assign n7145 = n7143 & n7144 ;
  assign n7146 = ~n7142 & n7145 ;
  assign n7148 = n3962 & ~n4032 ;
  assign n7149 = ~n4023 & ~n7148 ;
  assign n7150 = n7143 & ~n7149 ;
  assign n7147 = n3991 & n4025 ;
  assign n7151 = ~n4017 & ~n7147 ;
  assign n7152 = ~n7150 & n7151 ;
  assign n7153 = ~n7146 & n7152 ;
  assign n7154 = n3530 & ~n7153 ;
  assign n7155 = ~n3530 & n7153 ;
  assign n7156 = ~n7154 & ~n7155 ;
  assign n7157 = n6568 & ~n7156 ;
  assign n7158 = ~n7125 & ~n7157 ;
  assign n7159 = n6282 & ~n7158 ;
  assign n7160 = n6974 & ~n6981 ;
  assign n7161 = n6969 & ~n7160 ;
  assign n7162 = n6182 & ~n7161 ;
  assign n7163 = ~n3178 & ~n3550 ;
  assign n7164 = ~n3549 & ~n6972 ;
  assign n7165 = n7163 & ~n7164 ;
  assign n7166 = ~n7162 & n7165 ;
  assign n7167 = ~n3177 & ~n7166 ;
  assign n7168 = n7003 & n7005 ;
  assign n7169 = ~n6990 & n6993 ;
  assign n7170 = n6983 & n7000 ;
  assign n7171 = ~n7169 & n7170 ;
  assign n7172 = n6996 & n7000 ;
  assign n7173 = n7017 & ~n7172 ;
  assign n7174 = ~n7171 & n7173 ;
  assign n7175 = n6999 & n7006 ;
  assign n7176 = ~n7174 & n7175 ;
  assign n7177 = n7168 & n7176 ;
  assign n7178 = n7006 & ~n7020 ;
  assign n7179 = ~n7011 & ~n7178 ;
  assign n7180 = n7168 & ~n7179 ;
  assign n7181 = n7003 & n7014 ;
  assign n7182 = n6978 & ~n7181 ;
  assign n7183 = ~n7180 & n7182 ;
  assign n7184 = ~n7177 & n7183 ;
  assign n7185 = n6974 & n6976 ;
  assign n7186 = ~n3177 & n7185 ;
  assign n7187 = n6182 & n7186 ;
  assign n7188 = ~n7184 & n7187 ;
  assign n7189 = ~n7167 & ~n7188 ;
  assign n7190 = n3530 & n7189 ;
  assign n7191 = ~n3530 & ~n7189 ;
  assign n7192 = ~n7190 & ~n7191 ;
  assign n7193 = n6568 & ~n7192 ;
  assign n7194 = ~n7125 & ~n7193 ;
  assign n7195 = n6207 & ~n7194 ;
  assign n7196 = n2713 & ~n3176 ;
  assign n7197 = n3437 & ~n7099 ;
  assign n7198 = ~n2713 & ~n6312 ;
  assign n7199 = ~n7197 & n7198 ;
  assign n7200 = ~n7196 & ~n7199 ;
  assign n7201 = n4011 & ~n7200 ;
  assign n7202 = n3518 & ~n7108 ;
  assign n7203 = ~n6652 & ~n7202 ;
  assign n7204 = n6359 & n7203 ;
  assign n7205 = ~n7201 & ~n7204 ;
  assign n7206 = n6568 & ~n7205 ;
  assign n7207 = n3523 & ~n6668 ;
  assign n7208 = n3518 & ~n6649 ;
  assign n7209 = ~n7207 & ~n7208 ;
  assign n7210 = ~n7206 & n7209 ;
  assign n7211 = ~n7195 & n7210 ;
  assign n7212 = ~n7159 & n7211 ;
  assign n7213 = n6097 & ~n7212 ;
  assign n7214 = ~n7124 & ~n7213 ;
  assign n7215 = \P1_state_reg[0]/NET0131  & ~n7214 ;
  assign n7216 = \P1_reg3_reg[26]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7217 = n3523 & n4130 ;
  assign n7218 = ~n7216 & ~n7217 ;
  assign n7219 = ~n7215 & n7218 ;
  assign n7220 = \P3_reg2_reg[19]/NET0131  & ~n2143 ;
  assign n7221 = \P3_reg2_reg[19]/NET0131  & n2145 ;
  assign n7229 = \P3_reg2_reg[19]/NET0131  & ~n2427 ;
  assign n7230 = n2427 & n6552 ;
  assign n7231 = ~n7229 & ~n7230 ;
  assign n7232 = ~n2518 & ~n7231 ;
  assign n7222 = \P3_reg2_reg[19]/NET0131  & ~n2408 ;
  assign n7226 = n2408 & n6552 ;
  assign n7227 = ~n7222 & ~n7226 ;
  assign n7228 = n2425 & ~n7227 ;
  assign n7238 = ~n1110 & n2441 ;
  assign n7236 = \P3_reg2_reg[19]/NET0131  & ~n2429 ;
  assign n7237 = ~n1090 & n2283 ;
  assign n7239 = ~n7236 & ~n7237 ;
  assign n7240 = ~n7238 & n7239 ;
  assign n7241 = ~n7228 & n7240 ;
  assign n7242 = ~n7232 & n7241 ;
  assign n7223 = n2408 & ~n6546 ;
  assign n7224 = ~n7222 & ~n7223 ;
  assign n7225 = n737 & ~n7224 ;
  assign n7233 = n2427 & ~n6531 ;
  assign n7234 = ~n7229 & ~n7233 ;
  assign n7235 = n714 & ~n7234 ;
  assign n7243 = ~n7225 & ~n7235 ;
  assign n7244 = n7242 & n7243 ;
  assign n7245 = n2147 & ~n7244 ;
  assign n7246 = ~n7221 & ~n7245 ;
  assign n7247 = \P1_state_reg[0]/NET0131  & ~n7246 ;
  assign n7248 = ~n7220 & ~n7247 ;
  assign n7249 = \P3_reg2_reg[20]/NET0131  & ~n2143 ;
  assign n7250 = \P3_reg2_reg[20]/NET0131  & n2145 ;
  assign n7253 = \P3_reg2_reg[20]/NET0131  & ~n2427 ;
  assign n7254 = n2095 & n2489 ;
  assign n7255 = ~n2095 & ~n2489 ;
  assign n7256 = ~n7254 & ~n7255 ;
  assign n7257 = n2427 & ~n7256 ;
  assign n7258 = ~n7253 & ~n7257 ;
  assign n7259 = n714 & ~n7258 ;
  assign n7251 = n1063 & n2285 ;
  assign n7252 = n2427 & n7251 ;
  assign n7278 = ~n1068 & n2283 ;
  assign n7279 = \P3_reg2_reg[20]/NET0131  & ~n2429 ;
  assign n7280 = ~n7278 & ~n7279 ;
  assign n7281 = ~n7252 & n7280 ;
  assign n7282 = ~n7259 & n7281 ;
  assign n7269 = n2095 & ~n2413 ;
  assign n7270 = ~n2095 & n2413 ;
  assign n7271 = ~n7269 & ~n7270 ;
  assign n7275 = n2427 & ~n7271 ;
  assign n7276 = ~n7253 & ~n7275 ;
  assign n7277 = ~n2518 & ~n7276 ;
  assign n7260 = \P3_reg2_reg[20]/NET0131  & ~n2408 ;
  assign n7261 = ~n1095 & n2239 ;
  assign n7262 = n1038 & ~n6541 ;
  assign n7263 = ~n2239 & ~n2264 ;
  assign n7264 = ~n7262 & n7263 ;
  assign n7265 = ~n7261 & ~n7264 ;
  assign n7266 = n2408 & ~n7265 ;
  assign n7267 = ~n7260 & ~n7266 ;
  assign n7268 = n737 & ~n7267 ;
  assign n7272 = n2408 & ~n7271 ;
  assign n7273 = ~n7260 & ~n7272 ;
  assign n7274 = n2425 & ~n7273 ;
  assign n7283 = ~n7268 & ~n7274 ;
  assign n7284 = ~n7277 & n7283 ;
  assign n7285 = n7282 & n7284 ;
  assign n7286 = n2147 & ~n7285 ;
  assign n7287 = ~n7250 & ~n7286 ;
  assign n7288 = \P1_state_reg[0]/NET0131  & ~n7287 ;
  assign n7289 = ~n7249 & ~n7288 ;
  assign n7292 = ~n1034 & n2145 ;
  assign n7294 = ~n1034 & ~n2163 ;
  assign n7295 = n2087 & n2362 ;
  assign n7296 = ~n2087 & ~n2362 ;
  assign n7297 = ~n7295 & ~n7296 ;
  assign n7298 = n2163 & ~n7297 ;
  assign n7299 = ~n7294 & ~n7298 ;
  assign n7300 = n2393 & ~n7299 ;
  assign n7311 = n1000 & ~n2264 ;
  assign n7312 = ~n2239 & ~n5615 ;
  assign n7313 = ~n7311 & n7312 ;
  assign n7314 = ~n1072 & n2239 ;
  assign n7315 = ~n7313 & ~n7314 ;
  assign n7316 = n2163 & ~n7315 ;
  assign n7317 = ~n7294 & ~n7316 ;
  assign n7318 = n737 & ~n7317 ;
  assign n7293 = n1029 & n2580 ;
  assign n7319 = ~n1034 & ~n2583 ;
  assign n7320 = ~n7293 & ~n7319 ;
  assign n7321 = ~n7318 & n7320 ;
  assign n7322 = ~n7300 & n7321 ;
  assign n7301 = ~n1034 & ~n2236 ;
  assign n7302 = n2236 & ~n7297 ;
  assign n7303 = ~n7301 & ~n7302 ;
  assign n7304 = n2391 & ~n7303 ;
  assign n7305 = n2087 & ~n2209 ;
  assign n7306 = ~n2087 & n2209 ;
  assign n7307 = ~n7305 & ~n7306 ;
  assign n7308 = n2236 & ~n7307 ;
  assign n7309 = ~n7301 & ~n7308 ;
  assign n7310 = n2234 & ~n7309 ;
  assign n7323 = ~n7304 & ~n7310 ;
  assign n7324 = n7322 & n7323 ;
  assign n7325 = n2147 & ~n7324 ;
  assign n7326 = ~n7292 & ~n7325 ;
  assign n7327 = \P1_state_reg[0]/NET0131  & ~n7326 ;
  assign n7290 = n765 & ~n1034 ;
  assign n7291 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[21]/NET0131  ;
  assign n7328 = ~n7290 & ~n7291 ;
  assign n7329 = ~n7327 & n7328 ;
  assign n7332 = ~n996 & n2145 ;
  assign n7333 = ~n996 & ~n2236 ;
  assign n7336 = ~n5740 & ~n5745 ;
  assign n7334 = ~n2085 & n2351 ;
  assign n7337 = n5741 & n7334 ;
  assign n7338 = ~n7336 & n7337 ;
  assign n7335 = ~n5748 & n7334 ;
  assign n7339 = n5732 & ~n7335 ;
  assign n7340 = ~n7338 & n7339 ;
  assign n7341 = n2045 & n7340 ;
  assign n7342 = ~n2045 & ~n7340 ;
  assign n7343 = ~n7341 & ~n7342 ;
  assign n7344 = n2236 & ~n7343 ;
  assign n7345 = ~n7333 & ~n7344 ;
  assign n7346 = n2391 & ~n7345 ;
  assign n7347 = ~n996 & ~n2163 ;
  assign n7359 = n933 & ~n5615 ;
  assign n7360 = ~n2239 & ~n5616 ;
  assign n7361 = ~n7359 & n7360 ;
  assign n7362 = ~n1038 & n2239 ;
  assign n7363 = ~n7361 & ~n7362 ;
  assign n7364 = n2163 & ~n7363 ;
  assign n7365 = ~n7347 & ~n7364 ;
  assign n7366 = n737 & ~n7365 ;
  assign n7351 = ~n996 & ~n2583 ;
  assign n7367 = n991 & n2580 ;
  assign n7368 = ~n7351 & ~n7367 ;
  assign n7369 = ~n7366 & n7368 ;
  assign n7370 = ~n7346 & n7369 ;
  assign n7348 = n2163 & ~n7343 ;
  assign n7349 = ~n7347 & ~n7348 ;
  assign n7350 = n2393 & ~n7349 ;
  assign n7352 = ~n5715 & n5718 ;
  assign n7353 = n2045 & ~n7352 ;
  assign n7354 = ~n2045 & n7352 ;
  assign n7355 = ~n7353 & ~n7354 ;
  assign n7356 = n2236 & ~n7355 ;
  assign n7357 = ~n7333 & ~n7356 ;
  assign n7358 = n2234 & ~n7357 ;
  assign n7371 = ~n7350 & ~n7358 ;
  assign n7372 = n7370 & n7371 ;
  assign n7373 = n2147 & ~n7372 ;
  assign n7374 = ~n7332 & ~n7373 ;
  assign n7375 = \P1_state_reg[0]/NET0131  & ~n7374 ;
  assign n7330 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[22]/NET0131  ;
  assign n7331 = n765 & ~n996 ;
  assign n7376 = ~n7330 & ~n7331 ;
  assign n7377 = ~n7375 & n7376 ;
  assign n7380 = ~n929 & n2145 ;
  assign n7381 = ~n929 & ~n2236 ;
  assign n7402 = ~n2605 & n2608 ;
  assign n7403 = n2090 & ~n7402 ;
  assign n7404 = ~n2090 & n7402 ;
  assign n7405 = ~n7403 & ~n7404 ;
  assign n7406 = n2236 & ~n7405 ;
  assign n7407 = ~n7381 & ~n7406 ;
  assign n7408 = n2234 & ~n7407 ;
  assign n7390 = ~n929 & ~n2163 ;
  assign n7394 = n1236 & ~n5616 ;
  assign n7395 = ~n2239 & ~n5617 ;
  assign n7396 = ~n7394 & n7395 ;
  assign n7397 = ~n1000 & n2239 ;
  assign n7398 = ~n7396 & ~n7397 ;
  assign n7399 = n2163 & ~n7398 ;
  assign n7400 = ~n7390 & ~n7399 ;
  assign n7401 = n737 & ~n7400 ;
  assign n7409 = n886 & n2580 ;
  assign n7410 = ~n929 & ~n2583 ;
  assign n7411 = ~n7409 & ~n7410 ;
  assign n7412 = ~n7401 & n7411 ;
  assign n7413 = ~n7408 & n7412 ;
  assign n7382 = ~n2549 & n2551 ;
  assign n7383 = ~n2558 & ~n7382 ;
  assign n7384 = n2090 & n7383 ;
  assign n7385 = ~n2090 & ~n7383 ;
  assign n7386 = ~n7384 & ~n7385 ;
  assign n7387 = n2236 & ~n7386 ;
  assign n7388 = ~n7381 & ~n7387 ;
  assign n7389 = n2391 & ~n7388 ;
  assign n7391 = n2163 & ~n7386 ;
  assign n7392 = ~n7390 & ~n7391 ;
  assign n7393 = n2393 & ~n7392 ;
  assign n7414 = ~n7389 & ~n7393 ;
  assign n7415 = n7413 & n7414 ;
  assign n7416 = n2147 & ~n7415 ;
  assign n7417 = ~n7380 & ~n7416 ;
  assign n7418 = \P1_state_reg[0]/NET0131  & ~n7417 ;
  assign n7378 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[23]/NET0131  ;
  assign n7379 = n765 & ~n929 ;
  assign n7419 = ~n7378 & ~n7379 ;
  assign n7420 = ~n7418 & n7419 ;
  assign n7423 = ~n1068 & n2145 ;
  assign n7425 = ~n1068 & ~n2236 ;
  assign n7426 = n2236 & ~n7271 ;
  assign n7427 = ~n7425 & ~n7426 ;
  assign n7428 = n2234 & ~n7427 ;
  assign n7424 = n1063 & n2580 ;
  assign n7439 = ~n1068 & ~n2583 ;
  assign n7440 = ~n7424 & ~n7439 ;
  assign n7441 = ~n7428 & n7440 ;
  assign n7429 = ~n1068 & ~n2163 ;
  assign n7436 = n2163 & ~n7256 ;
  assign n7437 = ~n7429 & ~n7436 ;
  assign n7438 = n2393 & ~n7437 ;
  assign n7430 = n2163 & ~n7265 ;
  assign n7431 = ~n7429 & ~n7430 ;
  assign n7432 = n737 & ~n7431 ;
  assign n7433 = n2236 & ~n7256 ;
  assign n7434 = ~n7425 & ~n7433 ;
  assign n7435 = n2391 & ~n7434 ;
  assign n7442 = ~n7432 & ~n7435 ;
  assign n7443 = ~n7438 & n7442 ;
  assign n7444 = n7441 & n7443 ;
  assign n7445 = n2147 & ~n7444 ;
  assign n7446 = ~n7423 & ~n7445 ;
  assign n7447 = \P1_state_reg[0]/NET0131  & ~n7446 ;
  assign n7421 = n765 & ~n1068 ;
  assign n7422 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[20]/NET0131  ;
  assign n7448 = ~n7421 & ~n7422 ;
  assign n7449 = ~n7447 & n7448 ;
  assign n7452 = n4618 & n5585 ;
  assign n7453 = ~n4211 & n4218 ;
  assign n7454 = n4618 & ~n7453 ;
  assign n7455 = n4922 & n5268 ;
  assign n7456 = n4921 & ~n5031 ;
  assign n7457 = n5280 & ~n7456 ;
  assign n7458 = n4817 & ~n7457 ;
  assign n7459 = n5291 & ~n7458 ;
  assign n7460 = ~n7455 & n7459 ;
  assign n7461 = n5296 & ~n7460 ;
  assign n7462 = n4712 & ~n7461 ;
  assign n7463 = n5998 & n7462 ;
  assign n7464 = ~n5998 & ~n7462 ;
  assign n7465 = ~n7463 & ~n7464 ;
  assign n7466 = n7453 & ~n7465 ;
  assign n7467 = ~n7454 & ~n7466 ;
  assign n7468 = n5329 & ~n7467 ;
  assign n7486 = n4601 & ~n5371 ;
  assign n7487 = ~n4601 & n5371 ;
  assign n7488 = ~n7486 & ~n7487 ;
  assign n7489 = ~n4231 & ~n7488 ;
  assign n7490 = n4231 & n4647 ;
  assign n7491 = ~n7489 & ~n7490 ;
  assign n7492 = n7453 & n7491 ;
  assign n7493 = ~n7454 & ~n7492 ;
  assign n7494 = n5383 & ~n7493 ;
  assign n7472 = n5399 & n5454 ;
  assign n7469 = n5398 & n5412 ;
  assign n7470 = n5465 & ~n7469 ;
  assign n7471 = n5391 & ~n7470 ;
  assign n7473 = n5476 & ~n7471 ;
  assign n7474 = ~n7472 & n7473 ;
  assign n7475 = n5485 & ~n7474 ;
  assign n7476 = n5504 & ~n7475 ;
  assign n7477 = n5998 & ~n7476 ;
  assign n7478 = ~n5998 & n7476 ;
  assign n7479 = ~n7477 & ~n7478 ;
  assign n7480 = n7453 & ~n7479 ;
  assign n7481 = ~n7454 & ~n7480 ;
  assign n7482 = n5526 & ~n7481 ;
  assign n7495 = ~n4694 & n5547 ;
  assign n7496 = ~n4675 & n7495 ;
  assign n7497 = n5548 & n7496 ;
  assign n7498 = n4613 & ~n7497 ;
  assign n7499 = n5547 & n5551 ;
  assign n7500 = ~n7498 & ~n7499 ;
  assign n7501 = n5563 & n7500 ;
  assign n7502 = n7453 & n7501 ;
  assign n7483 = ~n6395 & ~n7453 ;
  assign n7484 = ~n5568 & ~n7483 ;
  assign n7485 = n4618 & ~n7484 ;
  assign n7503 = n5565 & n7453 ;
  assign n7504 = ~n5574 & ~n7503 ;
  assign n7505 = n4613 & ~n7504 ;
  assign n7506 = ~n7485 & ~n7505 ;
  assign n7507 = ~n7502 & n7506 ;
  assign n7508 = ~n7482 & n7507 ;
  assign n7509 = ~n7494 & n7508 ;
  assign n7510 = ~n7468 & n7509 ;
  assign n7511 = n5583 & ~n7510 ;
  assign n7512 = ~n7452 & ~n7511 ;
  assign n7513 = \P1_state_reg[0]/NET0131  & ~n7512 ;
  assign n7450 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[25]/NET0131  ;
  assign n7451 = n4618 & n5786 ;
  assign n7514 = ~n7450 & ~n7451 ;
  assign n7515 = ~n7513 & n7514 ;
  assign n7516 = n4548 & n5585 ;
  assign n7517 = n4548 & ~n7453 ;
  assign n7518 = ~n5430 & n5436 ;
  assign n7519 = ~n5442 & ~n7518 ;
  assign n7520 = ~n5405 & ~n5451 ;
  assign n7521 = n5433 & n7520 ;
  assign n7522 = ~n7519 & n7521 ;
  assign n7523 = n5447 & n7520 ;
  assign n7524 = ~n5409 & ~n7523 ;
  assign n7525 = ~n7522 & n7524 ;
  assign n7526 = ~n5404 & n5805 ;
  assign n7527 = ~n7525 & n7526 ;
  assign n7528 = ~n5403 & n5805 ;
  assign n7529 = ~n5935 & ~n7528 ;
  assign n7530 = ~n7527 & n7529 ;
  assign n7531 = n5390 & n5396 ;
  assign n7532 = ~n7530 & n7531 ;
  assign n7533 = n5390 & n5460 ;
  assign n7534 = ~n5470 & ~n7533 ;
  assign n7535 = ~n7532 & n7534 ;
  assign n7536 = n5387 & n5481 ;
  assign n7537 = n5484 & n5488 ;
  assign n7538 = n7536 & n7537 ;
  assign n7539 = ~n7535 & n7538 ;
  assign n7541 = n5475 & n5481 ;
  assign n7542 = ~n5498 & ~n7541 ;
  assign n7543 = n7537 & ~n7542 ;
  assign n7540 = n5488 & n5503 ;
  assign n7544 = ~n5509 & ~n7540 ;
  assign n7545 = ~n7543 & n7544 ;
  assign n7546 = ~n7539 & n7545 ;
  assign n7547 = n5982 & ~n7546 ;
  assign n7548 = ~n5982 & n7546 ;
  assign n7549 = ~n7547 & ~n7548 ;
  assign n7550 = n7453 & ~n7549 ;
  assign n7551 = ~n7517 & ~n7550 ;
  assign n7552 = n5526 & ~n7551 ;
  assign n7553 = ~n5252 & ~n5257 ;
  assign n7554 = n5083 & n5266 ;
  assign n7555 = ~n7553 & n7554 ;
  assign n7556 = ~n5262 & n5266 ;
  assign n7557 = n5025 & ~n7556 ;
  assign n7558 = ~n7555 & n7557 ;
  assign n7559 = n4869 & n4975 ;
  assign n7560 = n4816 & n4920 ;
  assign n7561 = n7559 & n7560 ;
  assign n7562 = ~n7558 & n7561 ;
  assign n7563 = n4869 & n5030 ;
  assign n7564 = ~n5274 & ~n7563 ;
  assign n7565 = n7560 & ~n7564 ;
  assign n7566 = n4816 & n5279 ;
  assign n7567 = ~n5285 & ~n7566 ;
  assign n7568 = ~n7565 & n7567 ;
  assign n7569 = ~n7562 & n7568 ;
  assign n7570 = ~n4626 & n4667 ;
  assign n7571 = n4765 & n5295 ;
  assign n7572 = ~n4602 & n7571 ;
  assign n7573 = n7570 & n7572 ;
  assign n7574 = ~n7569 & n7573 ;
  assign n7575 = ~n5290 & n5295 ;
  assign n7576 = n4706 & ~n7575 ;
  assign n7577 = n7570 & ~n7576 ;
  assign n7578 = ~n4626 & ~n4711 ;
  assign n7579 = n4624 & ~n7578 ;
  assign n7580 = ~n7577 & n7579 ;
  assign n7581 = ~n4602 & ~n7580 ;
  assign n7582 = ~n7574 & ~n7581 ;
  assign n7583 = n5982 & n7582 ;
  assign n7584 = ~n5982 & ~n7582 ;
  assign n7585 = ~n7583 & ~n7584 ;
  assign n7586 = n7453 & ~n7585 ;
  assign n7587 = ~n7517 & ~n7586 ;
  assign n7588 = n5329 & ~n7587 ;
  assign n7589 = ~n4728 & n5360 ;
  assign n7590 = n5363 & n7589 ;
  assign n7591 = n5357 & n7590 ;
  assign n7592 = ~n4763 & n5367 ;
  assign n7593 = n7591 & n7592 ;
  assign n7594 = ~n4601 & ~n4622 ;
  assign n7595 = ~n4647 & n7594 ;
  assign n7596 = ~n4552 & n7595 ;
  assign n7597 = n7593 & n7596 ;
  assign n7598 = ~n4500 & ~n7597 ;
  assign n7599 = n4500 & n7597 ;
  assign n7600 = ~n7598 & ~n7599 ;
  assign n7601 = ~n4231 & ~n7600 ;
  assign n7602 = n4231 & ~n4601 ;
  assign n7603 = ~n7601 & ~n7602 ;
  assign n7604 = n7453 & ~n7603 ;
  assign n7605 = ~n7517 & ~n7604 ;
  assign n7606 = n5383 & ~n7605 ;
  assign n7608 = n4543 & ~n5553 ;
  assign n7609 = ~n5554 & ~n7608 ;
  assign n7610 = n5563 & n7609 ;
  assign n7611 = n7453 & n7610 ;
  assign n7607 = n4548 & ~n7484 ;
  assign n7612 = n4543 & ~n7504 ;
  assign n7613 = ~n7607 & ~n7612 ;
  assign n7614 = ~n7611 & n7613 ;
  assign n7615 = ~n7606 & n7614 ;
  assign n7616 = ~n7588 & n7615 ;
  assign n7617 = ~n7552 & n7616 ;
  assign n7618 = n5583 & ~n7617 ;
  assign n7619 = ~n7516 & ~n7618 ;
  assign n7620 = \P1_state_reg[0]/NET0131  & ~n7619 ;
  assign n7621 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[27]/NET0131  ;
  assign n7622 = n4548 & n5786 ;
  assign n7623 = ~n7621 & ~n7622 ;
  assign n7624 = ~n7620 & n7623 ;
  assign n7625 = n4496 & n5585 ;
  assign n7626 = n4496 & ~n7453 ;
  assign n7627 = ~n6801 & n7453 ;
  assign n7628 = ~n7626 & ~n7627 ;
  assign n7629 = n5329 & ~n7628 ;
  assign n7630 = ~n6818 & n7453 ;
  assign n7631 = ~n7626 & ~n7630 ;
  assign n7632 = n5526 & ~n7631 ;
  assign n7633 = ~n6828 & n7453 ;
  assign n7634 = ~n7626 & ~n7633 ;
  assign n7635 = n5383 & ~n7634 ;
  assign n7637 = n6832 & n7453 ;
  assign n7638 = ~n7626 & ~n7637 ;
  assign n7639 = n5563 & ~n7638 ;
  assign n7636 = n4487 & ~n7504 ;
  assign n7640 = n5565 & ~n7453 ;
  assign n7641 = ~n5568 & ~n7640 ;
  assign n7642 = n4496 & ~n7641 ;
  assign n7643 = ~n7636 & ~n7642 ;
  assign n7644 = ~n7639 & n7643 ;
  assign n7645 = ~n7635 & n7644 ;
  assign n7646 = ~n7632 & n7645 ;
  assign n7647 = ~n7629 & n7646 ;
  assign n7648 = n5583 & ~n7647 ;
  assign n7649 = ~n7625 & ~n7648 ;
  assign n7650 = \P1_state_reg[0]/NET0131  & ~n7649 ;
  assign n7651 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[28]/NET0131  ;
  assign n7652 = n4496 & n5786 ;
  assign n7653 = ~n7651 & ~n7652 ;
  assign n7654 = ~n7650 & n7653 ;
  assign n7655 = n3030 & ~n6568 ;
  assign n7656 = n4027 & n4062 ;
  assign n7657 = ~n4059 & n7656 ;
  assign n7658 = ~n4026 & n4062 ;
  assign n7659 = ~n4020 & ~n7658 ;
  assign n7660 = ~n7657 & n7659 ;
  assign n7661 = n3037 & ~n7660 ;
  assign n7662 = ~n3037 & n7660 ;
  assign n7663 = ~n7661 & ~n7662 ;
  assign n7664 = n6568 & ~n7663 ;
  assign n7665 = ~n7655 & ~n7664 ;
  assign n7666 = n6282 & ~n7665 ;
  assign n7667 = n6628 & ~n6973 ;
  assign n7668 = n6178 & ~n7163 ;
  assign n7669 = ~n3438 & ~n3528 ;
  assign n7670 = ~n7668 & n7669 ;
  assign n7671 = ~n7667 & n7670 ;
  assign n7672 = ~n3439 & ~n7671 ;
  assign n7673 = ~n7002 & n7021 ;
  assign n7674 = n7008 & ~n7673 ;
  assign n7675 = n7004 & ~n7015 ;
  assign n7676 = n6982 & ~n7675 ;
  assign n7677 = ~n7674 & n7676 ;
  assign n7678 = ~n3439 & n6975 ;
  assign n7679 = n6628 & n7678 ;
  assign n7680 = ~n7677 & n7679 ;
  assign n7681 = ~n7672 & ~n7680 ;
  assign n7682 = n3037 & n7681 ;
  assign n7683 = ~n3037 & ~n7681 ;
  assign n7684 = ~n7682 & ~n7683 ;
  assign n7685 = n6568 & ~n7684 ;
  assign n7686 = ~n7655 & ~n7685 ;
  assign n7687 = n6207 & ~n7686 ;
  assign n7689 = n3410 & ~n6313 ;
  assign n7690 = ~n6314 & ~n7689 ;
  assign n7691 = ~n2713 & ~n7690 ;
  assign n7692 = n2713 & n3437 ;
  assign n7693 = n4011 & ~n7692 ;
  assign n7694 = ~n7691 & n7693 ;
  assign n7695 = n3019 & ~n6654 ;
  assign n7696 = ~n6353 & n6359 ;
  assign n7697 = ~n7695 & n7696 ;
  assign n7698 = ~n7694 & ~n7697 ;
  assign n7699 = n6568 & ~n7698 ;
  assign n7688 = n3030 & ~n6668 ;
  assign n7700 = n3019 & ~n6649 ;
  assign n7701 = ~n7688 & ~n7700 ;
  assign n7702 = ~n7699 & n7701 ;
  assign n7703 = ~n7687 & n7702 ;
  assign n7704 = ~n7666 & n7703 ;
  assign n7705 = n6097 & ~n7704 ;
  assign n7706 = n3030 & n6095 ;
  assign n7707 = ~n7705 & ~n7706 ;
  assign n7708 = \P1_state_reg[0]/NET0131  & ~n7707 ;
  assign n7709 = \P1_reg3_reg[28]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7710 = n3030 & n4130 ;
  assign n7711 = ~n7709 & ~n7710 ;
  assign n7712 = ~n7708 & n7711 ;
  assign n7715 = ~n1268 & n2145 ;
  assign n7716 = ~n1268 & ~n2236 ;
  assign n7717 = n2236 & ~n5657 ;
  assign n7718 = ~n7716 & ~n7717 ;
  assign n7719 = n2234 & ~n7718 ;
  assign n7720 = ~n1268 & ~n2163 ;
  assign n7728 = n2163 & ~n5679 ;
  assign n7729 = ~n7720 & ~n7728 ;
  assign n7730 = n737 & ~n7729 ;
  assign n7727 = n1262 & n2580 ;
  assign n7731 = ~n1268 & ~n2583 ;
  assign n7732 = ~n7727 & ~n7731 ;
  assign n7733 = ~n7730 & n7732 ;
  assign n7734 = ~n7719 & n7733 ;
  assign n7721 = n2163 & ~n5669 ;
  assign n7722 = ~n7720 & ~n7721 ;
  assign n7723 = n2393 & ~n7722 ;
  assign n7724 = n2236 & ~n5669 ;
  assign n7725 = ~n7716 & ~n7724 ;
  assign n7726 = n2391 & ~n7725 ;
  assign n7735 = ~n7723 & ~n7726 ;
  assign n7736 = n7734 & n7735 ;
  assign n7737 = n2147 & ~n7736 ;
  assign n7738 = ~n7715 & ~n7737 ;
  assign n7739 = \P1_state_reg[0]/NET0131  & ~n7738 ;
  assign n7713 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[25]/NET0131  ;
  assign n7714 = n765 & ~n1268 ;
  assign n7740 = ~n7713 & ~n7714 ;
  assign n7741 = ~n7739 & n7740 ;
  assign n7744 = ~n1470 & n2145 ;
  assign n7745 = ~n1470 & ~n2236 ;
  assign n7746 = n2236 & ~n5727 ;
  assign n7747 = ~n7745 & ~n7746 ;
  assign n7748 = n2234 & ~n7747 ;
  assign n7749 = ~n1470 & ~n2163 ;
  assign n7757 = n2163 & ~n5770 ;
  assign n7758 = ~n7749 & ~n7757 ;
  assign n7759 = n737 & ~n7758 ;
  assign n7756 = n1465 & n2580 ;
  assign n7760 = ~n1470 & ~n2583 ;
  assign n7761 = ~n7756 & ~n7760 ;
  assign n7762 = ~n7759 & n7761 ;
  assign n7763 = ~n7748 & n7762 ;
  assign n7750 = n2163 & ~n5757 ;
  assign n7751 = ~n7749 & ~n7750 ;
  assign n7752 = n2393 & ~n7751 ;
  assign n7753 = n2236 & ~n5757 ;
  assign n7754 = ~n7745 & ~n7753 ;
  assign n7755 = n2391 & ~n7754 ;
  assign n7764 = ~n7752 & ~n7755 ;
  assign n7765 = n7763 & n7764 ;
  assign n7766 = n2147 & ~n7765 ;
  assign n7767 = ~n7744 & ~n7766 ;
  assign n7768 = \P1_state_reg[0]/NET0131  & ~n7767 ;
  assign n7742 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[26]/NET0131  ;
  assign n7743 = n765 & ~n1470 ;
  assign n7769 = ~n7742 & ~n7743 ;
  assign n7770 = ~n7768 & n7769 ;
  assign n7771 = \P1_reg1_reg[25]/NET0131  & ~n6078 ;
  assign n7772 = \P1_reg1_reg[25]/NET0131  & n6095 ;
  assign n7780 = \P1_reg1_reg[25]/NET0131  & ~n6683 ;
  assign n7784 = n6683 & ~n7093 ;
  assign n7785 = ~n7780 & ~n7784 ;
  assign n7786 = n6207 & ~n7785 ;
  assign n7781 = n6683 & ~n7079 ;
  assign n7782 = ~n7780 & ~n7781 ;
  assign n7783 = n6282 & ~n7782 ;
  assign n7774 = n4011 & n7103 ;
  assign n7773 = n6359 & n7109 ;
  assign n7775 = n3165 & n6365 ;
  assign n7776 = ~n7773 & ~n7775 ;
  assign n7777 = ~n7774 & n7776 ;
  assign n7778 = n6683 & ~n7777 ;
  assign n7779 = \P1_reg1_reg[25]/NET0131  & ~n6696 ;
  assign n7787 = ~n7778 & ~n7779 ;
  assign n7788 = ~n7783 & n7787 ;
  assign n7789 = ~n7786 & n7788 ;
  assign n7790 = n6097 & ~n7789 ;
  assign n7791 = ~n7772 & ~n7790 ;
  assign n7792 = \P1_state_reg[0]/NET0131  & ~n7791 ;
  assign n7793 = ~n7771 & ~n7792 ;
  assign n7794 = \P1_reg1_reg[28]/NET0131  & ~n6683 ;
  assign n7795 = n6683 & ~n7663 ;
  assign n7796 = ~n7794 & ~n7795 ;
  assign n7797 = n6282 & ~n7796 ;
  assign n7798 = n6683 & ~n7684 ;
  assign n7799 = ~n7794 & ~n7798 ;
  assign n7800 = n6207 & ~n7799 ;
  assign n7801 = n3019 & n6365 ;
  assign n7802 = n7698 & ~n7801 ;
  assign n7803 = n6683 & ~n7802 ;
  assign n7804 = n6359 & ~n6683 ;
  assign n7805 = n6365 & ~n6683 ;
  assign n7806 = n6424 & ~n7805 ;
  assign n7807 = ~n7804 & n7806 ;
  assign n7808 = ~n6692 & n7807 ;
  assign n7809 = \P1_reg1_reg[28]/NET0131  & ~n7808 ;
  assign n7810 = ~n7803 & ~n7809 ;
  assign n7811 = ~n7800 & n7810 ;
  assign n7812 = ~n7797 & n7811 ;
  assign n7813 = n6097 & ~n7812 ;
  assign n7814 = \P1_reg1_reg[28]/NET0131  & n6095 ;
  assign n7815 = ~n7813 & ~n7814 ;
  assign n7816 = \P1_state_reg[0]/NET0131  & ~n7815 ;
  assign n7817 = \P1_reg1_reg[28]/NET0131  & ~n6078 ;
  assign n7818 = ~n7816 & ~n7817 ;
  assign n7819 = \P2_reg0_reg[24]/NET0131  & ~n5589 ;
  assign n7820 = \P2_reg0_reg[24]/NET0131  & n5585 ;
  assign n7836 = n4635 & n5565 ;
  assign n7837 = n5364 & n5365 ;
  assign n7838 = n5368 & n7837 ;
  assign n7839 = n4622 & ~n7838 ;
  assign n7840 = ~n5371 & ~n7839 ;
  assign n7841 = ~n4231 & ~n7840 ;
  assign n7842 = n4231 & n4665 ;
  assign n7843 = n5383 & ~n7842 ;
  assign n7844 = ~n7841 & n7843 ;
  assign n7845 = ~n4656 & n7496 ;
  assign n7846 = n4635 & ~n7845 ;
  assign n7847 = n5563 & ~n7497 ;
  assign n7848 = ~n7846 & n7847 ;
  assign n7849 = n5828 & n5836 ;
  assign n7850 = ~n5808 & n5835 ;
  assign n7851 = n5843 & ~n7850 ;
  assign n7852 = n5832 & ~n7851 ;
  assign n7853 = n5850 & ~n7852 ;
  assign n7854 = ~n7849 & n7853 ;
  assign n7856 = ~n5984 & ~n7854 ;
  assign n7855 = n5984 & n7854 ;
  assign n7857 = n5526 & ~n7855 ;
  assign n7858 = ~n7856 & n7857 ;
  assign n7859 = ~n7848 & ~n7858 ;
  assign n7860 = ~n7844 & n7859 ;
  assign n7861 = ~n7836 & n7860 ;
  assign n7862 = n6706 & ~n7861 ;
  assign n7821 = n6748 & n6762 ;
  assign n7822 = ~n6754 & n6758 ;
  assign n7823 = n6769 & ~n7822 ;
  assign n7824 = n6761 & ~n7823 ;
  assign n7825 = n6776 & ~n7824 ;
  assign n7826 = ~n7821 & n7825 ;
  assign n7827 = n6781 & ~n7826 ;
  assign n7828 = ~n6791 & ~n7827 ;
  assign n7829 = n5984 & n7828 ;
  assign n7830 = ~n5984 & ~n7828 ;
  assign n7831 = ~n7829 & ~n7830 ;
  assign n7832 = n6706 & n7831 ;
  assign n7833 = ~\P2_reg0_reg[24]/NET0131  & ~n6706 ;
  assign n7834 = n5329 & ~n7833 ;
  assign n7835 = ~n7832 & n7834 ;
  assign n7863 = n5565 & ~n6706 ;
  assign n7864 = n6394 & ~n7863 ;
  assign n7865 = ~n5526 & ~n5563 ;
  assign n7866 = ~n5383 & n7865 ;
  assign n7867 = ~n6706 & ~n7866 ;
  assign n7868 = n7864 & ~n7867 ;
  assign n7869 = \P2_reg0_reg[24]/NET0131  & ~n7868 ;
  assign n7870 = ~n7835 & ~n7869 ;
  assign n7871 = ~n7862 & n7870 ;
  assign n7872 = n5583 & ~n7871 ;
  assign n7873 = ~n7820 & ~n7872 ;
  assign n7874 = \P1_state_reg[0]/NET0131  & ~n7873 ;
  assign n7875 = ~n7819 & ~n7874 ;
  assign n7876 = \P2_reg0_reg[26]/NET0131  & ~n5589 ;
  assign n7877 = \P2_reg0_reg[26]/NET0131  & n5585 ;
  assign n7878 = \P2_reg0_reg[26]/NET0131  & ~n6706 ;
  assign n7913 = ~n5816 & ~n5819 ;
  assign n7914 = n5809 & n5825 ;
  assign n7915 = ~n7913 & n7914 ;
  assign n7916 = ~n5822 & n5825 ;
  assign n7917 = ~n5801 & ~n7916 ;
  assign n7918 = ~n7915 & n7917 ;
  assign n7919 = n5450 & n5804 ;
  assign n7920 = ~n7918 & n7919 ;
  assign n7921 = n5793 & n5834 ;
  assign n7922 = n7920 & n7921 ;
  assign n7923 = n5799 & n5804 ;
  assign n7924 = ~n5795 & ~n7923 ;
  assign n7925 = n7921 & ~n7924 ;
  assign n7926 = n5792 & n5834 ;
  assign n7927 = ~n5839 & ~n7926 ;
  assign n7928 = ~n7925 & n7927 ;
  assign n7929 = ~n7922 & n7928 ;
  assign n7930 = n5789 & n5830 ;
  assign n7931 = n5831 & n5833 ;
  assign n7932 = n7930 & n7931 ;
  assign n7933 = ~n7929 & n7932 ;
  assign n7935 = n5831 & n5842 ;
  assign n7936 = ~n5846 & ~n7935 ;
  assign n7937 = n7930 & ~n7936 ;
  assign n7934 = n5789 & n5849 ;
  assign n7938 = ~n5856 & ~n7934 ;
  assign n7939 = ~n7937 & n7938 ;
  assign n7940 = ~n7933 & n7939 ;
  assign n7941 = n5977 & n7940 ;
  assign n7942 = ~n5977 & ~n7940 ;
  assign n7943 = ~n7941 & ~n7942 ;
  assign n7944 = n6706 & n7943 ;
  assign n7945 = ~n7878 & ~n7944 ;
  assign n7946 = n5526 & ~n7945 ;
  assign n7879 = n6757 & n6760 ;
  assign n7880 = n6731 & n6745 ;
  assign n7881 = ~n6740 & n7880 ;
  assign n7882 = ~n6743 & n6745 ;
  assign n7883 = n6750 & ~n7882 ;
  assign n7884 = ~n7881 & n7883 ;
  assign n7885 = n6746 & n6756 ;
  assign n7886 = ~n7884 & n7885 ;
  assign n7887 = n7879 & n7886 ;
  assign n7888 = ~n6753 & n6756 ;
  assign n7889 = ~n6765 & ~n7888 ;
  assign n7890 = n7879 & ~n7889 ;
  assign n7891 = n6760 & n6768 ;
  assign n7892 = ~n6772 & ~n7891 ;
  assign n7893 = ~n7890 & n7892 ;
  assign n7894 = ~n7887 & n7893 ;
  assign n7895 = n6759 & n6779 ;
  assign n7896 = ~n4686 & n7570 ;
  assign n7897 = n7895 & n7896 ;
  assign n7898 = ~n7894 & n7897 ;
  assign n7899 = ~n6775 & n6779 ;
  assign n7900 = n6788 & ~n7899 ;
  assign n7901 = n7896 & ~n7900 ;
  assign n7902 = n4667 & ~n6786 ;
  assign n7903 = n6785 & ~n7902 ;
  assign n7904 = ~n4626 & ~n7903 ;
  assign n7905 = ~n7901 & ~n7904 ;
  assign n7906 = ~n7898 & n7905 ;
  assign n7907 = n5977 & n7906 ;
  assign n7908 = ~n5977 & ~n7906 ;
  assign n7909 = ~n7907 & ~n7908 ;
  assign n7910 = n6706 & ~n7909 ;
  assign n7911 = ~n7878 & ~n7910 ;
  assign n7912 = n5329 & ~n7911 ;
  assign n7948 = n7593 & n7595 ;
  assign n7949 = n4552 & ~n7948 ;
  assign n7950 = ~n7597 & ~n7949 ;
  assign n7951 = ~n4231 & ~n7950 ;
  assign n7952 = n4231 & n4622 ;
  assign n7953 = ~n7951 & ~n7952 ;
  assign n7954 = n6706 & n7953 ;
  assign n7955 = ~n7878 & ~n7954 ;
  assign n7956 = n5383 & ~n7955 ;
  assign n7947 = \P2_reg0_reg[26]/NET0131  & ~n6717 ;
  assign n7957 = n4592 & n5565 ;
  assign n7958 = n4592 & ~n7499 ;
  assign n7959 = ~n5553 & n5563 ;
  assign n7960 = ~n7958 & n7959 ;
  assign n7961 = ~n7957 & ~n7960 ;
  assign n7962 = n6706 & ~n7961 ;
  assign n7963 = ~n7947 & ~n7962 ;
  assign n7964 = ~n7956 & n7963 ;
  assign n7965 = ~n7912 & n7964 ;
  assign n7966 = ~n7946 & n7965 ;
  assign n7967 = n5583 & ~n7966 ;
  assign n7968 = ~n7877 & ~n7967 ;
  assign n7969 = \P1_state_reg[0]/NET0131  & ~n7968 ;
  assign n7970 = ~n7876 & ~n7969 ;
  assign n7971 = \P2_reg0_reg[27]/NET0131  & n5585 ;
  assign n7972 = \P2_reg0_reg[27]/NET0131  & ~n6706 ;
  assign n7973 = n6706 & ~n7549 ;
  assign n7974 = ~n7972 & ~n7973 ;
  assign n7975 = n5526 & ~n7974 ;
  assign n7976 = n6706 & ~n7585 ;
  assign n7977 = ~n7972 & ~n7976 ;
  assign n7978 = n5329 & ~n7977 ;
  assign n7979 = n5383 & ~n7603 ;
  assign n7980 = n4543 & n5565 ;
  assign n7981 = ~n7610 & ~n7980 ;
  assign n7982 = ~n7979 & n7981 ;
  assign n7983 = n6706 & ~n7982 ;
  assign n7984 = n5383 & ~n6706 ;
  assign n7985 = n6717 & ~n7984 ;
  assign n7986 = \P2_reg0_reg[27]/NET0131  & ~n7985 ;
  assign n7987 = ~n7983 & ~n7986 ;
  assign n7988 = ~n7978 & n7987 ;
  assign n7989 = ~n7975 & n7988 ;
  assign n7990 = n5583 & ~n7989 ;
  assign n7991 = ~n7971 & ~n7990 ;
  assign n7992 = \P1_state_reg[0]/NET0131  & ~n7991 ;
  assign n7993 = \P2_reg0_reg[27]/NET0131  & ~n5589 ;
  assign n7994 = ~n7992 & ~n7993 ;
  assign n7995 = \P2_reg1_reg[25]/NET0131  & ~n5589 ;
  assign n7996 = \P2_reg1_reg[25]/NET0131  & n5585 ;
  assign n8002 = n5383 & n7491 ;
  assign n8001 = n5526 & ~n7479 ;
  assign n8000 = n4613 & n5565 ;
  assign n8003 = ~n7501 & ~n8000 ;
  assign n8004 = ~n8001 & n8003 ;
  assign n8005 = ~n8002 & n8004 ;
  assign n8006 = n6380 & ~n8005 ;
  assign n7997 = n5383 & ~n6380 ;
  assign n7998 = n6398 & ~n7997 ;
  assign n7999 = \P2_reg1_reg[25]/NET0131  & ~n7998 ;
  assign n8008 = n6380 & n7465 ;
  assign n8007 = ~\P2_reg1_reg[25]/NET0131  & ~n6380 ;
  assign n8009 = n5329 & ~n8007 ;
  assign n8010 = ~n8008 & n8009 ;
  assign n8011 = ~n7999 & ~n8010 ;
  assign n8012 = ~n8006 & n8011 ;
  assign n8013 = n5583 & ~n8012 ;
  assign n8014 = ~n7996 & ~n8013 ;
  assign n8015 = \P1_state_reg[0]/NET0131  & ~n8014 ;
  assign n8016 = ~n7995 & ~n8015 ;
  assign n8017 = \P2_reg1_reg[27]/NET0131  & n5585 ;
  assign n8018 = \P2_reg1_reg[27]/NET0131  & ~n6380 ;
  assign n8019 = n6380 & ~n7549 ;
  assign n8020 = ~n8018 & ~n8019 ;
  assign n8021 = n5526 & ~n8020 ;
  assign n8022 = n6380 & ~n7585 ;
  assign n8023 = ~n8018 & ~n8022 ;
  assign n8024 = n5329 & ~n8023 ;
  assign n8025 = n6380 & ~n7982 ;
  assign n8026 = n6397 & ~n7997 ;
  assign n8027 = \P2_reg1_reg[27]/NET0131  & ~n8026 ;
  assign n8028 = ~n8025 & ~n8027 ;
  assign n8029 = ~n8024 & n8028 ;
  assign n8030 = ~n8021 & n8029 ;
  assign n8031 = n5583 & ~n8030 ;
  assign n8032 = ~n8017 & ~n8031 ;
  assign n8033 = \P1_state_reg[0]/NET0131  & ~n8032 ;
  assign n8034 = \P2_reg1_reg[27]/NET0131  & ~n5589 ;
  assign n8035 = ~n8033 & ~n8034 ;
  assign n8036 = \P2_reg1_reg[28]/NET0131  & ~n5589 ;
  assign n8037 = \P2_reg1_reg[28]/NET0131  & n5585 ;
  assign n8038 = \P2_reg1_reg[28]/NET0131  & ~n6380 ;
  assign n8039 = n6380 & ~n6801 ;
  assign n8040 = ~n8038 & ~n8039 ;
  assign n8041 = n5329 & ~n8040 ;
  assign n8042 = n6380 & ~n6818 ;
  assign n8043 = ~n8038 & ~n8042 ;
  assign n8044 = n5526 & ~n8043 ;
  assign n8045 = n6380 & ~n6835 ;
  assign n8046 = \P2_reg1_reg[28]/NET0131  & ~n8026 ;
  assign n8047 = ~n8045 & ~n8046 ;
  assign n8048 = ~n8044 & n8047 ;
  assign n8049 = ~n8041 & n8048 ;
  assign n8050 = n5583 & ~n8049 ;
  assign n8051 = ~n8037 & ~n8050 ;
  assign n8052 = \P1_state_reg[0]/NET0131  & ~n8051 ;
  assign n8053 = ~n8036 & ~n8052 ;
  assign n8054 = \P1_reg2_reg[28]/NET0131  & ~n6078 ;
  assign n8065 = n6113 & n7663 ;
  assign n8064 = ~\P1_reg2_reg[28]/NET0131  & ~n6113 ;
  assign n8066 = n6282 & ~n8064 ;
  assign n8067 = ~n8065 & n8066 ;
  assign n8055 = n6207 & ~n7684 ;
  assign n8056 = n7802 & ~n8055 ;
  assign n8057 = n6113 & ~n8056 ;
  assign n8058 = n3030 & n4112 ;
  assign n8059 = ~n4009 & ~n6426 ;
  assign n8060 = ~n6365 & n8059 ;
  assign n8061 = ~n6113 & ~n8060 ;
  assign n8062 = ~n6361 & ~n8061 ;
  assign n8063 = \P1_reg2_reg[28]/NET0131  & ~n8062 ;
  assign n8068 = ~n8058 & ~n8063 ;
  assign n8069 = ~n8057 & n8068 ;
  assign n8070 = ~n8067 & n8069 ;
  assign n8071 = n6097 & ~n8070 ;
  assign n8072 = \P1_reg2_reg[28]/NET0131  & n6095 ;
  assign n8073 = ~n8071 & ~n8072 ;
  assign n8074 = \P1_state_reg[0]/NET0131  & ~n8073 ;
  assign n8075 = ~n8054 & ~n8074 ;
  assign n8076 = \P2_reg2_reg[27]/NET0131  & n5585 ;
  assign n8077 = \P2_reg2_reg[27]/NET0131  & ~n4219 ;
  assign n8078 = n4219 & ~n7549 ;
  assign n8079 = ~n8077 & ~n8078 ;
  assign n8080 = n5526 & ~n8079 ;
  assign n8081 = n4219 & ~n7585 ;
  assign n8082 = ~n8077 & ~n8081 ;
  assign n8083 = n5329 & ~n8082 ;
  assign n8084 = n4219 & ~n7603 ;
  assign n8085 = ~n8077 & ~n8084 ;
  assign n8086 = n5383 & ~n8085 ;
  assign n8088 = n4219 & n7609 ;
  assign n8089 = ~n8077 & ~n8088 ;
  assign n8090 = n5563 & ~n8089 ;
  assign n8092 = n4219 & n7980 ;
  assign n8087 = \P2_reg2_reg[27]/NET0131  & ~n5570 ;
  assign n8091 = n4548 & n5574 ;
  assign n8093 = ~n8087 & ~n8091 ;
  assign n8094 = ~n8092 & n8093 ;
  assign n8095 = ~n8090 & n8094 ;
  assign n8096 = ~n8086 & n8095 ;
  assign n8097 = ~n8083 & n8096 ;
  assign n8098 = ~n8080 & n8097 ;
  assign n8099 = n5583 & ~n8098 ;
  assign n8100 = ~n8076 & ~n8099 ;
  assign n8101 = \P1_state_reg[0]/NET0131  & ~n8100 ;
  assign n8102 = \P2_reg2_reg[27]/NET0131  & ~n5589 ;
  assign n8103 = ~n8101 & ~n8102 ;
  assign n8104 = \P1_reg0_reg[26]/NET0131  & ~n6078 ;
  assign n8105 = \P1_reg0_reg[26]/NET0131  & n6095 ;
  assign n8106 = \P1_reg0_reg[26]/NET0131  & ~n6409 ;
  assign n8107 = n6409 & ~n7156 ;
  assign n8108 = ~n8106 & ~n8107 ;
  assign n8109 = n6282 & ~n8108 ;
  assign n8110 = n6409 & ~n7192 ;
  assign n8111 = ~n8106 & ~n8110 ;
  assign n8112 = n6207 & ~n8111 ;
  assign n8113 = \P1_reg0_reg[26]/NET0131  & ~n6429 ;
  assign n8114 = n3518 & n6365 ;
  assign n8115 = ~n7201 & ~n8114 ;
  assign n8116 = ~n7204 & n8115 ;
  assign n8117 = n6409 & ~n8116 ;
  assign n8118 = ~n8113 & ~n8117 ;
  assign n8119 = ~n8112 & n8118 ;
  assign n8120 = ~n8109 & n8119 ;
  assign n8121 = n6097 & ~n8120 ;
  assign n8122 = ~n8105 & ~n8121 ;
  assign n8123 = \P1_state_reg[0]/NET0131  & ~n8122 ;
  assign n8124 = ~n8104 & ~n8123 ;
  assign n8125 = \P1_reg0_reg[27]/NET0131  & ~n6409 ;
  assign n8126 = n6409 & ~n6603 ;
  assign n8127 = ~n8125 & ~n8126 ;
  assign n8128 = n6282 & ~n8127 ;
  assign n8129 = n6409 & ~n6644 ;
  assign n8130 = ~n8125 & ~n8129 ;
  assign n8131 = n6207 & ~n8130 ;
  assign n8132 = n3427 & n6365 ;
  assign n8133 = n6663 & ~n8132 ;
  assign n8134 = n6409 & ~n8133 ;
  assign n8135 = \P1_reg0_reg[27]/NET0131  & ~n6429 ;
  assign n8136 = ~n8134 & ~n8135 ;
  assign n8137 = ~n8131 & n8136 ;
  assign n8138 = ~n8128 & n8137 ;
  assign n8139 = n6097 & ~n8138 ;
  assign n8140 = \P1_reg0_reg[27]/NET0131  & n6095 ;
  assign n8141 = ~n8139 & ~n8140 ;
  assign n8142 = \P1_state_reg[0]/NET0131  & ~n8141 ;
  assign n8143 = \P1_reg0_reg[27]/NET0131  & ~n6078 ;
  assign n8144 = ~n8142 & ~n8143 ;
  assign n8145 = \P1_reg0_reg[24]/NET0131  & ~n6078 ;
  assign n8146 = \P1_reg0_reg[24]/NET0131  & n6095 ;
  assign n8153 = \P1_reg0_reg[24]/NET0131  & ~n6409 ;
  assign n8157 = n6409 & ~n7031 ;
  assign n8158 = ~n8153 & ~n8157 ;
  assign n8159 = n6207 & ~n8158 ;
  assign n8154 = n6409 & ~n6964 ;
  assign n8155 = ~n8153 & ~n8154 ;
  assign n8156 = n6282 & ~n8155 ;
  assign n8147 = \P1_reg0_reg[24]/NET0131  & ~n6429 ;
  assign n8149 = n4011 & n7044 ;
  assign n8148 = n3539 & n6365 ;
  assign n8150 = ~n7050 & ~n8148 ;
  assign n8151 = ~n8149 & n8150 ;
  assign n8152 = n6409 & ~n8151 ;
  assign n8160 = ~n8147 & ~n8152 ;
  assign n8161 = ~n8156 & n8160 ;
  assign n8162 = ~n8159 & n8161 ;
  assign n8163 = n6097 & ~n8162 ;
  assign n8164 = ~n8146 & ~n8163 ;
  assign n8165 = \P1_state_reg[0]/NET0131  & ~n8164 ;
  assign n8166 = ~n8145 & ~n8165 ;
  assign n8167 = \P3_reg0_reg[24]/NET0131  & ~n2143 ;
  assign n8168 = \P3_reg0_reg[24]/NET0131  & n2145 ;
  assign n8169 = \P3_reg0_reg[24]/NET0131  & ~n2163 ;
  assign n8178 = n2163 & ~n5634 ;
  assign n8179 = ~n8169 & ~n8178 ;
  assign n8180 = n2234 & ~n8179 ;
  assign n8172 = \P3_reg0_reg[24]/NET0131  & ~n2236 ;
  assign n8175 = n2236 & ~n5621 ;
  assign n8176 = ~n8172 & ~n8175 ;
  assign n8177 = n737 & ~n8176 ;
  assign n8181 = \P3_reg0_reg[24]/NET0131  & ~n2287 ;
  assign n8182 = n1223 & n2289 ;
  assign n8183 = ~n8181 & ~n8182 ;
  assign n8184 = ~n8177 & n8183 ;
  assign n8185 = ~n8180 & n8184 ;
  assign n8170 = ~n5611 & ~n8169 ;
  assign n8171 = n2391 & ~n8170 ;
  assign n8173 = ~n5607 & ~n8172 ;
  assign n8174 = n2393 & ~n8173 ;
  assign n8186 = ~n8171 & ~n8174 ;
  assign n8187 = n8185 & n8186 ;
  assign n8188 = n2147 & ~n8187 ;
  assign n8189 = ~n8168 & ~n8188 ;
  assign n8190 = \P1_state_reg[0]/NET0131  & ~n8189 ;
  assign n8191 = ~n8167 & ~n8190 ;
  assign n8192 = \P3_reg0_reg[25]/NET0131  & ~n2143 ;
  assign n8193 = \P3_reg0_reg[25]/NET0131  & n2145 ;
  assign n8194 = \P3_reg0_reg[25]/NET0131  & ~n2163 ;
  assign n8195 = n2163 & ~n5657 ;
  assign n8196 = ~n8194 & ~n8195 ;
  assign n8197 = n2234 & ~n8196 ;
  assign n8198 = \P3_reg0_reg[25]/NET0131  & ~n2236 ;
  assign n8204 = n2236 & ~n5679 ;
  assign n8205 = ~n8198 & ~n8204 ;
  assign n8206 = n737 & ~n8205 ;
  assign n8203 = \P3_reg0_reg[25]/NET0131  & ~n2287 ;
  assign n8207 = n1262 & n2289 ;
  assign n8208 = ~n8203 & ~n8207 ;
  assign n8209 = ~n8206 & n8208 ;
  assign n8210 = ~n8197 & n8209 ;
  assign n8199 = ~n7724 & ~n8198 ;
  assign n8200 = n2393 & ~n8199 ;
  assign n8201 = ~n7721 & ~n8194 ;
  assign n8202 = n2391 & ~n8201 ;
  assign n8211 = ~n8200 & ~n8202 ;
  assign n8212 = n8210 & n8211 ;
  assign n8213 = n2147 & ~n8212 ;
  assign n8214 = ~n8193 & ~n8213 ;
  assign n8215 = \P1_state_reg[0]/NET0131  & ~n8214 ;
  assign n8216 = ~n8192 & ~n8215 ;
  assign n8217 = \P1_reg0_reg[28]/NET0131  & ~n6409 ;
  assign n8218 = n6409 & ~n7663 ;
  assign n8219 = ~n8217 & ~n8218 ;
  assign n8220 = n6282 & ~n8219 ;
  assign n8221 = n6409 & ~n7684 ;
  assign n8222 = ~n8217 & ~n8221 ;
  assign n8223 = n6207 & ~n8222 ;
  assign n8224 = n6409 & ~n7802 ;
  assign n8225 = \P1_reg0_reg[28]/NET0131  & ~n6429 ;
  assign n8226 = ~n8224 & ~n8225 ;
  assign n8227 = ~n8223 & n8226 ;
  assign n8228 = ~n8220 & n8227 ;
  assign n8229 = n6097 & ~n8228 ;
  assign n8230 = \P1_reg0_reg[28]/NET0131  & n6095 ;
  assign n8231 = ~n8229 & ~n8230 ;
  assign n8232 = \P1_state_reg[0]/NET0131  & ~n8231 ;
  assign n8233 = \P1_reg0_reg[28]/NET0131  & ~n6078 ;
  assign n8234 = ~n8232 & ~n8233 ;
  assign n8235 = \P3_reg0_reg[26]/NET0131  & ~n2143 ;
  assign n8236 = \P3_reg0_reg[26]/NET0131  & n2145 ;
  assign n8237 = \P3_reg0_reg[26]/NET0131  & ~n2163 ;
  assign n8238 = n2163 & ~n5727 ;
  assign n8239 = ~n8237 & ~n8238 ;
  assign n8240 = n2234 & ~n8239 ;
  assign n8241 = \P3_reg0_reg[26]/NET0131  & ~n2236 ;
  assign n8247 = n2236 & ~n5770 ;
  assign n8248 = ~n8241 & ~n8247 ;
  assign n8249 = n737 & ~n8248 ;
  assign n8246 = n1465 & n2289 ;
  assign n8250 = \P3_reg0_reg[26]/NET0131  & ~n2287 ;
  assign n8251 = ~n8246 & ~n8250 ;
  assign n8252 = ~n8249 & n8251 ;
  assign n8253 = ~n8240 & n8252 ;
  assign n8242 = ~n7753 & ~n8241 ;
  assign n8243 = n2393 & ~n8242 ;
  assign n8244 = ~n7750 & ~n8237 ;
  assign n8245 = n2391 & ~n8244 ;
  assign n8254 = ~n8243 & ~n8245 ;
  assign n8255 = n8253 & n8254 ;
  assign n8256 = n2147 & ~n8255 ;
  assign n8257 = ~n8236 & ~n8256 ;
  assign n8258 = \P1_state_reg[0]/NET0131  & ~n8257 ;
  assign n8259 = ~n8235 & ~n8258 ;
  assign n8260 = \P3_reg1_reg[25]/NET0131  & ~n2143 ;
  assign n8261 = \P3_reg1_reg[25]/NET0131  & n2145 ;
  assign n8262 = \P3_reg1_reg[25]/NET0131  & ~n2427 ;
  assign n8263 = ~n5662 & ~n8262 ;
  assign n8264 = n2425 & ~n8263 ;
  assign n8272 = n2427 & ~n5679 ;
  assign n8273 = ~n8262 & ~n8272 ;
  assign n8274 = n737 & ~n8273 ;
  assign n8271 = \P3_reg1_reg[25]/NET0131  & ~n6449 ;
  assign n8275 = n1262 & n6451 ;
  assign n8276 = ~n8271 & ~n8275 ;
  assign n8277 = ~n8274 & n8276 ;
  assign n8278 = ~n8264 & n8277 ;
  assign n8265 = \P3_reg1_reg[25]/NET0131  & ~n2408 ;
  assign n8266 = ~n5658 & ~n8265 ;
  assign n8267 = ~n2518 & ~n8266 ;
  assign n8268 = n2408 & ~n5669 ;
  assign n8269 = ~n8265 & ~n8268 ;
  assign n8270 = n714 & ~n8269 ;
  assign n8279 = ~n8267 & ~n8270 ;
  assign n8280 = n8278 & n8279 ;
  assign n8281 = n2147 & ~n8280 ;
  assign n8282 = ~n8261 & ~n8281 ;
  assign n8283 = \P1_state_reg[0]/NET0131  & ~n8282 ;
  assign n8284 = ~n8260 & ~n8283 ;
  assign n8285 = \P3_reg1_reg[26]/NET0131  & ~n2143 ;
  assign n8286 = \P3_reg1_reg[26]/NET0131  & n2145 ;
  assign n8287 = \P3_reg1_reg[26]/NET0131  & ~n2408 ;
  assign n8288 = ~n5762 & ~n8287 ;
  assign n8289 = ~n2518 & ~n8288 ;
  assign n8293 = \P3_reg1_reg[26]/NET0131  & ~n2427 ;
  assign n8297 = n2427 & ~n5770 ;
  assign n8298 = ~n8293 & ~n8297 ;
  assign n8299 = n737 & ~n8298 ;
  assign n8296 = n1465 & n6451 ;
  assign n8300 = \P3_reg1_reg[26]/NET0131  & ~n6449 ;
  assign n8301 = ~n8296 & ~n8300 ;
  assign n8302 = ~n8299 & n8301 ;
  assign n8303 = ~n8289 & n8302 ;
  assign n8290 = n2408 & ~n5757 ;
  assign n8291 = ~n8287 & ~n8290 ;
  assign n8292 = n714 & ~n8291 ;
  assign n8294 = ~n5728 & ~n8293 ;
  assign n8295 = n2425 & ~n8294 ;
  assign n8304 = ~n8292 & ~n8295 ;
  assign n8305 = n8303 & n8304 ;
  assign n8306 = n2147 & ~n8305 ;
  assign n8307 = ~n8286 & ~n8306 ;
  assign n8308 = \P1_state_reg[0]/NET0131  & ~n8307 ;
  assign n8309 = ~n8285 & ~n8308 ;
  assign n8310 = \P3_reg1_reg[24]/NET0131  & ~n2143 ;
  assign n8311 = \P3_reg1_reg[24]/NET0131  & n2145 ;
  assign n8312 = \P3_reg1_reg[24]/NET0131  & ~n2408 ;
  assign n8313 = n2408 & ~n5606 ;
  assign n8314 = ~n8312 & ~n8313 ;
  assign n8315 = n714 & ~n8314 ;
  assign n8316 = \P3_reg1_reg[24]/NET0131  & ~n2427 ;
  assign n8317 = ~n6481 & ~n8316 ;
  assign n8318 = n2425 & ~n8317 ;
  assign n8319 = \P3_reg1_reg[24]/NET0131  & ~n6449 ;
  assign n8320 = n1223 & n6451 ;
  assign n8326 = ~n8319 & ~n8320 ;
  assign n8327 = ~n8318 & n8326 ;
  assign n8321 = ~n6475 & ~n8312 ;
  assign n8322 = ~n2518 & ~n8321 ;
  assign n8323 = n2427 & ~n5621 ;
  assign n8324 = ~n8316 & ~n8323 ;
  assign n8325 = n737 & ~n8324 ;
  assign n8328 = ~n8322 & ~n8325 ;
  assign n8329 = n8327 & n8328 ;
  assign n8330 = ~n8315 & n8329 ;
  assign n8331 = n2147 & ~n8330 ;
  assign n8332 = ~n8311 & ~n8331 ;
  assign n8333 = \P1_state_reg[0]/NET0131  & ~n8332 ;
  assign n8334 = ~n8310 & ~n8333 ;
  assign n8335 = \P3_reg2_reg[22]/NET0131  & ~n2143 ;
  assign n8336 = \P3_reg2_reg[22]/NET0131  & n2145 ;
  assign n8337 = \P3_reg2_reg[22]/NET0131  & ~n2427 ;
  assign n8338 = n2427 & ~n7343 ;
  assign n8339 = ~n8337 & ~n8338 ;
  assign n8340 = n714 & ~n8339 ;
  assign n8341 = \P3_reg2_reg[22]/NET0131  & ~n2408 ;
  assign n8349 = n2408 & ~n7363 ;
  assign n8350 = ~n8341 & ~n8349 ;
  assign n8351 = n737 & ~n8350 ;
  assign n8345 = n991 & n2441 ;
  assign n8352 = \P3_reg2_reg[22]/NET0131  & ~n2429 ;
  assign n8353 = ~n996 & n2283 ;
  assign n8354 = ~n8352 & ~n8353 ;
  assign n8355 = ~n8345 & n8354 ;
  assign n8356 = ~n8351 & n8355 ;
  assign n8357 = ~n8340 & n8356 ;
  assign n8342 = n2408 & ~n7355 ;
  assign n8343 = ~n8341 & ~n8342 ;
  assign n8344 = n2425 & ~n8343 ;
  assign n8346 = n2427 & ~n7355 ;
  assign n8347 = ~n8337 & ~n8346 ;
  assign n8348 = ~n2518 & ~n8347 ;
  assign n8358 = ~n8344 & ~n8348 ;
  assign n8359 = n8357 & n8358 ;
  assign n8360 = n2147 & ~n8359 ;
  assign n8361 = ~n8336 & ~n8360 ;
  assign n8362 = \P1_state_reg[0]/NET0131  & ~n8361 ;
  assign n8363 = ~n8335 & ~n8362 ;
  assign n8364 = \P3_reg2_reg[21]/NET0131  & ~n2143 ;
  assign n8365 = \P3_reg2_reg[21]/NET0131  & n2145 ;
  assign n8370 = \P3_reg2_reg[21]/NET0131  & ~n2427 ;
  assign n8371 = n2427 & ~n7297 ;
  assign n8372 = ~n8370 & ~n8371 ;
  assign n8373 = n714 & ~n8372 ;
  assign n8366 = \P3_reg2_reg[21]/NET0131  & ~n2408 ;
  assign n8367 = n2408 & ~n7315 ;
  assign n8368 = ~n8366 & ~n8367 ;
  assign n8369 = n737 & ~n8368 ;
  assign n8380 = n1029 & n2441 ;
  assign n8381 = \P3_reg2_reg[21]/NET0131  & ~n2429 ;
  assign n8382 = ~n1034 & n2283 ;
  assign n8383 = ~n8381 & ~n8382 ;
  assign n8384 = ~n8380 & n8383 ;
  assign n8385 = ~n8369 & n8384 ;
  assign n8386 = ~n8373 & n8385 ;
  assign n8374 = n2408 & ~n7307 ;
  assign n8375 = ~n8366 & ~n8374 ;
  assign n8376 = n2425 & ~n8375 ;
  assign n8377 = n2427 & ~n7307 ;
  assign n8378 = ~n8370 & ~n8377 ;
  assign n8379 = ~n2518 & ~n8378 ;
  assign n8387 = ~n8376 & ~n8379 ;
  assign n8388 = n8386 & n8387 ;
  assign n8389 = n2147 & ~n8388 ;
  assign n8390 = ~n8365 & ~n8389 ;
  assign n8391 = \P1_state_reg[0]/NET0131  & ~n8390 ;
  assign n8392 = ~n8364 & ~n8391 ;
  assign n8393 = \P3_reg2_reg[23]/NET0131  & ~n2143 ;
  assign n8394 = \P3_reg2_reg[23]/NET0131  & n2145 ;
  assign n8395 = \P3_reg2_reg[23]/NET0131  & ~n2427 ;
  assign n8396 = n2427 & ~n7386 ;
  assign n8397 = ~n8395 & ~n8396 ;
  assign n8398 = n714 & ~n8397 ;
  assign n8399 = n2427 & ~n7405 ;
  assign n8400 = ~n8395 & ~n8399 ;
  assign n8401 = ~n2518 & ~n8400 ;
  assign n8404 = n886 & n2441 ;
  assign n8402 = \P3_reg2_reg[23]/NET0131  & ~n2429 ;
  assign n8403 = ~n929 & n2283 ;
  assign n8412 = ~n8402 & ~n8403 ;
  assign n8413 = ~n8404 & n8412 ;
  assign n8414 = ~n8401 & n8413 ;
  assign n8405 = \P3_reg2_reg[23]/NET0131  & ~n2408 ;
  assign n8406 = n2408 & ~n7398 ;
  assign n8407 = ~n8405 & ~n8406 ;
  assign n8408 = n737 & ~n8407 ;
  assign n8409 = n2408 & ~n7405 ;
  assign n8410 = ~n8405 & ~n8409 ;
  assign n8411 = n2425 & ~n8410 ;
  assign n8415 = ~n8408 & ~n8411 ;
  assign n8416 = n8414 & n8415 ;
  assign n8417 = ~n8398 & n8416 ;
  assign n8418 = n2147 & ~n8417 ;
  assign n8419 = ~n8394 & ~n8418 ;
  assign n8420 = \P1_state_reg[0]/NET0131  & ~n8419 ;
  assign n8421 = ~n8393 & ~n8420 ;
  assign n8424 = n4793 & n5585 ;
  assign n8426 = n4793 & ~n7453 ;
  assign n8427 = n4728 & ~n5364 ;
  assign n8428 = ~n7591 & ~n8427 ;
  assign n8429 = ~n4231 & ~n8428 ;
  assign n8430 = n4231 & n4774 ;
  assign n8431 = ~n8429 & ~n8430 ;
  assign n8432 = n7453 & n8431 ;
  assign n8433 = ~n8426 & ~n8432 ;
  assign n8434 = n5383 & ~n8433 ;
  assign n8447 = ~n4789 & n5544 ;
  assign n8448 = n4814 & ~n8447 ;
  assign n8449 = ~n4814 & n8447 ;
  assign n8450 = ~n8448 & ~n8449 ;
  assign n8451 = n7453 & n8450 ;
  assign n8452 = ~n8426 & ~n8451 ;
  assign n8453 = n5563 & ~n8452 ;
  assign n8425 = n4814 & ~n7504 ;
  assign n8454 = n4793 & ~n7641 ;
  assign n8455 = ~n8425 & ~n8454 ;
  assign n8456 = ~n8453 & n8455 ;
  assign n8457 = ~n8434 & n8456 ;
  assign n8435 = n5990 & ~n7929 ;
  assign n8436 = ~n5990 & n7929 ;
  assign n8437 = ~n8435 & ~n8436 ;
  assign n8438 = n7453 & ~n8437 ;
  assign n8439 = ~n8426 & ~n8438 ;
  assign n8440 = n5526 & ~n8439 ;
  assign n8441 = n5990 & ~n7894 ;
  assign n8442 = ~n5990 & n7894 ;
  assign n8443 = ~n8441 & ~n8442 ;
  assign n8444 = n7453 & n8443 ;
  assign n8445 = ~n8426 & ~n8444 ;
  assign n8446 = n5329 & ~n8445 ;
  assign n8458 = ~n8440 & ~n8446 ;
  assign n8459 = n8457 & n8458 ;
  assign n8460 = n5583 & ~n8459 ;
  assign n8461 = ~n8424 & ~n8460 ;
  assign n8462 = \P1_state_reg[0]/NET0131  & ~n8461 ;
  assign n8422 = n4793 & n5786 ;
  assign n8423 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[18]/NET0131  ;
  assign n8463 = ~n8422 & ~n8423 ;
  assign n8464 = ~n8462 & n8463 ;
  assign n8467 = n4770 & n5585 ;
  assign n8469 = n4770 & ~n7453 ;
  assign n8470 = n4921 & ~n5269 ;
  assign n8471 = n5280 & ~n8470 ;
  assign n8472 = n5979 & n8471 ;
  assign n8473 = ~n5979 & ~n8471 ;
  assign n8474 = ~n8472 & ~n8473 ;
  assign n8475 = n7453 & ~n8474 ;
  assign n8476 = ~n8469 & ~n8475 ;
  assign n8477 = n5329 & ~n8476 ;
  assign n8478 = n5361 & n5362 ;
  assign n8479 = n4799 & ~n8478 ;
  assign n8480 = ~n5364 & ~n8479 ;
  assign n8481 = ~n4231 & ~n8480 ;
  assign n8482 = n4231 & n4879 ;
  assign n8483 = ~n8481 & ~n8482 ;
  assign n8484 = n7453 & n8483 ;
  assign n8485 = ~n8469 & ~n8484 ;
  assign n8486 = n5383 & ~n8485 ;
  assign n8487 = n5398 & ~n5455 ;
  assign n8488 = n5465 & ~n8487 ;
  assign n8489 = n5979 & n8488 ;
  assign n8490 = ~n5979 & ~n8488 ;
  assign n8491 = ~n8489 & ~n8490 ;
  assign n8492 = n7453 & n8491 ;
  assign n8493 = ~n8469 & ~n8492 ;
  assign n8494 = n5526 & ~n8493 ;
  assign n8495 = n4789 & ~n5544 ;
  assign n8496 = ~n8447 & ~n8495 ;
  assign n8497 = n7453 & n8496 ;
  assign n8498 = ~n8469 & ~n8497 ;
  assign n8499 = n5563 & ~n8498 ;
  assign n8468 = n4789 & ~n7504 ;
  assign n8500 = n4770 & ~n7641 ;
  assign n8501 = ~n8468 & ~n8500 ;
  assign n8502 = ~n8499 & n8501 ;
  assign n8503 = ~n8494 & n8502 ;
  assign n8504 = ~n8486 & n8503 ;
  assign n8505 = ~n8477 & n8504 ;
  assign n8506 = n5583 & ~n8505 ;
  assign n8507 = ~n8467 & ~n8506 ;
  assign n8508 = \P1_state_reg[0]/NET0131  & ~n8507 ;
  assign n8465 = n4770 & n5786 ;
  assign n8466 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[17]/NET0131  ;
  assign n8509 = ~n8465 & ~n8466 ;
  assign n8510 = ~n8508 & n8509 ;
  assign n8512 = n4722 & n5585 ;
  assign n8514 = n4722 & ~n7453 ;
  assign n8515 = n5987 & ~n7535 ;
  assign n8516 = ~n5987 & n7535 ;
  assign n8517 = ~n8515 & ~n8516 ;
  assign n8518 = n7453 & ~n8517 ;
  assign n8519 = ~n8514 & ~n8518 ;
  assign n8520 = n5526 & ~n8519 ;
  assign n8521 = n5987 & ~n7569 ;
  assign n8522 = ~n5987 & n7569 ;
  assign n8523 = ~n8521 & ~n8522 ;
  assign n8524 = n7453 & n8523 ;
  assign n8525 = ~n8514 & ~n8524 ;
  assign n8526 = n5329 & ~n8525 ;
  assign n8527 = n4763 & ~n7591 ;
  assign n8528 = ~n4763 & n7591 ;
  assign n8529 = ~n8527 & ~n8528 ;
  assign n8530 = ~n4231 & ~n8529 ;
  assign n8531 = n4231 & n4799 ;
  assign n8532 = ~n8530 & ~n8531 ;
  assign n8533 = n7453 & n8532 ;
  assign n8534 = ~n8514 & ~n8533 ;
  assign n8535 = n5383 & ~n8534 ;
  assign n8536 = n4745 & ~n8449 ;
  assign n8537 = n5528 & n8447 ;
  assign n8538 = ~n8536 & ~n8537 ;
  assign n8539 = n5563 & n8538 ;
  assign n8540 = n7453 & n8539 ;
  assign n8513 = n4722 & ~n7484 ;
  assign n8541 = n4745 & ~n7504 ;
  assign n8542 = ~n8513 & ~n8541 ;
  assign n8543 = ~n8540 & n8542 ;
  assign n8544 = ~n8535 & n8543 ;
  assign n8545 = ~n8526 & n8544 ;
  assign n8546 = ~n8520 & n8545 ;
  assign n8547 = n5583 & ~n8546 ;
  assign n8548 = ~n8512 & ~n8547 ;
  assign n8549 = \P1_state_reg[0]/NET0131  & ~n8548 ;
  assign n8511 = n4722 & n5786 ;
  assign n8550 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[19]/NET0131  ;
  assign n8551 = ~n8511 & ~n8550 ;
  assign n8552 = ~n8549 & n8551 ;
  assign n8555 = ~n1116 & n2145 ;
  assign n8556 = ~n1116 & ~n2163 ;
  assign n8570 = n1095 & ~n6539 ;
  assign n8571 = ~n2239 & ~n6540 ;
  assign n8572 = ~n8570 & n8571 ;
  assign n8573 = ~n1152 & n2239 ;
  assign n8574 = ~n8572 & ~n8573 ;
  assign n8575 = n2163 & ~n8574 ;
  assign n8576 = ~n8556 & ~n8575 ;
  assign n8577 = n737 & ~n8576 ;
  assign n8563 = ~n1116 & ~n2236 ;
  assign n8564 = n2074 & ~n5713 ;
  assign n8565 = ~n2074 & n5713 ;
  assign n8566 = ~n8564 & ~n8565 ;
  assign n8567 = n2236 & ~n8566 ;
  assign n8568 = ~n8563 & ~n8567 ;
  assign n8569 = n2234 & ~n8568 ;
  assign n8581 = ~n1137 & n2580 ;
  assign n8582 = ~n1116 & ~n2583 ;
  assign n8583 = ~n8581 & ~n8582 ;
  assign n8584 = ~n8569 & n8583 ;
  assign n8585 = ~n8577 & n8584 ;
  assign n8557 = n2074 & ~n5750 ;
  assign n8558 = ~n2074 & n5750 ;
  assign n8559 = ~n8557 & ~n8558 ;
  assign n8560 = n2163 & n8559 ;
  assign n8561 = ~n8556 & ~n8560 ;
  assign n8562 = n2393 & ~n8561 ;
  assign n8578 = n2236 & n8559 ;
  assign n8579 = ~n8563 & ~n8578 ;
  assign n8580 = n2391 & ~n8579 ;
  assign n8586 = ~n8562 & ~n8580 ;
  assign n8587 = n8585 & n8586 ;
  assign n8588 = n2147 & ~n8587 ;
  assign n8589 = ~n8555 & ~n8588 ;
  assign n8590 = \P1_state_reg[0]/NET0131  & ~n8589 ;
  assign n8553 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[18]/NET0131  ;
  assign n8554 = n765 & ~n1116 ;
  assign n8591 = ~n8553 & ~n8554 ;
  assign n8592 = ~n8590 & n8591 ;
  assign n8595 = ~n1146 & n2145 ;
  assign n8598 = ~n1146 & ~n2236 ;
  assign n8599 = n2078 & ~n2347 ;
  assign n8600 = ~n2078 & n2347 ;
  assign n8601 = ~n8599 & ~n8600 ;
  assign n8602 = n2236 & ~n8601 ;
  assign n8603 = ~n8598 & ~n8602 ;
  assign n8604 = n2391 & ~n8603 ;
  assign n8596 = ~n1166 & n2580 ;
  assign n8597 = ~n1146 & ~n2583 ;
  assign n8623 = ~n8596 & ~n8597 ;
  assign n8624 = ~n8604 & n8623 ;
  assign n8611 = ~n1146 & ~n2163 ;
  assign n8615 = n1121 & ~n2260 ;
  assign n8616 = ~n2239 & ~n6539 ;
  assign n8617 = ~n8615 & n8616 ;
  assign n8618 = ~n1197 & n2239 ;
  assign n8619 = ~n8617 & ~n8618 ;
  assign n8620 = n2163 & ~n8619 ;
  assign n8621 = ~n8611 & ~n8620 ;
  assign n8622 = n737 & ~n8621 ;
  assign n8605 = n2078 & ~n2199 ;
  assign n8606 = ~n2078 & n2199 ;
  assign n8607 = ~n8605 & ~n8606 ;
  assign n8608 = n2236 & n8607 ;
  assign n8609 = ~n8598 & ~n8608 ;
  assign n8610 = n2234 & ~n8609 ;
  assign n8612 = n2163 & ~n8601 ;
  assign n8613 = ~n8611 & ~n8612 ;
  assign n8614 = n2393 & ~n8613 ;
  assign n8625 = ~n8610 & ~n8614 ;
  assign n8626 = ~n8622 & n8625 ;
  assign n8627 = n8624 & n8626 ;
  assign n8628 = n2147 & ~n8627 ;
  assign n8629 = ~n8595 & ~n8628 ;
  assign n8630 = \P1_state_reg[0]/NET0131  & ~n8629 ;
  assign n8593 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[17]/NET0131  ;
  assign n8594 = n765 & ~n1146 ;
  assign n8631 = ~n8593 & ~n8594 ;
  assign n8632 = ~n8630 & n8631 ;
  assign n8633 = n4643 & n5585 ;
  assign n8643 = n7453 & ~n7860 ;
  assign n8635 = n7453 & n7831 ;
  assign n8634 = ~n4643 & ~n7453 ;
  assign n8636 = n5329 & ~n8634 ;
  assign n8637 = ~n8635 & n8636 ;
  assign n8638 = ~n7453 & ~n7865 ;
  assign n8639 = n7641 & ~n8638 ;
  assign n8640 = n5383 & ~n7453 ;
  assign n8641 = n8639 & ~n8640 ;
  assign n8642 = n4643 & ~n8641 ;
  assign n8644 = n4635 & ~n7504 ;
  assign n8645 = ~n8642 & ~n8644 ;
  assign n8646 = ~n8637 & n8645 ;
  assign n8647 = ~n8643 & n8646 ;
  assign n8648 = n5583 & ~n8647 ;
  assign n8649 = ~n8633 & ~n8648 ;
  assign n8650 = \P1_state_reg[0]/NET0131  & ~n8649 ;
  assign n8651 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[24]/NET0131  ;
  assign n8652 = n4643 & n5786 ;
  assign n8653 = ~n8651 & ~n8652 ;
  assign n8654 = ~n8650 & n8653 ;
  assign n8655 = n2883 & n6095 ;
  assign n8656 = ~n6207 & ~n6282 ;
  assign n8657 = n2883 & ~n8656 ;
  assign n8658 = ~n6568 & ~n8657 ;
  assign n8685 = ~n7142 & n7144 ;
  assign n8686 = n7149 & ~n8685 ;
  assign n8688 = ~n2890 & ~n8686 ;
  assign n8687 = n2890 & n8686 ;
  assign n8689 = n6282 & ~n8687 ;
  assign n8690 = ~n8688 & n8689 ;
  assign n8676 = ~n7176 & n7179 ;
  assign n8677 = n7168 & n7185 ;
  assign n8678 = ~n8676 & n8677 ;
  assign n8675 = ~n7182 & n7185 ;
  assign n8679 = n7161 & ~n8675 ;
  assign n8680 = ~n8678 & n8679 ;
  assign n8682 = ~n2890 & n8680 ;
  assign n8681 = n2890 & ~n8680 ;
  assign n8683 = n6207 & ~n8681 ;
  assign n8684 = ~n8682 & n8683 ;
  assign n8659 = ~n2942 & n6345 ;
  assign n8660 = ~n3588 & n8659 ;
  assign n8661 = ~n3294 & n8660 ;
  assign n8662 = n2830 & ~n8661 ;
  assign n8663 = n6346 & n8660 ;
  assign n8664 = n6359 & ~n8663 ;
  assign n8665 = ~n8662 & n8664 ;
  assign n8666 = n6303 & n6307 ;
  assign n8667 = n3283 & ~n8666 ;
  assign n8668 = n6303 & n6308 ;
  assign n8669 = ~n8667 & ~n8668 ;
  assign n8670 = ~n2713 & ~n8669 ;
  assign n8671 = n2713 & n3303 ;
  assign n8672 = n4011 & ~n8671 ;
  assign n8673 = ~n8670 & n8672 ;
  assign n8674 = ~n8665 & ~n8673 ;
  assign n8691 = n6568 & n8674 ;
  assign n8692 = ~n8684 & n8691 ;
  assign n8693 = ~n8690 & n8692 ;
  assign n8694 = ~n8658 & ~n8693 ;
  assign n8695 = n2883 & ~n6668 ;
  assign n8696 = n2830 & ~n6649 ;
  assign n8697 = ~n8695 & ~n8696 ;
  assign n8698 = ~n8694 & n8697 ;
  assign n8699 = n6097 & ~n8698 ;
  assign n8700 = ~n8655 & ~n8699 ;
  assign n8701 = \P1_state_reg[0]/NET0131  & ~n8700 ;
  assign n8702 = \P1_reg3_reg[22]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8703 = n2883 & n4130 ;
  assign n8704 = ~n8702 & ~n8703 ;
  assign n8705 = ~n8701 & n8704 ;
  assign n8706 = \P1_reg2_reg[31]/NET0131  & ~n6078 ;
  assign n8716 = ~n3500 & n6354 ;
  assign n8717 = n3467 & ~n8716 ;
  assign n8718 = ~n3467 & n8716 ;
  assign n8719 = ~n8717 & ~n8718 ;
  assign n8720 = n6113 & ~n8719 ;
  assign n8715 = ~\P1_reg2_reg[31]/NET0131  & ~n6113 ;
  assign n8721 = n6359 & ~n8715 ;
  assign n8722 = ~n8720 & n8721 ;
  assign n8712 = ~n3473 & n6320 ;
  assign n8713 = n4011 & n6113 ;
  assign n8714 = n8712 & n8713 ;
  assign n8707 = n6113 & n6365 ;
  assign n8708 = n3467 & n8707 ;
  assign n8709 = ~n4111 & ~n6113 ;
  assign n8710 = ~n6361 & ~n8709 ;
  assign n8711 = \P1_reg2_reg[31]/NET0131  & ~n8710 ;
  assign n8723 = ~n6367 & ~n8711 ;
  assign n8724 = ~n8708 & n8723 ;
  assign n8725 = ~n8714 & n8724 ;
  assign n8726 = ~n8722 & n8725 ;
  assign n8727 = n6097 & ~n8726 ;
  assign n8728 = \P1_reg2_reg[31]/NET0131  & n6095 ;
  assign n8729 = ~n8727 & ~n8728 ;
  assign n8730 = \P1_state_reg[0]/NET0131  & ~n8729 ;
  assign n8731 = ~n8706 & ~n8730 ;
  assign n8732 = n4680 & ~n7453 ;
  assign n8733 = ~n7886 & n7889 ;
  assign n8734 = n7879 & ~n8733 ;
  assign n8735 = n7892 & ~n8734 ;
  assign n8736 = n7895 & ~n8735 ;
  assign n8737 = n7900 & ~n8736 ;
  assign n8738 = n5983 & n8737 ;
  assign n8739 = ~n5983 & ~n8737 ;
  assign n8740 = ~n8738 & ~n8739 ;
  assign n8741 = n7453 & ~n8740 ;
  assign n8742 = ~n8732 & ~n8741 ;
  assign n8743 = n5329 & ~n8742 ;
  assign n8756 = n5366 & n8528 ;
  assign n8757 = n4665 & ~n8756 ;
  assign n8758 = ~n7593 & ~n8757 ;
  assign n8759 = ~n4231 & ~n8758 ;
  assign n8760 = n4231 & n4703 ;
  assign n8761 = ~n8759 & ~n8760 ;
  assign n8762 = n7453 & n8761 ;
  assign n8763 = ~n8732 & ~n8762 ;
  assign n8764 = n5383 & ~n8763 ;
  assign n8744 = ~n7920 & n7924 ;
  assign n8745 = n7921 & n7931 ;
  assign n8746 = ~n8744 & n8745 ;
  assign n8747 = ~n7927 & n7931 ;
  assign n8748 = n7936 & ~n8747 ;
  assign n8749 = ~n8746 & n8748 ;
  assign n8750 = n5983 & ~n8749 ;
  assign n8751 = ~n5983 & n8749 ;
  assign n8752 = ~n8750 & ~n8751 ;
  assign n8753 = n7453 & ~n8752 ;
  assign n8754 = ~n8732 & ~n8753 ;
  assign n8755 = n5526 & ~n8754 ;
  assign n8766 = n4675 & ~n7495 ;
  assign n8767 = ~n7496 & ~n8766 ;
  assign n8768 = n7453 & n8767 ;
  assign n8769 = ~n8732 & ~n8768 ;
  assign n8770 = n5563 & ~n8769 ;
  assign n8765 = n4675 & ~n7504 ;
  assign n8771 = n4680 & ~n7641 ;
  assign n8772 = ~n8765 & ~n8771 ;
  assign n8773 = ~n8770 & n8772 ;
  assign n8774 = ~n8755 & n8773 ;
  assign n8775 = ~n8764 & n8774 ;
  assign n8776 = ~n8743 & n8775 ;
  assign n8777 = n5583 & ~n8776 ;
  assign n8778 = n4680 & n5585 ;
  assign n8779 = ~n8777 & ~n8778 ;
  assign n8780 = \P1_state_reg[0]/NET0131  & ~n8779 ;
  assign n8781 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[22]/NET0131  ;
  assign n8782 = n4680 & n5786 ;
  assign n8783 = ~n8781 & ~n8782 ;
  assign n8784 = ~n8780 & n8783 ;
  assign n8787 = n4597 & n5585 ;
  assign n8788 = n4597 & ~n7453 ;
  assign n8792 = n7453 & ~n7909 ;
  assign n8793 = ~n8788 & ~n8792 ;
  assign n8794 = n5329 & ~n8793 ;
  assign n8789 = n7453 & n7943 ;
  assign n8790 = ~n8788 & ~n8789 ;
  assign n8791 = n5526 & ~n8790 ;
  assign n8796 = n7453 & n7953 ;
  assign n8797 = ~n8788 & ~n8796 ;
  assign n8798 = n5383 & ~n8797 ;
  assign n8799 = n7453 & n7960 ;
  assign n8795 = n4597 & ~n7484 ;
  assign n8800 = n4592 & ~n7504 ;
  assign n8801 = ~n8795 & ~n8800 ;
  assign n8802 = ~n8799 & n8801 ;
  assign n8803 = ~n8798 & n8802 ;
  assign n8804 = ~n8791 & n8803 ;
  assign n8805 = ~n8794 & n8804 ;
  assign n8806 = n5583 & ~n8805 ;
  assign n8807 = ~n8787 & ~n8806 ;
  assign n8808 = \P1_state_reg[0]/NET0131  & ~n8807 ;
  assign n8785 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[26]/NET0131  ;
  assign n8786 = n4597 & n5786 ;
  assign n8809 = ~n8785 & ~n8786 ;
  assign n8810 = ~n8808 & n8809 ;
  assign n8811 = \P2_reg2_reg[31]/NET0131  & ~n5589 ;
  assign n8812 = \P2_reg2_reg[31]/NET0131  & n5585 ;
  assign n8813 = \P2_reg2_reg[31]/NET0131  & ~n4219 ;
  assign n8814 = n5557 & ~n5895 ;
  assign n8815 = n5879 & ~n8814 ;
  assign n8816 = ~n5879 & n8814 ;
  assign n8817 = ~n8815 & ~n8816 ;
  assign n8818 = n4219 & n8817 ;
  assign n8819 = ~n8813 & ~n8818 ;
  assign n8820 = n5563 & ~n8819 ;
  assign n8821 = ~n5339 & n5373 ;
  assign n8822 = n7948 & n8821 ;
  assign n8823 = ~n5333 & ~n5345 ;
  assign n8824 = ~n8822 & n8823 ;
  assign n8825 = n4219 & n5383 ;
  assign n8826 = n8824 & n8825 ;
  assign n8827 = n4219 & n5879 ;
  assign n8828 = ~n8813 & ~n8827 ;
  assign n8829 = n5565 & ~n8828 ;
  assign n8830 = ~n4219 & ~n5562 ;
  assign n8831 = ~n5568 & ~n8830 ;
  assign n8832 = \P2_reg2_reg[31]/NET0131  & ~n8831 ;
  assign n8833 = ~n5575 & ~n8832 ;
  assign n8834 = ~n8829 & n8833 ;
  assign n8835 = ~n8826 & n8834 ;
  assign n8836 = ~n8820 & n8835 ;
  assign n8837 = n5583 & ~n8836 ;
  assign n8838 = ~n8812 & ~n8837 ;
  assign n8839 = \P1_state_reg[0]/NET0131  & ~n8838 ;
  assign n8840 = ~n8811 & ~n8839 ;
  assign n8841 = \P1_reg1_reg[24]/NET0131  & ~n6078 ;
  assign n8842 = \P1_reg1_reg[24]/NET0131  & n6095 ;
  assign n8845 = \P1_reg1_reg[24]/NET0131  & ~n6683 ;
  assign n8849 = n6683 & ~n7031 ;
  assign n8850 = ~n8845 & ~n8849 ;
  assign n8851 = n6207 & ~n8850 ;
  assign n8846 = n6683 & ~n6964 ;
  assign n8847 = ~n8845 & ~n8846 ;
  assign n8848 = n6282 & ~n8847 ;
  assign n8843 = \P1_reg1_reg[24]/NET0131  & ~n7808 ;
  assign n8844 = n6683 & ~n8151 ;
  assign n8852 = ~n8843 & ~n8844 ;
  assign n8853 = ~n8848 & n8852 ;
  assign n8854 = ~n8851 & n8853 ;
  assign n8855 = n6097 & ~n8854 ;
  assign n8856 = ~n8842 & ~n8855 ;
  assign n8857 = \P1_state_reg[0]/NET0131  & ~n8856 ;
  assign n8858 = ~n8841 & ~n8857 ;
  assign n8859 = \P1_reg1_reg[26]/NET0131  & ~n6078 ;
  assign n8860 = \P1_reg1_reg[26]/NET0131  & n6095 ;
  assign n8861 = \P1_reg1_reg[26]/NET0131  & ~n6683 ;
  assign n8862 = n6683 & ~n7156 ;
  assign n8863 = ~n8861 & ~n8862 ;
  assign n8864 = n6282 & ~n8863 ;
  assign n8865 = n6683 & ~n7192 ;
  assign n8866 = ~n8861 & ~n8865 ;
  assign n8867 = n6207 & ~n8866 ;
  assign n8868 = ~n7204 & ~n8114 ;
  assign n8869 = n6683 & ~n8868 ;
  assign n8870 = n6683 & ~n7200 ;
  assign n8871 = ~n8861 & ~n8870 ;
  assign n8872 = n4011 & ~n8871 ;
  assign n8873 = \P1_reg1_reg[26]/NET0131  & ~n6695 ;
  assign n8874 = ~n8872 & ~n8873 ;
  assign n8875 = ~n8869 & n8874 ;
  assign n8876 = ~n8867 & n8875 ;
  assign n8877 = ~n8864 & n8876 ;
  assign n8878 = n6097 & ~n8877 ;
  assign n8879 = ~n8860 & ~n8878 ;
  assign n8880 = \P1_state_reg[0]/NET0131  & ~n8879 ;
  assign n8881 = ~n8859 & ~n8880 ;
  assign n8882 = \P2_reg0_reg[25]/NET0131  & ~n5589 ;
  assign n8883 = \P2_reg0_reg[25]/NET0131  & n5585 ;
  assign n8889 = n6706 & ~n8005 ;
  assign n8884 = ~n5329 & ~n5526 ;
  assign n8885 = ~n6706 & ~n8884 ;
  assign n8886 = n6717 & ~n8885 ;
  assign n8887 = ~n7984 & n8886 ;
  assign n8888 = \P2_reg0_reg[25]/NET0131  & ~n8887 ;
  assign n8890 = n5329 & n6706 ;
  assign n8891 = ~n7465 & n8890 ;
  assign n8892 = ~n8888 & ~n8891 ;
  assign n8893 = ~n8889 & n8892 ;
  assign n8894 = n5583 & ~n8893 ;
  assign n8895 = ~n8883 & ~n8894 ;
  assign n8896 = \P1_state_reg[0]/NET0131  & ~n8895 ;
  assign n8897 = ~n8882 & ~n8896 ;
  assign n8898 = n5329 & ~n6380 ;
  assign n8899 = ~n5582 & n5589 ;
  assign n8900 = n6398 & n8899 ;
  assign n8901 = ~n8898 & n8900 ;
  assign n8902 = ~n7997 & n8901 ;
  assign n8903 = \P2_reg1_reg[22]/NET0131  & ~n8902 ;
  assign n8904 = n5329 & ~n8740 ;
  assign n8906 = n5383 & n8761 ;
  assign n8905 = n5526 & ~n8752 ;
  assign n8907 = n4675 & n5565 ;
  assign n8908 = n5563 & n8767 ;
  assign n8909 = ~n8907 & ~n8908 ;
  assign n8910 = ~n8905 & n8909 ;
  assign n8911 = ~n8906 & n8910 ;
  assign n8912 = ~n8904 & n8911 ;
  assign n8913 = n6380 & n8899 ;
  assign n8914 = ~n8912 & n8913 ;
  assign n8915 = ~n8903 & ~n8914 ;
  assign n8916 = \P2_reg1_reg[24]/NET0131  & ~n5589 ;
  assign n8917 = \P2_reg1_reg[24]/NET0131  & n5585 ;
  assign n8918 = n7998 & ~n8898 ;
  assign n8919 = \P2_reg1_reg[24]/NET0131  & ~n8918 ;
  assign n8920 = n5329 & ~n7831 ;
  assign n8921 = n7861 & ~n8920 ;
  assign n8922 = n6380 & ~n8921 ;
  assign n8923 = ~n8919 & ~n8922 ;
  assign n8924 = n5583 & ~n8923 ;
  assign n8925 = ~n8917 & ~n8924 ;
  assign n8926 = \P1_state_reg[0]/NET0131  & ~n8925 ;
  assign n8927 = ~n8916 & ~n8926 ;
  assign n8928 = \P2_reg1_reg[26]/NET0131  & ~n5589 ;
  assign n8929 = \P2_reg1_reg[26]/NET0131  & n5585 ;
  assign n8930 = \P2_reg1_reg[26]/NET0131  & ~n6380 ;
  assign n8934 = n6380 & n7943 ;
  assign n8935 = ~n8930 & ~n8934 ;
  assign n8936 = n5526 & ~n8935 ;
  assign n8931 = n6380 & ~n7909 ;
  assign n8932 = ~n8930 & ~n8931 ;
  assign n8933 = n5329 & ~n8932 ;
  assign n8938 = n6380 & n7953 ;
  assign n8939 = ~n8930 & ~n8938 ;
  assign n8940 = n5383 & ~n8939 ;
  assign n8937 = \P2_reg1_reg[26]/NET0131  & ~n6397 ;
  assign n8941 = n6380 & ~n7961 ;
  assign n8942 = ~n8937 & ~n8941 ;
  assign n8943 = ~n8940 & n8942 ;
  assign n8944 = ~n8933 & n8943 ;
  assign n8945 = ~n8936 & n8944 ;
  assign n8946 = n5583 & ~n8945 ;
  assign n8947 = ~n8929 & ~n8946 ;
  assign n8948 = \P1_state_reg[0]/NET0131  & ~n8947 ;
  assign n8949 = ~n8928 & ~n8948 ;
  assign n8950 = \P1_reg2_reg[25]/NET0131  & ~n6078 ;
  assign n8951 = \P1_reg2_reg[25]/NET0131  & n6095 ;
  assign n8959 = \P1_reg2_reg[25]/NET0131  & ~n6113 ;
  assign n8963 = n6113 & ~n7093 ;
  assign n8964 = ~n8959 & ~n8963 ;
  assign n8965 = n6207 & ~n8964 ;
  assign n8960 = n6113 & ~n7079 ;
  assign n8961 = ~n8959 & ~n8960 ;
  assign n8962 = n6282 & ~n8961 ;
  assign n8952 = n6113 & ~n7777 ;
  assign n8953 = n3172 & n4112 ;
  assign n8954 = ~n6113 & n6365 ;
  assign n8955 = ~n6361 & ~n8954 ;
  assign n8956 = ~n6113 & n6427 ;
  assign n8957 = n8955 & ~n8956 ;
  assign n8958 = \P1_reg2_reg[25]/NET0131  & ~n8957 ;
  assign n8966 = ~n8953 & ~n8958 ;
  assign n8967 = ~n8952 & n8966 ;
  assign n8968 = ~n8962 & n8967 ;
  assign n8969 = ~n8965 & n8968 ;
  assign n8970 = n6097 & ~n8969 ;
  assign n8971 = ~n8951 & ~n8970 ;
  assign n8972 = \P1_state_reg[0]/NET0131  & ~n8971 ;
  assign n8973 = ~n8950 & ~n8972 ;
  assign n8974 = \P2_reg2_reg[25]/NET0131  & ~n5589 ;
  assign n8975 = \P2_reg2_reg[25]/NET0131  & n5585 ;
  assign n8976 = \P2_reg2_reg[25]/NET0131  & ~n4219 ;
  assign n8977 = n4219 & ~n7465 ;
  assign n8978 = ~n8976 & ~n8977 ;
  assign n8979 = n5329 & ~n8978 ;
  assign n8984 = n4219 & n7491 ;
  assign n8985 = ~n8976 & ~n8984 ;
  assign n8986 = n5383 & ~n8985 ;
  assign n8980 = n4219 & ~n7479 ;
  assign n8981 = ~n8976 & ~n8980 ;
  assign n8982 = n5526 & ~n8981 ;
  assign n8987 = n4219 & n7500 ;
  assign n8988 = ~n8976 & ~n8987 ;
  assign n8989 = n5563 & ~n8988 ;
  assign n8991 = n4219 & n8000 ;
  assign n8983 = \P2_reg2_reg[25]/NET0131  & ~n5570 ;
  assign n8990 = n4618 & n5574 ;
  assign n8992 = ~n8983 & ~n8990 ;
  assign n8993 = ~n8991 & n8992 ;
  assign n8994 = ~n8989 & n8993 ;
  assign n8995 = ~n8982 & n8994 ;
  assign n8996 = ~n8986 & n8995 ;
  assign n8997 = ~n8979 & n8996 ;
  assign n8998 = n5583 & ~n8997 ;
  assign n8999 = ~n8975 & ~n8998 ;
  assign n9000 = \P1_state_reg[0]/NET0131  & ~n8999 ;
  assign n9001 = ~n8974 & ~n9000 ;
  assign n9002 = \P2_reg2_reg[26]/NET0131  & ~n5589 ;
  assign n9003 = \P2_reg2_reg[26]/NET0131  & n5585 ;
  assign n9004 = \P2_reg2_reg[26]/NET0131  & ~n4219 ;
  assign n9008 = n4219 & n7943 ;
  assign n9009 = ~n9004 & ~n9008 ;
  assign n9010 = n5526 & ~n9009 ;
  assign n9005 = n4219 & ~n7909 ;
  assign n9006 = ~n9004 & ~n9005 ;
  assign n9007 = n5329 & ~n9006 ;
  assign n9012 = n4219 & n7953 ;
  assign n9013 = ~n9004 & ~n9012 ;
  assign n9014 = n5383 & ~n9013 ;
  assign n9016 = n4219 & ~n7961 ;
  assign n9011 = \P2_reg2_reg[26]/NET0131  & ~n6839 ;
  assign n9015 = n4597 & n5574 ;
  assign n9017 = ~n9011 & ~n9015 ;
  assign n9018 = ~n9016 & n9017 ;
  assign n9019 = ~n9014 & n9018 ;
  assign n9020 = ~n9007 & n9019 ;
  assign n9021 = ~n9010 & n9020 ;
  assign n9022 = n5583 & ~n9021 ;
  assign n9023 = ~n9003 & ~n9022 ;
  assign n9024 = \P1_state_reg[0]/NET0131  & ~n9023 ;
  assign n9025 = ~n9002 & ~n9024 ;
  assign n9026 = \P1_reg0_reg[25]/NET0131  & ~n6078 ;
  assign n9027 = \P1_reg0_reg[25]/NET0131  & n6095 ;
  assign n9030 = \P1_reg0_reg[25]/NET0131  & ~n6409 ;
  assign n9034 = n6409 & ~n7093 ;
  assign n9035 = ~n9030 & ~n9034 ;
  assign n9036 = n6207 & ~n9035 ;
  assign n9031 = n6409 & ~n7079 ;
  assign n9032 = ~n9030 & ~n9031 ;
  assign n9033 = n6282 & ~n9032 ;
  assign n9028 = \P1_reg0_reg[25]/NET0131  & ~n6429 ;
  assign n9029 = n6409 & ~n7777 ;
  assign n9037 = ~n9028 & ~n9029 ;
  assign n9038 = ~n9033 & n9037 ;
  assign n9039 = ~n9036 & n9038 ;
  assign n9040 = n6097 & ~n9039 ;
  assign n9041 = ~n9027 & ~n9040 ;
  assign n9042 = \P1_state_reg[0]/NET0131  & ~n9041 ;
  assign n9043 = ~n9026 & ~n9042 ;
  assign n9044 = \P1_state_reg[0]/NET0131  & n6097 ;
  assign n9045 = n6683 & n9044 ;
  assign n9046 = n2830 & n6365 ;
  assign n9047 = n8674 & ~n9046 ;
  assign n9048 = ~n8684 & n9047 ;
  assign n9049 = ~n8690 & n9048 ;
  assign n9050 = n9045 & ~n9049 ;
  assign n9051 = ~n6683 & ~n8059 ;
  assign n9052 = n9044 & ~n9051 ;
  assign n9053 = n7806 & n9052 ;
  assign n9054 = \P1_reg1_reg[22]/NET0131  & ~n9053 ;
  assign n9055 = ~n9050 & ~n9054 ;
  assign n9057 = n3645 & n6095 ;
  assign n9063 = ~n3329 & n6293 ;
  assign n9064 = ~n3677 & n9063 ;
  assign n9065 = n6294 & n9064 ;
  assign n9066 = n3354 & ~n9065 ;
  assign n9067 = n6296 & n9063 ;
  assign n9068 = ~n9066 & ~n9067 ;
  assign n9069 = ~n2713 & ~n9068 ;
  assign n9070 = n2713 & n3255 ;
  assign n9071 = ~n9069 & ~n9070 ;
  assign n9072 = n4011 & n9071 ;
  assign n9059 = ~n3641 & n6338 ;
  assign n9060 = n3641 & ~n6338 ;
  assign n9061 = ~n9059 & ~n9060 ;
  assign n9062 = n6359 & n9061 ;
  assign n9074 = n3653 & n4055 ;
  assign n9073 = ~n3653 & ~n4055 ;
  assign n9075 = n6282 & ~n9073 ;
  assign n9076 = ~n9074 & n9075 ;
  assign n9078 = ~n3653 & n7673 ;
  assign n9077 = n3653 & ~n7673 ;
  assign n9079 = n6207 & ~n9077 ;
  assign n9080 = ~n9078 & n9079 ;
  assign n9081 = ~n9076 & ~n9080 ;
  assign n9082 = ~n9062 & n9081 ;
  assign n9083 = ~n9072 & n9082 ;
  assign n9084 = n6568 & ~n9083 ;
  assign n9058 = n3641 & ~n6649 ;
  assign n9085 = ~n6568 & ~n8060 ;
  assign n9086 = ~n6361 & ~n9085 ;
  assign n9087 = n3645 & ~n9086 ;
  assign n9088 = ~n9058 & ~n9087 ;
  assign n9089 = ~n9084 & n9088 ;
  assign n9090 = n6097 & ~n9089 ;
  assign n9091 = ~n9057 & ~n9090 ;
  assign n9092 = \P1_state_reg[0]/NET0131  & ~n9091 ;
  assign n9056 = n3645 & n4130 ;
  assign n9093 = \P1_reg3_reg[12]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9094 = ~n9056 & ~n9093 ;
  assign n9095 = ~n9092 & n9094 ;
  assign n9098 = n3199 & n6095 ;
  assign n9100 = n3199 & ~n6568 ;
  assign n9101 = n7007 & ~n7673 ;
  assign n9102 = n7015 & ~n9101 ;
  assign n9103 = n3206 & n9102 ;
  assign n9104 = ~n3206 & ~n9102 ;
  assign n9105 = ~n9103 & ~n9104 ;
  assign n9106 = n6568 & ~n9105 ;
  assign n9107 = ~n9100 & ~n9106 ;
  assign n9108 = n6207 & ~n9107 ;
  assign n9116 = n3206 & ~n4057 ;
  assign n9117 = ~n3206 & n4057 ;
  assign n9118 = ~n9116 & ~n9117 ;
  assign n9119 = n6568 & ~n9118 ;
  assign n9120 = ~n9100 & ~n9119 ;
  assign n9121 = n6282 & ~n9120 ;
  assign n9122 = ~n3081 & n6301 ;
  assign n9123 = n3081 & ~n6301 ;
  assign n9124 = ~n9122 & ~n9123 ;
  assign n9125 = ~n2713 & ~n9124 ;
  assign n9126 = n2713 & n3623 ;
  assign n9127 = ~n9125 & ~n9126 ;
  assign n9128 = n6568 & n9127 ;
  assign n9129 = ~n9100 & ~n9128 ;
  assign n9130 = n4011 & ~n9129 ;
  assign n9109 = ~n3614 & n6341 ;
  assign n9110 = ~n3194 & n9109 ;
  assign n9111 = n3194 & ~n9109 ;
  assign n9112 = ~n9110 & ~n9111 ;
  assign n9113 = n6568 & n9112 ;
  assign n9114 = ~n9100 & ~n9113 ;
  assign n9115 = n6359 & ~n9114 ;
  assign n9099 = n3194 & ~n6649 ;
  assign n9131 = n3199 & ~n6666 ;
  assign n9132 = ~n9099 & ~n9131 ;
  assign n9133 = ~n9115 & n9132 ;
  assign n9134 = ~n9130 & n9133 ;
  assign n9135 = ~n9121 & n9134 ;
  assign n9136 = ~n9108 & n9135 ;
  assign n9137 = n6097 & ~n9136 ;
  assign n9138 = ~n9098 & ~n9137 ;
  assign n9139 = \P1_state_reg[0]/NET0131  & ~n9138 ;
  assign n9096 = \P1_reg3_reg[16]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9097 = n3199 & n4130 ;
  assign n9140 = ~n9096 & ~n9097 ;
  assign n9141 = ~n9139 & n9140 ;
  assign n9144 = ~n1193 & n2145 ;
  assign n9158 = ~n1193 & ~n2236 ;
  assign n9170 = ~n2013 & n2061 ;
  assign n9171 = n2013 & ~n2061 ;
  assign n9172 = ~n9170 & ~n9171 ;
  assign n9173 = n2236 & ~n9172 ;
  assign n9174 = ~n9158 & ~n9173 ;
  assign n9175 = n2234 & ~n9174 ;
  assign n9146 = ~n1193 & ~n2163 ;
  assign n9147 = ~n1521 & n2239 ;
  assign n9148 = ~n1569 & n2255 ;
  assign n9149 = n2256 & n9148 ;
  assign n9150 = ~n1197 & n9149 ;
  assign n9151 = n1152 & ~n9150 ;
  assign n9152 = ~n2239 & ~n2260 ;
  assign n9153 = ~n9151 & n9152 ;
  assign n9154 = ~n9147 & ~n9153 ;
  assign n9155 = n2163 & ~n9154 ;
  assign n9156 = ~n9146 & ~n9155 ;
  assign n9157 = n737 & ~n9156 ;
  assign n9145 = ~n1185 & n2580 ;
  assign n9176 = ~n1193 & ~n2583 ;
  assign n9177 = ~n9145 & ~n9176 ;
  assign n9178 = ~n9157 & n9177 ;
  assign n9179 = ~n9175 & n9178 ;
  assign n9159 = ~n2468 & n2473 ;
  assign n9160 = n2480 & ~n9159 ;
  assign n9161 = n2061 & ~n9160 ;
  assign n9162 = ~n2061 & n9160 ;
  assign n9163 = ~n9161 & ~n9162 ;
  assign n9164 = n2236 & n9163 ;
  assign n9165 = ~n9158 & ~n9164 ;
  assign n9166 = n2391 & ~n9165 ;
  assign n9167 = n2163 & n9163 ;
  assign n9168 = ~n9146 & ~n9167 ;
  assign n9169 = n2393 & ~n9168 ;
  assign n9180 = ~n9166 & ~n9169 ;
  assign n9181 = n9179 & n9180 ;
  assign n9182 = n2147 & ~n9181 ;
  assign n9183 = ~n9144 & ~n9182 ;
  assign n9184 = \P1_state_reg[0]/NET0131  & ~n9183 ;
  assign n9142 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[16]/NET0131  ;
  assign n9143 = n765 & ~n1193 ;
  assign n9185 = ~n9142 & ~n9143 ;
  assign n9186 = ~n9184 & n9185 ;
  assign n9187 = \P1_reg3_reg[18]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9190 = n3102 & ~n6568 ;
  assign n9191 = n3112 & ~n7142 ;
  assign n9192 = ~n3112 & n7142 ;
  assign n9193 = ~n9191 & ~n9192 ;
  assign n9194 = n6568 & ~n9193 ;
  assign n9195 = ~n9190 & ~n9194 ;
  assign n9196 = n6282 & ~n9195 ;
  assign n9203 = n3112 & ~n7184 ;
  assign n9204 = ~n3112 & n7184 ;
  assign n9205 = ~n9203 & ~n9204 ;
  assign n9206 = n6568 & n9205 ;
  assign n9207 = ~n9190 & ~n9206 ;
  assign n9208 = n6207 & ~n9207 ;
  assign n9197 = ~n3072 & n9110 ;
  assign n9198 = n3100 & ~n9197 ;
  assign n9199 = ~n6345 & ~n9198 ;
  assign n9200 = n6568 & n9199 ;
  assign n9201 = ~n9190 & ~n9200 ;
  assign n9202 = n6359 & ~n9201 ;
  assign n9209 = ~n2952 & n6303 ;
  assign n9210 = n2952 & ~n6303 ;
  assign n9211 = ~n9209 & ~n9210 ;
  assign n9212 = ~n2713 & ~n9211 ;
  assign n9213 = n2713 & n3081 ;
  assign n9214 = ~n9212 & ~n9213 ;
  assign n9215 = n6568 & n9214 ;
  assign n9216 = ~n9190 & ~n9215 ;
  assign n9217 = n4011 & ~n9216 ;
  assign n9189 = n3100 & ~n6649 ;
  assign n9218 = n3102 & ~n6666 ;
  assign n9219 = n6097 & ~n9218 ;
  assign n9220 = ~n9189 & n9219 ;
  assign n9221 = ~n9217 & n9220 ;
  assign n9222 = ~n9202 & n9221 ;
  assign n9223 = ~n9208 & n9222 ;
  assign n9224 = ~n9196 & n9223 ;
  assign n9188 = ~n3102 & ~n6097 ;
  assign n9225 = \P1_state_reg[0]/NET0131  & ~n9188 ;
  assign n9226 = ~n9224 & n9225 ;
  assign n9227 = ~n9187 & ~n9226 ;
  assign n9228 = \P1_reg3_reg[19]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9235 = n2955 & ~n6589 ;
  assign n9236 = ~n2955 & n6589 ;
  assign n9237 = ~n9235 & ~n9236 ;
  assign n9238 = n6282 & ~n9237 ;
  assign n9232 = ~n2955 & n6627 ;
  assign n9231 = n2955 & ~n6627 ;
  assign n9233 = n6207 & ~n9231 ;
  assign n9234 = ~n9232 & n9233 ;
  assign n9239 = n3597 & ~n9209 ;
  assign n9240 = ~n3597 & n9209 ;
  assign n9241 = ~n9239 & ~n9240 ;
  assign n9242 = ~n2713 & ~n9241 ;
  assign n9243 = n2713 & n3109 ;
  assign n9244 = n4011 & ~n9243 ;
  assign n9245 = ~n9242 & n9244 ;
  assign n9246 = n2942 & ~n6345 ;
  assign n9247 = n6359 & ~n8659 ;
  assign n9248 = ~n9246 & n9247 ;
  assign n9249 = ~n9245 & ~n9248 ;
  assign n9250 = ~n9234 & n9249 ;
  assign n9251 = ~n9238 & n9250 ;
  assign n9252 = n6568 & ~n9251 ;
  assign n9230 = n2942 & ~n6649 ;
  assign n9253 = n2945 & ~n9086 ;
  assign n9254 = n6097 & ~n9253 ;
  assign n9255 = ~n9230 & n9254 ;
  assign n9256 = ~n9252 & n9255 ;
  assign n9229 = ~n2945 & ~n6097 ;
  assign n9257 = \P1_state_reg[0]/NET0131  & ~n9229 ;
  assign n9258 = ~n9256 & n9257 ;
  assign n9259 = ~n9228 & ~n9258 ;
  assign n9262 = n4757 & n5585 ;
  assign n9264 = n4757 & ~n7453 ;
  assign n9271 = ~n4703 & n7837 ;
  assign n9272 = n4703 & ~n7837 ;
  assign n9273 = ~n9271 & ~n9272 ;
  assign n9274 = ~n4231 & ~n9273 ;
  assign n9275 = n4231 & n4728 ;
  assign n9276 = ~n9274 & ~n9275 ;
  assign n9277 = n7453 & n9276 ;
  assign n9278 = ~n9264 & ~n9277 ;
  assign n9279 = n5383 & ~n9278 ;
  assign n9265 = n5978 & n6778 ;
  assign n9266 = ~n5978 & ~n6778 ;
  assign n9267 = ~n9265 & ~n9266 ;
  assign n9268 = n7453 & ~n9267 ;
  assign n9269 = ~n9264 & ~n9268 ;
  assign n9270 = n5329 & ~n9269 ;
  assign n9280 = n5978 & ~n6810 ;
  assign n9281 = ~n5978 & n6810 ;
  assign n9282 = ~n9280 & ~n9281 ;
  assign n9283 = n7453 & ~n9282 ;
  assign n9284 = ~n9264 & ~n9283 ;
  assign n9285 = n5526 & ~n9284 ;
  assign n9286 = n4754 & ~n8537 ;
  assign n9287 = ~n5547 & ~n9286 ;
  assign n9288 = n7453 & n9287 ;
  assign n9289 = ~n9264 & ~n9288 ;
  assign n9290 = n5563 & ~n9289 ;
  assign n9263 = n4754 & ~n7504 ;
  assign n9291 = n4757 & ~n7641 ;
  assign n9292 = ~n9263 & ~n9291 ;
  assign n9293 = ~n9290 & n9292 ;
  assign n9294 = ~n9285 & n9293 ;
  assign n9295 = ~n9270 & n9294 ;
  assign n9296 = ~n9279 & n9295 ;
  assign n9297 = n5583 & ~n9296 ;
  assign n9298 = ~n9262 & ~n9297 ;
  assign n9299 = \P1_state_reg[0]/NET0131  & ~n9298 ;
  assign n9260 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[20]/NET0131  ;
  assign n9261 = n4757 & n5786 ;
  assign n9300 = ~n9260 & ~n9261 ;
  assign n9301 = ~n9299 & n9300 ;
  assign n9304 = n3299 & n6095 ;
  assign n9306 = n3299 & ~n6568 ;
  assign n9328 = n3294 & ~n8660 ;
  assign n9329 = ~n8661 & ~n9328 ;
  assign n9330 = n6568 & n9329 ;
  assign n9331 = ~n9306 & ~n9330 ;
  assign n9332 = n6359 & ~n9331 ;
  assign n9316 = n3306 & ~n6255 ;
  assign n9317 = ~n3306 & n6255 ;
  assign n9318 = ~n9316 & ~n9317 ;
  assign n9319 = n6568 & ~n9318 ;
  assign n9320 = ~n9306 & ~n9319 ;
  assign n9321 = n6282 & ~n9320 ;
  assign n9305 = n3299 & ~n6666 ;
  assign n9333 = n3294 & ~n6649 ;
  assign n9334 = ~n9305 & ~n9333 ;
  assign n9335 = ~n9321 & n9334 ;
  assign n9336 = ~n9332 & n9335 ;
  assign n9307 = n6305 & n9209 ;
  assign n9308 = n2887 & ~n9307 ;
  assign n9309 = ~n8666 & ~n9308 ;
  assign n9310 = ~n2713 & ~n9309 ;
  assign n9311 = n2713 & n3597 ;
  assign n9312 = ~n9310 & ~n9311 ;
  assign n9313 = n6568 & n9312 ;
  assign n9314 = ~n9306 & ~n9313 ;
  assign n9315 = n4011 & ~n9314 ;
  assign n9322 = n3306 & n6177 ;
  assign n9323 = ~n3306 & ~n6177 ;
  assign n9324 = ~n9322 & ~n9323 ;
  assign n9325 = n6568 & ~n9324 ;
  assign n9326 = ~n9306 & ~n9325 ;
  assign n9327 = n6207 & ~n9326 ;
  assign n9337 = ~n9315 & ~n9327 ;
  assign n9338 = n9336 & n9337 ;
  assign n9339 = n6097 & ~n9338 ;
  assign n9340 = ~n9304 & ~n9339 ;
  assign n9341 = \P1_state_reg[0]/NET0131  & ~n9340 ;
  assign n9302 = \P1_reg3_reg[21]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9303 = n3299 & n4130 ;
  assign n9342 = ~n9302 & ~n9303 ;
  assign n9343 = ~n9341 & n9342 ;
  assign n9344 = \P1_reg2_reg[21]/NET0131  & ~n6078 ;
  assign n9345 = \P1_reg2_reg[21]/NET0131  & n6095 ;
  assign n9348 = \P1_reg2_reg[21]/NET0131  & ~n6113 ;
  assign n9358 = n6113 & n9329 ;
  assign n9359 = ~n9348 & ~n9358 ;
  assign n9360 = n6359 & ~n9359 ;
  assign n9352 = n6113 & ~n9318 ;
  assign n9353 = ~n9348 & ~n9352 ;
  assign n9354 = n6282 & ~n9353 ;
  assign n9346 = n3294 & n6365 ;
  assign n9347 = n6113 & n9346 ;
  assign n9361 = n3299 & n4112 ;
  assign n9362 = \P1_reg2_reg[21]/NET0131  & ~n8955 ;
  assign n9363 = ~n9361 & ~n9362 ;
  assign n9364 = ~n9347 & n9363 ;
  assign n9365 = ~n9354 & n9364 ;
  assign n9366 = ~n9360 & n9365 ;
  assign n9349 = n6113 & n9312 ;
  assign n9350 = ~n9348 & ~n9349 ;
  assign n9351 = n4011 & ~n9350 ;
  assign n9355 = n6113 & ~n9324 ;
  assign n9356 = ~n9348 & ~n9355 ;
  assign n9357 = n6207 & ~n9356 ;
  assign n9367 = ~n9351 & ~n9357 ;
  assign n9368 = n9366 & n9367 ;
  assign n9369 = n6097 & ~n9368 ;
  assign n9370 = ~n9345 & ~n9369 ;
  assign n9371 = \P1_state_reg[0]/NET0131  & ~n9370 ;
  assign n9372 = ~n9344 & ~n9371 ;
  assign n9374 = n4697 & n5585 ;
  assign n9393 = ~n5293 & n5989 ;
  assign n9392 = n5293 & ~n5989 ;
  assign n9394 = n5329 & ~n9392 ;
  assign n9395 = ~n9393 & n9394 ;
  assign n9385 = n4694 & ~n5547 ;
  assign n9386 = n5563 & ~n7495 ;
  assign n9387 = ~n9385 & n9386 ;
  assign n9389 = ~n5478 & ~n5989 ;
  assign n9388 = n5478 & n5989 ;
  assign n9390 = n5526 & ~n9388 ;
  assign n9391 = ~n9389 & n9390 ;
  assign n9396 = ~n9387 & ~n9391 ;
  assign n9397 = ~n9395 & n9396 ;
  assign n9398 = n7453 & ~n9397 ;
  assign n9375 = ~n4684 & ~n9271 ;
  assign n9376 = n4684 & n9271 ;
  assign n9377 = ~n9375 & ~n9376 ;
  assign n9378 = ~n4231 & ~n9377 ;
  assign n9379 = n4231 & ~n4763 ;
  assign n9380 = ~n9378 & ~n9379 ;
  assign n9381 = n7453 & n9380 ;
  assign n9382 = ~n4697 & ~n7453 ;
  assign n9383 = n5383 & ~n9382 ;
  assign n9384 = ~n9381 & n9383 ;
  assign n9399 = n4694 & ~n7504 ;
  assign n9400 = ~n7453 & ~n8884 ;
  assign n9401 = n7484 & ~n9400 ;
  assign n9402 = n4697 & ~n9401 ;
  assign n9403 = ~n9399 & ~n9402 ;
  assign n9404 = ~n9384 & n9403 ;
  assign n9405 = ~n9398 & n9404 ;
  assign n9406 = n5583 & ~n9405 ;
  assign n9407 = ~n9374 & ~n9406 ;
  assign n9408 = \P1_state_reg[0]/NET0131  & ~n9407 ;
  assign n9373 = n4697 & n5786 ;
  assign n9409 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[21]/NET0131  ;
  assign n9410 = ~n9373 & ~n9409 ;
  assign n9411 = ~n9408 & n9410 ;
  assign n9412 = \P1_reg2_reg[17]/NET0131  & ~n6078 ;
  assign n9413 = \P1_reg2_reg[17]/NET0131  & n6095 ;
  assign n9415 = \P1_reg2_reg[17]/NET0131  & ~n6113 ;
  assign n9416 = n6120 & ~n6161 ;
  assign n9417 = n6168 & ~n9416 ;
  assign n9418 = n3084 & n9417 ;
  assign n9419 = ~n3084 & ~n9417 ;
  assign n9420 = ~n9418 & ~n9419 ;
  assign n9421 = n6113 & ~n9420 ;
  assign n9422 = ~n9415 & ~n9421 ;
  assign n9423 = n6207 & ~n9422 ;
  assign n9429 = n6241 & n7068 ;
  assign n9430 = n7071 & ~n9429 ;
  assign n9431 = n3084 & n9430 ;
  assign n9432 = ~n3084 & ~n9430 ;
  assign n9433 = ~n9431 & ~n9432 ;
  assign n9434 = n6113 & n9433 ;
  assign n9435 = ~n9415 & ~n9434 ;
  assign n9436 = n6282 & ~n9435 ;
  assign n9437 = n3109 & ~n9122 ;
  assign n9438 = ~n6303 & ~n9437 ;
  assign n9439 = ~n2713 & ~n9438 ;
  assign n9440 = n2713 & n3203 ;
  assign n9441 = ~n9439 & ~n9440 ;
  assign n9442 = n6113 & n9441 ;
  assign n9443 = ~n9415 & ~n9442 ;
  assign n9444 = n4011 & ~n9443 ;
  assign n9424 = n3072 & ~n9110 ;
  assign n9425 = ~n9197 & ~n9424 ;
  assign n9426 = n6113 & n9425 ;
  assign n9427 = ~n9415 & ~n9426 ;
  assign n9428 = n6359 & ~n9427 ;
  assign n9446 = n3072 & n6365 ;
  assign n9447 = n6113 & n9446 ;
  assign n9414 = \P1_reg2_reg[17]/NET0131  & ~n8955 ;
  assign n9445 = n3077 & n4112 ;
  assign n9448 = ~n9414 & ~n9445 ;
  assign n9449 = ~n9447 & n9448 ;
  assign n9450 = ~n9428 & n9449 ;
  assign n9451 = ~n9444 & n9450 ;
  assign n9452 = ~n9436 & n9451 ;
  assign n9453 = ~n9423 & n9452 ;
  assign n9454 = n6097 & ~n9453 ;
  assign n9455 = ~n9413 & ~n9454 ;
  assign n9456 = \P1_state_reg[0]/NET0131  & ~n9455 ;
  assign n9457 = ~n9412 & ~n9456 ;
  assign n9458 = \P2_reg0_reg[17]/NET0131  & ~n5589 ;
  assign n9459 = \P2_reg0_reg[17]/NET0131  & n5585 ;
  assign n9467 = \P2_reg0_reg[17]/NET0131  & ~n6706 ;
  assign n9468 = n6706 & ~n8474 ;
  assign n9469 = ~n9467 & ~n9468 ;
  assign n9470 = n5329 & ~n9469 ;
  assign n9471 = n6706 & n8483 ;
  assign n9472 = ~n9467 & ~n9471 ;
  assign n9473 = n5383 & ~n9472 ;
  assign n9460 = n4789 & n5565 ;
  assign n9461 = n5563 & n8496 ;
  assign n9462 = ~n9460 & ~n9461 ;
  assign n9463 = n5526 & n8491 ;
  assign n9464 = n9462 & ~n9463 ;
  assign n9465 = n6706 & ~n9464 ;
  assign n9466 = \P2_reg0_reg[17]/NET0131  & ~n6718 ;
  assign n9474 = ~n9465 & ~n9466 ;
  assign n9475 = ~n9473 & n9474 ;
  assign n9476 = ~n9470 & n9475 ;
  assign n9477 = n5583 & ~n9476 ;
  assign n9478 = ~n9459 & ~n9477 ;
  assign n9479 = \P1_state_reg[0]/NET0131  & ~n9478 ;
  assign n9480 = ~n9458 & ~n9479 ;
  assign n9481 = \P2_reg0_reg[18]/NET0131  & ~n5589 ;
  assign n9482 = \P2_reg0_reg[18]/NET0131  & n5585 ;
  assign n9484 = \P2_reg0_reg[18]/NET0131  & ~n6706 ;
  assign n9485 = n6706 & n8431 ;
  assign n9486 = ~n9484 & ~n9485 ;
  assign n9487 = n5383 & ~n9486 ;
  assign n9483 = \P2_reg0_reg[18]/NET0131  & ~n6717 ;
  assign n9494 = n4814 & n5565 ;
  assign n9495 = n5563 & n8450 ;
  assign n9496 = ~n9494 & ~n9495 ;
  assign n9497 = n6706 & ~n9496 ;
  assign n9498 = ~n9483 & ~n9497 ;
  assign n9499 = ~n9487 & n9498 ;
  assign n9488 = n6706 & n8443 ;
  assign n9489 = ~n9484 & ~n9488 ;
  assign n9490 = n5329 & ~n9489 ;
  assign n9491 = n6706 & ~n8437 ;
  assign n9492 = ~n9484 & ~n9491 ;
  assign n9493 = n5526 & ~n9492 ;
  assign n9500 = ~n9490 & ~n9493 ;
  assign n9501 = n9499 & n9500 ;
  assign n9502 = n5583 & ~n9501 ;
  assign n9503 = ~n9482 & ~n9502 ;
  assign n9504 = \P1_state_reg[0]/NET0131  & ~n9503 ;
  assign n9505 = ~n9481 & ~n9504 ;
  assign n9506 = \P2_reg0_reg[19]/NET0131  & ~n5589 ;
  assign n9507 = \P2_reg0_reg[19]/NET0131  & n5585 ;
  assign n9513 = \P2_reg0_reg[19]/NET0131  & ~n6706 ;
  assign n9514 = n6706 & ~n8517 ;
  assign n9515 = ~n9513 & ~n9514 ;
  assign n9516 = n5526 & ~n9515 ;
  assign n9517 = n6706 & n8523 ;
  assign n9518 = ~n9513 & ~n9517 ;
  assign n9519 = n5329 & ~n9518 ;
  assign n9509 = n5383 & n8532 ;
  assign n9508 = n4745 & n5565 ;
  assign n9510 = ~n8539 & ~n9508 ;
  assign n9511 = ~n9509 & n9510 ;
  assign n9512 = n6706 & ~n9511 ;
  assign n9520 = \P2_reg0_reg[19]/NET0131  & ~n7985 ;
  assign n9521 = ~n9512 & ~n9520 ;
  assign n9522 = ~n9519 & n9521 ;
  assign n9523 = ~n9516 & n9522 ;
  assign n9524 = n5583 & ~n9523 ;
  assign n9525 = ~n9507 & ~n9524 ;
  assign n9526 = \P1_state_reg[0]/NET0131  & ~n9525 ;
  assign n9527 = ~n9506 & ~n9526 ;
  assign n9528 = ~n5562 & ~n6706 ;
  assign n9529 = n5525 & n9528 ;
  assign n9530 = n6718 & n8899 ;
  assign n9531 = ~n9529 & n9530 ;
  assign n9532 = \P2_reg0_reg[22]/NET0131  & ~n9531 ;
  assign n9533 = n6706 & n8899 ;
  assign n9534 = ~n8912 & n9533 ;
  assign n9535 = ~n9532 & ~n9534 ;
  assign n9536 = \P1_reg1_reg[31]/NET0131  & ~n6078 ;
  assign n9537 = \P1_reg1_reg[31]/NET0131  & n6095 ;
  assign n9538 = \P1_reg1_reg[31]/NET0131  & ~n6683 ;
  assign n9539 = n6683 & n8719 ;
  assign n9540 = ~n9538 & ~n9539 ;
  assign n9541 = n6359 & ~n9540 ;
  assign n9549 = n4011 & n6683 ;
  assign n9550 = n8712 & n9549 ;
  assign n9542 = n3467 & n6683 ;
  assign n9543 = ~n9538 & ~n9542 ;
  assign n9544 = n6365 & ~n9543 ;
  assign n9545 = ~n4010 & ~n6426 ;
  assign n9546 = ~n6683 & ~n9545 ;
  assign n9547 = n6424 & ~n9546 ;
  assign n9548 = \P1_reg1_reg[31]/NET0131  & ~n9547 ;
  assign n9551 = ~n9544 & ~n9548 ;
  assign n9552 = ~n9550 & n9551 ;
  assign n9553 = ~n9541 & n9552 ;
  assign n9554 = n6097 & ~n9553 ;
  assign n9555 = ~n9537 & ~n9554 ;
  assign n9556 = \P1_state_reg[0]/NET0131  & ~n9555 ;
  assign n9557 = ~n9536 & ~n9556 ;
  assign n9558 = \P2_reg0_reg[31]/NET0131  & ~n5589 ;
  assign n9559 = \P2_reg0_reg[31]/NET0131  & n5585 ;
  assign n9560 = \P2_reg0_reg[31]/NET0131  & ~n6706 ;
  assign n9561 = n6706 & n8817 ;
  assign n9562 = ~n9560 & ~n9561 ;
  assign n9563 = n5563 & ~n9562 ;
  assign n9569 = n5383 & n6706 ;
  assign n9570 = n8824 & n9569 ;
  assign n9564 = n5879 & n6706 ;
  assign n9565 = ~n9560 & ~n9564 ;
  assign n9566 = n5565 & ~n9565 ;
  assign n9567 = n6394 & ~n9528 ;
  assign n9568 = \P2_reg0_reg[31]/NET0131  & ~n9567 ;
  assign n9571 = ~n9566 & ~n9568 ;
  assign n9572 = ~n9570 & n9571 ;
  assign n9573 = ~n9563 & n9572 ;
  assign n9574 = n5583 & ~n9573 ;
  assign n9575 = ~n9559 & ~n9574 ;
  assign n9576 = \P1_state_reg[0]/NET0131  & ~n9575 ;
  assign n9577 = ~n9558 & ~n9576 ;
  assign n9578 = \P2_reg1_reg[17]/NET0131  & ~n5589 ;
  assign n9579 = \P2_reg1_reg[17]/NET0131  & n5585 ;
  assign n9582 = \P2_reg1_reg[17]/NET0131  & ~n6380 ;
  assign n9583 = n6380 & ~n8474 ;
  assign n9584 = ~n9582 & ~n9583 ;
  assign n9585 = n5329 & ~n9584 ;
  assign n9586 = n6380 & n8483 ;
  assign n9587 = ~n9582 & ~n9586 ;
  assign n9588 = n5383 & ~n9587 ;
  assign n9580 = \P2_reg1_reg[17]/NET0131  & ~n6398 ;
  assign n9581 = n6380 & ~n9464 ;
  assign n9589 = ~n9580 & ~n9581 ;
  assign n9590 = ~n9588 & n9589 ;
  assign n9591 = ~n9585 & n9590 ;
  assign n9592 = n5583 & ~n9591 ;
  assign n9593 = ~n9579 & ~n9592 ;
  assign n9594 = \P1_state_reg[0]/NET0131  & ~n9593 ;
  assign n9595 = ~n9578 & ~n9594 ;
  assign n9596 = \P2_reg1_reg[18]/NET0131  & ~n5589 ;
  assign n9597 = \P2_reg1_reg[18]/NET0131  & n5585 ;
  assign n9599 = \P2_reg1_reg[18]/NET0131  & ~n6380 ;
  assign n9600 = n6380 & n8443 ;
  assign n9601 = ~n9599 & ~n9600 ;
  assign n9602 = n5329 & ~n9601 ;
  assign n9598 = \P2_reg1_reg[18]/NET0131  & ~n6397 ;
  assign n9609 = n6380 & ~n9496 ;
  assign n9610 = ~n9598 & ~n9609 ;
  assign n9611 = ~n9602 & n9610 ;
  assign n9603 = n6380 & ~n8437 ;
  assign n9604 = ~n9599 & ~n9603 ;
  assign n9605 = n5526 & ~n9604 ;
  assign n9606 = n6380 & n8431 ;
  assign n9607 = ~n9599 & ~n9606 ;
  assign n9608 = n5383 & ~n9607 ;
  assign n9612 = ~n9605 & ~n9608 ;
  assign n9613 = n9611 & n9612 ;
  assign n9614 = n5583 & ~n9613 ;
  assign n9615 = ~n9597 & ~n9614 ;
  assign n9616 = \P1_state_reg[0]/NET0131  & ~n9615 ;
  assign n9617 = ~n9596 & ~n9616 ;
  assign n9618 = \P2_reg1_reg[19]/NET0131  & ~n5589 ;
  assign n9619 = \P2_reg1_reg[19]/NET0131  & n5585 ;
  assign n9621 = \P2_reg1_reg[19]/NET0131  & ~n6380 ;
  assign n9622 = n6380 & ~n8517 ;
  assign n9623 = ~n9621 & ~n9622 ;
  assign n9624 = n5526 & ~n9623 ;
  assign n9625 = n6380 & n8523 ;
  assign n9626 = ~n9621 & ~n9625 ;
  assign n9627 = n5329 & ~n9626 ;
  assign n9620 = n6380 & ~n9511 ;
  assign n9628 = \P2_reg1_reg[19]/NET0131  & ~n8026 ;
  assign n9629 = ~n9620 & ~n9628 ;
  assign n9630 = ~n9627 & n9629 ;
  assign n9631 = ~n9624 & n9630 ;
  assign n9632 = n5583 & ~n9631 ;
  assign n9633 = ~n9619 & ~n9632 ;
  assign n9634 = \P1_state_reg[0]/NET0131  & ~n9633 ;
  assign n9635 = ~n9618 & ~n9634 ;
  assign n9636 = \P2_reg1_reg[21]/NET0131  & ~n8902 ;
  assign n9638 = n5383 & ~n9380 ;
  assign n9637 = n4694 & n5565 ;
  assign n9639 = n9397 & ~n9637 ;
  assign n9640 = ~n9638 & n9639 ;
  assign n9641 = n8913 & ~n9640 ;
  assign n9642 = ~n9636 & ~n9641 ;
  assign n9643 = n2883 & n4112 ;
  assign n9644 = n6113 & ~n9049 ;
  assign n9645 = ~n9643 & ~n9644 ;
  assign n9646 = n9044 & ~n9645 ;
  assign n9647 = n8062 & n9044 ;
  assign n9648 = \P1_reg2_reg[22]/NET0131  & ~n9647 ;
  assign n9649 = ~n9646 & ~n9648 ;
  assign n9654 = \P2_reg1_reg[31]/NET0131  & ~n6380 ;
  assign n9655 = n8817 & n8913 ;
  assign n9656 = ~n9654 & ~n9655 ;
  assign n9657 = n5563 & ~n9656 ;
  assign n9650 = ~n5562 & ~n6380 ;
  assign n9651 = n6394 & n8899 ;
  assign n9652 = ~n9650 & n9651 ;
  assign n9653 = \P2_reg1_reg[31]/NET0131  & ~n9652 ;
  assign n9658 = n5879 & n6380 ;
  assign n9659 = ~n9654 & ~n9658 ;
  assign n9660 = n5565 & ~n9659 ;
  assign n9661 = n5383 & n6380 ;
  assign n9662 = n8824 & n9661 ;
  assign n9663 = ~n9660 & ~n9662 ;
  assign n9664 = n8899 & ~n9663 ;
  assign n9665 = ~n9653 & ~n9664 ;
  assign n9666 = ~n9657 & n9665 ;
  assign n9667 = \P2_reg2_reg[18]/NET0131  & ~n5589 ;
  assign n9668 = \P2_reg2_reg[18]/NET0131  & n5585 ;
  assign n9670 = \P2_reg2_reg[18]/NET0131  & ~n4219 ;
  assign n9671 = n4219 & ~n8437 ;
  assign n9672 = ~n9670 & ~n9671 ;
  assign n9673 = n5526 & ~n9672 ;
  assign n9681 = n4219 & ~n9496 ;
  assign n9669 = \P2_reg2_reg[18]/NET0131  & ~n6839 ;
  assign n9680 = n4793 & n5574 ;
  assign n9682 = ~n9669 & ~n9680 ;
  assign n9683 = ~n9681 & n9682 ;
  assign n9684 = ~n9673 & n9683 ;
  assign n9674 = n4219 & n8443 ;
  assign n9675 = ~n9670 & ~n9674 ;
  assign n9676 = n5329 & ~n9675 ;
  assign n9677 = n4219 & n8431 ;
  assign n9678 = ~n9670 & ~n9677 ;
  assign n9679 = n5383 & ~n9678 ;
  assign n9685 = ~n9676 & ~n9679 ;
  assign n9686 = n9684 & n9685 ;
  assign n9687 = n5583 & ~n9686 ;
  assign n9688 = ~n9668 & ~n9687 ;
  assign n9689 = \P1_state_reg[0]/NET0131  & ~n9688 ;
  assign n9690 = ~n9667 & ~n9689 ;
  assign n9691 = \P2_reg2_reg[17]/NET0131  & ~n5589 ;
  assign n9692 = \P2_reg2_reg[17]/NET0131  & n5585 ;
  assign n9694 = \P2_reg2_reg[17]/NET0131  & ~n4219 ;
  assign n9695 = n4219 & ~n8474 ;
  assign n9696 = ~n9694 & ~n9695 ;
  assign n9697 = n5329 & ~n9696 ;
  assign n9698 = n4219 & n8483 ;
  assign n9699 = ~n9694 & ~n9698 ;
  assign n9700 = n5383 & ~n9699 ;
  assign n9701 = n4219 & n8491 ;
  assign n9702 = ~n9694 & ~n9701 ;
  assign n9703 = n5526 & ~n9702 ;
  assign n9704 = n4219 & ~n9462 ;
  assign n9693 = \P2_reg2_reg[17]/NET0131  & ~n6839 ;
  assign n9705 = n4770 & n5574 ;
  assign n9706 = ~n9693 & ~n9705 ;
  assign n9707 = ~n9704 & n9706 ;
  assign n9708 = ~n9703 & n9707 ;
  assign n9709 = ~n9700 & n9708 ;
  assign n9710 = ~n9697 & n9709 ;
  assign n9711 = n5583 & ~n9710 ;
  assign n9712 = ~n9692 & ~n9711 ;
  assign n9713 = \P1_state_reg[0]/NET0131  & ~n9712 ;
  assign n9714 = ~n9691 & ~n9713 ;
  assign n9715 = \P2_reg2_reg[19]/NET0131  & ~n5589 ;
  assign n9716 = \P2_reg2_reg[19]/NET0131  & n5585 ;
  assign n9718 = \P2_reg2_reg[19]/NET0131  & ~n4219 ;
  assign n9719 = n4219 & ~n8517 ;
  assign n9720 = ~n9718 & ~n9719 ;
  assign n9721 = n5526 & ~n9720 ;
  assign n9722 = n4219 & n8523 ;
  assign n9723 = ~n9718 & ~n9722 ;
  assign n9724 = n5329 & ~n9723 ;
  assign n9725 = n4219 & n8532 ;
  assign n9726 = ~n9718 & ~n9725 ;
  assign n9727 = n5383 & ~n9726 ;
  assign n9728 = n4219 & n8538 ;
  assign n9729 = ~n9718 & ~n9728 ;
  assign n9730 = n5563 & ~n9729 ;
  assign n9732 = \P2_reg2_reg[19]/NET0131  & ~n5570 ;
  assign n9717 = n4219 & n9508 ;
  assign n9731 = n4722 & n5574 ;
  assign n9733 = ~n9717 & ~n9731 ;
  assign n9734 = ~n9732 & n9733 ;
  assign n9735 = ~n9730 & n9734 ;
  assign n9736 = ~n9727 & n9735 ;
  assign n9737 = ~n9724 & n9736 ;
  assign n9738 = ~n9721 & n9737 ;
  assign n9739 = n5583 & ~n9738 ;
  assign n9740 = ~n9716 & ~n9739 ;
  assign n9741 = \P1_state_reg[0]/NET0131  & ~n9740 ;
  assign n9742 = ~n9715 & ~n9741 ;
  assign n9743 = \P2_reg2_reg[20]/NET0131  & ~n5589 ;
  assign n9744 = \P2_reg2_reg[20]/NET0131  & n5585 ;
  assign n9746 = \P2_reg2_reg[20]/NET0131  & ~n4219 ;
  assign n9750 = n4219 & n9276 ;
  assign n9751 = ~n9746 & ~n9750 ;
  assign n9752 = n5383 & ~n9751 ;
  assign n9747 = n4219 & ~n9267 ;
  assign n9748 = ~n9746 & ~n9747 ;
  assign n9749 = n5329 & ~n9748 ;
  assign n9753 = n4219 & ~n9282 ;
  assign n9754 = ~n9746 & ~n9753 ;
  assign n9755 = n5526 & ~n9754 ;
  assign n9757 = n4754 & n5565 ;
  assign n9758 = n5563 & n9287 ;
  assign n9759 = ~n9757 & ~n9758 ;
  assign n9760 = n4219 & ~n9759 ;
  assign n9745 = \P2_reg2_reg[20]/NET0131  & ~n6839 ;
  assign n9756 = n4757 & n5574 ;
  assign n9761 = ~n9745 & ~n9756 ;
  assign n9762 = ~n9760 & n9761 ;
  assign n9763 = ~n9755 & n9762 ;
  assign n9764 = ~n9749 & n9763 ;
  assign n9765 = ~n9752 & n9764 ;
  assign n9766 = n5583 & ~n9765 ;
  assign n9767 = ~n9744 & ~n9766 ;
  assign n9768 = \P1_state_reg[0]/NET0131  & ~n9767 ;
  assign n9769 = ~n9743 & ~n9768 ;
  assign n9770 = ~n4219 & ~n8884 ;
  assign n9771 = n6839 & ~n9770 ;
  assign n9772 = ~n6840 & n9771 ;
  assign n9773 = n8899 & n9772 ;
  assign n9774 = \P2_reg2_reg[21]/NET0131  & ~n9773 ;
  assign n9775 = n4219 & ~n9640 ;
  assign n9776 = n4697 & n5574 ;
  assign n9777 = ~n9775 & ~n9776 ;
  assign n9778 = n8899 & ~n9777 ;
  assign n9779 = ~n9774 & ~n9778 ;
  assign n9780 = \P2_reg2_reg[22]/NET0131  & ~n5589 ;
  assign n9781 = \P2_reg2_reg[22]/NET0131  & n5585 ;
  assign n9788 = n4219 & n8740 ;
  assign n9787 = ~\P2_reg2_reg[22]/NET0131  & ~n4219 ;
  assign n9789 = n5329 & ~n9787 ;
  assign n9790 = ~n9788 & n9789 ;
  assign n9782 = n4219 & ~n8911 ;
  assign n9783 = n4680 & n5574 ;
  assign n9784 = ~n4219 & n5526 ;
  assign n9785 = n6841 & ~n9784 ;
  assign n9786 = \P2_reg2_reg[22]/NET0131  & ~n9785 ;
  assign n9791 = ~n9783 & ~n9786 ;
  assign n9792 = ~n9782 & n9791 ;
  assign n9793 = ~n9790 & n9792 ;
  assign n9794 = n5583 & ~n9793 ;
  assign n9795 = ~n9781 & ~n9794 ;
  assign n9796 = \P1_state_reg[0]/NET0131  & ~n9795 ;
  assign n9797 = ~n9780 & ~n9796 ;
  assign n9798 = \P1_reg0_reg[17]/NET0131  & ~n6078 ;
  assign n9799 = \P1_reg0_reg[17]/NET0131  & n6095 ;
  assign n9801 = \P1_reg0_reg[17]/NET0131  & ~n6409 ;
  assign n9802 = n6409 & ~n9420 ;
  assign n9803 = ~n9801 & ~n9802 ;
  assign n9804 = n6207 & ~n9803 ;
  assign n9808 = n6409 & n9433 ;
  assign n9809 = ~n9801 & ~n9808 ;
  assign n9810 = n6282 & ~n9809 ;
  assign n9811 = n6409 & n9441 ;
  assign n9812 = ~n9801 & ~n9811 ;
  assign n9813 = n4011 & ~n9812 ;
  assign n9805 = n6409 & n9425 ;
  assign n9806 = ~n9801 & ~n9805 ;
  assign n9807 = n6359 & ~n9806 ;
  assign n9800 = n6409 & n9446 ;
  assign n9814 = \P1_reg0_reg[17]/NET0131  & ~n6425 ;
  assign n9815 = ~n9800 & ~n9814 ;
  assign n9816 = ~n9807 & n9815 ;
  assign n9817 = ~n9813 & n9816 ;
  assign n9818 = ~n9810 & n9817 ;
  assign n9819 = ~n9804 & n9818 ;
  assign n9820 = n6097 & ~n9819 ;
  assign n9821 = ~n9799 & ~n9820 ;
  assign n9822 = \P1_state_reg[0]/NET0131  & ~n9821 ;
  assign n9823 = ~n9798 & ~n9822 ;
  assign n9824 = ~n6409 & ~n8060 ;
  assign n9825 = n6424 & ~n9824 ;
  assign n9826 = n9044 & n9825 ;
  assign n9827 = ~n8684 & n9826 ;
  assign n9828 = \P1_reg0_reg[22]/NET0131  & ~n9827 ;
  assign n9829 = n6409 & n9044 ;
  assign n9830 = ~n9049 & n9829 ;
  assign n9831 = ~n9828 & ~n9830 ;
  assign n9832 = \P3_reg0_reg[17]/NET0131  & ~n2143 ;
  assign n9833 = \P3_reg0_reg[17]/NET0131  & n2145 ;
  assign n9836 = \P3_reg0_reg[17]/NET0131  & ~n2236 ;
  assign n9837 = ~n8602 & ~n9836 ;
  assign n9838 = n2393 & ~n9837 ;
  assign n9834 = \P3_reg0_reg[17]/NET0131  & ~n2287 ;
  assign n9835 = ~n1166 & n2289 ;
  assign n9848 = ~n9834 & ~n9835 ;
  assign n9849 = ~n9838 & n9848 ;
  assign n9845 = n2236 & ~n8619 ;
  assign n9846 = ~n9836 & ~n9845 ;
  assign n9847 = n737 & ~n9846 ;
  assign n9839 = \P3_reg0_reg[17]/NET0131  & ~n2163 ;
  assign n9840 = n2163 & n8607 ;
  assign n9841 = ~n9839 & ~n9840 ;
  assign n9842 = n2234 & ~n9841 ;
  assign n9843 = ~n8612 & ~n9839 ;
  assign n9844 = n2391 & ~n9843 ;
  assign n9850 = ~n9842 & ~n9844 ;
  assign n9851 = ~n9847 & n9850 ;
  assign n9852 = n9849 & n9851 ;
  assign n9853 = n2147 & ~n9852 ;
  assign n9854 = ~n9833 & ~n9853 ;
  assign n9855 = \P1_state_reg[0]/NET0131  & ~n9854 ;
  assign n9856 = ~n9832 & ~n9855 ;
  assign n9857 = \P3_reg0_reg[18]/NET0131  & ~n2143 ;
  assign n9858 = \P3_reg0_reg[18]/NET0131  & n2145 ;
  assign n9859 = \P3_reg0_reg[18]/NET0131  & ~n2236 ;
  assign n9866 = n2236 & ~n8574 ;
  assign n9867 = ~n9859 & ~n9866 ;
  assign n9868 = n737 & ~n9867 ;
  assign n9862 = \P3_reg0_reg[18]/NET0131  & ~n2163 ;
  assign n9863 = n2163 & ~n8566 ;
  assign n9864 = ~n9862 & ~n9863 ;
  assign n9865 = n2234 & ~n9864 ;
  assign n9871 = \P3_reg0_reg[18]/NET0131  & ~n2287 ;
  assign n9872 = ~n1137 & n2285 ;
  assign n9873 = n2163 & n9872 ;
  assign n9874 = ~n9871 & ~n9873 ;
  assign n9875 = ~n9865 & n9874 ;
  assign n9876 = ~n9868 & n9875 ;
  assign n9860 = ~n8578 & ~n9859 ;
  assign n9861 = n2393 & ~n9860 ;
  assign n9869 = ~n8560 & ~n9862 ;
  assign n9870 = n2391 & ~n9869 ;
  assign n9877 = ~n9861 & ~n9870 ;
  assign n9878 = n9876 & n9877 ;
  assign n9879 = n2147 & ~n9878 ;
  assign n9880 = ~n9858 & ~n9879 ;
  assign n9881 = \P1_state_reg[0]/NET0131  & ~n9880 ;
  assign n9882 = ~n9857 & ~n9881 ;
  assign n9883 = \P3_reg0_reg[19]/NET0131  & ~n2143 ;
  assign n9884 = \P3_reg0_reg[19]/NET0131  & n2145 ;
  assign n9886 = \P3_reg0_reg[19]/NET0131  & ~n2236 ;
  assign n9887 = ~n6536 & ~n9886 ;
  assign n9888 = n2393 & ~n9887 ;
  assign n9889 = \P3_reg0_reg[19]/NET0131  & ~n2163 ;
  assign n9895 = n2163 & n6552 ;
  assign n9896 = ~n9889 & ~n9895 ;
  assign n9897 = n2234 & ~n9896 ;
  assign n9885 = \P3_reg0_reg[19]/NET0131  & ~n2287 ;
  assign n9898 = ~n1110 & n2289 ;
  assign n9899 = ~n9885 & ~n9898 ;
  assign n9900 = ~n9897 & n9899 ;
  assign n9901 = ~n9888 & n9900 ;
  assign n9890 = ~n6532 & ~n9889 ;
  assign n9891 = n2391 & ~n9890 ;
  assign n9892 = n2236 & ~n6546 ;
  assign n9893 = ~n9886 & ~n9892 ;
  assign n9894 = n737 & ~n9893 ;
  assign n9902 = ~n9891 & ~n9894 ;
  assign n9903 = n9901 & n9902 ;
  assign n9904 = n2147 & ~n9903 ;
  assign n9905 = ~n9884 & ~n9904 ;
  assign n9906 = \P1_state_reg[0]/NET0131  & ~n9905 ;
  assign n9907 = ~n9883 & ~n9906 ;
  assign n9908 = \P3_reg0_reg[20]/NET0131  & ~n2143 ;
  assign n9909 = \P3_reg0_reg[20]/NET0131  & n2145 ;
  assign n9911 = \P3_reg0_reg[20]/NET0131  & ~n2163 ;
  assign n9912 = n2163 & ~n7271 ;
  assign n9913 = ~n9911 & ~n9912 ;
  assign n9914 = n2234 & ~n9913 ;
  assign n9910 = n1063 & n2289 ;
  assign n9923 = \P3_reg0_reg[20]/NET0131  & ~n2287 ;
  assign n9924 = ~n9910 & ~n9923 ;
  assign n9925 = ~n9914 & n9924 ;
  assign n9915 = \P3_reg0_reg[20]/NET0131  & ~n2236 ;
  assign n9921 = ~n7433 & ~n9915 ;
  assign n9922 = n2393 & ~n9921 ;
  assign n9916 = n2236 & ~n7265 ;
  assign n9917 = ~n9915 & ~n9916 ;
  assign n9918 = n737 & ~n9917 ;
  assign n9919 = ~n7436 & ~n9911 ;
  assign n9920 = n2391 & ~n9919 ;
  assign n9926 = ~n9918 & ~n9920 ;
  assign n9927 = ~n9922 & n9926 ;
  assign n9928 = n9925 & n9927 ;
  assign n9929 = n2147 & ~n9928 ;
  assign n9930 = ~n9909 & ~n9929 ;
  assign n9931 = \P1_state_reg[0]/NET0131  & ~n9930 ;
  assign n9932 = ~n9908 & ~n9931 ;
  assign n9933 = \P3_reg0_reg[21]/NET0131  & ~n2143 ;
  assign n9934 = \P3_reg0_reg[21]/NET0131  & n2145 ;
  assign n9936 = \P3_reg0_reg[21]/NET0131  & ~n2236 ;
  assign n9937 = ~n7302 & ~n9936 ;
  assign n9938 = n2393 & ~n9937 ;
  assign n9945 = n2236 & ~n7315 ;
  assign n9946 = ~n9936 & ~n9945 ;
  assign n9947 = n737 & ~n9946 ;
  assign n9935 = \P3_reg0_reg[21]/NET0131  & ~n2287 ;
  assign n9948 = n1029 & n2289 ;
  assign n9949 = ~n9935 & ~n9948 ;
  assign n9950 = ~n9947 & n9949 ;
  assign n9951 = ~n9938 & n9950 ;
  assign n9939 = \P3_reg0_reg[21]/NET0131  & ~n2163 ;
  assign n9940 = ~n7298 & ~n9939 ;
  assign n9941 = n2391 & ~n9940 ;
  assign n9942 = n2163 & ~n7307 ;
  assign n9943 = ~n9939 & ~n9942 ;
  assign n9944 = n2234 & ~n9943 ;
  assign n9952 = ~n9941 & ~n9944 ;
  assign n9953 = n9951 & n9952 ;
  assign n9954 = n2147 & ~n9953 ;
  assign n9955 = ~n9934 & ~n9954 ;
  assign n9956 = \P1_state_reg[0]/NET0131  & ~n9955 ;
  assign n9957 = ~n9933 & ~n9956 ;
  assign n9958 = \P3_reg0_reg[22]/NET0131  & ~n2143 ;
  assign n9959 = \P3_reg0_reg[22]/NET0131  & n2145 ;
  assign n9960 = \P3_reg0_reg[22]/NET0131  & ~n2163 ;
  assign n9961 = ~n7348 & ~n9960 ;
  assign n9962 = n2391 & ~n9961 ;
  assign n9963 = \P3_reg0_reg[22]/NET0131  & ~n2236 ;
  assign n9970 = n2236 & ~n7363 ;
  assign n9971 = ~n9963 & ~n9970 ;
  assign n9972 = n737 & ~n9971 ;
  assign n9966 = n991 & n2289 ;
  assign n9973 = \P3_reg0_reg[22]/NET0131  & ~n2287 ;
  assign n9974 = ~n9966 & ~n9973 ;
  assign n9975 = ~n9972 & n9974 ;
  assign n9976 = ~n9962 & n9975 ;
  assign n9964 = ~n7344 & ~n9963 ;
  assign n9965 = n2393 & ~n9964 ;
  assign n9967 = n2163 & ~n7355 ;
  assign n9968 = ~n9960 & ~n9967 ;
  assign n9969 = n2234 & ~n9968 ;
  assign n9977 = ~n9965 & ~n9969 ;
  assign n9978 = n9976 & n9977 ;
  assign n9979 = n2147 & ~n9978 ;
  assign n9980 = ~n9959 & ~n9979 ;
  assign n9981 = \P1_state_reg[0]/NET0131  & ~n9980 ;
  assign n9982 = ~n9958 & ~n9981 ;
  assign n9983 = \P3_reg0_reg[23]/NET0131  & ~n2143 ;
  assign n9984 = \P3_reg0_reg[23]/NET0131  & n2145 ;
  assign n9985 = \P3_reg0_reg[23]/NET0131  & ~n2163 ;
  assign n9994 = n2163 & ~n7405 ;
  assign n9995 = ~n9985 & ~n9994 ;
  assign n9996 = n2234 & ~n9995 ;
  assign n9988 = \P3_reg0_reg[23]/NET0131  & ~n2236 ;
  assign n9991 = n2236 & ~n7398 ;
  assign n9992 = ~n9988 & ~n9991 ;
  assign n9993 = n737 & ~n9992 ;
  assign n9997 = \P3_reg0_reg[23]/NET0131  & ~n2287 ;
  assign n9998 = n886 & n2289 ;
  assign n9999 = ~n9997 & ~n9998 ;
  assign n10000 = ~n9993 & n9999 ;
  assign n10001 = ~n9996 & n10000 ;
  assign n9986 = ~n7391 & ~n9985 ;
  assign n9987 = n2391 & ~n9986 ;
  assign n9989 = ~n7387 & ~n9988 ;
  assign n9990 = n2393 & ~n9989 ;
  assign n10002 = ~n9987 & ~n9990 ;
  assign n10003 = n10001 & n10002 ;
  assign n10004 = n2147 & ~n10003 ;
  assign n10005 = ~n9984 & ~n10004 ;
  assign n10006 = \P1_state_reg[0]/NET0131  & ~n10005 ;
  assign n10007 = ~n9983 & ~n10006 ;
  assign n10012 = \P1_reg0_reg[31]/NET0131  & ~n6409 ;
  assign n10013 = n8719 & n9829 ;
  assign n10014 = ~n10012 & ~n10013 ;
  assign n10015 = n6359 & ~n10014 ;
  assign n10008 = ~n6409 & ~n9545 ;
  assign n10009 = n6424 & ~n10008 ;
  assign n10010 = n9044 & n10009 ;
  assign n10011 = \P1_reg0_reg[31]/NET0131  & ~n10010 ;
  assign n10016 = n4011 & n6409 ;
  assign n10017 = n8712 & n10016 ;
  assign n10018 = n3467 & n6409 ;
  assign n10019 = ~n10012 & ~n10018 ;
  assign n10020 = n6365 & ~n10019 ;
  assign n10021 = ~n10017 & ~n10020 ;
  assign n10022 = n9044 & ~n10021 ;
  assign n10023 = ~n10011 & ~n10022 ;
  assign n10024 = ~n10015 & n10023 ;
  assign n10025 = \P3_reg1_reg[18]/NET0131  & ~n2143 ;
  assign n10026 = \P3_reg1_reg[18]/NET0131  & n2145 ;
  assign n10034 = \P3_reg1_reg[18]/NET0131  & ~n2408 ;
  assign n10038 = n2408 & n8559 ;
  assign n10039 = ~n10034 & ~n10038 ;
  assign n10040 = n714 & ~n10039 ;
  assign n10027 = \P3_reg1_reg[18]/NET0131  & ~n2427 ;
  assign n10028 = n2427 & ~n8566 ;
  assign n10029 = ~n10027 & ~n10028 ;
  assign n10030 = n2425 & ~n10029 ;
  assign n10041 = \P3_reg1_reg[18]/NET0131  & ~n6449 ;
  assign n10042 = n2408 & n9872 ;
  assign n10043 = ~n10041 & ~n10042 ;
  assign n10044 = ~n10030 & n10043 ;
  assign n10031 = n2427 & ~n8574 ;
  assign n10032 = ~n10027 & ~n10031 ;
  assign n10033 = n737 & ~n10032 ;
  assign n10035 = n2408 & ~n8566 ;
  assign n10036 = ~n10034 & ~n10035 ;
  assign n10037 = ~n2518 & ~n10036 ;
  assign n10045 = ~n10033 & ~n10037 ;
  assign n10046 = n10044 & n10045 ;
  assign n10047 = ~n10040 & n10046 ;
  assign n10048 = n2147 & ~n10047 ;
  assign n10049 = ~n10026 & ~n10048 ;
  assign n10050 = \P1_state_reg[0]/NET0131  & ~n10049 ;
  assign n10051 = ~n10025 & ~n10050 ;
  assign n10052 = \P3_reg1_reg[19]/NET0131  & ~n2143 ;
  assign n10053 = \P3_reg1_reg[19]/NET0131  & n2145 ;
  assign n10054 = \P3_reg1_reg[19]/NET0131  & ~n2427 ;
  assign n10061 = ~n7230 & ~n10054 ;
  assign n10062 = n2425 & ~n10061 ;
  assign n10058 = \P3_reg1_reg[19]/NET0131  & ~n2408 ;
  assign n10059 = ~n7226 & ~n10058 ;
  assign n10060 = ~n2518 & ~n10059 ;
  assign n10066 = ~n1110 & n6451 ;
  assign n10067 = \P3_reg1_reg[19]/NET0131  & ~n6449 ;
  assign n10068 = ~n10066 & ~n10067 ;
  assign n10069 = ~n10060 & n10068 ;
  assign n10070 = ~n10062 & n10069 ;
  assign n10055 = n2427 & ~n6546 ;
  assign n10056 = ~n10054 & ~n10055 ;
  assign n10057 = n737 & ~n10056 ;
  assign n10063 = n2408 & ~n6531 ;
  assign n10064 = ~n10058 & ~n10063 ;
  assign n10065 = n714 & ~n10064 ;
  assign n10071 = ~n10057 & ~n10065 ;
  assign n10072 = n10070 & n10071 ;
  assign n10073 = n2147 & ~n10072 ;
  assign n10074 = ~n10053 & ~n10073 ;
  assign n10075 = \P1_state_reg[0]/NET0131  & ~n10074 ;
  assign n10076 = ~n10052 & ~n10075 ;
  assign n10077 = \P3_reg1_reg[17]/NET0131  & ~n2143 ;
  assign n10078 = \P3_reg1_reg[17]/NET0131  & n2145 ;
  assign n10081 = \P3_reg1_reg[17]/NET0131  & ~n2408 ;
  assign n10082 = n2408 & ~n8601 ;
  assign n10083 = ~n10081 & ~n10082 ;
  assign n10084 = n714 & ~n10083 ;
  assign n10079 = \P3_reg1_reg[17]/NET0131  & ~n6449 ;
  assign n10080 = ~n1166 & n6451 ;
  assign n10095 = ~n10079 & ~n10080 ;
  assign n10096 = ~n10084 & n10095 ;
  assign n10092 = n2408 & n8607 ;
  assign n10093 = ~n10081 & ~n10092 ;
  assign n10094 = ~n2518 & ~n10093 ;
  assign n10085 = \P3_reg1_reg[17]/NET0131  & ~n2427 ;
  assign n10086 = n2427 & n8607 ;
  assign n10087 = ~n10085 & ~n10086 ;
  assign n10088 = n2425 & ~n10087 ;
  assign n10089 = n2427 & ~n8619 ;
  assign n10090 = ~n10085 & ~n10089 ;
  assign n10091 = n737 & ~n10090 ;
  assign n10097 = ~n10088 & ~n10091 ;
  assign n10098 = ~n10094 & n10097 ;
  assign n10099 = n10096 & n10098 ;
  assign n10100 = n2147 & ~n10099 ;
  assign n10101 = ~n10078 & ~n10100 ;
  assign n10102 = \P1_state_reg[0]/NET0131  & ~n10101 ;
  assign n10103 = ~n10077 & ~n10102 ;
  assign n10104 = \P3_reg1_reg[21]/NET0131  & ~n2143 ;
  assign n10105 = \P3_reg1_reg[21]/NET0131  & n2145 ;
  assign n10107 = \P3_reg1_reg[21]/NET0131  & ~n2427 ;
  assign n10108 = ~n8377 & ~n10107 ;
  assign n10109 = n2425 & ~n10108 ;
  assign n10116 = n2427 & ~n7315 ;
  assign n10117 = ~n10107 & ~n10116 ;
  assign n10118 = n737 & ~n10117 ;
  assign n10106 = \P3_reg1_reg[21]/NET0131  & ~n6449 ;
  assign n10119 = n1029 & n6451 ;
  assign n10120 = ~n10106 & ~n10119 ;
  assign n10121 = ~n10118 & n10120 ;
  assign n10122 = ~n10109 & n10121 ;
  assign n10110 = \P3_reg1_reg[21]/NET0131  & ~n2408 ;
  assign n10111 = n2408 & ~n7297 ;
  assign n10112 = ~n10110 & ~n10111 ;
  assign n10113 = n714 & ~n10112 ;
  assign n10114 = ~n8374 & ~n10110 ;
  assign n10115 = ~n2518 & ~n10114 ;
  assign n10123 = ~n10113 & ~n10115 ;
  assign n10124 = n10122 & n10123 ;
  assign n10125 = n2147 & ~n10124 ;
  assign n10126 = ~n10105 & ~n10125 ;
  assign n10127 = \P1_state_reg[0]/NET0131  & ~n10126 ;
  assign n10128 = ~n10104 & ~n10127 ;
  assign n10129 = \P3_reg1_reg[20]/NET0131  & ~n2143 ;
  assign n10130 = \P3_reg1_reg[20]/NET0131  & n2145 ;
  assign n10132 = \P3_reg1_reg[20]/NET0131  & ~n2408 ;
  assign n10133 = n2408 & ~n7256 ;
  assign n10134 = ~n10132 & ~n10133 ;
  assign n10135 = n714 & ~n10134 ;
  assign n10131 = n2408 & n7251 ;
  assign n10144 = \P3_reg1_reg[20]/NET0131  & ~n6449 ;
  assign n10145 = ~n10131 & ~n10144 ;
  assign n10146 = ~n10135 & n10145 ;
  assign n10142 = ~n7272 & ~n10132 ;
  assign n10143 = ~n2518 & ~n10142 ;
  assign n10136 = \P3_reg1_reg[20]/NET0131  & ~n2427 ;
  assign n10137 = n2427 & ~n7265 ;
  assign n10138 = ~n10136 & ~n10137 ;
  assign n10139 = n737 & ~n10138 ;
  assign n10140 = ~n7275 & ~n10136 ;
  assign n10141 = n2425 & ~n10140 ;
  assign n10147 = ~n10139 & ~n10141 ;
  assign n10148 = ~n10143 & n10147 ;
  assign n10149 = n10146 & n10148 ;
  assign n10150 = n2147 & ~n10149 ;
  assign n10151 = ~n10130 & ~n10150 ;
  assign n10152 = \P1_state_reg[0]/NET0131  & ~n10151 ;
  assign n10153 = ~n10129 & ~n10152 ;
  assign n10154 = \P3_reg1_reg[22]/NET0131  & ~n2143 ;
  assign n10155 = \P3_reg1_reg[22]/NET0131  & n2145 ;
  assign n10156 = \P3_reg1_reg[22]/NET0131  & ~n2408 ;
  assign n10157 = n2408 & ~n7343 ;
  assign n10158 = ~n10156 & ~n10157 ;
  assign n10159 = n714 & ~n10158 ;
  assign n10160 = \P3_reg1_reg[22]/NET0131  & ~n2427 ;
  assign n10166 = n2427 & ~n7363 ;
  assign n10167 = ~n10160 & ~n10166 ;
  assign n10168 = n737 & ~n10167 ;
  assign n10163 = \P3_reg1_reg[22]/NET0131  & ~n6449 ;
  assign n10169 = n991 & n6451 ;
  assign n10170 = ~n10163 & ~n10169 ;
  assign n10171 = ~n10168 & n10170 ;
  assign n10172 = ~n10159 & n10171 ;
  assign n10161 = ~n8346 & ~n10160 ;
  assign n10162 = n2425 & ~n10161 ;
  assign n10164 = ~n8342 & ~n10156 ;
  assign n10165 = ~n2518 & ~n10164 ;
  assign n10173 = ~n10162 & ~n10165 ;
  assign n10174 = n10172 & n10173 ;
  assign n10175 = n2147 & ~n10174 ;
  assign n10176 = ~n10155 & ~n10175 ;
  assign n10177 = \P1_state_reg[0]/NET0131  & ~n10176 ;
  assign n10178 = ~n10154 & ~n10177 ;
  assign n10179 = \P3_reg1_reg[23]/NET0131  & ~n2143 ;
  assign n10180 = \P3_reg1_reg[23]/NET0131  & n2145 ;
  assign n10181 = \P3_reg1_reg[23]/NET0131  & ~n2408 ;
  assign n10182 = n2408 & ~n7386 ;
  assign n10183 = ~n10181 & ~n10182 ;
  assign n10184 = n714 & ~n10183 ;
  assign n10185 = ~n8409 & ~n10181 ;
  assign n10186 = ~n2518 & ~n10185 ;
  assign n10187 = n886 & n6451 ;
  assign n10188 = \P3_reg1_reg[23]/NET0131  & ~n6449 ;
  assign n10195 = ~n10187 & ~n10188 ;
  assign n10196 = ~n10186 & n10195 ;
  assign n10189 = \P3_reg1_reg[23]/NET0131  & ~n2427 ;
  assign n10190 = n2427 & ~n7398 ;
  assign n10191 = ~n10189 & ~n10190 ;
  assign n10192 = n737 & ~n10191 ;
  assign n10193 = ~n8399 & ~n10189 ;
  assign n10194 = n2425 & ~n10193 ;
  assign n10197 = ~n10192 & ~n10194 ;
  assign n10198 = n10196 & n10197 ;
  assign n10199 = ~n10184 & n10198 ;
  assign n10200 = n2147 & ~n10199 ;
  assign n10201 = ~n10180 & ~n10200 ;
  assign n10202 = \P1_state_reg[0]/NET0131  & ~n10201 ;
  assign n10203 = ~n10179 & ~n10202 ;
  assign n10204 = \P3_reg2_reg[17]/NET0131  & ~n2143 ;
  assign n10205 = \P3_reg2_reg[17]/NET0131  & n2145 ;
  assign n10207 = \P3_reg2_reg[17]/NET0131  & ~n2427 ;
  assign n10208 = n2427 & ~n8601 ;
  assign n10209 = ~n10207 & ~n10208 ;
  assign n10210 = n714 & ~n10209 ;
  assign n10220 = ~n1166 & n2441 ;
  assign n10206 = \P3_reg2_reg[17]/NET0131  & ~n2429 ;
  assign n10219 = ~n1146 & n2283 ;
  assign n10221 = ~n10206 & ~n10219 ;
  assign n10222 = ~n10220 & n10221 ;
  assign n10223 = ~n10210 & n10222 ;
  assign n10217 = ~n10086 & ~n10207 ;
  assign n10218 = ~n2518 & ~n10217 ;
  assign n10211 = \P3_reg2_reg[17]/NET0131  & ~n2408 ;
  assign n10212 = ~n10092 & ~n10211 ;
  assign n10213 = n2425 & ~n10212 ;
  assign n10214 = n2408 & ~n8619 ;
  assign n10215 = ~n10211 & ~n10214 ;
  assign n10216 = n737 & ~n10215 ;
  assign n10224 = ~n10213 & ~n10216 ;
  assign n10225 = ~n10218 & n10224 ;
  assign n10226 = n10223 & n10225 ;
  assign n10227 = n2147 & ~n10226 ;
  assign n10228 = ~n10205 & ~n10227 ;
  assign n10229 = \P1_state_reg[0]/NET0131  & ~n10228 ;
  assign n10230 = ~n10204 & ~n10229 ;
  assign n10231 = \P3_reg2_reg[18]/NET0131  & ~n2143 ;
  assign n10232 = \P3_reg2_reg[18]/NET0131  & n2145 ;
  assign n10239 = \P3_reg2_reg[18]/NET0131  & ~n2427 ;
  assign n10242 = n2427 & n8559 ;
  assign n10243 = ~n10239 & ~n10242 ;
  assign n10244 = n714 & ~n10243 ;
  assign n10233 = \P3_reg2_reg[18]/NET0131  & ~n2408 ;
  assign n10234 = n2408 & ~n8574 ;
  assign n10235 = ~n10233 & ~n10234 ;
  assign n10236 = n737 & ~n10235 ;
  assign n10245 = n2427 & n9872 ;
  assign n10246 = ~n1116 & n2283 ;
  assign n10247 = \P3_reg2_reg[18]/NET0131  & ~n2429 ;
  assign n10248 = ~n10246 & ~n10247 ;
  assign n10249 = ~n10245 & n10248 ;
  assign n10250 = ~n10236 & n10249 ;
  assign n10237 = ~n10035 & ~n10233 ;
  assign n10238 = n2425 & ~n10237 ;
  assign n10240 = ~n10028 & ~n10239 ;
  assign n10241 = ~n2518 & ~n10240 ;
  assign n10251 = ~n10238 & ~n10241 ;
  assign n10252 = n10250 & n10251 ;
  assign n10253 = ~n10244 & n10252 ;
  assign n10254 = n2147 & ~n10253 ;
  assign n10255 = ~n10232 & ~n10254 ;
  assign n10256 = \P1_state_reg[0]/NET0131  & ~n10255 ;
  assign n10257 = ~n10231 & ~n10256 ;
  assign n10258 = \P1_reg1_reg[17]/NET0131  & ~n6078 ;
  assign n10259 = \P1_reg1_reg[17]/NET0131  & n6095 ;
  assign n10261 = \P1_reg1_reg[17]/NET0131  & ~n6683 ;
  assign n10262 = n6683 & ~n9420 ;
  assign n10263 = ~n10261 & ~n10262 ;
  assign n10264 = n6207 & ~n10263 ;
  assign n10268 = n6683 & n9433 ;
  assign n10269 = ~n10261 & ~n10268 ;
  assign n10270 = n6282 & ~n10269 ;
  assign n10271 = n6683 & n9441 ;
  assign n10272 = ~n10261 & ~n10271 ;
  assign n10273 = n4011 & ~n10272 ;
  assign n10265 = n6683 & n9425 ;
  assign n10266 = ~n10261 & ~n10265 ;
  assign n10267 = n6359 & ~n10266 ;
  assign n10260 = n6683 & n9446 ;
  assign n10274 = \P1_reg1_reg[17]/NET0131  & ~n7806 ;
  assign n10275 = ~n10260 & ~n10274 ;
  assign n10276 = ~n10267 & n10275 ;
  assign n10277 = ~n10273 & n10276 ;
  assign n10278 = ~n10270 & n10277 ;
  assign n10279 = ~n10264 & n10278 ;
  assign n10280 = n6097 & ~n10279 ;
  assign n10281 = ~n10259 & ~n10280 ;
  assign n10282 = \P1_state_reg[0]/NET0131  & ~n10281 ;
  assign n10283 = ~n10258 & ~n10282 ;
  assign n10286 = ~n1657 & n2145 ;
  assign n10301 = ~n1657 & ~n2163 ;
  assign n10305 = ~n1687 & n2239 ;
  assign n10306 = ~n1663 & n2251 ;
  assign n10307 = n1637 & ~n10306 ;
  assign n10308 = ~n2239 & ~n2253 ;
  assign n10309 = ~n10307 & n10308 ;
  assign n10310 = ~n10305 & ~n10309 ;
  assign n10311 = n2163 & ~n10310 ;
  assign n10312 = ~n10301 & ~n10311 ;
  assign n10313 = n737 & ~n10312 ;
  assign n10288 = ~n1657 & ~n2236 ;
  assign n10289 = n2067 & ~n2331 ;
  assign n10290 = ~n2067 & n2331 ;
  assign n10291 = ~n10289 & ~n10290 ;
  assign n10292 = n2236 & n10291 ;
  assign n10293 = ~n10288 & ~n10292 ;
  assign n10294 = n2391 & ~n10293 ;
  assign n10287 = ~n1677 & n2580 ;
  assign n10314 = ~n1657 & ~n2583 ;
  assign n10315 = ~n10287 & ~n10314 ;
  assign n10316 = ~n10294 & n10315 ;
  assign n10295 = n2067 & ~n2179 ;
  assign n10296 = ~n2067 & n2179 ;
  assign n10297 = ~n10295 & ~n10296 ;
  assign n10298 = n2236 & ~n10297 ;
  assign n10299 = ~n10288 & ~n10298 ;
  assign n10300 = n2234 & ~n10299 ;
  assign n10302 = n2163 & n10291 ;
  assign n10303 = ~n10301 & ~n10302 ;
  assign n10304 = n2393 & ~n10303 ;
  assign n10317 = ~n10300 & ~n10304 ;
  assign n10318 = n10316 & n10317 ;
  assign n10319 = ~n10313 & n10318 ;
  assign n10320 = n2147 & ~n10319 ;
  assign n10321 = ~n10286 & ~n10320 ;
  assign n10322 = \P1_state_reg[0]/NET0131  & ~n10321 ;
  assign n10284 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[9]/NET0131  ;
  assign n10285 = n765 & ~n1657 ;
  assign n10323 = ~n10284 & ~n10285 ;
  assign n10324 = ~n10322 & n10323 ;
  assign n10327 = ~n4231 & ~n4931 ;
  assign n10328 = ~n5040 & n5353 ;
  assign n10329 = ~n5008 & n10328 ;
  assign n10330 = ~n4984 & n10329 ;
  assign n10331 = ~n10327 & ~n10330 ;
  assign n10332 = ~n5357 & ~n10331 ;
  assign n10333 = n4231 & ~n5008 ;
  assign n10334 = ~n10332 & ~n10333 ;
  assign n10335 = n5383 & ~n10334 ;
  assign n10337 = n5992 & ~n7918 ;
  assign n10336 = ~n5992 & n7918 ;
  assign n10338 = n5526 & ~n10336 ;
  assign n10339 = ~n10337 & n10338 ;
  assign n10341 = n5992 & n7884 ;
  assign n10340 = ~n5992 & ~n7884 ;
  assign n10342 = n5329 & ~n10340 ;
  assign n10343 = ~n10341 & n10342 ;
  assign n10344 = ~n10339 & ~n10343 ;
  assign n10345 = ~n10335 & n10344 ;
  assign n10346 = n7453 & ~n10345 ;
  assign n10349 = ~n5022 & n5536 ;
  assign n10350 = ~n4997 & ~n10349 ;
  assign n10351 = ~n5538 & ~n10350 ;
  assign n10352 = n7453 & ~n10351 ;
  assign n10353 = ~n4978 & ~n7453 ;
  assign n10354 = n5563 & ~n10353 ;
  assign n10355 = ~n10352 & n10354 ;
  assign n10326 = ~n4997 & ~n7504 ;
  assign n10347 = n7641 & ~n9400 ;
  assign n10348 = n4978 & ~n10347 ;
  assign n10356 = ~n10326 & ~n10348 ;
  assign n10357 = ~n10355 & n10356 ;
  assign n10358 = ~n10346 & n10357 ;
  assign n10359 = n5583 & ~n10358 ;
  assign n10360 = ~n5582 & ~n8640 ;
  assign n10361 = n4978 & ~n5316 ;
  assign n10362 = ~n10360 & n10361 ;
  assign n10363 = ~n10359 & ~n10362 ;
  assign n10364 = \P1_state_reg[0]/NET0131  & ~n10363 ;
  assign n10325 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[10]/NET0131  ;
  assign n10365 = n4978 & n5786 ;
  assign n10366 = ~n10325 & ~n10365 ;
  assign n10367 = ~n10364 & n10366 ;
  assign n10370 = n4952 & n5585 ;
  assign n10372 = n4952 & ~n7453 ;
  assign n10379 = ~n4958 & n5357 ;
  assign n10380 = n4854 & ~n10379 ;
  assign n10381 = ~n4854 & n10379 ;
  assign n10382 = ~n10380 & ~n10381 ;
  assign n10383 = ~n4231 & ~n10382 ;
  assign n10384 = n4231 & n4931 ;
  assign n10385 = ~n10383 & ~n10384 ;
  assign n10386 = n7453 & n10385 ;
  assign n10387 = ~n10372 & ~n10386 ;
  assign n10388 = n5383 & ~n10387 ;
  assign n10373 = n5996 & ~n6755 ;
  assign n10374 = ~n5996 & n6755 ;
  assign n10375 = ~n10373 & ~n10374 ;
  assign n10376 = n7453 & n10375 ;
  assign n10377 = ~n10372 & ~n10376 ;
  assign n10378 = n5329 & ~n10377 ;
  assign n10389 = n5996 & ~n6805 ;
  assign n10390 = ~n5996 & n6805 ;
  assign n10391 = ~n10389 & ~n10390 ;
  assign n10392 = n7453 & ~n10391 ;
  assign n10393 = ~n10372 & ~n10392 ;
  assign n10394 = n5526 & ~n10393 ;
  assign n10395 = ~n4948 & n5538 ;
  assign n10396 = n4973 & ~n10395 ;
  assign n10397 = ~n5540 & ~n10396 ;
  assign n10398 = n7453 & n10397 ;
  assign n10399 = ~n10372 & ~n10398 ;
  assign n10400 = n5563 & ~n10399 ;
  assign n10371 = n4973 & ~n7504 ;
  assign n10401 = n4952 & ~n7641 ;
  assign n10402 = ~n10371 & ~n10401 ;
  assign n10403 = ~n10400 & n10402 ;
  assign n10404 = ~n10394 & n10403 ;
  assign n10405 = ~n10378 & n10404 ;
  assign n10406 = ~n10388 & n10405 ;
  assign n10407 = n5583 & ~n10406 ;
  assign n10408 = ~n10370 & ~n10407 ;
  assign n10409 = \P1_state_reg[0]/NET0131  & ~n10408 ;
  assign n10368 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[12]/NET0131  ;
  assign n10369 = n4952 & n5786 ;
  assign n10410 = ~n10368 & ~n10369 ;
  assign n10411 = ~n10409 & n10410 ;
  assign n10413 = n4849 & n5585 ;
  assign n10433 = ~n5269 & n6000 ;
  assign n10432 = n5269 & ~n6000 ;
  assign n10434 = n5329 & ~n10432 ;
  assign n10435 = ~n10433 & n10434 ;
  assign n10417 = n4827 & ~n10381 ;
  assign n10418 = ~n4827 & n10381 ;
  assign n10419 = ~n10417 & ~n10418 ;
  assign n10420 = ~n4231 & ~n10419 ;
  assign n10421 = n4231 & n4958 ;
  assign n10422 = n5383 & ~n10421 ;
  assign n10423 = ~n10420 & n10422 ;
  assign n10425 = n4867 & ~n5540 ;
  assign n10424 = ~n4867 & n5540 ;
  assign n10426 = n5563 & ~n10424 ;
  assign n10427 = ~n10425 & n10426 ;
  assign n10429 = ~n5455 & ~n6000 ;
  assign n10428 = n5455 & n6000 ;
  assign n10430 = n5526 & ~n10428 ;
  assign n10431 = ~n10429 & n10430 ;
  assign n10436 = ~n10427 & ~n10431 ;
  assign n10437 = ~n10423 & n10436 ;
  assign n10438 = ~n10435 & n10437 ;
  assign n10439 = n7453 & ~n10438 ;
  assign n10414 = n7484 & ~n8640 ;
  assign n10415 = ~n9400 & n10414 ;
  assign n10416 = n4849 & ~n10415 ;
  assign n10440 = n4867 & ~n7504 ;
  assign n10441 = ~n10416 & ~n10440 ;
  assign n10442 = ~n10439 & n10441 ;
  assign n10443 = n5583 & ~n10442 ;
  assign n10444 = ~n10413 & ~n10443 ;
  assign n10445 = \P1_state_reg[0]/NET0131  & ~n10444 ;
  assign n10412 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[13]/NET0131  ;
  assign n10446 = n4849 & n5786 ;
  assign n10447 = ~n10412 & ~n10446 ;
  assign n10448 = ~n10445 & n10447 ;
  assign n10450 = n5003 & n5585 ;
  assign n10452 = n5003 & ~n7453 ;
  assign n10453 = n4984 & ~n10329 ;
  assign n10454 = ~n10330 & ~n10453 ;
  assign n10455 = ~n4231 & ~n10454 ;
  assign n10456 = n4231 & n5040 ;
  assign n10457 = ~n10455 & ~n10456 ;
  assign n10458 = n7453 & n10457 ;
  assign n10459 = ~n10452 & ~n10458 ;
  assign n10460 = n5383 & ~n10459 ;
  assign n10462 = n5449 & n5975 ;
  assign n10461 = ~n5449 & ~n5975 ;
  assign n10463 = n5526 & ~n10461 ;
  assign n10464 = ~n10462 & n10463 ;
  assign n10466 = ~n5264 & n5975 ;
  assign n10465 = n5264 & ~n5975 ;
  assign n10467 = n5329 & ~n10465 ;
  assign n10468 = ~n10466 & n10467 ;
  assign n10469 = ~n10464 & ~n10468 ;
  assign n10470 = n7453 & ~n10469 ;
  assign n10471 = n5022 & ~n5536 ;
  assign n10472 = ~n10349 & ~n10471 ;
  assign n10473 = n7453 & n10472 ;
  assign n10474 = ~n10452 & ~n10473 ;
  assign n10475 = n5563 & ~n10474 ;
  assign n10451 = n5022 & ~n7504 ;
  assign n10476 = n5003 & ~n10347 ;
  assign n10477 = ~n10451 & ~n10476 ;
  assign n10478 = ~n10475 & n10477 ;
  assign n10479 = ~n10470 & n10478 ;
  assign n10480 = ~n10460 & n10479 ;
  assign n10481 = n5583 & ~n10480 ;
  assign n10482 = ~n10450 & ~n10481 ;
  assign n10483 = \P1_state_reg[0]/NET0131  & ~n10482 ;
  assign n10449 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[9]/NET0131  ;
  assign n10484 = n5003 & n5786 ;
  assign n10485 = ~n10449 & ~n10484 ;
  assign n10486 = ~n10483 & n10485 ;
  assign n10489 = ~n1631 & n2145 ;
  assign n10498 = ~n1631 & ~n2236 ;
  assign n10492 = n2053 & ~n5738 ;
  assign n10493 = ~n2053 & n5738 ;
  assign n10494 = ~n10492 & ~n10493 ;
  assign n10499 = n2236 & n10494 ;
  assign n10500 = ~n10498 & ~n10499 ;
  assign n10501 = n2391 & ~n10500 ;
  assign n10491 = ~n1631 & ~n2163 ;
  assign n10495 = n2163 & n10494 ;
  assign n10496 = ~n10491 & ~n10495 ;
  assign n10497 = n2393 & ~n10496 ;
  assign n10503 = ~n1613 & n2253 ;
  assign n10502 = n1613 & ~n2253 ;
  assign n10504 = ~n2239 & ~n10502 ;
  assign n10505 = ~n10503 & n10504 ;
  assign n10506 = ~n1663 & n2239 ;
  assign n10507 = ~n10505 & ~n10506 ;
  assign n10508 = n2163 & ~n10507 ;
  assign n10509 = ~n10491 & ~n10508 ;
  assign n10510 = n737 & ~n10509 ;
  assign n10511 = n2053 & ~n5703 ;
  assign n10512 = ~n2053 & n5703 ;
  assign n10513 = ~n10511 & ~n10512 ;
  assign n10514 = n2236 & ~n10513 ;
  assign n10515 = ~n10498 & ~n10514 ;
  assign n10516 = n2234 & ~n10515 ;
  assign n10490 = ~n1651 & n2580 ;
  assign n10517 = ~n1631 & ~n2583 ;
  assign n10518 = ~n10490 & ~n10517 ;
  assign n10519 = ~n10516 & n10518 ;
  assign n10520 = ~n10510 & n10519 ;
  assign n10521 = ~n10497 & n10520 ;
  assign n10522 = ~n10501 & n10521 ;
  assign n10523 = n2147 & ~n10522 ;
  assign n10524 = ~n10489 & ~n10523 ;
  assign n10525 = \P1_state_reg[0]/NET0131  & ~n10524 ;
  assign n10487 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[10]/NET0131  ;
  assign n10488 = n765 & ~n1631 ;
  assign n10526 = ~n10487 & ~n10488 ;
  assign n10527 = ~n10525 & n10526 ;
  assign n10530 = ~n1608 & n2145 ;
  assign n10532 = ~n1608 & ~n2163 ;
  assign n10533 = n2050 & ~n2538 ;
  assign n10534 = ~n2050 & n2538 ;
  assign n10535 = ~n10533 & ~n10534 ;
  assign n10536 = n2163 & n10535 ;
  assign n10537 = ~n10532 & ~n10536 ;
  assign n10538 = n2393 & ~n10537 ;
  assign n10539 = ~n1608 & ~n2236 ;
  assign n10551 = n2050 & ~n2593 ;
  assign n10552 = ~n2050 & n2593 ;
  assign n10553 = ~n10551 & ~n10552 ;
  assign n10554 = n2236 & ~n10553 ;
  assign n10555 = ~n10539 & ~n10554 ;
  assign n10556 = n2234 & ~n10555 ;
  assign n10531 = ~n1627 & n2580 ;
  assign n10557 = ~n1608 & ~n2583 ;
  assign n10558 = ~n10531 & ~n10557 ;
  assign n10559 = ~n10556 & n10558 ;
  assign n10560 = ~n10538 & n10559 ;
  assign n10540 = n2236 & n10535 ;
  assign n10541 = ~n10539 & ~n10540 ;
  assign n10542 = n2391 & ~n10541 ;
  assign n10543 = ~n1637 & n2239 ;
  assign n10544 = n1594 & ~n10503 ;
  assign n10545 = ~n2239 & ~n2255 ;
  assign n10546 = ~n10544 & n10545 ;
  assign n10547 = ~n10543 & ~n10546 ;
  assign n10548 = n2163 & ~n10547 ;
  assign n10549 = ~n10532 & ~n10548 ;
  assign n10550 = n737 & ~n10549 ;
  assign n10561 = ~n10542 & ~n10550 ;
  assign n10562 = n10560 & n10561 ;
  assign n10563 = n2147 & ~n10562 ;
  assign n10564 = ~n10530 & ~n10563 ;
  assign n10565 = \P1_state_reg[0]/NET0131  & ~n10564 ;
  assign n10528 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[11]/NET0131  ;
  assign n10529 = n765 & ~n1608 ;
  assign n10566 = ~n10528 & ~n10529 ;
  assign n10567 = ~n10565 & n10566 ;
  assign n10570 = ~n1589 & n2145 ;
  assign n10572 = ~n1589 & ~n2163 ;
  assign n10586 = n1569 & ~n2255 ;
  assign n10587 = ~n2239 & ~n9148 ;
  assign n10588 = ~n10586 & n10587 ;
  assign n10589 = ~n1613 & n2239 ;
  assign n10590 = ~n10588 & ~n10589 ;
  assign n10591 = n2163 & ~n10590 ;
  assign n10592 = ~n10572 & ~n10591 ;
  assign n10593 = n737 & ~n10592 ;
  assign n10579 = ~n1589 & ~n2236 ;
  assign n10580 = ~n2011 & n2077 ;
  assign n10581 = n2011 & ~n2077 ;
  assign n10582 = ~n10580 & ~n10581 ;
  assign n10583 = n2236 & ~n10582 ;
  assign n10584 = ~n10579 & ~n10583 ;
  assign n10585 = n2234 & ~n10584 ;
  assign n10571 = n1584 & n2580 ;
  assign n10597 = ~n1589 & ~n2583 ;
  assign n10598 = ~n10571 & ~n10597 ;
  assign n10599 = ~n10585 & n10598 ;
  assign n10600 = ~n10593 & n10599 ;
  assign n10573 = n2077 & ~n2468 ;
  assign n10574 = ~n2077 & n2468 ;
  assign n10575 = ~n10573 & ~n10574 ;
  assign n10576 = n2163 & n10575 ;
  assign n10577 = ~n10572 & ~n10576 ;
  assign n10578 = n2393 & ~n10577 ;
  assign n10594 = n2236 & n10575 ;
  assign n10595 = ~n10579 & ~n10594 ;
  assign n10596 = n2391 & ~n10595 ;
  assign n10601 = ~n10578 & ~n10596 ;
  assign n10602 = n10600 & n10601 ;
  assign n10603 = n2147 & ~n10602 ;
  assign n10604 = ~n10570 & ~n10603 ;
  assign n10605 = \P1_state_reg[0]/NET0131  & ~n10604 ;
  assign n10568 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[12]/NET0131  ;
  assign n10569 = n765 & ~n1589 ;
  assign n10606 = ~n10568 & ~n10569 ;
  assign n10607 = ~n10605 & n10606 ;
  assign n10610 = ~n1564 & n2145 ;
  assign n10612 = ~n1564 & ~n2163 ;
  assign n10625 = n1531 & ~n9148 ;
  assign n10624 = ~n1531 & n9148 ;
  assign n10626 = ~n2239 & ~n10624 ;
  assign n10627 = ~n10625 & n10626 ;
  assign n10628 = ~n1594 & n2239 ;
  assign n10629 = ~n10627 & ~n10628 ;
  assign n10630 = n2163 & ~n10629 ;
  assign n10631 = ~n10612 & ~n10630 ;
  assign n10632 = n737 & ~n10631 ;
  assign n10613 = n2084 & ~n2342 ;
  assign n10614 = ~n2084 & n2342 ;
  assign n10615 = ~n10613 & ~n10614 ;
  assign n10616 = n2163 & n10615 ;
  assign n10617 = ~n10612 & ~n10616 ;
  assign n10618 = n2393 & ~n10617 ;
  assign n10611 = ~n1560 & n2580 ;
  assign n10619 = ~n1564 & ~n2583 ;
  assign n10639 = ~n10611 & ~n10619 ;
  assign n10640 = ~n10618 & n10639 ;
  assign n10620 = ~n1564 & ~n2236 ;
  assign n10621 = n2236 & n10615 ;
  assign n10622 = ~n10620 & ~n10621 ;
  assign n10623 = n2391 & ~n10622 ;
  assign n10633 = n2084 & ~n2189 ;
  assign n10634 = ~n2084 & n2189 ;
  assign n10635 = ~n10633 & ~n10634 ;
  assign n10636 = n2236 & ~n10635 ;
  assign n10637 = ~n10620 & ~n10636 ;
  assign n10638 = n2234 & ~n10637 ;
  assign n10641 = ~n10623 & ~n10638 ;
  assign n10642 = n10640 & n10641 ;
  assign n10643 = ~n10632 & n10642 ;
  assign n10644 = n2147 & ~n10643 ;
  assign n10645 = ~n10610 & ~n10644 ;
  assign n10646 = \P1_state_reg[0]/NET0131  & ~n10645 ;
  assign n10608 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[13]/NET0131  ;
  assign n10609 = n765 & ~n1564 ;
  assign n10647 = ~n10608 & ~n10609 ;
  assign n10648 = ~n10646 & n10647 ;
  assign n10651 = ~n1525 & n2145 ;
  assign n10653 = ~n1525 & ~n2163 ;
  assign n10663 = n2046 & ~n7336 ;
  assign n10664 = ~n2046 & n7336 ;
  assign n10665 = ~n10663 & ~n10664 ;
  assign n10669 = n2163 & ~n10665 ;
  assign n10670 = ~n10653 & ~n10669 ;
  assign n10671 = n2393 & ~n10670 ;
  assign n10662 = ~n1525 & ~n2236 ;
  assign n10666 = n2236 & ~n10665 ;
  assign n10667 = ~n10662 & ~n10666 ;
  assign n10668 = n2391 & ~n10667 ;
  assign n10654 = n1521 & ~n10624 ;
  assign n10655 = ~n2239 & ~n9149 ;
  assign n10656 = ~n10654 & n10655 ;
  assign n10657 = ~n1569 & n2239 ;
  assign n10658 = ~n10656 & ~n10657 ;
  assign n10659 = n2163 & ~n10658 ;
  assign n10660 = ~n10653 & ~n10659 ;
  assign n10661 = n737 & ~n10660 ;
  assign n10672 = n2046 & ~n5708 ;
  assign n10673 = ~n2046 & n5708 ;
  assign n10674 = ~n10672 & ~n10673 ;
  assign n10675 = n2236 & n10674 ;
  assign n10676 = ~n10662 & ~n10675 ;
  assign n10677 = n2234 & ~n10676 ;
  assign n10652 = ~n1544 & n2580 ;
  assign n10678 = ~n1525 & ~n2583 ;
  assign n10679 = ~n10652 & ~n10678 ;
  assign n10680 = ~n10677 & n10679 ;
  assign n10681 = ~n10661 & n10680 ;
  assign n10682 = ~n10668 & n10681 ;
  assign n10683 = ~n10671 & n10682 ;
  assign n10684 = n2147 & ~n10683 ;
  assign n10685 = ~n10651 & ~n10684 ;
  assign n10686 = \P1_state_reg[0]/NET0131  & ~n10685 ;
  assign n10649 = n765 & ~n1525 ;
  assign n10650 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[14]/NET0131  ;
  assign n10687 = ~n10649 & ~n10650 ;
  assign n10688 = ~n10686 & n10687 ;
  assign n10691 = n3593 & n6095 ;
  assign n10693 = n3593 & ~n6568 ;
  assign n10700 = n3303 & ~n9240 ;
  assign n10701 = ~n9307 & ~n10700 ;
  assign n10702 = ~n2713 & ~n10701 ;
  assign n10703 = n2713 & n2952 ;
  assign n10704 = ~n10702 & ~n10703 ;
  assign n10705 = n6568 & n10704 ;
  assign n10706 = ~n10693 & ~n10705 ;
  assign n10707 = n4011 & ~n10706 ;
  assign n10694 = n3600 & ~n4059 ;
  assign n10695 = ~n3600 & n4059 ;
  assign n10696 = ~n10694 & ~n10695 ;
  assign n10697 = n6568 & ~n10696 ;
  assign n10698 = ~n10693 & ~n10697 ;
  assign n10699 = n6282 & ~n10698 ;
  assign n10708 = n3600 & n7677 ;
  assign n10709 = ~n3600 & ~n7677 ;
  assign n10710 = ~n10708 & ~n10709 ;
  assign n10711 = n6568 & ~n10710 ;
  assign n10712 = ~n10693 & ~n10711 ;
  assign n10713 = n6207 & ~n10712 ;
  assign n10714 = n3588 & ~n8659 ;
  assign n10715 = ~n8660 & ~n10714 ;
  assign n10716 = n6359 & n10715 ;
  assign n10717 = n6568 & n10716 ;
  assign n10692 = n3593 & ~n7036 ;
  assign n10718 = n3588 & ~n6649 ;
  assign n10719 = ~n10692 & ~n10718 ;
  assign n10720 = ~n10717 & n10719 ;
  assign n10721 = ~n10713 & n10720 ;
  assign n10722 = ~n10699 & n10721 ;
  assign n10723 = ~n10707 & n10722 ;
  assign n10724 = n6097 & ~n10723 ;
  assign n10725 = ~n10691 & ~n10724 ;
  assign n10726 = \P1_state_reg[0]/NET0131  & ~n10725 ;
  assign n10689 = n3593 & n4130 ;
  assign n10690 = \P1_reg3_reg[20]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n10727 = ~n10689 & ~n10690 ;
  assign n10728 = ~n10726 & n10727 ;
  assign n10729 = n4661 & ~n7453 ;
  assign n10730 = ~n7535 & n7536 ;
  assign n10731 = n7542 & ~n10730 ;
  assign n10732 = n5986 & ~n10731 ;
  assign n10733 = ~n5986 & n10731 ;
  assign n10734 = ~n10732 & ~n10733 ;
  assign n10735 = n7453 & ~n10734 ;
  assign n10736 = ~n10729 & ~n10735 ;
  assign n10737 = n5526 & ~n10736 ;
  assign n10738 = ~n7558 & n7559 ;
  assign n10739 = n7564 & ~n10738 ;
  assign n10740 = n7560 & n7571 ;
  assign n10741 = ~n10739 & n10740 ;
  assign n10742 = ~n7567 & n7571 ;
  assign n10743 = n7576 & ~n10742 ;
  assign n10744 = ~n10741 & n10743 ;
  assign n10745 = n5986 & n10744 ;
  assign n10746 = ~n5986 & ~n10744 ;
  assign n10747 = ~n10745 & ~n10746 ;
  assign n10748 = n7453 & ~n10747 ;
  assign n10749 = ~n10729 & ~n10748 ;
  assign n10750 = n5329 & ~n10749 ;
  assign n10753 = ~n4647 & n7593 ;
  assign n10754 = n4647 & ~n7593 ;
  assign n10755 = ~n10753 & ~n10754 ;
  assign n10756 = ~n4231 & ~n10755 ;
  assign n10752 = n4231 & n4684 ;
  assign n10757 = n5383 & ~n10752 ;
  assign n10758 = ~n10756 & n10757 ;
  assign n10759 = n4656 & ~n7496 ;
  assign n10760 = n5563 & ~n7845 ;
  assign n10761 = ~n10759 & n10760 ;
  assign n10762 = ~n10758 & ~n10761 ;
  assign n10763 = n7453 & ~n10762 ;
  assign n10751 = n4661 & ~n10414 ;
  assign n10764 = n4656 & ~n7504 ;
  assign n10765 = ~n10751 & ~n10764 ;
  assign n10766 = ~n10763 & n10765 ;
  assign n10767 = ~n10750 & n10766 ;
  assign n10768 = ~n10737 & n10767 ;
  assign n10769 = n5583 & ~n10768 ;
  assign n10770 = n4661 & n5585 ;
  assign n10771 = ~n10769 & ~n10770 ;
  assign n10772 = \P1_state_reg[0]/NET0131  & ~n10771 ;
  assign n10773 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[23]/NET0131  ;
  assign n10774 = n4661 & n5786 ;
  assign n10775 = ~n10773 & ~n10774 ;
  assign n10776 = ~n10772 & n10775 ;
  assign n10777 = \P2_reg0_reg[20]/NET0131  & ~n5589 ;
  assign n10778 = \P2_reg0_reg[20]/NET0131  & n5585 ;
  assign n10780 = \P2_reg0_reg[20]/NET0131  & ~n6706 ;
  assign n10784 = n6706 & n9276 ;
  assign n10785 = ~n10780 & ~n10784 ;
  assign n10786 = n5383 & ~n10785 ;
  assign n10781 = n6706 & ~n9267 ;
  assign n10782 = ~n10780 & ~n10781 ;
  assign n10783 = n5329 & ~n10782 ;
  assign n10787 = n6706 & ~n9282 ;
  assign n10788 = ~n10780 & ~n10787 ;
  assign n10789 = n5526 & ~n10788 ;
  assign n10779 = \P2_reg0_reg[20]/NET0131  & ~n6717 ;
  assign n10790 = n6706 & ~n9759 ;
  assign n10791 = ~n10779 & ~n10790 ;
  assign n10792 = ~n10789 & n10791 ;
  assign n10793 = ~n10783 & n10792 ;
  assign n10794 = ~n10786 & n10793 ;
  assign n10795 = n5583 & ~n10794 ;
  assign n10796 = ~n10778 & ~n10795 ;
  assign n10797 = \P1_state_reg[0]/NET0131  & ~n10796 ;
  assign n10798 = ~n10777 & ~n10797 ;
  assign n10799 = \P2_reg0_reg[21]/NET0131  & ~n9531 ;
  assign n10800 = n9533 & ~n9640 ;
  assign n10801 = ~n10799 & ~n10800 ;
  assign n10802 = \P1_reg1_reg[30]/NET0131  & ~n6078 ;
  assign n10803 = \P1_reg1_reg[30]/NET0131  & n6095 ;
  assign n10804 = \P1_reg1_reg[30]/NET0131  & ~n6683 ;
  assign n10809 = n3500 & ~n6354 ;
  assign n10810 = ~n8716 & ~n10809 ;
  assign n10811 = n6683 & n10810 ;
  assign n10812 = ~n10804 & ~n10811 ;
  assign n10813 = n6359 & ~n10812 ;
  assign n10805 = n3500 & n6683 ;
  assign n10806 = ~n10804 & ~n10805 ;
  assign n10807 = n6365 & ~n10806 ;
  assign n10808 = \P1_reg1_reg[30]/NET0131  & ~n9547 ;
  assign n10814 = ~n10807 & ~n10808 ;
  assign n10815 = ~n9550 & n10814 ;
  assign n10816 = ~n10813 & n10815 ;
  assign n10817 = n6097 & ~n10816 ;
  assign n10818 = ~n10803 & ~n10817 ;
  assign n10819 = \P1_state_reg[0]/NET0131  & ~n10818 ;
  assign n10820 = ~n10802 & ~n10819 ;
  assign n10821 = \P1_reg2_reg[12]/NET0131  & ~n6078 ;
  assign n10822 = \P1_reg2_reg[12]/NET0131  & n6095 ;
  assign n10824 = \P1_reg2_reg[12]/NET0131  & ~n6113 ;
  assign n10825 = n6113 & n9071 ;
  assign n10826 = ~n10824 & ~n10825 ;
  assign n10827 = n4011 & ~n10826 ;
  assign n10828 = n3641 & n6365 ;
  assign n10829 = n9081 & ~n10828 ;
  assign n10830 = n6113 & ~n10829 ;
  assign n10831 = n6113 & n9061 ;
  assign n10832 = ~n10824 & ~n10831 ;
  assign n10833 = n6359 & ~n10832 ;
  assign n10823 = n3645 & n4112 ;
  assign n10834 = ~n6113 & ~n8656 ;
  assign n10835 = n8955 & ~n10834 ;
  assign n10836 = \P1_reg2_reg[12]/NET0131  & ~n10835 ;
  assign n10837 = ~n10823 & ~n10836 ;
  assign n10838 = ~n10833 & n10837 ;
  assign n10839 = ~n10830 & n10838 ;
  assign n10840 = ~n10827 & n10839 ;
  assign n10841 = n6097 & ~n10840 ;
  assign n10842 = ~n10822 & ~n10841 ;
  assign n10843 = \P1_state_reg[0]/NET0131  & ~n10842 ;
  assign n10844 = ~n10821 & ~n10843 ;
  assign n10845 = \P1_reg2_reg[16]/NET0131  & ~n6078 ;
  assign n10846 = \P1_reg2_reg[16]/NET0131  & n6095 ;
  assign n10849 = \P1_reg2_reg[16]/NET0131  & ~n6113 ;
  assign n10850 = n6113 & ~n9105 ;
  assign n10851 = ~n10849 & ~n10850 ;
  assign n10852 = n6207 & ~n10851 ;
  assign n10856 = n6113 & ~n9118 ;
  assign n10857 = ~n10849 & ~n10856 ;
  assign n10858 = n6282 & ~n10857 ;
  assign n10859 = n6113 & n9112 ;
  assign n10860 = ~n10849 & ~n10859 ;
  assign n10861 = n6359 & ~n10860 ;
  assign n10853 = n6113 & n9127 ;
  assign n10854 = ~n10849 & ~n10853 ;
  assign n10855 = n4011 & ~n10854 ;
  assign n10847 = n3194 & n6365 ;
  assign n10848 = n6113 & n10847 ;
  assign n10862 = n3199 & n4112 ;
  assign n10863 = \P1_reg2_reg[16]/NET0131  & ~n8955 ;
  assign n10864 = ~n10862 & ~n10863 ;
  assign n10865 = ~n10848 & n10864 ;
  assign n10866 = ~n10855 & n10865 ;
  assign n10867 = ~n10861 & n10866 ;
  assign n10868 = ~n10858 & n10867 ;
  assign n10869 = ~n10852 & n10868 ;
  assign n10870 = n6097 & ~n10869 ;
  assign n10871 = ~n10846 & ~n10870 ;
  assign n10872 = \P1_state_reg[0]/NET0131  & ~n10871 ;
  assign n10873 = ~n10845 & ~n10872 ;
  assign n10874 = \P1_reg2_reg[18]/NET0131  & ~n6078 ;
  assign n10875 = \P1_reg2_reg[18]/NET0131  & n6095 ;
  assign n10878 = \P1_reg2_reg[18]/NET0131  & ~n6113 ;
  assign n10879 = n6113 & ~n9193 ;
  assign n10880 = ~n10878 & ~n10879 ;
  assign n10881 = n6282 & ~n10880 ;
  assign n10885 = n6113 & n9199 ;
  assign n10886 = ~n10878 & ~n10885 ;
  assign n10887 = n6359 & ~n10886 ;
  assign n10882 = n6113 & n9205 ;
  assign n10883 = ~n10878 & ~n10882 ;
  assign n10884 = n6207 & ~n10883 ;
  assign n10888 = n6113 & n9214 ;
  assign n10889 = ~n10878 & ~n10888 ;
  assign n10890 = n4011 & ~n10889 ;
  assign n10876 = n3100 & n6365 ;
  assign n10877 = n6113 & n10876 ;
  assign n10891 = n3102 & n4112 ;
  assign n10892 = \P1_reg2_reg[18]/NET0131  & ~n8955 ;
  assign n10893 = ~n10891 & ~n10892 ;
  assign n10894 = ~n10877 & n10893 ;
  assign n10895 = ~n10890 & n10894 ;
  assign n10896 = ~n10884 & n10895 ;
  assign n10897 = ~n10887 & n10896 ;
  assign n10898 = ~n10881 & n10897 ;
  assign n10899 = n6097 & ~n10898 ;
  assign n10900 = ~n10875 & ~n10899 ;
  assign n10901 = \P1_state_reg[0]/NET0131  & ~n10900 ;
  assign n10902 = ~n10874 & ~n10901 ;
  assign n10903 = \P1_reg2_reg[20]/NET0131  & ~n6078 ;
  assign n10904 = \P1_reg2_reg[20]/NET0131  & n6095 ;
  assign n10907 = \P1_reg2_reg[20]/NET0131  & ~n6113 ;
  assign n10911 = n6113 & n10704 ;
  assign n10912 = ~n10907 & ~n10911 ;
  assign n10913 = n4011 & ~n10912 ;
  assign n10908 = n6113 & ~n10696 ;
  assign n10909 = ~n10907 & ~n10908 ;
  assign n10910 = n6282 & ~n10909 ;
  assign n10914 = n6113 & ~n10710 ;
  assign n10915 = ~n10907 & ~n10914 ;
  assign n10916 = n6207 & ~n10915 ;
  assign n10917 = n6113 & n10715 ;
  assign n10918 = ~n10907 & ~n10917 ;
  assign n10919 = n6359 & ~n10918 ;
  assign n10905 = n3588 & n6365 ;
  assign n10906 = n6113 & n10905 ;
  assign n10920 = n3593 & n4112 ;
  assign n10921 = \P1_reg2_reg[20]/NET0131  & ~n8955 ;
  assign n10922 = ~n10920 & ~n10921 ;
  assign n10923 = ~n10906 & n10922 ;
  assign n10924 = ~n10919 & n10923 ;
  assign n10925 = ~n10916 & n10924 ;
  assign n10926 = ~n10910 & n10925 ;
  assign n10927 = ~n10913 & n10926 ;
  assign n10928 = n6097 & ~n10927 ;
  assign n10929 = ~n10904 & ~n10928 ;
  assign n10930 = \P1_state_reg[0]/NET0131  & ~n10929 ;
  assign n10931 = ~n10903 & ~n10930 ;
  assign n10932 = \P2_reg1_reg[20]/NET0131  & ~n5589 ;
  assign n10933 = \P2_reg1_reg[20]/NET0131  & n5585 ;
  assign n10935 = \P2_reg1_reg[20]/NET0131  & ~n6380 ;
  assign n10939 = n6380 & n9276 ;
  assign n10940 = ~n10935 & ~n10939 ;
  assign n10941 = n5383 & ~n10940 ;
  assign n10936 = n6380 & ~n9267 ;
  assign n10937 = ~n10935 & ~n10936 ;
  assign n10938 = n5329 & ~n10937 ;
  assign n10942 = n6380 & ~n9282 ;
  assign n10943 = ~n10935 & ~n10942 ;
  assign n10944 = n5526 & ~n10943 ;
  assign n10934 = \P2_reg1_reg[20]/NET0131  & ~n6397 ;
  assign n10945 = n6380 & ~n9759 ;
  assign n10946 = ~n10934 & ~n10945 ;
  assign n10947 = ~n10944 & n10946 ;
  assign n10948 = ~n10938 & n10947 ;
  assign n10949 = ~n10941 & n10948 ;
  assign n10950 = n5583 & ~n10949 ;
  assign n10951 = ~n10933 & ~n10950 ;
  assign n10952 = \P1_state_reg[0]/NET0131  & ~n10951 ;
  assign n10953 = ~n10932 & ~n10952 ;
  assign n10954 = n2942 & n6365 ;
  assign n10955 = n9251 & ~n10954 ;
  assign n10956 = n6113 & ~n10955 ;
  assign n10957 = n2945 & n4112 ;
  assign n10958 = ~n10956 & ~n10957 ;
  assign n10959 = n9044 & ~n10958 ;
  assign n10962 = ~n6113 & n6693 ;
  assign n10960 = ~n6361 & n9044 ;
  assign n10961 = ~n6113 & ~n9545 ;
  assign n10963 = n10960 & ~n10961 ;
  assign n10964 = ~n10962 & n10963 ;
  assign n10965 = \P1_reg2_reg[19]/NET0131  & ~n10964 ;
  assign n10966 = ~n10959 & ~n10965 ;
  assign n10967 = \P1_reg2_reg[23]/NET0131  & ~n6078 ;
  assign n10968 = \P1_reg2_reg[23]/NET0131  & n6095 ;
  assign n10969 = \P1_reg2_reg[23]/NET0131  & ~n6113 ;
  assign n10970 = ~n6589 & n6590 ;
  assign n10971 = n6596 & ~n10970 ;
  assign n10972 = n3286 & ~n10971 ;
  assign n10973 = ~n3286 & n10971 ;
  assign n10974 = ~n10972 & ~n10973 ;
  assign n10975 = n6113 & ~n10974 ;
  assign n10976 = ~n10969 & ~n10975 ;
  assign n10977 = n6282 & ~n10976 ;
  assign n10978 = n3273 & n6365 ;
  assign n10988 = ~n6619 & n6622 ;
  assign n10989 = n6607 & n6631 ;
  assign n10990 = ~n10988 & n10989 ;
  assign n10991 = ~n6625 & n6631 ;
  assign n10992 = ~n6636 & ~n10991 ;
  assign n10993 = ~n10990 & n10992 ;
  assign n10995 = n3286 & ~n10993 ;
  assign n10994 = ~n3286 & n10993 ;
  assign n10996 = n6207 & ~n10994 ;
  assign n10997 = ~n10995 & n10996 ;
  assign n10979 = n2713 & ~n2887 ;
  assign n10980 = n3548 & ~n8668 ;
  assign n10981 = ~n2713 & ~n7038 ;
  assign n10982 = ~n10980 & n10981 ;
  assign n10983 = ~n10979 & ~n10982 ;
  assign n10984 = n4011 & ~n10983 ;
  assign n10985 = n3273 & ~n8663 ;
  assign n10986 = ~n6350 & n6359 ;
  assign n10987 = ~n10985 & n10986 ;
  assign n10998 = ~n10984 & ~n10987 ;
  assign n10999 = ~n10997 & n10998 ;
  assign n11000 = ~n10978 & n10999 ;
  assign n11001 = n6113 & ~n11000 ;
  assign n11003 = \P1_reg2_reg[23]/NET0131  & ~n8957 ;
  assign n11002 = n3279 & n4112 ;
  assign n11004 = n6207 & n10969 ;
  assign n11005 = ~n11002 & ~n11004 ;
  assign n11006 = ~n11003 & n11005 ;
  assign n11007 = ~n11001 & n11006 ;
  assign n11008 = ~n10977 & n11007 ;
  assign n11009 = n6097 & ~n11008 ;
  assign n11010 = ~n10968 & ~n11009 ;
  assign n11011 = \P1_state_reg[0]/NET0131  & ~n11010 ;
  assign n11012 = ~n10967 & ~n11011 ;
  assign n11013 = \P1_reg2_reg[30]/NET0131  & ~n6078 ;
  assign n11014 = \P1_reg2_reg[30]/NET0131  & n6095 ;
  assign n11015 = \P1_reg2_reg[30]/NET0131  & ~n6113 ;
  assign n11016 = n6113 & n10810 ;
  assign n11017 = ~n11015 & ~n11016 ;
  assign n11018 = n6359 & ~n11017 ;
  assign n11019 = n3500 & n6113 ;
  assign n11020 = ~n11015 & ~n11019 ;
  assign n11021 = n6365 & ~n11020 ;
  assign n11022 = ~n6361 & ~n10961 ;
  assign n11023 = \P1_reg2_reg[30]/NET0131  & ~n11022 ;
  assign n11024 = ~n6367 & ~n11023 ;
  assign n11025 = ~n11021 & n11024 ;
  assign n11026 = ~n8714 & n11025 ;
  assign n11027 = ~n11018 & n11026 ;
  assign n11028 = n6097 & ~n11027 ;
  assign n11029 = ~n11014 & ~n11028 ;
  assign n11030 = \P1_state_reg[0]/NET0131  & ~n11029 ;
  assign n11031 = ~n11013 & ~n11030 ;
  assign n11032 = \P2_reg2_reg[23]/NET0131  & n5585 ;
  assign n11033 = \P2_reg2_reg[23]/NET0131  & ~n4219 ;
  assign n11034 = n4219 & ~n10734 ;
  assign n11035 = ~n11033 & ~n11034 ;
  assign n11036 = n5526 & ~n11035 ;
  assign n11037 = n4219 & ~n10747 ;
  assign n11038 = ~n11033 & ~n11037 ;
  assign n11039 = n5329 & ~n11038 ;
  assign n11040 = n4656 & n5565 ;
  assign n11041 = n10762 & ~n11040 ;
  assign n11042 = n4219 & ~n11041 ;
  assign n11043 = n4661 & n5574 ;
  assign n11044 = \P2_reg2_reg[23]/NET0131  & ~n6841 ;
  assign n11045 = ~n11043 & ~n11044 ;
  assign n11046 = ~n11042 & n11045 ;
  assign n11047 = ~n11039 & n11046 ;
  assign n11048 = ~n11036 & n11047 ;
  assign n11049 = n5583 & ~n11048 ;
  assign n11050 = ~n11032 & ~n11049 ;
  assign n11051 = \P1_state_reg[0]/NET0131  & ~n11050 ;
  assign n11052 = \P2_reg2_reg[23]/NET0131  & ~n5589 ;
  assign n11053 = ~n11051 & ~n11052 ;
  assign n11054 = \P1_reg0_reg[12]/NET0131  & ~n6078 ;
  assign n11055 = \P1_reg0_reg[12]/NET0131  & n6095 ;
  assign n11056 = \P1_reg0_reg[12]/NET0131  & ~n9825 ;
  assign n11057 = n9083 & ~n10828 ;
  assign n11058 = n6409 & ~n11057 ;
  assign n11059 = ~n11056 & ~n11058 ;
  assign n11060 = n6097 & ~n11059 ;
  assign n11061 = ~n11055 & ~n11060 ;
  assign n11062 = \P1_state_reg[0]/NET0131  & ~n11061 ;
  assign n11063 = ~n11054 & ~n11062 ;
  assign n11064 = \P1_reg0_reg[16]/NET0131  & ~n6078 ;
  assign n11065 = \P1_reg0_reg[16]/NET0131  & n6095 ;
  assign n11067 = \P1_reg0_reg[16]/NET0131  & ~n6409 ;
  assign n11068 = n6409 & ~n9105 ;
  assign n11069 = ~n11067 & ~n11068 ;
  assign n11070 = n6207 & ~n11069 ;
  assign n11074 = n6409 & ~n9118 ;
  assign n11075 = ~n11067 & ~n11074 ;
  assign n11076 = n6282 & ~n11075 ;
  assign n11077 = n6409 & n9127 ;
  assign n11078 = ~n11067 & ~n11077 ;
  assign n11079 = n4011 & ~n11078 ;
  assign n11071 = n6409 & n9112 ;
  assign n11072 = ~n11067 & ~n11071 ;
  assign n11073 = n6359 & ~n11072 ;
  assign n11066 = \P1_reg0_reg[16]/NET0131  & ~n6425 ;
  assign n11080 = n6409 & n10847 ;
  assign n11081 = ~n11066 & ~n11080 ;
  assign n11082 = ~n11073 & n11081 ;
  assign n11083 = ~n11079 & n11082 ;
  assign n11084 = ~n11076 & n11083 ;
  assign n11085 = ~n11070 & n11084 ;
  assign n11086 = n6097 & ~n11085 ;
  assign n11087 = ~n11065 & ~n11086 ;
  assign n11088 = \P1_state_reg[0]/NET0131  & ~n11087 ;
  assign n11089 = ~n11064 & ~n11088 ;
  assign n11090 = \P1_reg0_reg[18]/NET0131  & ~n6078 ;
  assign n11091 = \P1_reg0_reg[18]/NET0131  & n6095 ;
  assign n11093 = \P1_reg0_reg[18]/NET0131  & ~n6409 ;
  assign n11094 = n6409 & ~n9193 ;
  assign n11095 = ~n11093 & ~n11094 ;
  assign n11096 = n6282 & ~n11095 ;
  assign n11100 = n6409 & n9199 ;
  assign n11101 = ~n11093 & ~n11100 ;
  assign n11102 = n6359 & ~n11101 ;
  assign n11097 = n6409 & n9205 ;
  assign n11098 = ~n11093 & ~n11097 ;
  assign n11099 = n6207 & ~n11098 ;
  assign n11103 = n6409 & n9214 ;
  assign n11104 = ~n11093 & ~n11103 ;
  assign n11105 = n4011 & ~n11104 ;
  assign n11092 = \P1_reg0_reg[18]/NET0131  & ~n6425 ;
  assign n11106 = n6409 & n10876 ;
  assign n11107 = ~n11092 & ~n11106 ;
  assign n11108 = ~n11105 & n11107 ;
  assign n11109 = ~n11099 & n11108 ;
  assign n11110 = ~n11102 & n11109 ;
  assign n11111 = ~n11096 & n11110 ;
  assign n11112 = n6097 & ~n11111 ;
  assign n11113 = ~n11091 & ~n11112 ;
  assign n11114 = \P1_state_reg[0]/NET0131  & ~n11113 ;
  assign n11115 = ~n11090 & ~n11114 ;
  assign n11116 = n9829 & ~n10955 ;
  assign n11120 = n6409 & n9237 ;
  assign n11121 = n6282 & ~n11120 ;
  assign n11117 = ~n6409 & n6693 ;
  assign n11118 = n6424 & ~n11117 ;
  assign n11119 = n9044 & n11118 ;
  assign n11122 = n6206 & ~n6409 ;
  assign n11123 = n11119 & ~n11122 ;
  assign n11124 = ~n11121 & n11123 ;
  assign n11125 = \P1_reg0_reg[19]/NET0131  & ~n11124 ;
  assign n11126 = ~n11116 & ~n11125 ;
  assign n11127 = \P1_reg0_reg[20]/NET0131  & ~n6078 ;
  assign n11128 = \P1_reg0_reg[20]/NET0131  & n6095 ;
  assign n11131 = \P1_reg0_reg[20]/NET0131  & ~n6409 ;
  assign n11135 = n6409 & n10704 ;
  assign n11136 = ~n11131 & ~n11135 ;
  assign n11137 = n4011 & ~n11136 ;
  assign n11132 = n6409 & ~n10696 ;
  assign n11133 = ~n11131 & ~n11132 ;
  assign n11134 = n6282 & ~n11133 ;
  assign n11138 = n6409 & ~n10710 ;
  assign n11139 = ~n11131 & ~n11138 ;
  assign n11140 = n6207 & ~n11139 ;
  assign n11129 = ~n10716 & ~n10905 ;
  assign n11130 = n6409 & ~n11129 ;
  assign n11141 = n6359 & ~n6409 ;
  assign n11142 = n6425 & ~n11141 ;
  assign n11143 = \P1_reg0_reg[20]/NET0131  & ~n11142 ;
  assign n11144 = ~n11130 & ~n11143 ;
  assign n11145 = ~n11140 & n11144 ;
  assign n11146 = ~n11134 & n11145 ;
  assign n11147 = ~n11137 & n11146 ;
  assign n11148 = n6097 & ~n11147 ;
  assign n11149 = ~n11128 & ~n11148 ;
  assign n11150 = \P1_state_reg[0]/NET0131  & ~n11149 ;
  assign n11151 = ~n11127 & ~n11150 ;
  assign n11152 = \P1_reg0_reg[21]/NET0131  & ~n6078 ;
  assign n11153 = \P1_reg0_reg[21]/NET0131  & n6095 ;
  assign n11155 = \P1_reg0_reg[21]/NET0131  & ~n6409 ;
  assign n11165 = n6409 & n9329 ;
  assign n11166 = ~n11155 & ~n11165 ;
  assign n11167 = n6359 & ~n11166 ;
  assign n11159 = n6409 & ~n9318 ;
  assign n11160 = ~n11155 & ~n11159 ;
  assign n11161 = n6282 & ~n11160 ;
  assign n11154 = \P1_reg0_reg[21]/NET0131  & ~n6425 ;
  assign n11168 = n6409 & n9346 ;
  assign n11169 = ~n11154 & ~n11168 ;
  assign n11170 = ~n11161 & n11169 ;
  assign n11171 = ~n11167 & n11170 ;
  assign n11156 = n6409 & n9312 ;
  assign n11157 = ~n11155 & ~n11156 ;
  assign n11158 = n4011 & ~n11157 ;
  assign n11162 = n6409 & ~n9324 ;
  assign n11163 = ~n11155 & ~n11162 ;
  assign n11164 = n6207 & ~n11163 ;
  assign n11172 = ~n11158 & ~n11164 ;
  assign n11173 = n11171 & n11172 ;
  assign n11174 = n6097 & ~n11173 ;
  assign n11175 = ~n11153 & ~n11174 ;
  assign n11176 = \P1_state_reg[0]/NET0131  & ~n11175 ;
  assign n11177 = ~n11152 & ~n11176 ;
  assign n11178 = \P1_reg0_reg[30]/NET0131  & ~n6078 ;
  assign n11179 = \P1_reg0_reg[30]/NET0131  & n6095 ;
  assign n11180 = \P1_reg0_reg[30]/NET0131  & ~n6409 ;
  assign n11185 = n6409 & n10810 ;
  assign n11186 = ~n11180 & ~n11185 ;
  assign n11187 = n6359 & ~n11186 ;
  assign n11181 = n3500 & n6409 ;
  assign n11182 = ~n11180 & ~n11181 ;
  assign n11183 = n6365 & ~n11182 ;
  assign n11184 = \P1_reg0_reg[30]/NET0131  & ~n10009 ;
  assign n11188 = ~n11183 & ~n11184 ;
  assign n11189 = ~n10017 & n11188 ;
  assign n11190 = ~n11187 & n11189 ;
  assign n11191 = n6097 & ~n11190 ;
  assign n11192 = ~n11179 & ~n11191 ;
  assign n11193 = \P1_state_reg[0]/NET0131  & ~n11192 ;
  assign n11194 = ~n11178 & ~n11193 ;
  assign n11195 = \P1_reg1_reg[12]/NET0131  & ~n6078 ;
  assign n11196 = \P1_reg1_reg[12]/NET0131  & n6095 ;
  assign n11197 = ~n6683 & ~n8656 ;
  assign n11198 = n7808 & ~n11197 ;
  assign n11199 = \P1_reg1_reg[12]/NET0131  & ~n11198 ;
  assign n11200 = n6683 & ~n11057 ;
  assign n11201 = ~n11199 & ~n11200 ;
  assign n11202 = n6097 & ~n11201 ;
  assign n11203 = ~n11196 & ~n11202 ;
  assign n11204 = \P1_state_reg[0]/NET0131  & ~n11203 ;
  assign n11205 = ~n11195 & ~n11204 ;
  assign n11206 = \P1_reg1_reg[16]/NET0131  & ~n6078 ;
  assign n11207 = \P1_reg1_reg[16]/NET0131  & n6095 ;
  assign n11209 = \P1_reg1_reg[16]/NET0131  & ~n6683 ;
  assign n11210 = n6683 & ~n9105 ;
  assign n11211 = ~n11209 & ~n11210 ;
  assign n11212 = n6207 & ~n11211 ;
  assign n11216 = n6683 & ~n9118 ;
  assign n11217 = ~n11209 & ~n11216 ;
  assign n11218 = n6282 & ~n11217 ;
  assign n11219 = n6683 & n9127 ;
  assign n11220 = ~n11209 & ~n11219 ;
  assign n11221 = n4011 & ~n11220 ;
  assign n11213 = n6683 & n9112 ;
  assign n11214 = ~n11209 & ~n11213 ;
  assign n11215 = n6359 & ~n11214 ;
  assign n11208 = \P1_reg1_reg[16]/NET0131  & ~n7806 ;
  assign n11222 = n6683 & n10847 ;
  assign n11223 = ~n11208 & ~n11222 ;
  assign n11224 = ~n11215 & n11223 ;
  assign n11225 = ~n11221 & n11224 ;
  assign n11226 = ~n11218 & n11225 ;
  assign n11227 = ~n11212 & n11226 ;
  assign n11228 = n6097 & ~n11227 ;
  assign n11229 = ~n11207 & ~n11228 ;
  assign n11230 = \P1_state_reg[0]/NET0131  & ~n11229 ;
  assign n11231 = ~n11206 & ~n11230 ;
  assign n11232 = \P1_reg1_reg[18]/NET0131  & ~n6078 ;
  assign n11233 = \P1_reg1_reg[18]/NET0131  & n6095 ;
  assign n11235 = \P1_reg1_reg[18]/NET0131  & ~n6683 ;
  assign n11236 = n6683 & ~n9193 ;
  assign n11237 = ~n11235 & ~n11236 ;
  assign n11238 = n6282 & ~n11237 ;
  assign n11242 = n6683 & n9205 ;
  assign n11243 = ~n11235 & ~n11242 ;
  assign n11244 = n6207 & ~n11243 ;
  assign n11239 = n6683 & n9199 ;
  assign n11240 = ~n11235 & ~n11239 ;
  assign n11241 = n6359 & ~n11240 ;
  assign n11245 = n6683 & n9214 ;
  assign n11246 = ~n11235 & ~n11245 ;
  assign n11247 = n4011 & ~n11246 ;
  assign n11234 = \P1_reg1_reg[18]/NET0131  & ~n7806 ;
  assign n11248 = n6683 & n10876 ;
  assign n11249 = ~n11234 & ~n11248 ;
  assign n11250 = ~n11247 & n11249 ;
  assign n11251 = ~n11241 & n11250 ;
  assign n11252 = ~n11244 & n11251 ;
  assign n11253 = ~n11238 & n11252 ;
  assign n11254 = n6097 & ~n11253 ;
  assign n11255 = ~n11233 & ~n11254 ;
  assign n11256 = \P1_state_reg[0]/NET0131  & ~n11255 ;
  assign n11257 = ~n11232 & ~n11256 ;
  assign n11258 = n6696 & n9044 ;
  assign n11259 = ~n11197 & n11258 ;
  assign n11260 = \P1_reg1_reg[19]/NET0131  & ~n11259 ;
  assign n11261 = n9045 & ~n10955 ;
  assign n11262 = ~n11260 & ~n11261 ;
  assign n11263 = \P1_reg1_reg[20]/NET0131  & ~n6078 ;
  assign n11264 = \P1_reg1_reg[20]/NET0131  & n6095 ;
  assign n11266 = \P1_reg1_reg[20]/NET0131  & ~n6683 ;
  assign n11270 = n6683 & n10704 ;
  assign n11271 = ~n11266 & ~n11270 ;
  assign n11272 = n4011 & ~n11271 ;
  assign n11267 = n6683 & ~n10696 ;
  assign n11268 = ~n11266 & ~n11267 ;
  assign n11269 = n6282 & ~n11268 ;
  assign n11273 = n6683 & ~n10710 ;
  assign n11274 = ~n11266 & ~n11273 ;
  assign n11275 = n6207 & ~n11274 ;
  assign n11265 = n6683 & ~n11129 ;
  assign n11276 = \P1_reg1_reg[20]/NET0131  & ~n7807 ;
  assign n11277 = ~n11265 & ~n11276 ;
  assign n11278 = ~n11275 & n11277 ;
  assign n11279 = ~n11269 & n11278 ;
  assign n11280 = ~n11272 & n11279 ;
  assign n11281 = n6097 & ~n11280 ;
  assign n11282 = ~n11264 & ~n11281 ;
  assign n11283 = \P1_state_reg[0]/NET0131  & ~n11282 ;
  assign n11284 = ~n11263 & ~n11283 ;
  assign n11286 = n3250 & n6095 ;
  assign n11288 = ~n3255 & n9064 ;
  assign n11289 = n3650 & ~n11288 ;
  assign n11290 = ~n9065 & ~n11289 ;
  assign n11291 = ~n2713 & ~n11290 ;
  assign n11292 = n2713 & n3677 ;
  assign n11293 = ~n11291 & ~n11292 ;
  assign n11294 = n6568 & ~n11293 ;
  assign n11295 = ~n3250 & ~n6568 ;
  assign n11296 = n4011 & ~n11295 ;
  assign n11297 = ~n11294 & n11296 ;
  assign n11307 = ~n3258 & ~n6579 ;
  assign n11306 = n3258 & n6579 ;
  assign n11308 = n6282 & ~n11306 ;
  assign n11309 = ~n11307 & n11308 ;
  assign n11298 = ~n3668 & n6336 ;
  assign n11299 = n3246 & ~n11298 ;
  assign n11300 = ~n6338 & n6359 ;
  assign n11301 = ~n11299 & n11300 ;
  assign n11303 = ~n3258 & n6617 ;
  assign n11302 = n3258 & ~n6617 ;
  assign n11304 = n6207 & ~n11302 ;
  assign n11305 = ~n11303 & n11304 ;
  assign n11310 = ~n11301 & ~n11305 ;
  assign n11311 = ~n11309 & n11310 ;
  assign n11312 = n6568 & ~n11311 ;
  assign n11287 = n3246 & ~n6649 ;
  assign n11313 = ~n6568 & ~n8656 ;
  assign n11314 = n7036 & ~n11313 ;
  assign n11315 = n3250 & ~n11314 ;
  assign n11316 = ~n11287 & ~n11315 ;
  assign n11317 = ~n11312 & n11316 ;
  assign n11318 = ~n11297 & n11317 ;
  assign n11319 = n6097 & ~n11318 ;
  assign n11320 = ~n11286 & ~n11319 ;
  assign n11321 = \P1_state_reg[0]/NET0131  & ~n11320 ;
  assign n11285 = n3250 & n4130 ;
  assign n11322 = \P1_reg3_reg[11]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11323 = ~n11285 & ~n11322 ;
  assign n11324 = ~n11321 & n11323 ;
  assign n11327 = n4926 & n5585 ;
  assign n11329 = n4926 & ~n7453 ;
  assign n11336 = n4958 & ~n5357 ;
  assign n11337 = ~n10379 & ~n11336 ;
  assign n11338 = ~n4231 & ~n11337 ;
  assign n11339 = n4231 & n4984 ;
  assign n11340 = ~n11338 & ~n11339 ;
  assign n11341 = n7453 & n11340 ;
  assign n11342 = ~n11329 & ~n11341 ;
  assign n11343 = n5383 & ~n11342 ;
  assign n11330 = n5991 & ~n7558 ;
  assign n11331 = ~n5991 & n7558 ;
  assign n11332 = ~n11330 & ~n11331 ;
  assign n11333 = n7453 & n11332 ;
  assign n11334 = ~n11329 & ~n11333 ;
  assign n11335 = n5329 & ~n11334 ;
  assign n11344 = n5991 & ~n7525 ;
  assign n11345 = ~n5991 & n7525 ;
  assign n11346 = ~n11344 & ~n11345 ;
  assign n11347 = n7453 & ~n11346 ;
  assign n11348 = ~n11329 & ~n11347 ;
  assign n11349 = n5526 & ~n11348 ;
  assign n11350 = n4948 & ~n5538 ;
  assign n11351 = ~n10395 & ~n11350 ;
  assign n11352 = n7453 & n11351 ;
  assign n11353 = ~n11329 & ~n11352 ;
  assign n11354 = n5563 & ~n11353 ;
  assign n11328 = n4948 & ~n7504 ;
  assign n11355 = n4926 & ~n7641 ;
  assign n11356 = ~n11328 & ~n11355 ;
  assign n11357 = ~n11354 & n11356 ;
  assign n11358 = ~n11349 & n11357 ;
  assign n11359 = ~n11335 & n11358 ;
  assign n11360 = ~n11343 & n11359 ;
  assign n11361 = n5583 & ~n11360 ;
  assign n11362 = ~n11327 & ~n11361 ;
  assign n11363 = \P1_state_reg[0]/NET0131  & ~n11362 ;
  assign n11325 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[11]/NET0131  ;
  assign n11326 = n4926 & n5786 ;
  assign n11364 = ~n11325 & ~n11326 ;
  assign n11365 = ~n11363 & n11364 ;
  assign n11368 = n3618 & n6095 ;
  assign n11372 = n3618 & n6427 ;
  assign n11373 = ~n6568 & ~n11372 ;
  assign n11383 = n2713 & ~n3229 ;
  assign n11384 = ~n3229 & n9067 ;
  assign n11385 = ~n3623 & n11384 ;
  assign n11386 = n3203 & ~n11385 ;
  assign n11387 = ~n2713 & ~n6301 ;
  assign n11388 = ~n11386 & n11387 ;
  assign n11389 = ~n11383 & ~n11388 ;
  assign n11390 = n4011 & ~n11389 ;
  assign n11375 = n3626 & n6584 ;
  assign n11374 = ~n3626 & ~n6584 ;
  assign n11376 = n6282 & ~n11374 ;
  assign n11377 = ~n11375 & n11376 ;
  assign n11379 = ~n3626 & n10988 ;
  assign n11378 = n3626 & ~n10988 ;
  assign n11380 = n6207 & ~n11378 ;
  assign n11381 = ~n11379 & n11380 ;
  assign n11382 = ~n11377 & ~n11381 ;
  assign n11391 = n3614 & ~n6341 ;
  assign n11392 = n6359 & ~n9109 ;
  assign n11393 = ~n11391 & n11392 ;
  assign n11394 = n6568 & ~n11393 ;
  assign n11395 = n11382 & n11394 ;
  assign n11396 = ~n11390 & n11395 ;
  assign n11397 = ~n11373 & ~n11396 ;
  assign n11369 = n3614 & ~n6649 ;
  assign n11370 = n6666 & ~n11313 ;
  assign n11371 = n3618 & ~n11370 ;
  assign n11398 = ~n11369 & ~n11371 ;
  assign n11399 = ~n11397 & n11398 ;
  assign n11400 = n6097 & ~n11399 ;
  assign n11401 = ~n11368 & ~n11400 ;
  assign n11402 = \P1_state_reg[0]/NET0131  & ~n11401 ;
  assign n11366 = \P1_reg3_reg[15]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11367 = n3618 & n4130 ;
  assign n11403 = ~n11366 & ~n11367 ;
  assign n11404 = ~n11402 & n11403 ;
  assign n11407 = n4821 & n5585 ;
  assign n11408 = n4821 & ~n7453 ;
  assign n11415 = n4902 & ~n10418 ;
  assign n11416 = ~n5361 & ~n11415 ;
  assign n11417 = ~n4231 & ~n11416 ;
  assign n11418 = n4231 & n4854 ;
  assign n11419 = ~n11417 & ~n11418 ;
  assign n11420 = n7453 & n11419 ;
  assign n11421 = ~n11408 & ~n11420 ;
  assign n11422 = n5383 & ~n11421 ;
  assign n11424 = ~n4843 & n10424 ;
  assign n11423 = n4843 & ~n10424 ;
  assign n11425 = n5563 & ~n11423 ;
  assign n11426 = ~n11424 & n11425 ;
  assign n11428 = n5999 & ~n8733 ;
  assign n11427 = ~n5999 & n8733 ;
  assign n11429 = n5329 & ~n11427 ;
  assign n11430 = ~n11428 & n11429 ;
  assign n11431 = ~n11426 & ~n11430 ;
  assign n11432 = n7453 & ~n11431 ;
  assign n11409 = n5999 & ~n8744 ;
  assign n11410 = ~n5999 & n8744 ;
  assign n11411 = ~n11409 & ~n11410 ;
  assign n11412 = n7453 & ~n11411 ;
  assign n11413 = ~n11408 & ~n11412 ;
  assign n11414 = n5526 & ~n11413 ;
  assign n11433 = n4843 & ~n7504 ;
  assign n11434 = n5329 & ~n7453 ;
  assign n11435 = n7484 & ~n11434 ;
  assign n11436 = n4821 & ~n11435 ;
  assign n11437 = ~n11433 & ~n11436 ;
  assign n11438 = ~n11414 & n11437 ;
  assign n11439 = ~n11432 & n11438 ;
  assign n11440 = ~n11422 & n11439 ;
  assign n11441 = n5583 & ~n11440 ;
  assign n11442 = ~n11407 & ~n11441 ;
  assign n11443 = \P1_state_reg[0]/NET0131  & ~n11442 ;
  assign n11405 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[14]/NET0131  ;
  assign n11406 = n4821 & n5786 ;
  assign n11444 = ~n11405 & ~n11406 ;
  assign n11445 = ~n11443 & n11444 ;
  assign n11448 = n4898 & n5585 ;
  assign n11450 = n4898 & ~n7453 ;
  assign n11451 = n5988 & ~n10739 ;
  assign n11452 = ~n5988 & n10739 ;
  assign n11453 = ~n11451 & ~n11452 ;
  assign n11454 = n7453 & n11453 ;
  assign n11455 = ~n11450 & ~n11454 ;
  assign n11456 = n5329 & ~n11455 ;
  assign n11463 = ~n4879 & n5361 ;
  assign n11464 = n4879 & ~n5361 ;
  assign n11465 = ~n11463 & ~n11464 ;
  assign n11466 = ~n4231 & ~n11465 ;
  assign n11467 = n4231 & n4827 ;
  assign n11468 = ~n11466 & ~n11467 ;
  assign n11469 = n7453 & n11468 ;
  assign n11470 = ~n11450 & ~n11469 ;
  assign n11471 = n5383 & ~n11470 ;
  assign n11457 = n5988 & ~n7530 ;
  assign n11458 = ~n5988 & n7530 ;
  assign n11459 = ~n11457 & ~n11458 ;
  assign n11460 = n7453 & ~n11459 ;
  assign n11461 = ~n11450 & ~n11460 ;
  assign n11462 = n5526 & ~n11461 ;
  assign n11472 = n4918 & ~n11424 ;
  assign n11473 = n5541 & n10424 ;
  assign n11474 = ~n11472 & ~n11473 ;
  assign n11475 = n7453 & n11474 ;
  assign n11476 = ~n11450 & ~n11475 ;
  assign n11477 = n5563 & ~n11476 ;
  assign n11449 = n4918 & ~n7504 ;
  assign n11478 = n4898 & ~n7641 ;
  assign n11479 = ~n11449 & ~n11478 ;
  assign n11480 = ~n11477 & n11479 ;
  assign n11481 = ~n11462 & n11480 ;
  assign n11482 = ~n11471 & n11481 ;
  assign n11483 = ~n11456 & n11482 ;
  assign n11484 = n5583 & ~n11483 ;
  assign n11485 = ~n11448 & ~n11484 ;
  assign n11486 = \P1_state_reg[0]/NET0131  & ~n11485 ;
  assign n11446 = n4898 & n5786 ;
  assign n11447 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[15]/NET0131  ;
  assign n11487 = ~n11446 & ~n11447 ;
  assign n11488 = ~n11486 & n11487 ;
  assign n11490 = n4875 & n5585 ;
  assign n11492 = n4875 & ~n7453 ;
  assign n11493 = ~n6755 & n6758 ;
  assign n11494 = n6769 & ~n11493 ;
  assign n11495 = n5997 & n11494 ;
  assign n11496 = ~n5997 & ~n11494 ;
  assign n11497 = ~n11495 & ~n11496 ;
  assign n11498 = n7453 & ~n11497 ;
  assign n11499 = ~n11492 & ~n11498 ;
  assign n11500 = n5329 & ~n11499 ;
  assign n11501 = n4774 & ~n11463 ;
  assign n11502 = ~n8478 & ~n11501 ;
  assign n11503 = ~n4231 & ~n11502 ;
  assign n11504 = n4231 & n4902 ;
  assign n11505 = ~n11503 & ~n11504 ;
  assign n11506 = n7453 & n11505 ;
  assign n11507 = ~n11492 & ~n11506 ;
  assign n11508 = n5383 & ~n11507 ;
  assign n11509 = ~n5829 & n5997 ;
  assign n11510 = n5829 & ~n5997 ;
  assign n11511 = ~n11509 & ~n11510 ;
  assign n11512 = n7453 & ~n11511 ;
  assign n11513 = ~n11492 & ~n11512 ;
  assign n11514 = n5526 & ~n11513 ;
  assign n11515 = n4892 & ~n11473 ;
  assign n11516 = ~n5544 & ~n11515 ;
  assign n11517 = n7453 & n11516 ;
  assign n11518 = ~n11492 & ~n11517 ;
  assign n11519 = n5563 & ~n11518 ;
  assign n11491 = n4892 & ~n7504 ;
  assign n11520 = n4875 & ~n7641 ;
  assign n11521 = ~n11491 & ~n11520 ;
  assign n11522 = ~n11519 & n11521 ;
  assign n11523 = ~n11514 & n11522 ;
  assign n11524 = ~n11508 & n11523 ;
  assign n11525 = ~n11500 & n11524 ;
  assign n11526 = n5583 & ~n11525 ;
  assign n11527 = ~n11490 & ~n11526 ;
  assign n11528 = \P1_state_reg[0]/NET0131  & ~n11527 ;
  assign n11489 = n4875 & n5786 ;
  assign n11529 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[16]/NET0131  ;
  assign n11530 = ~n11489 & ~n11529 ;
  assign n11531 = ~n11528 & n11530 ;
  assign n11533 = n3818 & n6095 ;
  assign n11535 = n3818 & ~n6568 ;
  assign n11536 = n3329 & ~n6293 ;
  assign n11537 = ~n9063 & ~n11536 ;
  assign n11538 = ~n2713 & ~n11537 ;
  assign n11539 = n2713 & n3577 ;
  assign n11540 = ~n11538 & ~n11539 ;
  assign n11541 = n6568 & n11540 ;
  assign n11542 = ~n11535 & ~n11541 ;
  assign n11543 = n4011 & ~n11542 ;
  assign n11544 = n3825 & ~n6998 ;
  assign n11545 = ~n3825 & n6998 ;
  assign n11546 = ~n11544 & ~n11545 ;
  assign n11547 = n6568 & n11546 ;
  assign n11548 = ~n11535 & ~n11547 ;
  assign n11549 = n6207 & ~n11548 ;
  assign n11550 = n3825 & ~n4052 ;
  assign n11551 = ~n3825 & n4052 ;
  assign n11552 = ~n11550 & ~n11551 ;
  assign n11553 = n6568 & ~n11552 ;
  assign n11554 = ~n11535 & ~n11553 ;
  assign n11555 = n6282 & ~n11554 ;
  assign n11556 = n3813 & ~n6334 ;
  assign n11557 = ~n6335 & ~n11556 ;
  assign n11558 = n6568 & n11557 ;
  assign n11559 = ~n11535 & ~n11558 ;
  assign n11560 = n6359 & ~n11559 ;
  assign n11534 = n3813 & ~n6649 ;
  assign n11561 = n3818 & ~n6666 ;
  assign n11562 = ~n11534 & ~n11561 ;
  assign n11563 = ~n11560 & n11562 ;
  assign n11564 = ~n11555 & n11563 ;
  assign n11565 = ~n11549 & n11564 ;
  assign n11566 = ~n11543 & n11565 ;
  assign n11567 = n6097 & ~n11566 ;
  assign n11568 = ~n11533 & ~n11567 ;
  assign n11569 = \P1_state_reg[0]/NET0131  & ~n11568 ;
  assign n11532 = \P1_reg3_reg[8]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11570 = n3818 & n4130 ;
  assign n11571 = ~n11532 & ~n11570 ;
  assign n11572 = ~n11569 & n11571 ;
  assign n11575 = ~n1514 & n2145 ;
  assign n11584 = ~n1514 & ~n2163 ;
  assign n11588 = n1197 & ~n9149 ;
  assign n11589 = ~n2239 & ~n9150 ;
  assign n11590 = ~n11588 & n11589 ;
  assign n11591 = ~n1531 & n2239 ;
  assign n11592 = ~n11590 & ~n11591 ;
  assign n11593 = n2163 & ~n11592 ;
  assign n11594 = ~n11584 & ~n11593 ;
  assign n11595 = n737 & ~n11594 ;
  assign n11578 = n2036 & ~n2544 ;
  assign n11579 = ~n2036 & n2544 ;
  assign n11580 = ~n11578 & ~n11579 ;
  assign n11585 = n2163 & ~n11580 ;
  assign n11586 = ~n11584 & ~n11585 ;
  assign n11587 = n2393 & ~n11586 ;
  assign n11577 = ~n1514 & ~n2236 ;
  assign n11581 = n2236 & ~n11580 ;
  assign n11582 = ~n11577 & ~n11581 ;
  assign n11583 = n2391 & ~n11582 ;
  assign n11596 = n2036 & ~n2598 ;
  assign n11597 = ~n2036 & n2598 ;
  assign n11598 = ~n11596 & ~n11597 ;
  assign n11599 = n2236 & n11598 ;
  assign n11600 = ~n11577 & ~n11599 ;
  assign n11601 = n2234 & ~n11600 ;
  assign n11576 = ~n1512 & n2580 ;
  assign n11602 = ~n1514 & ~n2583 ;
  assign n11603 = ~n11576 & ~n11602 ;
  assign n11604 = ~n11601 & n11603 ;
  assign n11605 = ~n11583 & n11604 ;
  assign n11606 = ~n11587 & n11605 ;
  assign n11607 = ~n11595 & n11606 ;
  assign n11608 = n2147 & ~n11607 ;
  assign n11609 = ~n11575 & ~n11608 ;
  assign n11610 = \P1_state_reg[0]/NET0131  & ~n11609 ;
  assign n11573 = n765 & ~n1514 ;
  assign n11574 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[15]/NET0131  ;
  assign n11611 = ~n11573 & ~n11574 ;
  assign n11612 = ~n11610 & n11611 ;
  assign n11615 = ~n1681 & n2145 ;
  assign n11618 = ~n1681 & ~n2163 ;
  assign n11619 = n2064 & ~n2464 ;
  assign n11620 = ~n2064 & n2464 ;
  assign n11621 = ~n11619 & ~n11620 ;
  assign n11622 = n2163 & n11621 ;
  assign n11623 = ~n11618 & ~n11622 ;
  assign n11624 = n2393 & ~n11623 ;
  assign n11616 = ~n1704 & n2580 ;
  assign n11617 = ~n1681 & ~n2583 ;
  assign n11643 = ~n11616 & ~n11617 ;
  assign n11644 = ~n11624 & n11643 ;
  assign n11635 = n1663 & ~n2251 ;
  assign n11636 = ~n2239 & ~n10306 ;
  assign n11637 = ~n11635 & n11636 ;
  assign n11638 = ~n1729 & n2239 ;
  assign n11639 = ~n11637 & ~n11638 ;
  assign n11640 = n2163 & ~n11639 ;
  assign n11641 = ~n11618 & ~n11640 ;
  assign n11642 = n737 & ~n11641 ;
  assign n11625 = ~n1681 & ~n2236 ;
  assign n11626 = ~n1979 & n2064 ;
  assign n11627 = n1979 & ~n2064 ;
  assign n11628 = ~n11626 & ~n11627 ;
  assign n11629 = n2236 & ~n11628 ;
  assign n11630 = ~n11625 & ~n11629 ;
  assign n11631 = n2234 & ~n11630 ;
  assign n11632 = n2236 & n11621 ;
  assign n11633 = ~n11625 & ~n11632 ;
  assign n11634 = n2391 & ~n11633 ;
  assign n11645 = ~n11631 & ~n11634 ;
  assign n11646 = ~n11642 & n11645 ;
  assign n11647 = n11644 & n11646 ;
  assign n11648 = n2147 & ~n11647 ;
  assign n11649 = ~n11615 & ~n11648 ;
  assign n11650 = \P1_state_reg[0]/NET0131  & ~n11649 ;
  assign n11613 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[8]/NET0131  ;
  assign n11614 = n765 & ~n1681 ;
  assign n11651 = ~n11613 & ~n11614 ;
  assign n11652 = ~n11650 & n11651 ;
  assign n11653 = \P1_reg3_reg[10]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11656 = n3672 & ~n6568 ;
  assign n11657 = n3255 & ~n9064 ;
  assign n11658 = ~n11288 & ~n11657 ;
  assign n11659 = ~n2713 & ~n11658 ;
  assign n11660 = n2713 & n3329 ;
  assign n11661 = ~n11659 & ~n11660 ;
  assign n11662 = n6568 & n11661 ;
  assign n11663 = ~n11656 & ~n11662 ;
  assign n11664 = n4011 & ~n11663 ;
  assign n11671 = n3680 & ~n7132 ;
  assign n11672 = ~n3680 & n7132 ;
  assign n11673 = ~n11671 & ~n11672 ;
  assign n11674 = n6568 & ~n11673 ;
  assign n11675 = ~n11656 & ~n11674 ;
  assign n11676 = n6282 & ~n11675 ;
  assign n11665 = n3680 & ~n7174 ;
  assign n11666 = ~n3680 & n7174 ;
  assign n11667 = ~n11665 & ~n11666 ;
  assign n11668 = n6568 & n11667 ;
  assign n11669 = ~n11656 & ~n11668 ;
  assign n11670 = n6207 & ~n11669 ;
  assign n11677 = n3668 & ~n6336 ;
  assign n11678 = ~n11298 & ~n11677 ;
  assign n11679 = n6568 & n11678 ;
  assign n11680 = ~n11656 & ~n11679 ;
  assign n11681 = n6359 & ~n11680 ;
  assign n11682 = n3668 & ~n6649 ;
  assign n11655 = n3672 & ~n6666 ;
  assign n11683 = n6097 & ~n11655 ;
  assign n11684 = ~n11682 & n11683 ;
  assign n11685 = ~n11681 & n11684 ;
  assign n11686 = ~n11670 & n11685 ;
  assign n11687 = ~n11676 & n11686 ;
  assign n11688 = ~n11664 & n11687 ;
  assign n11654 = ~n3672 & ~n6097 ;
  assign n11689 = \P1_state_reg[0]/NET0131  & ~n11654 ;
  assign n11690 = ~n11688 & n11689 ;
  assign n11691 = ~n11653 & ~n11690 ;
  assign n11692 = \P1_reg3_reg[13]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11710 = ~n3357 & n6161 ;
  assign n11709 = n3357 & ~n6161 ;
  assign n11711 = n6207 & ~n11709 ;
  assign n11712 = ~n11710 & n11711 ;
  assign n11706 = ~n3357 & ~n6235 ;
  assign n11705 = n3357 & n6235 ;
  assign n11707 = n6282 & ~n11705 ;
  assign n11708 = ~n11706 & n11707 ;
  assign n11695 = n3229 & ~n9067 ;
  assign n11696 = ~n11384 & ~n11695 ;
  assign n11697 = ~n2713 & ~n11696 ;
  assign n11698 = n2713 & n3650 ;
  assign n11699 = n4011 & ~n11698 ;
  assign n11700 = ~n11697 & n11699 ;
  assign n11702 = n3345 & ~n9059 ;
  assign n11701 = ~n3345 & n9059 ;
  assign n11703 = n6359 & ~n11701 ;
  assign n11704 = ~n11702 & n11703 ;
  assign n11713 = ~n11700 & ~n11704 ;
  assign n11714 = ~n11708 & n11713 ;
  assign n11715 = ~n11712 & n11714 ;
  assign n11716 = n6568 & ~n11715 ;
  assign n11717 = n6668 & ~n11313 ;
  assign n11718 = n3349 & ~n11717 ;
  assign n11694 = n3345 & ~n6649 ;
  assign n11719 = n6097 & ~n11694 ;
  assign n11720 = ~n11718 & n11719 ;
  assign n11721 = ~n11716 & n11720 ;
  assign n11693 = ~n3349 & ~n6097 ;
  assign n11722 = \P1_state_reg[0]/NET0131  & ~n11693 ;
  assign n11723 = ~n11721 & n11722 ;
  assign n11724 = ~n11692 & ~n11723 ;
  assign n11725 = \P1_reg3_reg[9]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11728 = n3324 & ~n6568 ;
  assign n11729 = n3677 & ~n9063 ;
  assign n11730 = ~n9064 & ~n11729 ;
  assign n11731 = ~n2713 & ~n11730 ;
  assign n11732 = n2713 & n3822 ;
  assign n11733 = ~n11731 & ~n11732 ;
  assign n11734 = n6568 & n11733 ;
  assign n11735 = ~n11728 & ~n11734 ;
  assign n11736 = n4011 & ~n11735 ;
  assign n11743 = n3332 & ~n7067 ;
  assign n11744 = ~n3332 & n7067 ;
  assign n11745 = ~n11743 & ~n11744 ;
  assign n11746 = n6568 & ~n11745 ;
  assign n11747 = ~n11728 & ~n11746 ;
  assign n11748 = n6282 & ~n11747 ;
  assign n11737 = n3332 & ~n6157 ;
  assign n11738 = ~n3332 & n6157 ;
  assign n11739 = ~n11737 & ~n11738 ;
  assign n11740 = n6568 & n11739 ;
  assign n11741 = ~n11728 & ~n11740 ;
  assign n11742 = n6207 & ~n11741 ;
  assign n11749 = n3320 & ~n6335 ;
  assign n11750 = ~n6336 & ~n11749 ;
  assign n11751 = n6568 & n11750 ;
  assign n11752 = ~n11728 & ~n11751 ;
  assign n11753 = n6359 & ~n11752 ;
  assign n11754 = n3320 & n6568 ;
  assign n11755 = ~n11728 & ~n11754 ;
  assign n11756 = n6365 & ~n11755 ;
  assign n11727 = n3320 & n4112 ;
  assign n11757 = n3324 & n6361 ;
  assign n11758 = n6097 & ~n11757 ;
  assign n11759 = ~n11727 & n11758 ;
  assign n11760 = ~n11756 & n11759 ;
  assign n11761 = ~n11753 & n11760 ;
  assign n11762 = ~n11742 & n11761 ;
  assign n11763 = ~n11748 & n11762 ;
  assign n11764 = ~n11736 & n11763 ;
  assign n11726 = ~n3324 & ~n6097 ;
  assign n11765 = \P1_state_reg[0]/NET0131  & ~n11726 ;
  assign n11766 = ~n11764 & n11765 ;
  assign n11767 = ~n11725 & ~n11766 ;
  assign n11768 = n3279 & n6095 ;
  assign n11774 = n6568 & n10974 ;
  assign n11775 = ~n3279 & ~n6568 ;
  assign n11776 = n6282 & ~n11775 ;
  assign n11777 = ~n11774 & n11776 ;
  assign n11770 = n6568 & ~n10999 ;
  assign n11769 = n3273 & ~n6649 ;
  assign n11771 = n6207 & ~n6568 ;
  assign n11772 = n6668 & ~n11771 ;
  assign n11773 = n3279 & ~n11772 ;
  assign n11778 = ~n11769 & ~n11773 ;
  assign n11779 = ~n11770 & n11778 ;
  assign n11780 = ~n11777 & n11779 ;
  assign n11781 = n6097 & ~n11780 ;
  assign n11782 = ~n11768 & ~n11781 ;
  assign n11783 = \P1_state_reg[0]/NET0131  & ~n11782 ;
  assign n11784 = \P1_reg3_reg[23]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11785 = n3279 & n4130 ;
  assign n11786 = ~n11784 & ~n11785 ;
  assign n11787 = ~n11783 & n11786 ;
  assign n11788 = \P1_reg2_reg[10]/NET0131  & ~n6078 ;
  assign n11789 = \P1_reg2_reg[10]/NET0131  & n6095 ;
  assign n11792 = \P1_reg2_reg[10]/NET0131  & ~n6113 ;
  assign n11799 = n6113 & n11661 ;
  assign n11800 = ~n11792 & ~n11799 ;
  assign n11801 = n4011 & ~n11800 ;
  assign n11796 = n6113 & ~n11673 ;
  assign n11797 = ~n11792 & ~n11796 ;
  assign n11798 = n6282 & ~n11797 ;
  assign n11793 = n6113 & n11667 ;
  assign n11794 = ~n11792 & ~n11793 ;
  assign n11795 = n6207 & ~n11794 ;
  assign n11802 = n6113 & n11678 ;
  assign n11803 = ~n11792 & ~n11802 ;
  assign n11804 = n6359 & ~n11803 ;
  assign n11806 = \P1_reg2_reg[10]/NET0131  & ~n8955 ;
  assign n11790 = n3668 & n6365 ;
  assign n11791 = n6113 & n11790 ;
  assign n11805 = n3672 & n4112 ;
  assign n11807 = ~n11791 & ~n11805 ;
  assign n11808 = ~n11806 & n11807 ;
  assign n11809 = ~n11804 & n11808 ;
  assign n11810 = ~n11795 & n11809 ;
  assign n11811 = ~n11798 & n11810 ;
  assign n11812 = ~n11801 & n11811 ;
  assign n11813 = n6097 & ~n11812 ;
  assign n11814 = ~n11789 & ~n11813 ;
  assign n11815 = \P1_state_reg[0]/NET0131  & ~n11814 ;
  assign n11816 = ~n11788 & ~n11815 ;
  assign n11817 = \P1_reg2_reg[9]/NET0131  & ~n6078 ;
  assign n11818 = \P1_reg2_reg[9]/NET0131  & n6095 ;
  assign n11823 = \P1_reg2_reg[9]/NET0131  & ~n6113 ;
  assign n11824 = n6113 & n11733 ;
  assign n11825 = ~n11823 & ~n11824 ;
  assign n11826 = n4011 & ~n11825 ;
  assign n11830 = n6113 & n11739 ;
  assign n11831 = ~n11823 & ~n11830 ;
  assign n11832 = n6207 & ~n11831 ;
  assign n11827 = n6113 & ~n11745 ;
  assign n11828 = ~n11823 & ~n11827 ;
  assign n11829 = n6282 & ~n11828 ;
  assign n11819 = n3320 & n6365 ;
  assign n11820 = n6359 & n11750 ;
  assign n11821 = ~n11819 & ~n11820 ;
  assign n11822 = n6113 & ~n11821 ;
  assign n11833 = n3324 & n4112 ;
  assign n11834 = ~n6361 & ~n10962 ;
  assign n11835 = \P1_reg2_reg[9]/NET0131  & ~n11834 ;
  assign n11836 = ~n11833 & ~n11835 ;
  assign n11837 = ~n11822 & n11836 ;
  assign n11838 = ~n11829 & n11837 ;
  assign n11839 = ~n11832 & n11838 ;
  assign n11840 = ~n11826 & n11839 ;
  assign n11841 = n6097 & ~n11840 ;
  assign n11842 = ~n11818 & ~n11841 ;
  assign n11843 = \P1_state_reg[0]/NET0131  & ~n11842 ;
  assign n11844 = ~n11817 & ~n11843 ;
  assign n11845 = \P1_reg1_reg[23]/NET0131  & ~n11259 ;
  assign n11846 = n6282 & ~n10974 ;
  assign n11847 = n11000 & ~n11846 ;
  assign n11848 = n9045 & ~n11847 ;
  assign n11849 = ~n11845 & ~n11848 ;
  assign n11850 = \P2_reg0_reg[23]/NET0131  & ~n6706 ;
  assign n11851 = n6706 & ~n10734 ;
  assign n11852 = ~n11850 & ~n11851 ;
  assign n11853 = n5526 & ~n11852 ;
  assign n11854 = n6706 & ~n10747 ;
  assign n11855 = ~n11850 & ~n11854 ;
  assign n11856 = n5329 & ~n11855 ;
  assign n11857 = n6706 & ~n11041 ;
  assign n11858 = \P2_reg0_reg[23]/NET0131  & ~n7985 ;
  assign n11859 = ~n11857 & ~n11858 ;
  assign n11860 = ~n11856 & n11859 ;
  assign n11861 = ~n11853 & n11860 ;
  assign n11862 = n5583 & ~n11861 ;
  assign n11863 = \P2_reg0_reg[23]/NET0131  & n5585 ;
  assign n11864 = ~n11862 & ~n11863 ;
  assign n11865 = \P1_state_reg[0]/NET0131  & ~n11864 ;
  assign n11866 = \P2_reg0_reg[23]/NET0131  & ~n5589 ;
  assign n11867 = ~n11865 & ~n11866 ;
  assign n11868 = \P2_reg0_reg[30]/NET0131  & ~n6706 ;
  assign n11869 = ~n5557 & n5895 ;
  assign n11870 = ~n8814 & ~n11869 ;
  assign n11871 = n9533 & n11870 ;
  assign n11872 = ~n11868 & ~n11871 ;
  assign n11873 = n5563 & ~n11872 ;
  assign n11874 = n5895 & n6706 ;
  assign n11875 = ~n11868 & ~n11874 ;
  assign n11876 = n5565 & ~n11875 ;
  assign n11877 = ~n9570 & ~n11876 ;
  assign n11878 = n8899 & ~n11877 ;
  assign n11879 = ~n9528 & n9651 ;
  assign n11880 = \P2_reg0_reg[30]/NET0131  & ~n11879 ;
  assign n11881 = ~n11878 & ~n11880 ;
  assign n11882 = ~n11873 & n11881 ;
  assign n11883 = \P1_reg1_reg[9]/NET0131  & ~n6078 ;
  assign n11884 = \P1_reg1_reg[9]/NET0131  & n6095 ;
  assign n11886 = \P1_reg1_reg[9]/NET0131  & ~n6683 ;
  assign n11887 = n6683 & n11733 ;
  assign n11888 = ~n11886 & ~n11887 ;
  assign n11889 = n4011 & ~n11888 ;
  assign n11893 = n6683 & n11739 ;
  assign n11894 = ~n11886 & ~n11893 ;
  assign n11895 = n6207 & ~n11894 ;
  assign n11890 = n6683 & ~n11745 ;
  assign n11891 = ~n11886 & ~n11890 ;
  assign n11892 = n6282 & ~n11891 ;
  assign n11885 = n6683 & ~n11821 ;
  assign n11896 = \P1_reg1_reg[9]/NET0131  & ~n6695 ;
  assign n11897 = ~n11885 & ~n11896 ;
  assign n11898 = ~n11892 & n11897 ;
  assign n11899 = ~n11895 & n11898 ;
  assign n11900 = ~n11889 & n11899 ;
  assign n11901 = n6097 & ~n11900 ;
  assign n11902 = ~n11884 & ~n11901 ;
  assign n11903 = \P1_state_reg[0]/NET0131  & ~n11902 ;
  assign n11904 = ~n11883 & ~n11903 ;
  assign n11905 = \P2_reg0_reg[9]/NET0131  & ~n9531 ;
  assign n11907 = n5383 & n10457 ;
  assign n11906 = n5563 & n10472 ;
  assign n11908 = n5022 & n5565 ;
  assign n11909 = ~n11906 & ~n11908 ;
  assign n11910 = n10469 & n11909 ;
  assign n11911 = ~n11907 & n11910 ;
  assign n11912 = n9533 & ~n11911 ;
  assign n11913 = ~n11905 & ~n11912 ;
  assign n11914 = \P2_reg1_reg[10]/NET0131  & ~n8902 ;
  assign n11915 = ~n4997 & n5565 ;
  assign n11916 = n5563 & n10351 ;
  assign n11917 = ~n11915 & ~n11916 ;
  assign n11918 = n10345 & n11917 ;
  assign n11919 = n8913 & ~n11918 ;
  assign n11920 = ~n11914 & ~n11919 ;
  assign n11921 = \P2_reg1_reg[13]/NET0131  & ~n8902 ;
  assign n11922 = n4867 & n5565 ;
  assign n11923 = n10438 & ~n11922 ;
  assign n11924 = n8913 & ~n11923 ;
  assign n11925 = ~n11921 & ~n11924 ;
  assign n11926 = \P2_reg1_reg[23]/NET0131  & ~n5589 ;
  assign n11927 = \P2_reg1_reg[23]/NET0131  & ~n6380 ;
  assign n11928 = n6380 & ~n10734 ;
  assign n11929 = ~n11927 & ~n11928 ;
  assign n11930 = n5526 & ~n11929 ;
  assign n11931 = n6380 & ~n10747 ;
  assign n11932 = ~n11927 & ~n11931 ;
  assign n11933 = n5329 & ~n11932 ;
  assign n11934 = n6380 & ~n11041 ;
  assign n11935 = \P2_reg1_reg[23]/NET0131  & ~n8026 ;
  assign n11936 = ~n11934 & ~n11935 ;
  assign n11937 = ~n11933 & n11936 ;
  assign n11938 = ~n11930 & n11937 ;
  assign n11939 = n5583 & ~n11938 ;
  assign n11940 = \P2_reg1_reg[23]/NET0131  & n5585 ;
  assign n11941 = ~n11939 & ~n11940 ;
  assign n11942 = \P1_state_reg[0]/NET0131  & ~n11941 ;
  assign n11943 = ~n11926 & ~n11942 ;
  assign n11945 = \P2_reg1_reg[30]/NET0131  & ~n6380 ;
  assign n11946 = n8913 & n11870 ;
  assign n11947 = ~n11945 & ~n11946 ;
  assign n11948 = n5563 & ~n11947 ;
  assign n11944 = \P2_reg1_reg[30]/NET0131  & ~n9652 ;
  assign n11949 = n5895 & n6380 ;
  assign n11950 = ~n11945 & ~n11949 ;
  assign n11951 = n5565 & ~n11950 ;
  assign n11952 = ~n9662 & ~n11951 ;
  assign n11953 = n8899 & ~n11952 ;
  assign n11954 = ~n11944 & ~n11953 ;
  assign n11955 = ~n11948 & n11954 ;
  assign n11956 = \P2_reg1_reg[9]/NET0131  & ~n8902 ;
  assign n11957 = n8913 & ~n11911 ;
  assign n11958 = ~n11956 & ~n11957 ;
  assign n11959 = n4978 & n5574 ;
  assign n11960 = n4219 & ~n11918 ;
  assign n11961 = ~n11959 & ~n11960 ;
  assign n11962 = n8899 & ~n11961 ;
  assign n11963 = \P2_reg2_reg[10]/NET0131  & ~n9773 ;
  assign n11964 = ~n11962 & ~n11963 ;
  assign n11965 = \P2_reg2_reg[12]/NET0131  & ~n5589 ;
  assign n11966 = \P2_reg2_reg[12]/NET0131  & n5585 ;
  assign n11968 = \P2_reg2_reg[12]/NET0131  & ~n4219 ;
  assign n11972 = n4219 & n10385 ;
  assign n11973 = ~n11968 & ~n11972 ;
  assign n11974 = n5383 & ~n11973 ;
  assign n11969 = n4219 & n10375 ;
  assign n11970 = ~n11968 & ~n11969 ;
  assign n11971 = n5329 & ~n11970 ;
  assign n11975 = n4219 & ~n10391 ;
  assign n11976 = ~n11968 & ~n11975 ;
  assign n11977 = n5526 & ~n11976 ;
  assign n11979 = n4973 & n5565 ;
  assign n11980 = n5563 & n10397 ;
  assign n11981 = ~n11979 & ~n11980 ;
  assign n11982 = n4219 & ~n11981 ;
  assign n11967 = \P2_reg2_reg[12]/NET0131  & ~n6839 ;
  assign n11978 = n4952 & n5574 ;
  assign n11983 = ~n11967 & ~n11978 ;
  assign n11984 = ~n11982 & n11983 ;
  assign n11985 = ~n11977 & n11984 ;
  assign n11986 = ~n11971 & n11985 ;
  assign n11987 = ~n11974 & n11986 ;
  assign n11988 = n5583 & ~n11987 ;
  assign n11989 = ~n11966 & ~n11988 ;
  assign n11990 = \P1_state_reg[0]/NET0131  & ~n11989 ;
  assign n11991 = ~n11965 & ~n11990 ;
  assign n11992 = n4219 & ~n11923 ;
  assign n11993 = n4849 & n5574 ;
  assign n11994 = ~n11992 & ~n11993 ;
  assign n11995 = n8899 & ~n11994 ;
  assign n11996 = \P2_reg2_reg[13]/NET0131  & ~n9773 ;
  assign n11997 = ~n11995 & ~n11996 ;
  assign n11998 = \P2_reg2_reg[30]/NET0131  & ~n5589 ;
  assign n11999 = \P2_reg2_reg[30]/NET0131  & n5585 ;
  assign n12000 = \P2_reg2_reg[30]/NET0131  & ~n4219 ;
  assign n12001 = n4219 & n11870 ;
  assign n12002 = ~n12000 & ~n12001 ;
  assign n12003 = n5563 & ~n12002 ;
  assign n12004 = n4219 & n5895 ;
  assign n12005 = ~n12000 & ~n12004 ;
  assign n12006 = n5565 & ~n12005 ;
  assign n12007 = \P2_reg2_reg[30]/NET0131  & ~n8831 ;
  assign n12008 = ~n5575 & ~n12007 ;
  assign n12009 = ~n12006 & n12008 ;
  assign n12010 = ~n8826 & n12009 ;
  assign n12011 = ~n12003 & n12010 ;
  assign n12012 = n5583 & ~n12011 ;
  assign n12013 = ~n11999 & ~n12012 ;
  assign n12014 = \P1_state_reg[0]/NET0131  & ~n12013 ;
  assign n12015 = ~n11998 & ~n12014 ;
  assign n12016 = \P2_reg2_reg[9]/NET0131  & ~n9773 ;
  assign n12017 = n5003 & n5574 ;
  assign n12018 = n4219 & ~n11911 ;
  assign n12019 = ~n12017 & ~n12018 ;
  assign n12020 = n8899 & ~n12019 ;
  assign n12021 = ~n12016 & ~n12020 ;
  assign n12022 = \P1_reg0_reg[10]/NET0131  & ~n6078 ;
  assign n12023 = \P1_reg0_reg[10]/NET0131  & n6095 ;
  assign n12025 = \P1_reg0_reg[10]/NET0131  & ~n6409 ;
  assign n12032 = n6409 & n11661 ;
  assign n12033 = ~n12025 & ~n12032 ;
  assign n12034 = n4011 & ~n12033 ;
  assign n12029 = n6409 & ~n11673 ;
  assign n12030 = ~n12025 & ~n12029 ;
  assign n12031 = n6282 & ~n12030 ;
  assign n12026 = n6409 & n11667 ;
  assign n12027 = ~n12025 & ~n12026 ;
  assign n12028 = n6207 & ~n12027 ;
  assign n12035 = n6409 & n11678 ;
  assign n12036 = ~n12025 & ~n12035 ;
  assign n12037 = n6359 & ~n12036 ;
  assign n12024 = \P1_reg0_reg[10]/NET0131  & ~n6425 ;
  assign n12038 = n6409 & n11790 ;
  assign n12039 = ~n12024 & ~n12038 ;
  assign n12040 = ~n12037 & n12039 ;
  assign n12041 = ~n12028 & n12040 ;
  assign n12042 = ~n12031 & n12041 ;
  assign n12043 = ~n12034 & n12042 ;
  assign n12044 = n6097 & ~n12043 ;
  assign n12045 = ~n12023 & ~n12044 ;
  assign n12046 = \P1_state_reg[0]/NET0131  & ~n12045 ;
  assign n12047 = ~n12022 & ~n12046 ;
  assign n12048 = \P1_reg0_reg[13]/NET0131  & ~n9826 ;
  assign n12049 = n3345 & n6365 ;
  assign n12050 = n11715 & ~n12049 ;
  assign n12051 = n9829 & ~n12050 ;
  assign n12052 = ~n12048 & ~n12051 ;
  assign n12053 = ~n10008 & n11119 ;
  assign n12054 = \P1_reg0_reg[23]/NET0131  & ~n12053 ;
  assign n12055 = n9829 & ~n11847 ;
  assign n12056 = ~n12054 & ~n12055 ;
  assign n12057 = \P3_reg0_reg[10]/NET0131  & ~n2143 ;
  assign n12058 = \P3_reg0_reg[10]/NET0131  & n2145 ;
  assign n12064 = \P3_reg0_reg[10]/NET0131  & ~n2163 ;
  assign n12065 = ~n10495 & ~n12064 ;
  assign n12066 = n2391 & ~n12065 ;
  assign n12061 = \P3_reg0_reg[10]/NET0131  & ~n2236 ;
  assign n12062 = ~n10499 & ~n12061 ;
  assign n12063 = n2393 & ~n12062 ;
  assign n12067 = n2236 & ~n10507 ;
  assign n12068 = ~n12061 & ~n12067 ;
  assign n12069 = n737 & ~n12068 ;
  assign n12070 = n2163 & ~n10513 ;
  assign n12071 = ~n12064 & ~n12070 ;
  assign n12072 = n2234 & ~n12071 ;
  assign n12059 = ~n1651 & n2285 ;
  assign n12060 = n2163 & n12059 ;
  assign n12073 = \P3_reg0_reg[10]/NET0131  & ~n2287 ;
  assign n12074 = ~n12060 & ~n12073 ;
  assign n12075 = ~n12072 & n12074 ;
  assign n12076 = ~n12069 & n12075 ;
  assign n12077 = ~n12063 & n12076 ;
  assign n12078 = ~n12066 & n12077 ;
  assign n12079 = n2147 & ~n12078 ;
  assign n12080 = ~n12058 & ~n12079 ;
  assign n12081 = \P1_state_reg[0]/NET0131  & ~n12080 ;
  assign n12082 = ~n12057 & ~n12081 ;
  assign n12083 = \P3_reg0_reg[11]/NET0131  & ~n2143 ;
  assign n12084 = \P3_reg0_reg[11]/NET0131  & n2145 ;
  assign n12086 = \P3_reg0_reg[11]/NET0131  & ~n2236 ;
  assign n12087 = ~n10540 & ~n12086 ;
  assign n12088 = n2393 & ~n12087 ;
  assign n12089 = \P3_reg0_reg[11]/NET0131  & ~n2163 ;
  assign n12095 = n2163 & ~n10553 ;
  assign n12096 = ~n12089 & ~n12095 ;
  assign n12097 = n2234 & ~n12096 ;
  assign n12085 = \P3_reg0_reg[11]/NET0131  & ~n2287 ;
  assign n12098 = ~n1627 & n2289 ;
  assign n12099 = ~n12085 & ~n12098 ;
  assign n12100 = ~n12097 & n12099 ;
  assign n12101 = ~n12088 & n12100 ;
  assign n12090 = ~n10536 & ~n12089 ;
  assign n12091 = n2391 & ~n12090 ;
  assign n12092 = n2236 & ~n10547 ;
  assign n12093 = ~n12086 & ~n12092 ;
  assign n12094 = n737 & ~n12093 ;
  assign n12102 = ~n12091 & ~n12094 ;
  assign n12103 = n12101 & n12102 ;
  assign n12104 = n2147 & ~n12103 ;
  assign n12105 = ~n12084 & ~n12104 ;
  assign n12106 = \P1_state_reg[0]/NET0131  & ~n12105 ;
  assign n12107 = ~n12083 & ~n12106 ;
  assign n12108 = \P3_reg0_reg[12]/NET0131  & ~n2143 ;
  assign n12109 = \P3_reg0_reg[12]/NET0131  & n2145 ;
  assign n12111 = \P3_reg0_reg[12]/NET0131  & ~n2236 ;
  assign n12118 = n2236 & ~n10590 ;
  assign n12119 = ~n12111 & ~n12118 ;
  assign n12120 = n737 & ~n12119 ;
  assign n12114 = \P3_reg0_reg[12]/NET0131  & ~n2163 ;
  assign n12115 = n2163 & ~n10582 ;
  assign n12116 = ~n12114 & ~n12115 ;
  assign n12117 = n2234 & ~n12116 ;
  assign n12110 = \P3_reg0_reg[12]/NET0131  & ~n2287 ;
  assign n12123 = n1584 & n2289 ;
  assign n12124 = ~n12110 & ~n12123 ;
  assign n12125 = ~n12117 & n12124 ;
  assign n12126 = ~n12120 & n12125 ;
  assign n12112 = ~n10594 & ~n12111 ;
  assign n12113 = n2393 & ~n12112 ;
  assign n12121 = ~n10576 & ~n12114 ;
  assign n12122 = n2391 & ~n12121 ;
  assign n12127 = ~n12113 & ~n12122 ;
  assign n12128 = n12126 & n12127 ;
  assign n12129 = n2147 & ~n12128 ;
  assign n12130 = ~n12109 & ~n12129 ;
  assign n12131 = \P1_state_reg[0]/NET0131  & ~n12130 ;
  assign n12132 = ~n12108 & ~n12131 ;
  assign n12133 = \P3_reg0_reg[13]/NET0131  & ~n2143 ;
  assign n12134 = \P3_reg0_reg[13]/NET0131  & n2145 ;
  assign n12137 = \P3_reg0_reg[13]/NET0131  & ~n2236 ;
  assign n12145 = n2236 & ~n10629 ;
  assign n12146 = ~n12137 & ~n12145 ;
  assign n12147 = n737 & ~n12146 ;
  assign n12138 = ~n10621 & ~n12137 ;
  assign n12139 = n2393 & ~n12138 ;
  assign n12135 = ~n1560 & n2285 ;
  assign n12136 = n2163 & n12135 ;
  assign n12140 = \P3_reg0_reg[13]/NET0131  & ~n2287 ;
  assign n12150 = ~n12136 & ~n12140 ;
  assign n12151 = ~n12139 & n12150 ;
  assign n12141 = \P3_reg0_reg[13]/NET0131  & ~n2163 ;
  assign n12142 = n2163 & ~n10635 ;
  assign n12143 = ~n12141 & ~n12142 ;
  assign n12144 = n2234 & ~n12143 ;
  assign n12148 = ~n10616 & ~n12141 ;
  assign n12149 = n2391 & ~n12148 ;
  assign n12152 = ~n12144 & ~n12149 ;
  assign n12153 = n12151 & n12152 ;
  assign n12154 = ~n12147 & n12153 ;
  assign n12155 = n2147 & ~n12154 ;
  assign n12156 = ~n12134 & ~n12155 ;
  assign n12157 = \P1_state_reg[0]/NET0131  & ~n12156 ;
  assign n12158 = ~n12133 & ~n12157 ;
  assign n12159 = \P3_reg0_reg[14]/NET0131  & ~n2143 ;
  assign n12160 = \P3_reg0_reg[14]/NET0131  & n2145 ;
  assign n12169 = \P3_reg0_reg[14]/NET0131  & ~n2163 ;
  assign n12170 = ~n10669 & ~n12169 ;
  assign n12171 = n2391 & ~n12170 ;
  assign n12163 = \P3_reg0_reg[14]/NET0131  & ~n2236 ;
  assign n12167 = ~n10666 & ~n12163 ;
  assign n12168 = n2393 & ~n12167 ;
  assign n12164 = n2236 & ~n10658 ;
  assign n12165 = ~n12163 & ~n12164 ;
  assign n12166 = n737 & ~n12165 ;
  assign n12172 = n2163 & n10674 ;
  assign n12173 = ~n12169 & ~n12172 ;
  assign n12174 = n2234 & ~n12173 ;
  assign n12161 = ~n1544 & n2285 ;
  assign n12162 = n2163 & n12161 ;
  assign n12175 = \P3_reg0_reg[14]/NET0131  & ~n2287 ;
  assign n12176 = ~n12162 & ~n12175 ;
  assign n12177 = ~n12174 & n12176 ;
  assign n12178 = ~n12166 & n12177 ;
  assign n12179 = ~n12168 & n12178 ;
  assign n12180 = ~n12171 & n12179 ;
  assign n12181 = n2147 & ~n12180 ;
  assign n12182 = ~n12160 & ~n12181 ;
  assign n12183 = \P1_state_reg[0]/NET0131  & ~n12182 ;
  assign n12184 = ~n12159 & ~n12183 ;
  assign n12185 = \P3_reg0_reg[16]/NET0131  & ~n2143 ;
  assign n12186 = \P3_reg0_reg[16]/NET0131  & n2145 ;
  assign n12192 = \P3_reg0_reg[16]/NET0131  & ~n2163 ;
  assign n12197 = n2163 & ~n9172 ;
  assign n12198 = ~n12192 & ~n12197 ;
  assign n12199 = n2234 & ~n12198 ;
  assign n12188 = \P3_reg0_reg[16]/NET0131  & ~n2236 ;
  assign n12189 = n2236 & ~n9154 ;
  assign n12190 = ~n12188 & ~n12189 ;
  assign n12191 = n737 & ~n12190 ;
  assign n12187 = \P3_reg0_reg[16]/NET0131  & ~n2287 ;
  assign n12200 = ~n1185 & n2289 ;
  assign n12201 = ~n12187 & ~n12200 ;
  assign n12202 = ~n12191 & n12201 ;
  assign n12203 = ~n12199 & n12202 ;
  assign n12193 = ~n9167 & ~n12192 ;
  assign n12194 = n2391 & ~n12193 ;
  assign n12195 = ~n9164 & ~n12188 ;
  assign n12196 = n2393 & ~n12195 ;
  assign n12204 = ~n12194 & ~n12196 ;
  assign n12205 = n12203 & n12204 ;
  assign n12206 = n2147 & ~n12205 ;
  assign n12207 = ~n12186 & ~n12206 ;
  assign n12208 = \P1_state_reg[0]/NET0131  & ~n12207 ;
  assign n12209 = ~n12185 & ~n12208 ;
  assign n12210 = \P3_reg0_reg[9]/NET0131  & ~n2143 ;
  assign n12211 = \P3_reg0_reg[9]/NET0131  & n2145 ;
  assign n12222 = n2234 & ~n10297 ;
  assign n12220 = n2391 & n10291 ;
  assign n12221 = ~n1677 & n2285 ;
  assign n12223 = ~n12220 & ~n12221 ;
  assign n12224 = ~n12222 & n12223 ;
  assign n12225 = n2163 & ~n12224 ;
  assign n12216 = \P3_reg0_reg[9]/NET0131  & ~n2236 ;
  assign n12217 = n2236 & ~n10310 ;
  assign n12218 = ~n12216 & ~n12217 ;
  assign n12219 = n737 & ~n12218 ;
  assign n12212 = ~n2234 & ~n2391 ;
  assign n12213 = ~n2163 & ~n12212 ;
  assign n12214 = n2287 & ~n12213 ;
  assign n12215 = \P3_reg0_reg[9]/NET0131  & ~n12214 ;
  assign n12226 = ~n10292 & ~n12216 ;
  assign n12227 = n2393 & ~n12226 ;
  assign n12228 = ~n12215 & ~n12227 ;
  assign n12229 = ~n12219 & n12228 ;
  assign n12230 = ~n12225 & n12229 ;
  assign n12231 = n2147 & ~n12230 ;
  assign n12232 = ~n12211 & ~n12231 ;
  assign n12233 = \P1_state_reg[0]/NET0131  & ~n12232 ;
  assign n12234 = ~n12210 & ~n12233 ;
  assign n12235 = \P3_reg1_reg[10]/NET0131  & ~n2143 ;
  assign n12236 = \P3_reg1_reg[10]/NET0131  & n2145 ;
  assign n12238 = \P3_reg1_reg[10]/NET0131  & ~n2408 ;
  assign n12239 = n2408 & n10494 ;
  assign n12240 = ~n12238 & ~n12239 ;
  assign n12241 = n714 & ~n12240 ;
  assign n12242 = \P3_reg1_reg[10]/NET0131  & ~n2427 ;
  assign n12243 = n2427 & ~n10507 ;
  assign n12244 = ~n12242 & ~n12243 ;
  assign n12245 = n737 & ~n12244 ;
  assign n12250 = n2427 & ~n10513 ;
  assign n12251 = ~n12242 & ~n12250 ;
  assign n12252 = n2425 & ~n12251 ;
  assign n12247 = n2408 & ~n10513 ;
  assign n12248 = ~n12238 & ~n12247 ;
  assign n12249 = ~n2518 & ~n12248 ;
  assign n12237 = n2408 & n12059 ;
  assign n12246 = \P3_reg1_reg[10]/NET0131  & ~n6449 ;
  assign n12253 = ~n12237 & ~n12246 ;
  assign n12254 = ~n12249 & n12253 ;
  assign n12255 = ~n12252 & n12254 ;
  assign n12256 = ~n12245 & n12255 ;
  assign n12257 = ~n12241 & n12256 ;
  assign n12258 = n2147 & ~n12257 ;
  assign n12259 = ~n12236 & ~n12258 ;
  assign n12260 = \P1_state_reg[0]/NET0131  & ~n12259 ;
  assign n12261 = ~n12235 & ~n12260 ;
  assign n12262 = \P3_reg1_reg[11]/NET0131  & ~n2143 ;
  assign n12263 = \P3_reg1_reg[11]/NET0131  & n2145 ;
  assign n12272 = \P3_reg1_reg[11]/NET0131  & ~n2408 ;
  assign n12273 = n2408 & ~n10553 ;
  assign n12274 = ~n12272 & ~n12273 ;
  assign n12275 = ~n2518 & ~n12274 ;
  assign n12265 = \P3_reg1_reg[11]/NET0131  & ~n2427 ;
  assign n12269 = n2427 & ~n10553 ;
  assign n12270 = ~n12265 & ~n12269 ;
  assign n12271 = n2425 & ~n12270 ;
  assign n12264 = \P3_reg1_reg[11]/NET0131  & ~n6449 ;
  assign n12279 = ~n1627 & n6451 ;
  assign n12280 = ~n12264 & ~n12279 ;
  assign n12281 = ~n12271 & n12280 ;
  assign n12282 = ~n12275 & n12281 ;
  assign n12266 = n2427 & ~n10547 ;
  assign n12267 = ~n12265 & ~n12266 ;
  assign n12268 = n737 & ~n12267 ;
  assign n12276 = n2408 & n10535 ;
  assign n12277 = ~n12272 & ~n12276 ;
  assign n12278 = n714 & ~n12277 ;
  assign n12283 = ~n12268 & ~n12278 ;
  assign n12284 = n12282 & n12283 ;
  assign n12285 = n2147 & ~n12284 ;
  assign n12286 = ~n12263 & ~n12285 ;
  assign n12287 = \P1_state_reg[0]/NET0131  & ~n12286 ;
  assign n12288 = ~n12262 & ~n12287 ;
  assign n12289 = \P3_reg1_reg[12]/NET0131  & ~n2143 ;
  assign n12290 = \P3_reg1_reg[12]/NET0131  & n2145 ;
  assign n12296 = \P3_reg1_reg[12]/NET0131  & ~n2408 ;
  assign n12303 = n2408 & n10575 ;
  assign n12304 = ~n12296 & ~n12303 ;
  assign n12305 = n714 & ~n12304 ;
  assign n12292 = \P3_reg1_reg[12]/NET0131  & ~n2427 ;
  assign n12293 = n2427 & ~n10582 ;
  assign n12294 = ~n12292 & ~n12293 ;
  assign n12295 = n2425 & ~n12294 ;
  assign n12291 = \P3_reg1_reg[12]/NET0131  & ~n6449 ;
  assign n12306 = n1584 & n6451 ;
  assign n12307 = ~n12291 & ~n12306 ;
  assign n12308 = ~n12295 & n12307 ;
  assign n12297 = n2408 & ~n10582 ;
  assign n12298 = ~n12296 & ~n12297 ;
  assign n12299 = ~n2518 & ~n12298 ;
  assign n12300 = n2427 & ~n10590 ;
  assign n12301 = ~n12292 & ~n12300 ;
  assign n12302 = n737 & ~n12301 ;
  assign n12309 = ~n12299 & ~n12302 ;
  assign n12310 = n12308 & n12309 ;
  assign n12311 = ~n12305 & n12310 ;
  assign n12312 = n2147 & ~n12311 ;
  assign n12313 = ~n12290 & ~n12312 ;
  assign n12314 = \P1_state_reg[0]/NET0131  & ~n12313 ;
  assign n12315 = ~n12289 & ~n12314 ;
  assign n12316 = \P3_reg1_reg[13]/NET0131  & ~n2143 ;
  assign n12317 = \P3_reg1_reg[13]/NET0131  & n2145 ;
  assign n12327 = \P3_reg1_reg[13]/NET0131  & ~n2427 ;
  assign n12328 = n2427 & ~n10629 ;
  assign n12329 = ~n12327 & ~n12328 ;
  assign n12330 = n737 & ~n12329 ;
  assign n12319 = \P3_reg1_reg[13]/NET0131  & ~n2408 ;
  assign n12320 = n2408 & n10615 ;
  assign n12321 = ~n12319 & ~n12320 ;
  assign n12322 = n714 & ~n12321 ;
  assign n12318 = n2408 & n12135 ;
  assign n12323 = \P3_reg1_reg[13]/NET0131  & ~n6449 ;
  assign n12334 = ~n12318 & ~n12323 ;
  assign n12335 = ~n12322 & n12334 ;
  assign n12324 = n2408 & ~n10635 ;
  assign n12325 = ~n12319 & ~n12324 ;
  assign n12326 = ~n2518 & ~n12325 ;
  assign n12331 = n2427 & ~n10635 ;
  assign n12332 = ~n12327 & ~n12331 ;
  assign n12333 = n2425 & ~n12332 ;
  assign n12336 = ~n12326 & ~n12333 ;
  assign n12337 = n12335 & n12336 ;
  assign n12338 = ~n12330 & n12337 ;
  assign n12339 = n2147 & ~n12338 ;
  assign n12340 = ~n12317 & ~n12339 ;
  assign n12341 = \P1_state_reg[0]/NET0131  & ~n12340 ;
  assign n12342 = ~n12316 & ~n12341 ;
  assign n12343 = \P3_reg1_reg[14]/NET0131  & ~n2143 ;
  assign n12344 = \P3_reg1_reg[14]/NET0131  & n2145 ;
  assign n12346 = \P3_reg1_reg[14]/NET0131  & ~n2408 ;
  assign n12347 = n2408 & ~n10665 ;
  assign n12348 = ~n12346 & ~n12347 ;
  assign n12349 = n714 & ~n12348 ;
  assign n12350 = \P3_reg1_reg[14]/NET0131  & ~n2427 ;
  assign n12351 = n2427 & ~n10658 ;
  assign n12352 = ~n12350 & ~n12351 ;
  assign n12353 = n737 & ~n12352 ;
  assign n12358 = n2427 & n10674 ;
  assign n12359 = ~n12350 & ~n12358 ;
  assign n12360 = n2425 & ~n12359 ;
  assign n12355 = n2408 & n10674 ;
  assign n12356 = ~n12346 & ~n12355 ;
  assign n12357 = ~n2518 & ~n12356 ;
  assign n12345 = n2408 & n12161 ;
  assign n12354 = \P3_reg1_reg[14]/NET0131  & ~n6449 ;
  assign n12361 = ~n12345 & ~n12354 ;
  assign n12362 = ~n12357 & n12361 ;
  assign n12363 = ~n12360 & n12362 ;
  assign n12364 = ~n12353 & n12363 ;
  assign n12365 = ~n12349 & n12364 ;
  assign n12366 = n2147 & ~n12365 ;
  assign n12367 = ~n12344 & ~n12366 ;
  assign n12368 = \P1_state_reg[0]/NET0131  & ~n12367 ;
  assign n12369 = ~n12343 & ~n12368 ;
  assign n12370 = \P3_reg1_reg[16]/NET0131  & ~n2143 ;
  assign n12371 = \P3_reg1_reg[16]/NET0131  & n2145 ;
  assign n12377 = \P3_reg1_reg[16]/NET0131  & ~n2408 ;
  assign n12378 = n2408 & n9163 ;
  assign n12379 = ~n12377 & ~n12378 ;
  assign n12380 = n714 & ~n12379 ;
  assign n12373 = \P3_reg1_reg[16]/NET0131  & ~n2427 ;
  assign n12374 = n2427 & ~n9154 ;
  assign n12375 = ~n12373 & ~n12374 ;
  assign n12376 = n737 & ~n12375 ;
  assign n12372 = \P3_reg1_reg[16]/NET0131  & ~n6449 ;
  assign n12387 = ~n1185 & n6451 ;
  assign n12388 = ~n12372 & ~n12387 ;
  assign n12389 = ~n12376 & n12388 ;
  assign n12381 = n2427 & ~n9172 ;
  assign n12382 = ~n12373 & ~n12381 ;
  assign n12383 = n2425 & ~n12382 ;
  assign n12384 = n2408 & ~n9172 ;
  assign n12385 = ~n12377 & ~n12384 ;
  assign n12386 = ~n2518 & ~n12385 ;
  assign n12390 = ~n12383 & ~n12386 ;
  assign n12391 = n12389 & n12390 ;
  assign n12392 = ~n12380 & n12391 ;
  assign n12393 = n2147 & ~n12392 ;
  assign n12394 = ~n12371 & ~n12393 ;
  assign n12395 = \P1_state_reg[0]/NET0131  & ~n12394 ;
  assign n12396 = ~n12370 & ~n12395 ;
  assign n12397 = \P3_reg1_reg[9]/NET0131  & ~n2143 ;
  assign n12398 = \P3_reg1_reg[9]/NET0131  & n2145 ;
  assign n12404 = \P3_reg1_reg[9]/NET0131  & ~n2427 ;
  assign n12411 = n2427 & ~n10310 ;
  assign n12412 = ~n12404 & ~n12411 ;
  assign n12413 = n737 & ~n12412 ;
  assign n12400 = \P3_reg1_reg[9]/NET0131  & ~n2408 ;
  assign n12401 = n2408 & n10291 ;
  assign n12402 = ~n12400 & ~n12401 ;
  assign n12403 = n714 & ~n12402 ;
  assign n12399 = n2408 & n12221 ;
  assign n12414 = \P3_reg1_reg[9]/NET0131  & ~n6449 ;
  assign n12415 = ~n12399 & ~n12414 ;
  assign n12416 = ~n12403 & n12415 ;
  assign n12405 = n2427 & ~n10297 ;
  assign n12406 = ~n12404 & ~n12405 ;
  assign n12407 = n2425 & ~n12406 ;
  assign n12408 = n2408 & ~n10297 ;
  assign n12409 = ~n12400 & ~n12408 ;
  assign n12410 = ~n2518 & ~n12409 ;
  assign n12417 = ~n12407 & ~n12410 ;
  assign n12418 = n12416 & n12417 ;
  assign n12419 = ~n12413 & n12418 ;
  assign n12420 = n2147 & ~n12419 ;
  assign n12421 = ~n12398 & ~n12420 ;
  assign n12422 = \P1_state_reg[0]/NET0131  & ~n12421 ;
  assign n12423 = ~n12397 & ~n12422 ;
  assign n12424 = \P3_reg2_reg[10]/NET0131  & ~n2143 ;
  assign n12425 = \P3_reg2_reg[10]/NET0131  & n2145 ;
  assign n12427 = \P3_reg2_reg[10]/NET0131  & ~n2427 ;
  assign n12428 = n2427 & n10494 ;
  assign n12429 = ~n12427 & ~n12428 ;
  assign n12430 = n714 & ~n12429 ;
  assign n12431 = \P3_reg2_reg[10]/NET0131  & ~n2408 ;
  assign n12432 = n2408 & ~n10507 ;
  assign n12433 = ~n12431 & ~n12432 ;
  assign n12434 = n737 & ~n12433 ;
  assign n12437 = ~n12247 & ~n12431 ;
  assign n12438 = n2425 & ~n12437 ;
  assign n12435 = ~n12250 & ~n12427 ;
  assign n12436 = ~n2518 & ~n12435 ;
  assign n12426 = n2427 & n12059 ;
  assign n12439 = ~n1631 & n2283 ;
  assign n12440 = \P3_reg2_reg[10]/NET0131  & ~n2429 ;
  assign n12441 = ~n12439 & ~n12440 ;
  assign n12442 = ~n12426 & n12441 ;
  assign n12443 = ~n12436 & n12442 ;
  assign n12444 = ~n12438 & n12443 ;
  assign n12445 = ~n12434 & n12444 ;
  assign n12446 = ~n12430 & n12445 ;
  assign n12447 = n2147 & ~n12446 ;
  assign n12448 = ~n12425 & ~n12447 ;
  assign n12449 = \P1_state_reg[0]/NET0131  & ~n12448 ;
  assign n12450 = ~n12424 & ~n12449 ;
  assign n12451 = \P3_reg2_reg[11]/NET0131  & ~n2143 ;
  assign n12452 = \P3_reg2_reg[11]/NET0131  & n2145 ;
  assign n12460 = \P3_reg2_reg[11]/NET0131  & ~n2427 ;
  assign n12461 = ~n12269 & ~n12460 ;
  assign n12462 = ~n2518 & ~n12461 ;
  assign n12454 = \P3_reg2_reg[11]/NET0131  & ~n2408 ;
  assign n12458 = ~n12273 & ~n12454 ;
  assign n12459 = n2425 & ~n12458 ;
  assign n12467 = ~n1627 & n2441 ;
  assign n12453 = \P3_reg2_reg[11]/NET0131  & ~n2429 ;
  assign n12466 = ~n1608 & n2283 ;
  assign n12468 = ~n12453 & ~n12466 ;
  assign n12469 = ~n12467 & n12468 ;
  assign n12470 = ~n12459 & n12469 ;
  assign n12471 = ~n12462 & n12470 ;
  assign n12455 = n2408 & ~n10547 ;
  assign n12456 = ~n12454 & ~n12455 ;
  assign n12457 = n737 & ~n12456 ;
  assign n12463 = n2427 & n10535 ;
  assign n12464 = ~n12460 & ~n12463 ;
  assign n12465 = n714 & ~n12464 ;
  assign n12472 = ~n12457 & ~n12465 ;
  assign n12473 = n12471 & n12472 ;
  assign n12474 = n2147 & ~n12473 ;
  assign n12475 = ~n12452 & ~n12474 ;
  assign n12476 = \P1_state_reg[0]/NET0131  & ~n12475 ;
  assign n12477 = ~n12451 & ~n12476 ;
  assign n12478 = \P3_reg2_reg[12]/NET0131  & ~n2143 ;
  assign n12479 = \P3_reg2_reg[12]/NET0131  & n2145 ;
  assign n12484 = \P3_reg2_reg[12]/NET0131  & ~n2427 ;
  assign n12490 = n2427 & n10575 ;
  assign n12491 = ~n12484 & ~n12490 ;
  assign n12492 = n714 & ~n12491 ;
  assign n12481 = \P3_reg2_reg[12]/NET0131  & ~n2408 ;
  assign n12482 = ~n12297 & ~n12481 ;
  assign n12483 = n2425 & ~n12482 ;
  assign n12494 = n1584 & n2441 ;
  assign n12480 = \P3_reg2_reg[12]/NET0131  & ~n2429 ;
  assign n12493 = ~n1589 & n2283 ;
  assign n12495 = ~n12480 & ~n12493 ;
  assign n12496 = ~n12494 & n12495 ;
  assign n12497 = ~n12483 & n12496 ;
  assign n12485 = ~n12293 & ~n12484 ;
  assign n12486 = ~n2518 & ~n12485 ;
  assign n12487 = n2408 & ~n10590 ;
  assign n12488 = ~n12481 & ~n12487 ;
  assign n12489 = n737 & ~n12488 ;
  assign n12498 = ~n12486 & ~n12489 ;
  assign n12499 = n12497 & n12498 ;
  assign n12500 = ~n12492 & n12499 ;
  assign n12501 = n2147 & ~n12500 ;
  assign n12502 = ~n12479 & ~n12501 ;
  assign n12503 = \P1_state_reg[0]/NET0131  & ~n12502 ;
  assign n12504 = ~n12478 & ~n12503 ;
  assign n12505 = \P3_reg2_reg[13]/NET0131  & ~n2143 ;
  assign n12506 = \P3_reg2_reg[13]/NET0131  & n2145 ;
  assign n12514 = \P3_reg2_reg[13]/NET0131  & ~n2408 ;
  assign n12515 = n2408 & ~n10629 ;
  assign n12516 = ~n12514 & ~n12515 ;
  assign n12517 = n737 & ~n12516 ;
  assign n12508 = \P3_reg2_reg[13]/NET0131  & ~n2427 ;
  assign n12509 = n2427 & n10615 ;
  assign n12510 = ~n12508 & ~n12509 ;
  assign n12511 = n714 & ~n12510 ;
  assign n12507 = n2427 & n12135 ;
  assign n12520 = ~n1564 & n2283 ;
  assign n12521 = \P3_reg2_reg[13]/NET0131  & ~n2429 ;
  assign n12522 = ~n12520 & ~n12521 ;
  assign n12523 = ~n12507 & n12522 ;
  assign n12524 = ~n12511 & n12523 ;
  assign n12512 = ~n12331 & ~n12508 ;
  assign n12513 = ~n2518 & ~n12512 ;
  assign n12518 = ~n12324 & ~n12514 ;
  assign n12519 = n2425 & ~n12518 ;
  assign n12525 = ~n12513 & ~n12519 ;
  assign n12526 = n12524 & n12525 ;
  assign n12527 = ~n12517 & n12526 ;
  assign n12528 = n2147 & ~n12527 ;
  assign n12529 = ~n12506 & ~n12528 ;
  assign n12530 = \P1_state_reg[0]/NET0131  & ~n12529 ;
  assign n12531 = ~n12505 & ~n12530 ;
  assign n12532 = \P3_reg2_reg[14]/NET0131  & ~n2143 ;
  assign n12533 = \P3_reg2_reg[14]/NET0131  & n2145 ;
  assign n12535 = \P3_reg2_reg[14]/NET0131  & ~n2427 ;
  assign n12536 = n2427 & ~n10665 ;
  assign n12537 = ~n12535 & ~n12536 ;
  assign n12538 = n714 & ~n12537 ;
  assign n12539 = \P3_reg2_reg[14]/NET0131  & ~n2408 ;
  assign n12540 = n2408 & ~n10658 ;
  assign n12541 = ~n12539 & ~n12540 ;
  assign n12542 = n737 & ~n12541 ;
  assign n12545 = ~n12358 & ~n12535 ;
  assign n12546 = ~n2518 & ~n12545 ;
  assign n12543 = ~n12355 & ~n12539 ;
  assign n12544 = n2425 & ~n12543 ;
  assign n12534 = n2427 & n12161 ;
  assign n12547 = ~n1525 & n2283 ;
  assign n12548 = \P3_reg2_reg[14]/NET0131  & ~n2429 ;
  assign n12549 = ~n12547 & ~n12548 ;
  assign n12550 = ~n12534 & n12549 ;
  assign n12551 = ~n12544 & n12550 ;
  assign n12552 = ~n12546 & n12551 ;
  assign n12553 = ~n12542 & n12552 ;
  assign n12554 = ~n12538 & n12553 ;
  assign n12555 = n2147 & ~n12554 ;
  assign n12556 = ~n12533 & ~n12555 ;
  assign n12557 = \P1_state_reg[0]/NET0131  & ~n12556 ;
  assign n12558 = ~n12532 & ~n12557 ;
  assign n12559 = \P3_reg2_reg[16]/NET0131  & ~n2143 ;
  assign n12560 = \P3_reg2_reg[16]/NET0131  & n2145 ;
  assign n12566 = \P3_reg2_reg[16]/NET0131  & ~n2427 ;
  assign n12567 = n2427 & n9163 ;
  assign n12568 = ~n12566 & ~n12567 ;
  assign n12569 = n714 & ~n12568 ;
  assign n12562 = \P3_reg2_reg[16]/NET0131  & ~n2408 ;
  assign n12563 = n2408 & ~n9154 ;
  assign n12564 = ~n12562 & ~n12563 ;
  assign n12565 = n737 & ~n12564 ;
  assign n12575 = ~n1185 & n2441 ;
  assign n12561 = \P3_reg2_reg[16]/NET0131  & ~n2429 ;
  assign n12574 = ~n1193 & n2283 ;
  assign n12576 = ~n12561 & ~n12574 ;
  assign n12577 = ~n12575 & n12576 ;
  assign n12578 = ~n12565 & n12577 ;
  assign n12570 = ~n12384 & ~n12562 ;
  assign n12571 = n2425 & ~n12570 ;
  assign n12572 = ~n12381 & ~n12566 ;
  assign n12573 = ~n2518 & ~n12572 ;
  assign n12579 = ~n12571 & ~n12573 ;
  assign n12580 = n12578 & n12579 ;
  assign n12581 = ~n12569 & n12580 ;
  assign n12582 = n2147 & ~n12581 ;
  assign n12583 = ~n12560 & ~n12582 ;
  assign n12584 = \P1_state_reg[0]/NET0131  & ~n12583 ;
  assign n12585 = ~n12559 & ~n12584 ;
  assign n12586 = \P1_reg0_reg[8]/NET0131  & ~n6078 ;
  assign n12587 = \P1_reg0_reg[8]/NET0131  & n6095 ;
  assign n12594 = \P1_reg0_reg[8]/NET0131  & ~n6409 ;
  assign n12595 = n6409 & n11540 ;
  assign n12596 = ~n12594 & ~n12595 ;
  assign n12597 = n4011 & ~n12596 ;
  assign n12598 = n6409 & n11546 ;
  assign n12599 = ~n12594 & ~n12598 ;
  assign n12600 = n6207 & ~n12599 ;
  assign n12589 = n6282 & ~n11552 ;
  assign n12588 = n6359 & n11557 ;
  assign n12590 = n3813 & n6365 ;
  assign n12591 = ~n12588 & ~n12590 ;
  assign n12592 = ~n12589 & n12591 ;
  assign n12593 = n6409 & ~n12592 ;
  assign n12601 = n6282 & ~n6409 ;
  assign n12602 = n11142 & ~n12601 ;
  assign n12603 = \P1_reg0_reg[8]/NET0131  & ~n12602 ;
  assign n12604 = ~n12593 & ~n12603 ;
  assign n12605 = ~n12600 & n12604 ;
  assign n12606 = ~n12597 & n12605 ;
  assign n12607 = n6097 & ~n12606 ;
  assign n12608 = ~n12587 & ~n12607 ;
  assign n12609 = \P1_state_reg[0]/NET0131  & ~n12608 ;
  assign n12610 = ~n12586 & ~n12609 ;
  assign n12611 = n9044 & ~n9546 ;
  assign n12612 = n7807 & n12611 ;
  assign n12613 = \P1_reg1_reg[13]/NET0131  & ~n12612 ;
  assign n12614 = n9045 & ~n12050 ;
  assign n12615 = ~n12613 & ~n12614 ;
  assign n12616 = \P2_reg0_reg[10]/NET0131  & ~n9531 ;
  assign n12617 = n9533 & ~n11918 ;
  assign n12618 = ~n12616 & ~n12617 ;
  assign n12619 = \P3_reg2_reg[9]/NET0131  & ~n2143 ;
  assign n12620 = \P3_reg2_reg[9]/NET0131  & n2145 ;
  assign n12626 = \P3_reg2_reg[9]/NET0131  & ~n2408 ;
  assign n12631 = n2408 & ~n10310 ;
  assign n12632 = ~n12626 & ~n12631 ;
  assign n12633 = n737 & ~n12632 ;
  assign n12622 = \P3_reg2_reg[9]/NET0131  & ~n2427 ;
  assign n12623 = n2427 & n10291 ;
  assign n12624 = ~n12622 & ~n12623 ;
  assign n12625 = n714 & ~n12624 ;
  assign n12635 = \P3_reg2_reg[9]/NET0131  & ~n2429 ;
  assign n12621 = n2427 & n12221 ;
  assign n12634 = ~n1657 & n2283 ;
  assign n12636 = ~n12621 & ~n12634 ;
  assign n12637 = ~n12635 & n12636 ;
  assign n12638 = ~n12625 & n12637 ;
  assign n12627 = ~n12408 & ~n12626 ;
  assign n12628 = n2425 & ~n12627 ;
  assign n12629 = ~n12405 & ~n12622 ;
  assign n12630 = ~n2518 & ~n12629 ;
  assign n12639 = ~n12628 & ~n12630 ;
  assign n12640 = n12638 & n12639 ;
  assign n12641 = ~n12633 & n12640 ;
  assign n12642 = n2147 & ~n12641 ;
  assign n12643 = ~n12620 & ~n12642 ;
  assign n12644 = \P1_state_reg[0]/NET0131  & ~n12643 ;
  assign n12645 = ~n12619 & ~n12644 ;
  assign n12646 = n5327 & ~n5524 ;
  assign n12647 = ~n6706 & n12646 ;
  assign n12648 = n9530 & ~n12647 ;
  assign n12649 = \P2_reg0_reg[13]/NET0131  & ~n12648 ;
  assign n12650 = n9533 & ~n11923 ;
  assign n12651 = ~n12649 & ~n12650 ;
  assign n12653 = n3223 & n6095 ;
  assign n12672 = ~n3232 & n8676 ;
  assign n12671 = n3232 & ~n8676 ;
  assign n12673 = n6207 & ~n12671 ;
  assign n12674 = ~n12672 & n12673 ;
  assign n12665 = n3232 & n7137 ;
  assign n12664 = ~n3232 & ~n7137 ;
  assign n12666 = n6282 & ~n12664 ;
  assign n12667 = ~n12665 & n12666 ;
  assign n12668 = n3219 & ~n11701 ;
  assign n12669 = ~n6341 & n6359 ;
  assign n12670 = ~n12668 & n12669 ;
  assign n12675 = ~n12667 & ~n12670 ;
  assign n12676 = ~n12674 & n12675 ;
  assign n12677 = n6568 & ~n12676 ;
  assign n12655 = n3623 & ~n11384 ;
  assign n12656 = ~n11385 & ~n12655 ;
  assign n12657 = ~n2713 & ~n12656 ;
  assign n12658 = n2713 & n3354 ;
  assign n12659 = ~n12657 & ~n12658 ;
  assign n12660 = n6568 & ~n12659 ;
  assign n12661 = ~n3223 & ~n6568 ;
  assign n12662 = n4011 & ~n12661 ;
  assign n12663 = ~n12660 & n12662 ;
  assign n12654 = n3223 & ~n11314 ;
  assign n12678 = n3219 & ~n6649 ;
  assign n12679 = ~n12654 & ~n12678 ;
  assign n12680 = ~n12663 & n12679 ;
  assign n12681 = ~n12677 & n12680 ;
  assign n12682 = n6097 & ~n12681 ;
  assign n12683 = ~n12653 & ~n12682 ;
  assign n12684 = \P1_state_reg[0]/NET0131  & ~n12683 ;
  assign n12652 = \P1_reg3_reg[14]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n12685 = n3223 & n4130 ;
  assign n12686 = ~n12652 & ~n12685 ;
  assign n12687 = ~n12684 & n12686 ;
  assign n12689 = n5110 & n5585 ;
  assign n12693 = n5092 & ~n5351 ;
  assign n12694 = ~n5352 & ~n12693 ;
  assign n12695 = ~n4231 & ~n12694 ;
  assign n12696 = n4231 & n5203 ;
  assign n12697 = ~n12695 & ~n12696 ;
  assign n12698 = n5383 & n12697 ;
  assign n12708 = ~n5250 & n5976 ;
  assign n12707 = n5250 & ~n5976 ;
  assign n12709 = n5329 & ~n12707 ;
  assign n12710 = ~n12708 & n12709 ;
  assign n12700 = n5131 & ~n5532 ;
  assign n12699 = ~n5131 & n5532 ;
  assign n12701 = n5563 & ~n12699 ;
  assign n12702 = ~n12700 & n12701 ;
  assign n12704 = ~n5430 & ~n5976 ;
  assign n12703 = n5430 & n5976 ;
  assign n12705 = n5526 & ~n12703 ;
  assign n12706 = ~n12704 & n12705 ;
  assign n12711 = ~n12702 & ~n12706 ;
  assign n12712 = ~n12710 & n12711 ;
  assign n12713 = ~n12698 & n12712 ;
  assign n12714 = n7453 & ~n12713 ;
  assign n12690 = n8639 & ~n11434 ;
  assign n12691 = ~n8640 & n12690 ;
  assign n12692 = n5110 & ~n12691 ;
  assign n12715 = n5131 & ~n7504 ;
  assign n12716 = ~n12692 & ~n12715 ;
  assign n12717 = ~n12714 & n12716 ;
  assign n12718 = n5583 & ~n12717 ;
  assign n12719 = ~n12689 & ~n12718 ;
  assign n12720 = \P1_state_reg[0]/NET0131  & ~n12719 ;
  assign n12688 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[5]/NET0131  ;
  assign n12721 = n5110 & n5786 ;
  assign n12722 = ~n12688 & ~n12721 ;
  assign n12723 = ~n12720 & n12722 ;
  assign n12726 = n3791 & n6095 ;
  assign n12733 = n3791 & ~n6568 ;
  assign n12734 = n2713 & ~n3756 ;
  assign n12735 = ~n3795 & n6288 ;
  assign n12736 = n3137 & ~n12735 ;
  assign n12737 = ~n2713 & ~n6290 ;
  assign n12738 = ~n12736 & n12737 ;
  assign n12739 = ~n12734 & ~n12738 ;
  assign n12740 = n6568 & ~n12739 ;
  assign n12741 = ~n12733 & ~n12740 ;
  assign n12742 = n4011 & ~n12741 ;
  assign n12749 = ~n3798 & n4045 ;
  assign n12750 = n3798 & ~n4045 ;
  assign n12751 = ~n12749 & ~n12750 ;
  assign n12752 = n6568 & n12751 ;
  assign n12753 = ~n12733 & ~n12752 ;
  assign n12754 = n6282 & ~n12753 ;
  assign n12743 = n3798 & ~n6988 ;
  assign n12744 = ~n3798 & n6988 ;
  assign n12745 = ~n12743 & ~n12744 ;
  assign n12746 = n6568 & ~n12745 ;
  assign n12747 = ~n12733 & ~n12746 ;
  assign n12748 = n6207 & ~n12747 ;
  assign n12727 = ~n3786 & n6365 ;
  assign n12728 = ~n3786 & ~n6330 ;
  assign n12729 = ~n6331 & n6359 ;
  assign n12730 = ~n12728 & n12729 ;
  assign n12731 = ~n12727 & ~n12730 ;
  assign n12732 = n6568 & ~n12731 ;
  assign n12755 = ~n3786 & n4112 ;
  assign n12756 = ~n6568 & n6693 ;
  assign n12757 = ~n6361 & ~n12756 ;
  assign n12758 = n3791 & ~n12757 ;
  assign n12759 = ~n12755 & ~n12758 ;
  assign n12760 = ~n12732 & n12759 ;
  assign n12761 = ~n12748 & n12760 ;
  assign n12762 = ~n12754 & n12761 ;
  assign n12763 = ~n12742 & n12762 ;
  assign n12764 = n6097 & ~n12763 ;
  assign n12765 = ~n12726 & ~n12764 ;
  assign n12766 = \P1_state_reg[0]/NET0131  & ~n12765 ;
  assign n12724 = \P1_reg3_reg[4]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n12725 = n3791 & n4130 ;
  assign n12767 = ~n12724 & ~n12725 ;
  assign n12768 = ~n12766 & n12767 ;
  assign n12771 = n3133 & n6095 ;
  assign n12778 = n3133 & ~n6568 ;
  assign n12779 = n3140 & ~n6146 ;
  assign n12780 = ~n3140 & n6146 ;
  assign n12781 = ~n12779 & ~n12780 ;
  assign n12782 = n6568 & n12781 ;
  assign n12783 = ~n12778 & ~n12782 ;
  assign n12784 = n6207 & ~n12783 ;
  assign n12772 = ~n3128 & n6365 ;
  assign n12773 = ~n3128 & ~n6331 ;
  assign n12774 = ~n6332 & ~n12773 ;
  assign n12775 = n6359 & n12774 ;
  assign n12776 = ~n12772 & ~n12775 ;
  assign n12777 = n6568 & ~n12776 ;
  assign n12799 = ~n3128 & n4112 ;
  assign n12800 = n3133 & ~n12757 ;
  assign n12801 = ~n12799 & ~n12800 ;
  assign n12802 = ~n12777 & n12801 ;
  assign n12803 = ~n12784 & n12802 ;
  assign n12785 = n3746 & ~n6290 ;
  assign n12786 = ~n6291 & ~n12785 ;
  assign n12787 = ~n2713 & ~n12786 ;
  assign n12788 = n2713 & n3795 ;
  assign n12789 = ~n12787 & ~n12788 ;
  assign n12790 = n6568 & n12789 ;
  assign n12791 = ~n12778 & ~n12790 ;
  assign n12792 = n4011 & ~n12791 ;
  assign n12793 = n3140 & ~n6218 ;
  assign n12794 = ~n3140 & n6218 ;
  assign n12795 = ~n12793 & ~n12794 ;
  assign n12796 = n6568 & ~n12795 ;
  assign n12797 = ~n12778 & ~n12796 ;
  assign n12798 = n6282 & ~n12797 ;
  assign n12804 = ~n12792 & ~n12798 ;
  assign n12805 = n12803 & n12804 ;
  assign n12806 = n6097 & ~n12805 ;
  assign n12807 = ~n12771 & ~n12806 ;
  assign n12808 = \P1_state_reg[0]/NET0131  & ~n12807 ;
  assign n12769 = \P1_reg3_reg[5]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n12770 = n3133 & n4130 ;
  assign n12809 = ~n12769 & ~n12770 ;
  assign n12810 = ~n12808 & n12809 ;
  assign n12813 = ~n1774 & n2145 ;
  assign n12823 = ~n1774 & ~n2163 ;
  assign n12828 = n1755 & ~n2248 ;
  assign n12827 = ~n1755 & n2248 ;
  assign n12829 = ~n2239 & ~n12827 ;
  assign n12830 = ~n12828 & n12829 ;
  assign n12831 = ~n1806 & n2239 ;
  assign n12832 = ~n12830 & ~n12831 ;
  assign n12833 = n2163 & ~n12832 ;
  assign n12834 = ~n12823 & ~n12833 ;
  assign n12835 = n737 & ~n12834 ;
  assign n12816 = ~n1795 & ~n1822 ;
  assign n12817 = ~n2320 & n12816 ;
  assign n12818 = n2320 & ~n12816 ;
  assign n12819 = ~n12817 & ~n12818 ;
  assign n12824 = n2163 & ~n12819 ;
  assign n12825 = ~n12823 & ~n12824 ;
  assign n12826 = n2393 & ~n12825 ;
  assign n12815 = ~n1774 & ~n2236 ;
  assign n12820 = n2236 & ~n12819 ;
  assign n12821 = ~n12815 & ~n12820 ;
  assign n12822 = n2391 & ~n12821 ;
  assign n12836 = ~n2170 & n12816 ;
  assign n12837 = n2170 & ~n12816 ;
  assign n12838 = ~n12836 & ~n12837 ;
  assign n12839 = n2236 & n12838 ;
  assign n12840 = ~n12815 & ~n12839 ;
  assign n12841 = n2234 & ~n12840 ;
  assign n12814 = ~n1794 & n2580 ;
  assign n12842 = ~n1774 & ~n2583 ;
  assign n12843 = ~n12814 & ~n12842 ;
  assign n12844 = ~n12841 & n12843 ;
  assign n12845 = ~n12822 & n12844 ;
  assign n12846 = ~n12826 & n12845 ;
  assign n12847 = ~n12835 & n12846 ;
  assign n12848 = n2147 & ~n12847 ;
  assign n12849 = ~n12813 & ~n12848 ;
  assign n12850 = \P1_state_reg[0]/NET0131  & ~n12849 ;
  assign n12811 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[5]/NET0131  ;
  assign n12812 = n765 & ~n1774 ;
  assign n12851 = ~n12811 & ~n12812 ;
  assign n12852 = ~n12850 & n12851 ;
  assign n12855 = ~n1750 & n2145 ;
  assign n12857 = ~n1750 & ~n2163 ;
  assign n12873 = n1729 & ~n12827 ;
  assign n12872 = ~n1729 & n12827 ;
  assign n12874 = ~n2239 & ~n12872 ;
  assign n12875 = ~n12873 & n12874 ;
  assign n12876 = ~n1779 & n2239 ;
  assign n12877 = ~n12875 & ~n12876 ;
  assign n12878 = n2163 & ~n12877 ;
  assign n12879 = ~n12857 & ~n12878 ;
  assign n12880 = n737 & ~n12879 ;
  assign n12858 = n2068 & ~n2459 ;
  assign n12859 = ~n2068 & n2459 ;
  assign n12860 = ~n12858 & ~n12859 ;
  assign n12861 = n2163 & ~n12860 ;
  assign n12862 = ~n12857 & ~n12861 ;
  assign n12863 = n2393 & ~n12862 ;
  assign n12856 = ~n1768 & n2580 ;
  assign n12864 = ~n1750 & ~n2583 ;
  assign n12884 = ~n12856 & ~n12864 ;
  assign n12885 = ~n12863 & n12884 ;
  assign n12865 = ~n1750 & ~n2236 ;
  assign n12866 = ~n1975 & n2068 ;
  assign n12867 = n1975 & ~n2068 ;
  assign n12868 = ~n12866 & ~n12867 ;
  assign n12869 = n2236 & n12868 ;
  assign n12870 = ~n12865 & ~n12869 ;
  assign n12871 = n2234 & ~n12870 ;
  assign n12881 = n2236 & ~n12860 ;
  assign n12882 = ~n12865 & ~n12881 ;
  assign n12883 = n2391 & ~n12882 ;
  assign n12886 = ~n12871 & ~n12883 ;
  assign n12887 = n12885 & n12886 ;
  assign n12888 = ~n12880 & n12887 ;
  assign n12889 = n2147 & ~n12888 ;
  assign n12890 = ~n12855 & ~n12889 ;
  assign n12891 = \P1_state_reg[0]/NET0131  & ~n12890 ;
  assign n12853 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[6]/NET0131  ;
  assign n12854 = n765 & ~n1750 ;
  assign n12892 = ~n12853 & ~n12854 ;
  assign n12893 = ~n12891 & n12892 ;
  assign n12896 = ~n1724 & n2145 ;
  assign n12905 = ~n1724 & ~n2163 ;
  assign n12909 = ~n1755 & n2239 ;
  assign n12910 = n1687 & ~n12872 ;
  assign n12911 = ~n2239 & ~n2251 ;
  assign n12912 = ~n12910 & n12911 ;
  assign n12913 = ~n12909 & ~n12912 ;
  assign n12914 = n2163 & ~n12913 ;
  assign n12915 = ~n12905 & ~n12914 ;
  assign n12916 = n737 & ~n12915 ;
  assign n12899 = n2035 & ~n2533 ;
  assign n12900 = ~n2035 & n2533 ;
  assign n12901 = ~n12899 & ~n12900 ;
  assign n12906 = n2163 & n12901 ;
  assign n12907 = ~n12905 & ~n12906 ;
  assign n12908 = n2393 & ~n12907 ;
  assign n12898 = ~n1724 & ~n2236 ;
  assign n12902 = n2236 & n12901 ;
  assign n12903 = ~n12898 & ~n12902 ;
  assign n12904 = n2391 & ~n12903 ;
  assign n12917 = n2035 & ~n2588 ;
  assign n12918 = ~n2035 & n2588 ;
  assign n12919 = ~n12917 & ~n12918 ;
  assign n12920 = n2236 & ~n12919 ;
  assign n12921 = ~n12898 & ~n12920 ;
  assign n12922 = n2234 & ~n12921 ;
  assign n12897 = ~n1744 & n2580 ;
  assign n12923 = ~n1724 & ~n2583 ;
  assign n12924 = ~n12897 & ~n12923 ;
  assign n12925 = ~n12922 & n12924 ;
  assign n12926 = ~n12904 & n12925 ;
  assign n12927 = ~n12908 & n12926 ;
  assign n12928 = ~n12916 & n12927 ;
  assign n12929 = n2147 & ~n12928 ;
  assign n12930 = ~n12896 & ~n12929 ;
  assign n12931 = \P1_state_reg[0]/NET0131  & ~n12930 ;
  assign n12894 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[7]/NET0131  ;
  assign n12895 = n765 & ~n1724 ;
  assign n12932 = ~n12894 & ~n12895 ;
  assign n12933 = ~n12931 & n12932 ;
  assign n12934 = \P1_reg1_reg[8]/NET0131  & ~n6078 ;
  assign n12935 = \P1_reg1_reg[8]/NET0131  & n6095 ;
  assign n12937 = \P1_reg1_reg[8]/NET0131  & ~n6683 ;
  assign n12938 = n6683 & n11540 ;
  assign n12939 = ~n12937 & ~n12938 ;
  assign n12940 = n4011 & ~n12939 ;
  assign n12941 = n6683 & n11546 ;
  assign n12942 = ~n12937 & ~n12941 ;
  assign n12943 = n6207 & ~n12942 ;
  assign n12936 = n6683 & ~n12592 ;
  assign n12944 = n6282 & ~n6683 ;
  assign n12945 = n7807 & ~n12944 ;
  assign n12946 = \P1_reg1_reg[8]/NET0131  & ~n12945 ;
  assign n12947 = ~n12936 & ~n12946 ;
  assign n12948 = ~n12943 & n12947 ;
  assign n12949 = ~n12940 & n12948 ;
  assign n12950 = n6097 & ~n12949 ;
  assign n12951 = ~n12935 & ~n12950 ;
  assign n12952 = \P1_state_reg[0]/NET0131  & ~n12951 ;
  assign n12953 = ~n12934 & ~n12952 ;
  assign n12954 = n4011 & n11293 ;
  assign n12955 = n9647 & ~n12954 ;
  assign n12956 = \P1_reg2_reg[11]/NET0131  & ~n12955 ;
  assign n12957 = n3250 & n4112 ;
  assign n12958 = n3246 & n6365 ;
  assign n12959 = n11311 & ~n12958 ;
  assign n12960 = ~n12954 & n12959 ;
  assign n12961 = n6113 & ~n12960 ;
  assign n12962 = ~n12957 & ~n12961 ;
  assign n12963 = n9044 & ~n12962 ;
  assign n12964 = ~n12956 & ~n12963 ;
  assign n12965 = n6113 & ~n12050 ;
  assign n12966 = n3349 & n4112 ;
  assign n12967 = ~n12965 & ~n12966 ;
  assign n12968 = n9044 & ~n12967 ;
  assign n12969 = \P1_reg2_reg[13]/NET0131  & ~n9647 ;
  assign n12970 = ~n12968 & ~n12969 ;
  assign n12971 = \P1_reg2_reg[15]/NET0131  & ~n6078 ;
  assign n12972 = \P1_reg2_reg[15]/NET0131  & n6095 ;
  assign n12974 = n3614 & n6365 ;
  assign n12975 = ~n11393 & ~n12974 ;
  assign n12976 = n11382 & n12975 ;
  assign n12977 = n6113 & ~n12976 ;
  assign n12978 = n6113 & n11389 ;
  assign n12979 = ~\P1_reg2_reg[15]/NET0131  & ~n6113 ;
  assign n12980 = n4011 & ~n12979 ;
  assign n12981 = ~n12978 & n12980 ;
  assign n12973 = n3618 & n4112 ;
  assign n12982 = ~n6113 & n6359 ;
  assign n12983 = n8955 & ~n12982 ;
  assign n12984 = ~n10834 & n12983 ;
  assign n12985 = \P1_reg2_reg[15]/NET0131  & ~n12984 ;
  assign n12986 = ~n12973 & ~n12985 ;
  assign n12987 = ~n12981 & n12986 ;
  assign n12988 = ~n12977 & n12987 ;
  assign n12989 = n6097 & ~n12988 ;
  assign n12990 = ~n12972 & ~n12989 ;
  assign n12991 = \P1_state_reg[0]/NET0131  & ~n12990 ;
  assign n12992 = ~n12971 & ~n12991 ;
  assign n12993 = \P2_reg1_reg[12]/NET0131  & ~n5589 ;
  assign n12994 = \P2_reg1_reg[12]/NET0131  & n5585 ;
  assign n12996 = \P2_reg1_reg[12]/NET0131  & ~n6380 ;
  assign n13000 = n6380 & n10385 ;
  assign n13001 = ~n12996 & ~n13000 ;
  assign n13002 = n5383 & ~n13001 ;
  assign n12997 = n6380 & n10375 ;
  assign n12998 = ~n12996 & ~n12997 ;
  assign n12999 = n5329 & ~n12998 ;
  assign n13003 = n6380 & ~n10391 ;
  assign n13004 = ~n12996 & ~n13003 ;
  assign n13005 = n5526 & ~n13004 ;
  assign n12995 = \P2_reg1_reg[12]/NET0131  & ~n6397 ;
  assign n13006 = n6380 & ~n11981 ;
  assign n13007 = ~n12995 & ~n13006 ;
  assign n13008 = ~n13005 & n13007 ;
  assign n13009 = ~n12999 & n13008 ;
  assign n13010 = ~n13002 & n13009 ;
  assign n13011 = n5583 & ~n13010 ;
  assign n13012 = ~n12994 & ~n13011 ;
  assign n13013 = \P1_state_reg[0]/NET0131  & ~n13012 ;
  assign n13014 = ~n12993 & ~n13013 ;
  assign n13015 = \P2_reg1_reg[15]/NET0131  & ~n5589 ;
  assign n13016 = \P2_reg1_reg[15]/NET0131  & n5585 ;
  assign n13019 = \P2_reg1_reg[15]/NET0131  & ~n6380 ;
  assign n13020 = n6380 & n11453 ;
  assign n13021 = ~n13019 & ~n13020 ;
  assign n13022 = n5329 & ~n13021 ;
  assign n13026 = n6380 & n11468 ;
  assign n13027 = ~n13019 & ~n13026 ;
  assign n13028 = n5383 & ~n13027 ;
  assign n13023 = n6380 & ~n11459 ;
  assign n13024 = ~n13019 & ~n13023 ;
  assign n13025 = n5526 & ~n13024 ;
  assign n13029 = n6380 & n11474 ;
  assign n13030 = ~n13019 & ~n13029 ;
  assign n13031 = n5563 & ~n13030 ;
  assign n13017 = n4918 & n5565 ;
  assign n13018 = n6380 & n13017 ;
  assign n13032 = n5565 & ~n6380 ;
  assign n13033 = n6394 & ~n13032 ;
  assign n13034 = \P2_reg1_reg[15]/NET0131  & ~n13033 ;
  assign n13035 = ~n13018 & ~n13034 ;
  assign n13036 = ~n13031 & n13035 ;
  assign n13037 = ~n13025 & n13036 ;
  assign n13038 = ~n13028 & n13037 ;
  assign n13039 = ~n13022 & n13038 ;
  assign n13040 = n5583 & ~n13039 ;
  assign n13041 = ~n13016 & ~n13040 ;
  assign n13042 = \P1_state_reg[0]/NET0131  & ~n13041 ;
  assign n13043 = ~n13015 & ~n13042 ;
  assign n13044 = \P2_reg1_reg[16]/NET0131  & ~n5589 ;
  assign n13045 = \P2_reg1_reg[16]/NET0131  & n5585 ;
  assign n13047 = \P2_reg1_reg[16]/NET0131  & ~n6380 ;
  assign n13048 = n6380 & ~n11497 ;
  assign n13049 = ~n13047 & ~n13048 ;
  assign n13050 = n5329 & ~n13049 ;
  assign n13051 = n6380 & n11505 ;
  assign n13052 = ~n13047 & ~n13051 ;
  assign n13053 = n5383 & ~n13052 ;
  assign n13046 = \P2_reg1_reg[16]/NET0131  & ~n6398 ;
  assign n13055 = n5526 & ~n11511 ;
  assign n13054 = n5563 & n11516 ;
  assign n13056 = n4892 & n5565 ;
  assign n13057 = ~n13054 & ~n13056 ;
  assign n13058 = ~n13055 & n13057 ;
  assign n13059 = n6380 & ~n13058 ;
  assign n13060 = ~n13046 & ~n13059 ;
  assign n13061 = ~n13053 & n13060 ;
  assign n13062 = ~n13050 & n13061 ;
  assign n13063 = n5583 & ~n13062 ;
  assign n13064 = ~n13045 & ~n13063 ;
  assign n13065 = \P1_state_reg[0]/NET0131  & ~n13064 ;
  assign n13066 = ~n13044 & ~n13065 ;
  assign n13067 = \P2_reg2_reg[11]/NET0131  & ~n5589 ;
  assign n13068 = \P2_reg2_reg[11]/NET0131  & n5585 ;
  assign n13070 = \P2_reg2_reg[11]/NET0131  & ~n4219 ;
  assign n13074 = n4219 & n11340 ;
  assign n13075 = ~n13070 & ~n13074 ;
  assign n13076 = n5383 & ~n13075 ;
  assign n13071 = n4219 & n11332 ;
  assign n13072 = ~n13070 & ~n13071 ;
  assign n13073 = n5329 & ~n13072 ;
  assign n13077 = n4219 & ~n11346 ;
  assign n13078 = ~n13070 & ~n13077 ;
  assign n13079 = n5526 & ~n13078 ;
  assign n13081 = n4948 & n5565 ;
  assign n13082 = n5563 & n11351 ;
  assign n13083 = ~n13081 & ~n13082 ;
  assign n13084 = n4219 & ~n13083 ;
  assign n13069 = \P2_reg2_reg[11]/NET0131  & ~n6839 ;
  assign n13080 = n4926 & n5574 ;
  assign n13085 = ~n13069 & ~n13080 ;
  assign n13086 = ~n13084 & n13085 ;
  assign n13087 = ~n13079 & n13086 ;
  assign n13088 = ~n13073 & n13087 ;
  assign n13089 = ~n13076 & n13088 ;
  assign n13090 = n5583 & ~n13089 ;
  assign n13091 = ~n13068 & ~n13090 ;
  assign n13092 = \P1_state_reg[0]/NET0131  & ~n13091 ;
  assign n13093 = ~n13067 & ~n13092 ;
  assign n13094 = \P2_reg2_reg[14]/NET0131  & ~n9773 ;
  assign n13096 = n5383 & n11419 ;
  assign n13095 = n5526 & ~n11411 ;
  assign n13097 = n4843 & n5565 ;
  assign n13098 = ~n13095 & ~n13097 ;
  assign n13099 = n11431 & n13098 ;
  assign n13100 = ~n13096 & n13099 ;
  assign n13101 = n4219 & ~n13100 ;
  assign n13102 = n4821 & n5574 ;
  assign n13103 = ~n13101 & ~n13102 ;
  assign n13104 = n8899 & ~n13103 ;
  assign n13105 = ~n13094 & ~n13104 ;
  assign n13106 = \P2_reg2_reg[15]/NET0131  & ~n5589 ;
  assign n13107 = \P2_reg2_reg[15]/NET0131  & n5585 ;
  assign n13109 = \P2_reg2_reg[15]/NET0131  & ~n4219 ;
  assign n13110 = n4219 & n11453 ;
  assign n13111 = ~n13109 & ~n13110 ;
  assign n13112 = n5329 & ~n13111 ;
  assign n13116 = n4219 & n11468 ;
  assign n13117 = ~n13109 & ~n13116 ;
  assign n13118 = n5383 & ~n13117 ;
  assign n13113 = n4219 & ~n11459 ;
  assign n13114 = ~n13109 & ~n13113 ;
  assign n13115 = n5526 & ~n13114 ;
  assign n13119 = n4219 & n11474 ;
  assign n13120 = ~n13109 & ~n13119 ;
  assign n13121 = n5563 & ~n13120 ;
  assign n13123 = \P2_reg2_reg[15]/NET0131  & ~n5570 ;
  assign n13108 = n4219 & n13017 ;
  assign n13122 = n4898 & n5574 ;
  assign n13124 = ~n13108 & ~n13122 ;
  assign n13125 = ~n13123 & n13124 ;
  assign n13126 = ~n13121 & n13125 ;
  assign n13127 = ~n13115 & n13126 ;
  assign n13128 = ~n13118 & n13127 ;
  assign n13129 = ~n13112 & n13128 ;
  assign n13130 = n5583 & ~n13129 ;
  assign n13131 = ~n13107 & ~n13130 ;
  assign n13132 = \P1_state_reg[0]/NET0131  & ~n13131 ;
  assign n13133 = ~n13106 & ~n13132 ;
  assign n13134 = \P2_reg2_reg[16]/NET0131  & ~n5589 ;
  assign n13135 = \P2_reg2_reg[16]/NET0131  & n5585 ;
  assign n13139 = \P2_reg2_reg[16]/NET0131  & ~n4219 ;
  assign n13140 = n4219 & ~n11497 ;
  assign n13141 = ~n13139 & ~n13140 ;
  assign n13142 = n5329 & ~n13141 ;
  assign n13143 = n4219 & n11505 ;
  assign n13144 = ~n13139 & ~n13143 ;
  assign n13145 = n5383 & ~n13144 ;
  assign n13146 = n4219 & ~n13058 ;
  assign n13136 = n4875 & n5574 ;
  assign n13137 = n6839 & ~n9784 ;
  assign n13138 = \P2_reg2_reg[16]/NET0131  & ~n13137 ;
  assign n13147 = ~n13136 & ~n13138 ;
  assign n13148 = ~n13146 & n13147 ;
  assign n13149 = ~n13145 & n13148 ;
  assign n13150 = ~n13142 & n13149 ;
  assign n13151 = n5583 & ~n13150 ;
  assign n13152 = ~n13135 & ~n13151 ;
  assign n13153 = \P1_state_reg[0]/NET0131  & ~n13152 ;
  assign n13154 = ~n13134 & ~n13153 ;
  assign n13155 = \P1_reg2_reg[8]/NET0131  & ~n6078 ;
  assign n13156 = \P1_reg2_reg[8]/NET0131  & n6095 ;
  assign n13158 = \P1_reg2_reg[8]/NET0131  & ~n6113 ;
  assign n13159 = n6113 & n11540 ;
  assign n13160 = ~n13158 & ~n13159 ;
  assign n13161 = n4011 & ~n13160 ;
  assign n13162 = n6113 & n11546 ;
  assign n13163 = ~n13158 & ~n13162 ;
  assign n13164 = n6207 & ~n13163 ;
  assign n13165 = n6113 & ~n12592 ;
  assign n13157 = n3818 & n4112 ;
  assign n13166 = ~n6113 & n6282 ;
  assign n13167 = n12983 & ~n13166 ;
  assign n13168 = \P1_reg2_reg[8]/NET0131  & ~n13167 ;
  assign n13169 = ~n13157 & ~n13168 ;
  assign n13170 = ~n13165 & n13169 ;
  assign n13171 = ~n13164 & n13170 ;
  assign n13172 = ~n13161 & n13171 ;
  assign n13173 = n6097 & ~n13172 ;
  assign n13174 = ~n13156 & ~n13173 ;
  assign n13175 = \P1_state_reg[0]/NET0131  & ~n13174 ;
  assign n13176 = ~n13155 & ~n13175 ;
  assign n13177 = ~n10008 & n11142 ;
  assign n13178 = n9044 & n13177 ;
  assign n13179 = \P1_reg0_reg[15]/NET0131  & ~n13178 ;
  assign n13180 = ~n11390 & n12976 ;
  assign n13181 = n9829 & ~n13180 ;
  assign n13182 = ~n13179 & ~n13181 ;
  assign n13183 = \P3_reg0_reg[15]/NET0131  & ~n2143 ;
  assign n13184 = \P3_reg0_reg[15]/NET0131  & n2145 ;
  assign n13189 = \P3_reg0_reg[15]/NET0131  & ~n2236 ;
  assign n13192 = n2236 & ~n11592 ;
  assign n13193 = ~n13189 & ~n13192 ;
  assign n13194 = n737 & ~n13193 ;
  assign n13190 = ~n11581 & ~n13189 ;
  assign n13191 = n2393 & ~n13190 ;
  assign n13186 = \P3_reg0_reg[15]/NET0131  & ~n2163 ;
  assign n13187 = ~n11585 & ~n13186 ;
  assign n13188 = n2391 & ~n13187 ;
  assign n13195 = n2163 & n11598 ;
  assign n13196 = ~n13186 & ~n13195 ;
  assign n13197 = n2234 & ~n13196 ;
  assign n13185 = \P3_reg0_reg[15]/NET0131  & ~n2287 ;
  assign n13198 = ~n1512 & n2289 ;
  assign n13199 = ~n13185 & ~n13198 ;
  assign n13200 = ~n13197 & n13199 ;
  assign n13201 = ~n13188 & n13200 ;
  assign n13202 = ~n13191 & n13201 ;
  assign n13203 = ~n13194 & n13202 ;
  assign n13204 = n2147 & ~n13203 ;
  assign n13205 = ~n13184 & ~n13204 ;
  assign n13206 = \P1_state_reg[0]/NET0131  & ~n13205 ;
  assign n13207 = ~n13183 & ~n13206 ;
  assign n13208 = \P3_reg1_reg[15]/NET0131  & ~n2143 ;
  assign n13209 = \P3_reg1_reg[15]/NET0131  & n2145 ;
  assign n13216 = \P3_reg1_reg[15]/NET0131  & ~n2427 ;
  assign n13220 = n2427 & ~n11592 ;
  assign n13221 = ~n13216 & ~n13220 ;
  assign n13222 = n737 & ~n13221 ;
  assign n13211 = \P3_reg1_reg[15]/NET0131  & ~n2408 ;
  assign n13212 = n2408 & ~n11580 ;
  assign n13213 = ~n13211 & ~n13212 ;
  assign n13214 = n714 & ~n13213 ;
  assign n13223 = n2408 & n11598 ;
  assign n13224 = ~n13211 & ~n13223 ;
  assign n13225 = ~n2518 & ~n13224 ;
  assign n13217 = n2427 & n11598 ;
  assign n13218 = ~n13216 & ~n13217 ;
  assign n13219 = n2425 & ~n13218 ;
  assign n13210 = ~n1512 & n6451 ;
  assign n13215 = \P3_reg1_reg[15]/NET0131  & ~n6449 ;
  assign n13226 = ~n13210 & ~n13215 ;
  assign n13227 = ~n13219 & n13226 ;
  assign n13228 = ~n13225 & n13227 ;
  assign n13229 = ~n13214 & n13228 ;
  assign n13230 = ~n13222 & n13229 ;
  assign n13231 = n2147 & ~n13230 ;
  assign n13232 = ~n13209 & ~n13231 ;
  assign n13233 = \P1_state_reg[0]/NET0131  & ~n13232 ;
  assign n13234 = ~n13208 & ~n13233 ;
  assign n13235 = \P1_reg0_reg[9]/NET0131  & ~n6078 ;
  assign n13236 = \P1_reg0_reg[9]/NET0131  & n6095 ;
  assign n13238 = \P1_reg0_reg[9]/NET0131  & ~n6409 ;
  assign n13239 = n6409 & n11733 ;
  assign n13240 = ~n13238 & ~n13239 ;
  assign n13241 = n4011 & ~n13240 ;
  assign n13245 = n6409 & n11739 ;
  assign n13246 = ~n13238 & ~n13245 ;
  assign n13247 = n6207 & ~n13246 ;
  assign n13242 = n6409 & ~n11745 ;
  assign n13243 = ~n13238 & ~n13242 ;
  assign n13244 = n6282 & ~n13243 ;
  assign n13237 = n6409 & ~n11821 ;
  assign n13248 = \P1_reg0_reg[9]/NET0131  & ~n11118 ;
  assign n13249 = ~n13237 & ~n13248 ;
  assign n13250 = ~n13244 & n13249 ;
  assign n13251 = ~n13247 & n13250 ;
  assign n13252 = ~n13241 & n13251 ;
  assign n13253 = n6097 & ~n13252 ;
  assign n13254 = ~n13236 & ~n13253 ;
  assign n13255 = \P1_state_reg[0]/NET0131  & ~n13254 ;
  assign n13256 = ~n13235 & ~n13255 ;
  assign n13257 = \P3_reg2_reg[15]/NET0131  & ~n2143 ;
  assign n13258 = \P3_reg2_reg[15]/NET0131  & n2145 ;
  assign n13264 = \P3_reg2_reg[15]/NET0131  & ~n2408 ;
  assign n13267 = n2408 & ~n11592 ;
  assign n13268 = ~n13264 & ~n13267 ;
  assign n13269 = n737 & ~n13268 ;
  assign n13260 = \P3_reg2_reg[15]/NET0131  & ~n2427 ;
  assign n13261 = n2427 & ~n11580 ;
  assign n13262 = ~n13260 & ~n13261 ;
  assign n13263 = n714 & ~n13262 ;
  assign n13270 = ~n13217 & ~n13260 ;
  assign n13271 = ~n2518 & ~n13270 ;
  assign n13265 = ~n13223 & ~n13264 ;
  assign n13266 = n2425 & ~n13265 ;
  assign n13259 = ~n1512 & n2441 ;
  assign n13272 = ~n1514 & n2283 ;
  assign n13273 = \P3_reg2_reg[15]/NET0131  & ~n2429 ;
  assign n13274 = ~n13272 & ~n13273 ;
  assign n13275 = ~n13259 & n13274 ;
  assign n13276 = ~n13266 & n13275 ;
  assign n13277 = ~n13271 & n13276 ;
  assign n13278 = ~n13263 & n13277 ;
  assign n13279 = ~n13269 & n13278 ;
  assign n13280 = n2147 & ~n13279 ;
  assign n13281 = ~n13258 & ~n13280 ;
  assign n13282 = \P1_state_reg[0]/NET0131  & ~n13281 ;
  assign n13283 = ~n13257 & ~n13282 ;
  assign n13284 = \P1_reg1_reg[10]/NET0131  & ~n6078 ;
  assign n13285 = \P1_reg1_reg[10]/NET0131  & n6095 ;
  assign n13287 = \P1_reg1_reg[10]/NET0131  & ~n6683 ;
  assign n13294 = n6683 & n11661 ;
  assign n13295 = ~n13287 & ~n13294 ;
  assign n13296 = n4011 & ~n13295 ;
  assign n13291 = n6683 & n11667 ;
  assign n13292 = ~n13287 & ~n13291 ;
  assign n13293 = n6207 & ~n13292 ;
  assign n13288 = n6683 & ~n11673 ;
  assign n13289 = ~n13287 & ~n13288 ;
  assign n13290 = n6282 & ~n13289 ;
  assign n13297 = n6683 & n11678 ;
  assign n13298 = ~n13287 & ~n13297 ;
  assign n13299 = n6359 & ~n13298 ;
  assign n13286 = \P1_reg1_reg[10]/NET0131  & ~n7806 ;
  assign n13300 = n6683 & n11790 ;
  assign n13301 = ~n13286 & ~n13300 ;
  assign n13302 = ~n13299 & n13301 ;
  assign n13303 = ~n13290 & n13302 ;
  assign n13304 = ~n13293 & n13303 ;
  assign n13305 = ~n13296 & n13304 ;
  assign n13306 = n6097 & ~n13305 ;
  assign n13307 = ~n13285 & ~n13306 ;
  assign n13308 = \P1_state_reg[0]/NET0131  & ~n13307 ;
  assign n13309 = ~n13284 & ~n13308 ;
  assign n13310 = n9045 & ~n13180 ;
  assign n13311 = n6695 & n12611 ;
  assign n13312 = \P1_reg1_reg[15]/NET0131  & ~n13311 ;
  assign n13313 = ~n13310 & ~n13312 ;
  assign n13314 = \P2_reg0_reg[12]/NET0131  & ~n5589 ;
  assign n13315 = \P2_reg0_reg[12]/NET0131  & n5585 ;
  assign n13317 = \P2_reg0_reg[12]/NET0131  & ~n6706 ;
  assign n13321 = n6706 & n10385 ;
  assign n13322 = ~n13317 & ~n13321 ;
  assign n13323 = n5383 & ~n13322 ;
  assign n13318 = n6706 & n10375 ;
  assign n13319 = ~n13317 & ~n13318 ;
  assign n13320 = n5329 & ~n13319 ;
  assign n13324 = n6706 & ~n10391 ;
  assign n13325 = ~n13317 & ~n13324 ;
  assign n13326 = n5526 & ~n13325 ;
  assign n13316 = \P2_reg0_reg[12]/NET0131  & ~n6717 ;
  assign n13327 = n6706 & ~n11981 ;
  assign n13328 = ~n13316 & ~n13327 ;
  assign n13329 = ~n13326 & n13328 ;
  assign n13330 = ~n13320 & n13329 ;
  assign n13331 = ~n13323 & n13330 ;
  assign n13332 = n5583 & ~n13331 ;
  assign n13333 = ~n13315 & ~n13332 ;
  assign n13334 = \P1_state_reg[0]/NET0131  & ~n13333 ;
  assign n13335 = ~n13314 & ~n13334 ;
  assign n13336 = \P2_reg0_reg[15]/NET0131  & ~n5589 ;
  assign n13337 = \P2_reg0_reg[15]/NET0131  & n5585 ;
  assign n13339 = \P2_reg0_reg[15]/NET0131  & ~n6706 ;
  assign n13340 = n6706 & n11453 ;
  assign n13341 = ~n13339 & ~n13340 ;
  assign n13342 = n5329 & ~n13341 ;
  assign n13346 = n6706 & n11468 ;
  assign n13347 = ~n13339 & ~n13346 ;
  assign n13348 = n5383 & ~n13347 ;
  assign n13343 = n6706 & ~n11459 ;
  assign n13344 = ~n13339 & ~n13343 ;
  assign n13345 = n5526 & ~n13344 ;
  assign n13349 = n6706 & n11474 ;
  assign n13350 = ~n13339 & ~n13349 ;
  assign n13351 = n5563 & ~n13350 ;
  assign n13338 = n6706 & n13017 ;
  assign n13352 = \P2_reg0_reg[15]/NET0131  & ~n7864 ;
  assign n13353 = ~n13338 & ~n13352 ;
  assign n13354 = ~n13351 & n13353 ;
  assign n13355 = ~n13345 & n13354 ;
  assign n13356 = ~n13348 & n13355 ;
  assign n13357 = ~n13342 & n13356 ;
  assign n13358 = n5583 & ~n13357 ;
  assign n13359 = ~n13337 & ~n13358 ;
  assign n13360 = \P1_state_reg[0]/NET0131  & ~n13359 ;
  assign n13361 = ~n13336 & ~n13360 ;
  assign n13362 = \P2_reg0_reg[16]/NET0131  & ~n5589 ;
  assign n13363 = \P2_reg0_reg[16]/NET0131  & n5585 ;
  assign n13365 = \P2_reg0_reg[16]/NET0131  & ~n6706 ;
  assign n13366 = n6706 & ~n11497 ;
  assign n13367 = ~n13365 & ~n13366 ;
  assign n13368 = n5329 & ~n13367 ;
  assign n13369 = n6706 & n11505 ;
  assign n13370 = ~n13365 & ~n13369 ;
  assign n13371 = n5383 & ~n13370 ;
  assign n13364 = \P2_reg0_reg[16]/NET0131  & ~n6718 ;
  assign n13372 = n6706 & ~n13058 ;
  assign n13373 = ~n13364 & ~n13372 ;
  assign n13374 = ~n13371 & n13373 ;
  assign n13375 = ~n13368 & n13374 ;
  assign n13376 = n5583 & ~n13375 ;
  assign n13377 = ~n13363 & ~n13376 ;
  assign n13378 = \P1_state_reg[0]/NET0131  & ~n13377 ;
  assign n13379 = ~n13362 & ~n13378 ;
  assign n13382 = n5088 & n5585 ;
  assign n13384 = n5088 & ~n7453 ;
  assign n13385 = n5068 & ~n5352 ;
  assign n13386 = ~n5353 & ~n13385 ;
  assign n13387 = ~n4231 & ~n13386 ;
  assign n13388 = n4231 & n5117 ;
  assign n13389 = ~n13387 & ~n13388 ;
  assign n13390 = n7453 & n13389 ;
  assign n13391 = ~n13384 & ~n13390 ;
  assign n13392 = n5383 & ~n13391 ;
  assign n13399 = n5981 & ~n6740 ;
  assign n13400 = ~n5981 & n6740 ;
  assign n13401 = ~n13399 & ~n13400 ;
  assign n13402 = n7453 & ~n13401 ;
  assign n13403 = ~n13384 & ~n13402 ;
  assign n13404 = n5329 & ~n13403 ;
  assign n13393 = n5981 & ~n7913 ;
  assign n13394 = ~n5981 & n7913 ;
  assign n13395 = ~n13393 & ~n13394 ;
  assign n13396 = n7453 & n13395 ;
  assign n13397 = ~n13384 & ~n13396 ;
  assign n13398 = n5526 & ~n13397 ;
  assign n13405 = ~n5107 & ~n12699 ;
  assign n13406 = ~n5534 & n5563 ;
  assign n13407 = ~n13405 & n13406 ;
  assign n13408 = n7453 & n13407 ;
  assign n13383 = n5088 & ~n7484 ;
  assign n13409 = ~n5107 & ~n7504 ;
  assign n13410 = ~n13383 & ~n13409 ;
  assign n13411 = ~n13408 & n13410 ;
  assign n13412 = ~n13398 & n13411 ;
  assign n13413 = ~n13404 & n13412 ;
  assign n13414 = ~n13392 & n13413 ;
  assign n13415 = n5583 & ~n13414 ;
  assign n13416 = ~n13382 & ~n13415 ;
  assign n13417 = \P1_state_reg[0]/NET0131  & ~n13416 ;
  assign n13380 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[6]/NET0131  ;
  assign n13381 = n5088 & n5786 ;
  assign n13418 = ~n13380 & ~n13381 ;
  assign n13419 = ~n13417 & n13418 ;
  assign n13421 = n5063 & n5585 ;
  assign n13423 = n5040 & ~n5353 ;
  assign n13424 = ~n10328 & ~n13423 ;
  assign n13425 = ~n4231 & ~n13424 ;
  assign n13426 = n4231 & n5092 ;
  assign n13427 = n5383 & ~n13426 ;
  assign n13428 = ~n13425 & n13427 ;
  assign n13438 = n5980 & ~n7553 ;
  assign n13437 = ~n5980 & n7553 ;
  assign n13439 = n5329 & ~n13437 ;
  assign n13440 = ~n13438 & n13439 ;
  assign n13430 = n5980 & n7519 ;
  assign n13429 = ~n5980 & ~n7519 ;
  assign n13431 = n5526 & ~n13429 ;
  assign n13432 = ~n13430 & n13431 ;
  assign n13434 = ~n5081 & ~n5534 ;
  assign n13433 = n5081 & n5534 ;
  assign n13435 = n5563 & ~n13433 ;
  assign n13436 = ~n13434 & n13435 ;
  assign n13441 = ~n13432 & ~n13436 ;
  assign n13442 = ~n13440 & n13441 ;
  assign n13443 = ~n13428 & n13442 ;
  assign n13444 = n7453 & ~n13443 ;
  assign n13422 = ~n5081 & ~n7504 ;
  assign n13445 = ~n5329 & n7866 ;
  assign n13446 = ~n7453 & ~n13445 ;
  assign n13447 = n7641 & ~n13446 ;
  assign n13448 = n5063 & ~n13447 ;
  assign n13449 = ~n13422 & ~n13448 ;
  assign n13450 = ~n13444 & n13449 ;
  assign n13451 = n5583 & ~n13450 ;
  assign n13452 = ~n13421 & ~n13451 ;
  assign n13453 = \P1_state_reg[0]/NET0131  & ~n13452 ;
  assign n13420 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[7]/NET0131  ;
  assign n13454 = n5063 & n5786 ;
  assign n13455 = ~n13420 & ~n13454 ;
  assign n13456 = ~n13453 & n13455 ;
  assign n13459 = n5033 & n5585 ;
  assign n13462 = n5033 & ~n13445 ;
  assign n13463 = ~n7453 & ~n13462 ;
  assign n13472 = n5008 & ~n10328 ;
  assign n13473 = ~n10329 & ~n13472 ;
  assign n13474 = ~n4231 & ~n13473 ;
  assign n13475 = n4231 & n5068 ;
  assign n13476 = ~n13474 & ~n13475 ;
  assign n13477 = n5383 & n13476 ;
  assign n13464 = ~n5058 & ~n13433 ;
  assign n13465 = ~n5536 & n5563 ;
  assign n13466 = ~n13464 & n13465 ;
  assign n13468 = n5993 & ~n6744 ;
  assign n13467 = ~n5993 & n6744 ;
  assign n13469 = n5329 & ~n13467 ;
  assign n13470 = ~n13468 & n13469 ;
  assign n13471 = ~n13466 & ~n13470 ;
  assign n13479 = n5824 & n5993 ;
  assign n13478 = ~n5824 & ~n5993 ;
  assign n13480 = n5526 & ~n13478 ;
  assign n13481 = ~n13479 & n13480 ;
  assign n13482 = n7453 & ~n13481 ;
  assign n13483 = n13471 & n13482 ;
  assign n13484 = ~n13477 & n13483 ;
  assign n13485 = ~n13463 & ~n13484 ;
  assign n13460 = ~n5058 & ~n7504 ;
  assign n13461 = n5033 & ~n7641 ;
  assign n13486 = ~n13460 & ~n13461 ;
  assign n13487 = ~n13485 & n13486 ;
  assign n13488 = n5583 & ~n13487 ;
  assign n13489 = ~n13459 & ~n13488 ;
  assign n13490 = \P1_state_reg[0]/NET0131  & ~n13489 ;
  assign n13457 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[8]/NET0131  ;
  assign n13458 = n5033 & n5786 ;
  assign n13491 = ~n13457 & ~n13458 ;
  assign n13492 = ~n13490 & n13491 ;
  assign n13495 = ~\P1_reg3_reg[3]/NET0131  & n6095 ;
  assign n13502 = ~\P1_reg3_reg[3]/NET0131  & ~n6568 ;
  assign n13503 = n3795 & ~n6288 ;
  assign n13504 = ~n12735 & ~n13503 ;
  assign n13505 = ~n2713 & ~n13504 ;
  assign n13506 = n2713 & n3364 ;
  assign n13507 = ~n13505 & ~n13506 ;
  assign n13508 = n6568 & n13507 ;
  assign n13509 = ~n13502 & ~n13508 ;
  assign n13510 = n4011 & ~n13509 ;
  assign n13517 = n3773 & ~n6214 ;
  assign n13518 = ~n3773 & n6214 ;
  assign n13519 = ~n13517 & ~n13518 ;
  assign n13520 = n6568 & n13519 ;
  assign n13521 = ~n13502 & ~n13520 ;
  assign n13522 = n6282 & ~n13521 ;
  assign n13511 = n3773 & n6140 ;
  assign n13512 = ~n3773 & ~n6140 ;
  assign n13513 = ~n13511 & ~n13512 ;
  assign n13514 = n6568 & n13513 ;
  assign n13515 = ~n13502 & ~n13514 ;
  assign n13516 = n6207 & ~n13515 ;
  assign n13496 = ~n3770 & n6365 ;
  assign n13497 = ~n3770 & ~n6329 ;
  assign n13498 = ~n6330 & n6359 ;
  assign n13499 = ~n13497 & n13498 ;
  assign n13500 = ~n13496 & ~n13499 ;
  assign n13501 = n6568 & ~n13500 ;
  assign n13523 = ~n3770 & n4112 ;
  assign n13524 = ~\P1_reg3_reg[3]/NET0131  & ~n12757 ;
  assign n13525 = ~n13523 & ~n13524 ;
  assign n13526 = ~n13501 & n13525 ;
  assign n13527 = ~n13516 & n13526 ;
  assign n13528 = ~n13522 & n13527 ;
  assign n13529 = ~n13510 & n13528 ;
  assign n13530 = n6097 & ~n13529 ;
  assign n13531 = ~n13495 & ~n13530 ;
  assign n13532 = \P1_state_reg[0]/NET0131  & ~n13531 ;
  assign n13493 = \P1_reg3_reg[3]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n13494 = ~\P1_reg3_reg[3]/NET0131  & n4130 ;
  assign n13533 = ~n13493 & ~n13494 ;
  assign n13534 = ~n13532 & n13533 ;
  assign n13537 = n3739 & n6095 ;
  assign n13544 = n3739 & ~n6568 ;
  assign n13545 = n3577 & ~n6291 ;
  assign n13546 = ~n3577 & n6291 ;
  assign n13547 = ~n13545 & ~n13546 ;
  assign n13548 = ~n2713 & ~n13547 ;
  assign n13549 = n2713 & n3137 ;
  assign n13550 = ~n13548 & ~n13549 ;
  assign n13551 = n6568 & n13550 ;
  assign n13552 = ~n13544 & ~n13551 ;
  assign n13553 = n4011 & ~n13552 ;
  assign n13560 = n3749 & ~n7127 ;
  assign n13561 = ~n3749 & n7127 ;
  assign n13562 = ~n13560 & ~n13561 ;
  assign n13563 = n6568 & ~n13562 ;
  assign n13564 = ~n13544 & ~n13563 ;
  assign n13565 = n6282 & ~n13564 ;
  assign n13554 = n3749 & ~n7169 ;
  assign n13555 = ~n3749 & n7169 ;
  assign n13556 = ~n13554 & ~n13555 ;
  assign n13557 = n6568 & n13556 ;
  assign n13558 = ~n13544 & ~n13557 ;
  assign n13559 = n6207 & ~n13558 ;
  assign n13538 = n3737 & n6365 ;
  assign n13539 = n3737 & ~n6332 ;
  assign n13540 = ~n6333 & ~n13539 ;
  assign n13541 = n6359 & n13540 ;
  assign n13542 = ~n13538 & ~n13541 ;
  assign n13543 = n6568 & ~n13542 ;
  assign n13566 = n3737 & n4112 ;
  assign n13567 = n3739 & ~n12757 ;
  assign n13568 = ~n13566 & ~n13567 ;
  assign n13569 = ~n13543 & n13568 ;
  assign n13570 = ~n13559 & n13569 ;
  assign n13571 = ~n13565 & n13570 ;
  assign n13572 = ~n13553 & n13571 ;
  assign n13573 = n6097 & ~n13572 ;
  assign n13574 = ~n13537 & ~n13573 ;
  assign n13575 = \P1_state_reg[0]/NET0131  & ~n13574 ;
  assign n13535 = \P1_reg3_reg[6]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n13536 = n3739 & n4130 ;
  assign n13576 = ~n13535 & ~n13536 ;
  assign n13577 = ~n13575 & n13576 ;
  assign n13580 = n3573 & n6095 ;
  assign n13587 = n3573 & ~n6568 ;
  assign n13588 = n2713 & ~n3746 ;
  assign n13589 = n3822 & ~n13546 ;
  assign n13590 = ~n2713 & ~n6293 ;
  assign n13591 = ~n13589 & n13590 ;
  assign n13592 = ~n13588 & ~n13591 ;
  assign n13593 = n6568 & ~n13592 ;
  assign n13594 = ~n13587 & ~n13593 ;
  assign n13595 = n4011 & ~n13594 ;
  assign n13602 = n3580 & ~n6574 ;
  assign n13603 = ~n3580 & n6574 ;
  assign n13604 = ~n13602 & ~n13603 ;
  assign n13605 = n6568 & ~n13604 ;
  assign n13606 = ~n13587 & ~n13605 ;
  assign n13607 = n6282 & ~n13606 ;
  assign n13596 = n3580 & ~n6612 ;
  assign n13597 = ~n3580 & n6612 ;
  assign n13598 = ~n13596 & ~n13597 ;
  assign n13599 = n6568 & n13598 ;
  assign n13600 = ~n13587 & ~n13599 ;
  assign n13601 = n6207 & ~n13600 ;
  assign n13581 = n3568 & n6365 ;
  assign n13582 = n3568 & ~n6333 ;
  assign n13583 = ~n6334 & ~n13582 ;
  assign n13584 = n6359 & n13583 ;
  assign n13585 = ~n13581 & ~n13584 ;
  assign n13586 = n6568 & ~n13585 ;
  assign n13608 = n3568 & n4112 ;
  assign n13609 = n3573 & ~n12757 ;
  assign n13610 = ~n13608 & ~n13609 ;
  assign n13611 = ~n13586 & n13610 ;
  assign n13612 = ~n13601 & n13611 ;
  assign n13613 = ~n13607 & n13612 ;
  assign n13614 = ~n13595 & n13613 ;
  assign n13615 = n6097 & ~n13614 ;
  assign n13616 = ~n13580 & ~n13615 ;
  assign n13617 = \P1_state_reg[0]/NET0131  & ~n13616 ;
  assign n13578 = \P1_reg3_reg[7]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n13579 = n3573 & n4130 ;
  assign n13618 = ~n13578 & ~n13579 ;
  assign n13619 = ~n13617 & n13618 ;
  assign n13622 = ~n1801 & n2145 ;
  assign n13624 = ~n1801 & ~n2163 ;
  assign n13639 = ~n1852 & n2239 ;
  assign n13640 = ~n1806 & n2246 ;
  assign n13641 = n1779 & ~n13640 ;
  assign n13642 = ~n2239 & ~n2248 ;
  assign n13643 = ~n13641 & n13642 ;
  assign n13644 = ~n13639 & ~n13643 ;
  assign n13645 = n2163 & ~n13644 ;
  assign n13646 = ~n13624 & ~n13645 ;
  assign n13647 = n737 & ~n13646 ;
  assign n13625 = ~n1821 & ~n1916 ;
  assign n13626 = ~n2454 & n13625 ;
  assign n13627 = n2454 & ~n13625 ;
  assign n13628 = ~n13626 & ~n13627 ;
  assign n13632 = n2391 & ~n13628 ;
  assign n13633 = ~n1971 & n13625 ;
  assign n13634 = n1971 & ~n13625 ;
  assign n13635 = ~n13633 & ~n13634 ;
  assign n13636 = n2234 & n13635 ;
  assign n13637 = ~n13632 & ~n13636 ;
  assign n13638 = n2236 & ~n13637 ;
  assign n13629 = n2163 & ~n13628 ;
  assign n13630 = ~n13624 & ~n13629 ;
  assign n13631 = n2393 & ~n13630 ;
  assign n13623 = ~n1820 & n2580 ;
  assign n13648 = ~n2236 & ~n12212 ;
  assign n13649 = n2583 & ~n13648 ;
  assign n13650 = ~n1801 & ~n13649 ;
  assign n13651 = ~n13623 & ~n13650 ;
  assign n13652 = ~n13631 & n13651 ;
  assign n13653 = ~n13638 & n13652 ;
  assign n13654 = ~n13647 & n13653 ;
  assign n13655 = n2147 & ~n13654 ;
  assign n13656 = ~n13622 & ~n13655 ;
  assign n13657 = \P1_state_reg[0]/NET0131  & ~n13656 ;
  assign n13620 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[4]/NET0131  ;
  assign n13621 = n765 & ~n1801 ;
  assign n13658 = ~n13620 & ~n13621 ;
  assign n13659 = ~n13657 & n13658 ;
  assign n13660 = \P1_reg2_reg[5]/NET0131  & ~n6078 ;
  assign n13661 = \P1_reg2_reg[5]/NET0131  & n6095 ;
  assign n13663 = \P1_reg2_reg[5]/NET0131  & ~n6113 ;
  assign n13664 = n6113 & n12781 ;
  assign n13665 = ~n13663 & ~n13664 ;
  assign n13666 = n6207 & ~n13665 ;
  assign n13662 = n6113 & ~n12776 ;
  assign n13673 = n3133 & n4112 ;
  assign n13674 = \P1_reg2_reg[5]/NET0131  & ~n11834 ;
  assign n13675 = ~n13673 & ~n13674 ;
  assign n13676 = ~n13662 & n13675 ;
  assign n13677 = ~n13666 & n13676 ;
  assign n13667 = n6113 & n12789 ;
  assign n13668 = ~n13663 & ~n13667 ;
  assign n13669 = n4011 & ~n13668 ;
  assign n13670 = n6113 & ~n12795 ;
  assign n13671 = ~n13663 & ~n13670 ;
  assign n13672 = n6282 & ~n13671 ;
  assign n13678 = ~n13669 & ~n13672 ;
  assign n13679 = n13677 & n13678 ;
  assign n13680 = n6097 & ~n13679 ;
  assign n13681 = ~n13661 & ~n13680 ;
  assign n13682 = \P1_state_reg[0]/NET0131  & ~n13681 ;
  assign n13683 = ~n13660 & ~n13682 ;
  assign n13684 = \P1_reg1_reg[4]/NET0131  & ~n6078 ;
  assign n13685 = \P1_reg1_reg[4]/NET0131  & n6095 ;
  assign n13687 = \P1_reg1_reg[4]/NET0131  & ~n6683 ;
  assign n13688 = n6683 & ~n12739 ;
  assign n13689 = ~n13687 & ~n13688 ;
  assign n13690 = n4011 & ~n13689 ;
  assign n13694 = n6683 & ~n12745 ;
  assign n13695 = ~n13687 & ~n13694 ;
  assign n13696 = n6207 & ~n13695 ;
  assign n13691 = n6683 & n12751 ;
  assign n13692 = ~n13687 & ~n13691 ;
  assign n13693 = n6282 & ~n13692 ;
  assign n13686 = n6683 & ~n12731 ;
  assign n13697 = \P1_reg1_reg[4]/NET0131  & ~n6695 ;
  assign n13698 = ~n13686 & ~n13697 ;
  assign n13699 = ~n13693 & n13698 ;
  assign n13700 = ~n13696 & n13699 ;
  assign n13701 = ~n13690 & n13700 ;
  assign n13702 = n6097 & ~n13701 ;
  assign n13703 = ~n13685 & ~n13702 ;
  assign n13704 = \P1_state_reg[0]/NET0131  & ~n13703 ;
  assign n13705 = ~n13684 & ~n13704 ;
  assign n13706 = \P1_reg1_reg[5]/NET0131  & ~n6078 ;
  assign n13707 = \P1_reg1_reg[5]/NET0131  & n6095 ;
  assign n13709 = \P1_reg1_reg[5]/NET0131  & ~n6683 ;
  assign n13710 = n6683 & n12781 ;
  assign n13711 = ~n13709 & ~n13710 ;
  assign n13712 = n6207 & ~n13711 ;
  assign n13708 = n6683 & ~n12776 ;
  assign n13719 = \P1_reg1_reg[5]/NET0131  & ~n6695 ;
  assign n13720 = ~n13708 & ~n13719 ;
  assign n13721 = ~n13712 & n13720 ;
  assign n13713 = n6683 & n12789 ;
  assign n13714 = ~n13709 & ~n13713 ;
  assign n13715 = n4011 & ~n13714 ;
  assign n13716 = n6683 & ~n12795 ;
  assign n13717 = ~n13709 & ~n13716 ;
  assign n13718 = n6282 & ~n13717 ;
  assign n13722 = ~n13715 & ~n13718 ;
  assign n13723 = n13721 & n13722 ;
  assign n13724 = n6097 & ~n13723 ;
  assign n13725 = ~n13707 & ~n13724 ;
  assign n13726 = \P1_state_reg[0]/NET0131  & ~n13725 ;
  assign n13727 = ~n13706 & ~n13726 ;
  assign n13728 = n5131 & n5565 ;
  assign n13729 = n12712 & ~n13728 ;
  assign n13730 = ~n12698 & n13729 ;
  assign n13731 = n9533 & ~n13730 ;
  assign n13732 = n8887 & n8899 ;
  assign n13733 = \P2_reg0_reg[5]/NET0131  & ~n13732 ;
  assign n13734 = ~n13731 & ~n13733 ;
  assign n13735 = n4011 & n12659 ;
  assign n13736 = n3219 & n6365 ;
  assign n13737 = ~n13735 & ~n13736 ;
  assign n13738 = n12676 & n13737 ;
  assign n13739 = n6113 & ~n13738 ;
  assign n13740 = n3223 & n4112 ;
  assign n13741 = ~n13739 & ~n13740 ;
  assign n13742 = n9044 & ~n13741 ;
  assign n13743 = \P1_reg2_reg[14]/NET0131  & ~n9647 ;
  assign n13744 = ~n13742 & ~n13743 ;
  assign n13745 = \P2_reg1_reg[11]/NET0131  & ~n5589 ;
  assign n13746 = \P2_reg1_reg[11]/NET0131  & n5585 ;
  assign n13748 = \P2_reg1_reg[11]/NET0131  & ~n6380 ;
  assign n13752 = n6380 & n11340 ;
  assign n13753 = ~n13748 & ~n13752 ;
  assign n13754 = n5383 & ~n13753 ;
  assign n13749 = n6380 & n11332 ;
  assign n13750 = ~n13748 & ~n13749 ;
  assign n13751 = n5329 & ~n13750 ;
  assign n13755 = n6380 & ~n11346 ;
  assign n13756 = ~n13748 & ~n13755 ;
  assign n13757 = n5526 & ~n13756 ;
  assign n13747 = \P2_reg1_reg[11]/NET0131  & ~n6397 ;
  assign n13758 = n6380 & ~n13083 ;
  assign n13759 = ~n13747 & ~n13758 ;
  assign n13760 = ~n13757 & n13759 ;
  assign n13761 = ~n13751 & n13760 ;
  assign n13762 = ~n13754 & n13761 ;
  assign n13763 = n5583 & ~n13762 ;
  assign n13764 = ~n13746 & ~n13763 ;
  assign n13765 = \P1_state_reg[0]/NET0131  & ~n13764 ;
  assign n13766 = ~n13745 & ~n13765 ;
  assign n13767 = \P2_reg1_reg[14]/NET0131  & ~n8902 ;
  assign n13768 = n8913 & ~n13100 ;
  assign n13769 = ~n13767 & ~n13768 ;
  assign n13772 = \P2_reg1_reg[5]/NET0131  & ~n6380 ;
  assign n13773 = n8913 & n12697 ;
  assign n13774 = ~n13772 & ~n13773 ;
  assign n13775 = n5383 & ~n13774 ;
  assign n13770 = \P2_reg1_reg[5]/NET0131  & ~n8901 ;
  assign n13771 = n8913 & ~n13729 ;
  assign n13776 = ~n13770 & ~n13771 ;
  assign n13777 = ~n13775 & n13776 ;
  assign n13778 = \P1_reg2_reg[4]/NET0131  & ~n6078 ;
  assign n13779 = \P1_reg2_reg[4]/NET0131  & n6095 ;
  assign n13781 = \P1_reg2_reg[4]/NET0131  & ~n6113 ;
  assign n13782 = n6113 & ~n12739 ;
  assign n13783 = ~n13781 & ~n13782 ;
  assign n13784 = n4011 & ~n13783 ;
  assign n13788 = n6113 & n12751 ;
  assign n13789 = ~n13781 & ~n13788 ;
  assign n13790 = n6282 & ~n13789 ;
  assign n13785 = n6113 & ~n12745 ;
  assign n13786 = ~n13781 & ~n13785 ;
  assign n13787 = n6207 & ~n13786 ;
  assign n13780 = n6113 & ~n12731 ;
  assign n13791 = n3791 & n4112 ;
  assign n13792 = \P1_reg2_reg[4]/NET0131  & ~n11834 ;
  assign n13793 = ~n13791 & ~n13792 ;
  assign n13794 = ~n13780 & n13793 ;
  assign n13795 = ~n13787 & n13794 ;
  assign n13796 = ~n13790 & n13795 ;
  assign n13797 = ~n13784 & n13796 ;
  assign n13798 = n6097 & ~n13797 ;
  assign n13799 = ~n13779 & ~n13798 ;
  assign n13800 = \P1_state_reg[0]/NET0131  & ~n13799 ;
  assign n13801 = ~n13778 & ~n13800 ;
  assign n13802 = ~\P2_reg2_reg[5]/NET0131  & ~n8899 ;
  assign n13805 = n4219 & ~n12697 ;
  assign n13806 = n5383 & ~n13805 ;
  assign n13807 = n8899 & n9771 ;
  assign n13808 = ~n13806 & n13807 ;
  assign n13809 = \P2_reg2_reg[5]/NET0131  & ~n13808 ;
  assign n13803 = n5110 & n5574 ;
  assign n13804 = n4219 & ~n13730 ;
  assign n13810 = ~n13803 & ~n13804 ;
  assign n13811 = ~n13809 & n13810 ;
  assign n13812 = ~n13802 & ~n13811 ;
  assign n13813 = \P1_reg0_reg[11]/NET0131  & ~n9826 ;
  assign n13814 = n9829 & ~n12960 ;
  assign n13815 = ~n13813 & ~n13814 ;
  assign n13816 = \P1_reg0_reg[14]/NET0131  & ~n9826 ;
  assign n13817 = n9829 & ~n13738 ;
  assign n13818 = ~n13816 & ~n13817 ;
  assign n13819 = \P3_reg0_reg[5]/NET0131  & ~n2143 ;
  assign n13820 = \P3_reg0_reg[5]/NET0131  & n2145 ;
  assign n13822 = \P3_reg0_reg[5]/NET0131  & ~n2236 ;
  assign n13823 = n2236 & ~n12832 ;
  assign n13824 = ~n13822 & ~n13823 ;
  assign n13825 = n737 & ~n13824 ;
  assign n13828 = n2391 & ~n12819 ;
  assign n13829 = n2234 & n12838 ;
  assign n13830 = ~n1794 & n2285 ;
  assign n13831 = ~n13829 & ~n13830 ;
  assign n13832 = ~n13828 & n13831 ;
  assign n13833 = n2163 & ~n13832 ;
  assign n13821 = \P3_reg0_reg[5]/NET0131  & ~n12214 ;
  assign n13826 = ~n12820 & ~n13822 ;
  assign n13827 = n2393 & ~n13826 ;
  assign n13834 = ~n13821 & ~n13827 ;
  assign n13835 = ~n13833 & n13834 ;
  assign n13836 = ~n13825 & n13835 ;
  assign n13837 = n2147 & ~n13836 ;
  assign n13838 = ~n13820 & ~n13837 ;
  assign n13839 = \P1_state_reg[0]/NET0131  & ~n13838 ;
  assign n13840 = ~n13819 & ~n13839 ;
  assign n13841 = \P3_reg0_reg[6]/NET0131  & ~n2143 ;
  assign n13842 = \P3_reg0_reg[6]/NET0131  & n2145 ;
  assign n13844 = \P3_reg0_reg[6]/NET0131  & ~n2236 ;
  assign n13845 = n2236 & ~n12877 ;
  assign n13846 = ~n13844 & ~n13845 ;
  assign n13847 = n737 & ~n13846 ;
  assign n13851 = n2234 & n12868 ;
  assign n13850 = n2391 & ~n12860 ;
  assign n13852 = ~n1768 & n2285 ;
  assign n13853 = ~n13850 & ~n13852 ;
  assign n13854 = ~n13851 & n13853 ;
  assign n13855 = n2163 & ~n13854 ;
  assign n13843 = \P3_reg0_reg[6]/NET0131  & ~n12214 ;
  assign n13848 = ~n12881 & ~n13844 ;
  assign n13849 = n2393 & ~n13848 ;
  assign n13856 = ~n13843 & ~n13849 ;
  assign n13857 = ~n13855 & n13856 ;
  assign n13858 = ~n13847 & n13857 ;
  assign n13859 = n2147 & ~n13858 ;
  assign n13860 = ~n13842 & ~n13859 ;
  assign n13861 = \P1_state_reg[0]/NET0131  & ~n13860 ;
  assign n13862 = ~n13841 & ~n13861 ;
  assign n13863 = \P3_reg0_reg[7]/NET0131  & ~n2143 ;
  assign n13864 = \P3_reg0_reg[7]/NET0131  & n2145 ;
  assign n13867 = \P3_reg0_reg[7]/NET0131  & ~n2236 ;
  assign n13873 = n2236 & ~n12913 ;
  assign n13874 = ~n13867 & ~n13873 ;
  assign n13875 = n737 & ~n13874 ;
  assign n13870 = \P3_reg0_reg[7]/NET0131  & ~n2163 ;
  assign n13871 = ~n12906 & ~n13870 ;
  assign n13872 = n2391 & ~n13871 ;
  assign n13868 = ~n12902 & ~n13867 ;
  assign n13869 = n2393 & ~n13868 ;
  assign n13876 = n2163 & ~n12919 ;
  assign n13877 = ~n13870 & ~n13876 ;
  assign n13878 = n2234 & ~n13877 ;
  assign n13865 = ~n1744 & n2285 ;
  assign n13866 = n2163 & n13865 ;
  assign n13879 = \P3_reg0_reg[7]/NET0131  & ~n2287 ;
  assign n13880 = ~n13866 & ~n13879 ;
  assign n13881 = ~n13878 & n13880 ;
  assign n13882 = ~n13869 & n13881 ;
  assign n13883 = ~n13872 & n13882 ;
  assign n13884 = ~n13875 & n13883 ;
  assign n13885 = n2147 & ~n13884 ;
  assign n13886 = ~n13864 & ~n13885 ;
  assign n13887 = \P1_state_reg[0]/NET0131  & ~n13886 ;
  assign n13888 = ~n13863 & ~n13887 ;
  assign n13889 = \P3_reg0_reg[8]/NET0131  & ~n2143 ;
  assign n13890 = \P3_reg0_reg[8]/NET0131  & n2145 ;
  assign n13900 = n2234 & ~n11628 ;
  assign n13898 = n2391 & n11621 ;
  assign n13899 = ~n1704 & n2285 ;
  assign n13901 = ~n13898 & ~n13899 ;
  assign n13902 = ~n13900 & n13901 ;
  assign n13903 = n2163 & ~n13902 ;
  assign n13892 = \P3_reg0_reg[8]/NET0131  & ~n2236 ;
  assign n13896 = ~n11632 & ~n13892 ;
  assign n13897 = n2393 & ~n13896 ;
  assign n13891 = \P3_reg0_reg[8]/NET0131  & ~n12214 ;
  assign n13893 = n2236 & ~n11639 ;
  assign n13894 = ~n13892 & ~n13893 ;
  assign n13895 = n737 & ~n13894 ;
  assign n13904 = ~n13891 & ~n13895 ;
  assign n13905 = ~n13897 & n13904 ;
  assign n13906 = ~n13903 & n13905 ;
  assign n13907 = n2147 & ~n13906 ;
  assign n13908 = ~n13890 & ~n13907 ;
  assign n13909 = \P1_state_reg[0]/NET0131  & ~n13908 ;
  assign n13910 = ~n13889 & ~n13909 ;
  assign n13911 = \P1_reg0_reg[4]/NET0131  & ~n6078 ;
  assign n13912 = \P1_reg0_reg[4]/NET0131  & n6095 ;
  assign n13914 = \P1_reg0_reg[4]/NET0131  & ~n6409 ;
  assign n13915 = n6409 & ~n12739 ;
  assign n13916 = ~n13914 & ~n13915 ;
  assign n13917 = n4011 & ~n13916 ;
  assign n13921 = n6409 & n12751 ;
  assign n13922 = ~n13914 & ~n13921 ;
  assign n13923 = n6282 & ~n13922 ;
  assign n13918 = n6409 & ~n12745 ;
  assign n13919 = ~n13914 & ~n13918 ;
  assign n13920 = n6207 & ~n13919 ;
  assign n13913 = \P1_reg0_reg[4]/NET0131  & ~n11142 ;
  assign n13924 = n6409 & ~n12731 ;
  assign n13925 = ~n13913 & ~n13924 ;
  assign n13926 = ~n13920 & n13925 ;
  assign n13927 = ~n13923 & n13926 ;
  assign n13928 = ~n13917 & n13927 ;
  assign n13929 = n6097 & ~n13928 ;
  assign n13930 = ~n13912 & ~n13929 ;
  assign n13931 = \P1_state_reg[0]/NET0131  & ~n13930 ;
  assign n13932 = ~n13911 & ~n13931 ;
  assign n13933 = \P1_reg0_reg[5]/NET0131  & ~n6078 ;
  assign n13934 = \P1_reg0_reg[5]/NET0131  & n6095 ;
  assign n13936 = \P1_reg0_reg[5]/NET0131  & ~n6409 ;
  assign n13937 = n6409 & ~n12795 ;
  assign n13938 = ~n13936 & ~n13937 ;
  assign n13939 = n6282 & ~n13938 ;
  assign n13946 = n6409 & n12774 ;
  assign n13947 = ~n13936 & ~n13946 ;
  assign n13948 = n6359 & ~n13947 ;
  assign n13935 = \P1_reg0_reg[5]/NET0131  & ~n6424 ;
  assign n13949 = ~n3128 & n6409 ;
  assign n13950 = ~n13936 & ~n13949 ;
  assign n13951 = n6365 & ~n13950 ;
  assign n13952 = ~n13935 & ~n13951 ;
  assign n13953 = ~n13948 & n13952 ;
  assign n13954 = ~n13939 & n13953 ;
  assign n13940 = n6409 & n12781 ;
  assign n13941 = ~n13936 & ~n13940 ;
  assign n13942 = n6207 & ~n13941 ;
  assign n13943 = n6409 & n12789 ;
  assign n13944 = ~n13936 & ~n13943 ;
  assign n13945 = n4011 & ~n13944 ;
  assign n13955 = ~n13942 & ~n13945 ;
  assign n13956 = n13954 & n13955 ;
  assign n13957 = n6097 & ~n13956 ;
  assign n13958 = ~n13934 & ~n13957 ;
  assign n13959 = \P1_state_reg[0]/NET0131  & ~n13958 ;
  assign n13960 = ~n13933 & ~n13959 ;
  assign n13961 = \P3_reg1_reg[5]/NET0131  & ~n2143 ;
  assign n13962 = \P3_reg1_reg[5]/NET0131  & n2145 ;
  assign n13969 = \P3_reg1_reg[5]/NET0131  & ~n2427 ;
  assign n13973 = n2427 & ~n12832 ;
  assign n13974 = ~n13969 & ~n13973 ;
  assign n13975 = n737 & ~n13974 ;
  assign n13964 = \P3_reg1_reg[5]/NET0131  & ~n2408 ;
  assign n13965 = n2408 & ~n12819 ;
  assign n13966 = ~n13964 & ~n13965 ;
  assign n13967 = n714 & ~n13966 ;
  assign n13976 = n2408 & n12838 ;
  assign n13977 = ~n13964 & ~n13976 ;
  assign n13978 = ~n2518 & ~n13977 ;
  assign n13970 = n2427 & n12838 ;
  assign n13971 = ~n13969 & ~n13970 ;
  assign n13972 = n2425 & ~n13971 ;
  assign n13963 = n2408 & n13830 ;
  assign n13968 = \P3_reg1_reg[5]/NET0131  & ~n6449 ;
  assign n13979 = ~n13963 & ~n13968 ;
  assign n13980 = ~n13972 & n13979 ;
  assign n13981 = ~n13978 & n13980 ;
  assign n13982 = ~n13967 & n13981 ;
  assign n13983 = ~n13975 & n13982 ;
  assign n13984 = n2147 & ~n13983 ;
  assign n13985 = ~n13962 & ~n13984 ;
  assign n13986 = \P1_state_reg[0]/NET0131  & ~n13985 ;
  assign n13987 = ~n13961 & ~n13986 ;
  assign n13988 = \P3_reg1_reg[6]/NET0131  & ~n2143 ;
  assign n13989 = \P3_reg1_reg[6]/NET0131  & n2145 ;
  assign n13999 = \P3_reg1_reg[6]/NET0131  & ~n2427 ;
  assign n14000 = n2427 & ~n12877 ;
  assign n14001 = ~n13999 & ~n14000 ;
  assign n14002 = n737 & ~n14001 ;
  assign n13991 = \P3_reg1_reg[6]/NET0131  & ~n2408 ;
  assign n13992 = n2408 & n12868 ;
  assign n13993 = ~n13991 & ~n13992 ;
  assign n13994 = ~n2518 & ~n13993 ;
  assign n13990 = n2408 & n13852 ;
  assign n13995 = \P3_reg1_reg[6]/NET0131  & ~n6449 ;
  assign n14006 = ~n13990 & ~n13995 ;
  assign n14007 = ~n13994 & n14006 ;
  assign n13996 = n2408 & ~n12860 ;
  assign n13997 = ~n13991 & ~n13996 ;
  assign n13998 = n714 & ~n13997 ;
  assign n14003 = n2427 & n12868 ;
  assign n14004 = ~n13999 & ~n14003 ;
  assign n14005 = n2425 & ~n14004 ;
  assign n14008 = ~n13998 & ~n14005 ;
  assign n14009 = n14007 & n14008 ;
  assign n14010 = ~n14002 & n14009 ;
  assign n14011 = n2147 & ~n14010 ;
  assign n14012 = ~n13989 & ~n14011 ;
  assign n14013 = \P1_state_reg[0]/NET0131  & ~n14012 ;
  assign n14014 = ~n13988 & ~n14013 ;
  assign n14015 = \P3_reg1_reg[7]/NET0131  & ~n2143 ;
  assign n14016 = \P3_reg1_reg[7]/NET0131  & n2145 ;
  assign n14023 = \P3_reg1_reg[7]/NET0131  & ~n2427 ;
  assign n14027 = n2427 & ~n12913 ;
  assign n14028 = ~n14023 & ~n14027 ;
  assign n14029 = n737 & ~n14028 ;
  assign n14018 = \P3_reg1_reg[7]/NET0131  & ~n2408 ;
  assign n14019 = n2408 & n12901 ;
  assign n14020 = ~n14018 & ~n14019 ;
  assign n14021 = n714 & ~n14020 ;
  assign n14030 = n2408 & ~n12919 ;
  assign n14031 = ~n14018 & ~n14030 ;
  assign n14032 = ~n2518 & ~n14031 ;
  assign n14024 = n2427 & ~n12919 ;
  assign n14025 = ~n14023 & ~n14024 ;
  assign n14026 = n2425 & ~n14025 ;
  assign n14017 = n2408 & n13865 ;
  assign n14022 = \P3_reg1_reg[7]/NET0131  & ~n6449 ;
  assign n14033 = ~n14017 & ~n14022 ;
  assign n14034 = ~n14026 & n14033 ;
  assign n14035 = ~n14032 & n14034 ;
  assign n14036 = ~n14021 & n14035 ;
  assign n14037 = ~n14029 & n14036 ;
  assign n14038 = n2147 & ~n14037 ;
  assign n14039 = ~n14016 & ~n14038 ;
  assign n14040 = \P1_state_reg[0]/NET0131  & ~n14039 ;
  assign n14041 = ~n14015 & ~n14040 ;
  assign n14042 = \P3_reg1_reg[8]/NET0131  & ~n2143 ;
  assign n14043 = \P3_reg1_reg[8]/NET0131  & n2145 ;
  assign n14046 = \P3_reg1_reg[8]/NET0131  & ~n2427 ;
  assign n14047 = n2427 & ~n11639 ;
  assign n14048 = ~n14046 & ~n14047 ;
  assign n14049 = n737 & ~n14048 ;
  assign n14044 = n2408 & n13899 ;
  assign n14045 = \P3_reg1_reg[8]/NET0131  & ~n6449 ;
  assign n14060 = ~n14044 & ~n14045 ;
  assign n14061 = ~n14049 & n14060 ;
  assign n14057 = n2427 & ~n11628 ;
  assign n14058 = ~n14046 & ~n14057 ;
  assign n14059 = n2425 & ~n14058 ;
  assign n14050 = \P3_reg1_reg[8]/NET0131  & ~n2408 ;
  assign n14051 = n2408 & ~n11628 ;
  assign n14052 = ~n14050 & ~n14051 ;
  assign n14053 = ~n2518 & ~n14052 ;
  assign n14054 = n2408 & n11621 ;
  assign n14055 = ~n14050 & ~n14054 ;
  assign n14056 = n714 & ~n14055 ;
  assign n14062 = ~n14053 & ~n14056 ;
  assign n14063 = ~n14059 & n14062 ;
  assign n14064 = n14061 & n14063 ;
  assign n14065 = n2147 & ~n14064 ;
  assign n14066 = ~n14043 & ~n14065 ;
  assign n14067 = \P1_state_reg[0]/NET0131  & ~n14066 ;
  assign n14068 = ~n14042 & ~n14067 ;
  assign n14069 = \P1_reg1_reg[11]/NET0131  & ~n12612 ;
  assign n14070 = n9045 & ~n12960 ;
  assign n14071 = ~n14069 & ~n14070 ;
  assign n14072 = \P3_reg2_reg[5]/NET0131  & ~n2143 ;
  assign n14073 = \P3_reg2_reg[5]/NET0131  & n2145 ;
  assign n14079 = \P3_reg2_reg[5]/NET0131  & ~n2408 ;
  assign n14082 = n2408 & ~n12832 ;
  assign n14083 = ~n14079 & ~n14082 ;
  assign n14084 = n737 & ~n14083 ;
  assign n14075 = \P3_reg2_reg[5]/NET0131  & ~n2427 ;
  assign n14076 = n2427 & ~n12819 ;
  assign n14077 = ~n14075 & ~n14076 ;
  assign n14078 = n714 & ~n14077 ;
  assign n14085 = ~n13970 & ~n14075 ;
  assign n14086 = ~n2518 & ~n14085 ;
  assign n14080 = ~n13976 & ~n14079 ;
  assign n14081 = n2425 & ~n14080 ;
  assign n14088 = \P3_reg2_reg[5]/NET0131  & ~n2429 ;
  assign n14074 = n2427 & n13830 ;
  assign n14087 = ~n1774 & n2283 ;
  assign n14089 = ~n14074 & ~n14087 ;
  assign n14090 = ~n14088 & n14089 ;
  assign n14091 = ~n14081 & n14090 ;
  assign n14092 = ~n14086 & n14091 ;
  assign n14093 = ~n14078 & n14092 ;
  assign n14094 = ~n14084 & n14093 ;
  assign n14095 = n2147 & ~n14094 ;
  assign n14096 = ~n14073 & ~n14095 ;
  assign n14097 = \P1_state_reg[0]/NET0131  & ~n14096 ;
  assign n14098 = ~n14072 & ~n14097 ;
  assign n14099 = \P3_reg2_reg[6]/NET0131  & ~n2143 ;
  assign n14100 = \P3_reg2_reg[6]/NET0131  & n2145 ;
  assign n14108 = \P3_reg2_reg[6]/NET0131  & ~n2408 ;
  assign n14109 = n2408 & ~n12877 ;
  assign n14110 = ~n14108 & ~n14109 ;
  assign n14111 = n737 & ~n14110 ;
  assign n14102 = \P3_reg2_reg[6]/NET0131  & ~n2427 ;
  assign n14103 = ~n14003 & ~n14102 ;
  assign n14104 = ~n2518 & ~n14103 ;
  assign n14115 = \P3_reg2_reg[6]/NET0131  & ~n2429 ;
  assign n14101 = n2427 & n13852 ;
  assign n14114 = ~n1750 & n2283 ;
  assign n14116 = ~n14101 & ~n14114 ;
  assign n14117 = ~n14115 & n14116 ;
  assign n14118 = ~n14104 & n14117 ;
  assign n14105 = n2427 & ~n12860 ;
  assign n14106 = ~n14102 & ~n14105 ;
  assign n14107 = n714 & ~n14106 ;
  assign n14112 = ~n13992 & ~n14108 ;
  assign n14113 = n2425 & ~n14112 ;
  assign n14119 = ~n14107 & ~n14113 ;
  assign n14120 = n14118 & n14119 ;
  assign n14121 = ~n14111 & n14120 ;
  assign n14122 = n2147 & ~n14121 ;
  assign n14123 = ~n14100 & ~n14122 ;
  assign n14124 = \P1_state_reg[0]/NET0131  & ~n14123 ;
  assign n14125 = ~n14099 & ~n14124 ;
  assign n14126 = \P1_reg1_reg[14]/NET0131  & ~n9053 ;
  assign n14127 = n9045 & ~n13738 ;
  assign n14128 = ~n14126 & ~n14127 ;
  assign n14129 = \P3_reg2_reg[7]/NET0131  & ~n2143 ;
  assign n14130 = \P3_reg2_reg[7]/NET0131  & n2145 ;
  assign n14136 = \P3_reg2_reg[7]/NET0131  & ~n2408 ;
  assign n14139 = n2408 & ~n12913 ;
  assign n14140 = ~n14136 & ~n14139 ;
  assign n14141 = n737 & ~n14140 ;
  assign n14132 = \P3_reg2_reg[7]/NET0131  & ~n2427 ;
  assign n14133 = n2427 & n12901 ;
  assign n14134 = ~n14132 & ~n14133 ;
  assign n14135 = n714 & ~n14134 ;
  assign n14142 = ~n14024 & ~n14132 ;
  assign n14143 = ~n2518 & ~n14142 ;
  assign n14137 = ~n14030 & ~n14136 ;
  assign n14138 = n2425 & ~n14137 ;
  assign n14145 = \P3_reg2_reg[7]/NET0131  & ~n2429 ;
  assign n14131 = n2427 & n13865 ;
  assign n14144 = ~n1724 & n2283 ;
  assign n14146 = ~n14131 & ~n14144 ;
  assign n14147 = ~n14145 & n14146 ;
  assign n14148 = ~n14138 & n14147 ;
  assign n14149 = ~n14143 & n14148 ;
  assign n14150 = ~n14135 & n14149 ;
  assign n14151 = ~n14141 & n14150 ;
  assign n14152 = n2147 & ~n14151 ;
  assign n14153 = ~n14130 & ~n14152 ;
  assign n14154 = \P1_state_reg[0]/NET0131  & ~n14153 ;
  assign n14155 = ~n14129 & ~n14154 ;
  assign n14156 = \P3_reg2_reg[8]/NET0131  & ~n2143 ;
  assign n14157 = \P3_reg2_reg[8]/NET0131  & n2145 ;
  assign n14159 = \P3_reg2_reg[8]/NET0131  & ~n2408 ;
  assign n14160 = n2408 & ~n11639 ;
  assign n14161 = ~n14159 & ~n14160 ;
  assign n14162 = n737 & ~n14161 ;
  assign n14172 = \P3_reg2_reg[8]/NET0131  & ~n2429 ;
  assign n14158 = n2427 & n13899 ;
  assign n14171 = ~n1681 & n2283 ;
  assign n14173 = ~n14158 & ~n14171 ;
  assign n14174 = ~n14172 & n14173 ;
  assign n14175 = ~n14162 & n14174 ;
  assign n14169 = ~n14051 & ~n14159 ;
  assign n14170 = n2425 & ~n14169 ;
  assign n14163 = \P3_reg2_reg[8]/NET0131  & ~n2427 ;
  assign n14164 = ~n14057 & ~n14163 ;
  assign n14165 = ~n2518 & ~n14164 ;
  assign n14166 = n2427 & n11621 ;
  assign n14167 = ~n14163 & ~n14166 ;
  assign n14168 = n714 & ~n14167 ;
  assign n14176 = ~n14165 & ~n14168 ;
  assign n14177 = ~n14170 & n14176 ;
  assign n14178 = n14175 & n14177 ;
  assign n14179 = n2147 & ~n14178 ;
  assign n14180 = ~n14157 & ~n14179 ;
  assign n14181 = \P1_state_reg[0]/NET0131  & ~n14180 ;
  assign n14182 = ~n14156 & ~n14181 ;
  assign n14183 = \P2_reg0_reg[11]/NET0131  & ~n5589 ;
  assign n14184 = \P2_reg0_reg[11]/NET0131  & n5585 ;
  assign n14186 = \P2_reg0_reg[11]/NET0131  & ~n6706 ;
  assign n14190 = n6706 & n11340 ;
  assign n14191 = ~n14186 & ~n14190 ;
  assign n14192 = n5383 & ~n14191 ;
  assign n14187 = n6706 & n11332 ;
  assign n14188 = ~n14186 & ~n14187 ;
  assign n14189 = n5329 & ~n14188 ;
  assign n14193 = n6706 & ~n11346 ;
  assign n14194 = ~n14186 & ~n14193 ;
  assign n14195 = n5526 & ~n14194 ;
  assign n14185 = \P2_reg0_reg[11]/NET0131  & ~n6717 ;
  assign n14196 = n6706 & ~n13083 ;
  assign n14197 = ~n14185 & ~n14196 ;
  assign n14198 = ~n14195 & n14197 ;
  assign n14199 = ~n14189 & n14198 ;
  assign n14200 = ~n14192 & n14199 ;
  assign n14201 = n5583 & ~n14200 ;
  assign n14202 = ~n14184 & ~n14201 ;
  assign n14203 = \P1_state_reg[0]/NET0131  & ~n14202 ;
  assign n14204 = ~n14183 & ~n14203 ;
  assign n14205 = \P2_reg0_reg[14]/NET0131  & ~n9531 ;
  assign n14206 = n9533 & ~n13100 ;
  assign n14207 = ~n14205 & ~n14206 ;
  assign n14209 = ~\P2_reg3_reg[3]/NET0131  & n5585 ;
  assign n14228 = n5203 & ~n5349 ;
  assign n14229 = ~n5203 & n5349 ;
  assign n14230 = ~n14228 & ~n14229 ;
  assign n14231 = ~n4231 & ~n14230 ;
  assign n14232 = n4231 & n5139 ;
  assign n14233 = ~n14231 & ~n14232 ;
  assign n14234 = n7453 & ~n14233 ;
  assign n14235 = \P2_reg3_reg[3]/NET0131  & ~n7453 ;
  assign n14236 = n5383 & ~n14235 ;
  assign n14237 = ~n14234 & n14236 ;
  assign n14219 = ~n5194 & ~n5242 ;
  assign n14221 = n5995 & n14219 ;
  assign n14220 = ~n5995 & ~n14219 ;
  assign n14222 = n5329 & ~n14220 ;
  assign n14223 = ~n14221 & n14222 ;
  assign n14211 = ~n5424 & ~n5426 ;
  assign n14213 = n5995 & ~n14211 ;
  assign n14212 = ~n5995 & n14211 ;
  assign n14214 = n5526 & ~n14212 ;
  assign n14215 = ~n14213 & n14214 ;
  assign n14216 = ~n5240 & ~n5530 ;
  assign n14217 = ~n5531 & n5563 ;
  assign n14218 = ~n14216 & n14217 ;
  assign n14224 = ~n14215 & ~n14218 ;
  assign n14225 = ~n14223 & n14224 ;
  assign n14226 = n7453 & ~n14225 ;
  assign n14210 = ~\P2_reg3_reg[3]/NET0131  & ~n12690 ;
  assign n14227 = ~n5240 & ~n7504 ;
  assign n14238 = ~n14210 & ~n14227 ;
  assign n14239 = ~n14226 & n14238 ;
  assign n14240 = ~n14237 & n14239 ;
  assign n14241 = n5583 & ~n14240 ;
  assign n14242 = ~n14209 & ~n14241 ;
  assign n14243 = \P1_state_reg[0]/NET0131  & ~n14242 ;
  assign n14208 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[3]/NET0131  ;
  assign n14244 = ~\P2_reg3_reg[3]/NET0131  & n5786 ;
  assign n14245 = ~n14208 & ~n14244 ;
  assign n14246 = ~n14243 & n14245 ;
  assign n14249 = ~\P3_reg3_reg[3]/NET0131  & n2145 ;
  assign n14259 = ~\P3_reg3_reg[3]/NET0131  & ~n2163 ;
  assign n14263 = n1806 & ~n2246 ;
  assign n14264 = ~n2239 & ~n13640 ;
  assign n14265 = ~n14263 & n14264 ;
  assign n14266 = ~n1830 & n2239 ;
  assign n14267 = ~n14265 & ~n14266 ;
  assign n14268 = n2163 & ~n14267 ;
  assign n14269 = ~n14259 & ~n14268 ;
  assign n14270 = n737 & ~n14269 ;
  assign n14252 = ~n2311 & ~n2313 ;
  assign n14253 = n2039 & ~n14252 ;
  assign n14254 = ~n2039 & n14252 ;
  assign n14255 = ~n14253 & ~n14254 ;
  assign n14260 = n2163 & ~n14255 ;
  assign n14261 = ~n14259 & ~n14260 ;
  assign n14262 = n2393 & ~n14261 ;
  assign n14251 = ~\P3_reg3_reg[3]/NET0131  & ~n2236 ;
  assign n14256 = n2236 & ~n14255 ;
  assign n14257 = ~n14251 & ~n14256 ;
  assign n14258 = n2391 & ~n14257 ;
  assign n14271 = ~n1845 & ~n2167 ;
  assign n14272 = n2039 & ~n14271 ;
  assign n14273 = ~n2039 & n14271 ;
  assign n14274 = ~n14272 & ~n14273 ;
  assign n14275 = n2236 & n14274 ;
  assign n14276 = ~n14251 & ~n14275 ;
  assign n14277 = n2234 & ~n14276 ;
  assign n14250 = ~n1868 & n2580 ;
  assign n14278 = ~\P3_reg3_reg[3]/NET0131  & ~n2583 ;
  assign n14279 = ~n14250 & ~n14278 ;
  assign n14280 = ~n14277 & n14279 ;
  assign n14281 = ~n14258 & n14280 ;
  assign n14282 = ~n14262 & n14281 ;
  assign n14283 = ~n14270 & n14282 ;
  assign n14284 = n2147 & ~n14283 ;
  assign n14285 = ~n14249 & ~n14284 ;
  assign n14286 = \P1_state_reg[0]/NET0131  & ~n14285 ;
  assign n14247 = ~\P1_state_reg[0]/NET0131  & \P3_reg3_reg[3]/NET0131  ;
  assign n14248 = ~\P3_reg3_reg[3]/NET0131  & n765 ;
  assign n14287 = ~n14247 & ~n14248 ;
  assign n14288 = ~n14286 & n14287 ;
  assign n14289 = \P1_reg1_reg[3]/NET0131  & ~n6078 ;
  assign n14290 = \P1_reg1_reg[3]/NET0131  & n6095 ;
  assign n14292 = \P1_reg1_reg[3]/NET0131  & ~n6683 ;
  assign n14293 = n6683 & n13507 ;
  assign n14294 = ~n14292 & ~n14293 ;
  assign n14295 = n4011 & ~n14294 ;
  assign n14299 = n6683 & n13519 ;
  assign n14300 = ~n14292 & ~n14299 ;
  assign n14301 = n6282 & ~n14300 ;
  assign n14296 = n6683 & n13513 ;
  assign n14297 = ~n14292 & ~n14296 ;
  assign n14298 = n6207 & ~n14297 ;
  assign n14291 = n6683 & ~n13500 ;
  assign n14302 = \P1_reg1_reg[3]/NET0131  & ~n6695 ;
  assign n14303 = ~n14291 & ~n14302 ;
  assign n14304 = ~n14298 & n14303 ;
  assign n14305 = ~n14301 & n14304 ;
  assign n14306 = ~n14295 & n14305 ;
  assign n14307 = n6097 & ~n14306 ;
  assign n14308 = ~n14290 & ~n14307 ;
  assign n14309 = \P1_state_reg[0]/NET0131  & ~n14308 ;
  assign n14310 = ~n14289 & ~n14309 ;
  assign n14311 = \P1_reg1_reg[7]/NET0131  & ~n6078 ;
  assign n14312 = \P1_reg1_reg[7]/NET0131  & n6095 ;
  assign n14314 = \P1_reg1_reg[7]/NET0131  & ~n6683 ;
  assign n14315 = n6683 & ~n13592 ;
  assign n14316 = ~n14314 & ~n14315 ;
  assign n14317 = n4011 & ~n14316 ;
  assign n14321 = n6683 & ~n13604 ;
  assign n14322 = ~n14314 & ~n14321 ;
  assign n14323 = n6282 & ~n14322 ;
  assign n14318 = n6683 & n13598 ;
  assign n14319 = ~n14314 & ~n14318 ;
  assign n14320 = n6207 & ~n14319 ;
  assign n14313 = n6683 & ~n13585 ;
  assign n14324 = \P1_reg1_reg[7]/NET0131  & ~n6695 ;
  assign n14325 = ~n14313 & ~n14324 ;
  assign n14326 = ~n14320 & n14325 ;
  assign n14327 = ~n14323 & n14326 ;
  assign n14328 = ~n14317 & n14327 ;
  assign n14329 = n6097 & ~n14328 ;
  assign n14330 = ~n14312 & ~n14329 ;
  assign n14331 = \P1_state_reg[0]/NET0131  & ~n14330 ;
  assign n14332 = ~n14311 & ~n14331 ;
  assign n14333 = \P2_reg0_reg[7]/NET0131  & ~n9531 ;
  assign n14334 = ~n5081 & n5565 ;
  assign n14335 = n13443 & ~n14334 ;
  assign n14336 = n9533 & ~n14335 ;
  assign n14337 = ~n14333 & ~n14336 ;
  assign n14338 = ~n5058 & n5565 ;
  assign n14339 = ~n13481 & ~n14338 ;
  assign n14340 = n13471 & n14339 ;
  assign n14341 = ~n13477 & n14340 ;
  assign n14342 = n9533 & ~n14341 ;
  assign n14343 = \P2_reg0_reg[8]/NET0131  & ~n9531 ;
  assign n14344 = ~n14342 & ~n14343 ;
  assign n14345 = \P2_reg1_reg[7]/NET0131  & ~n5589 ;
  assign n14346 = \P2_reg1_reg[7]/NET0131  & n5585 ;
  assign n14347 = \P2_reg1_reg[7]/NET0131  & ~n8918 ;
  assign n14348 = n6380 & ~n14335 ;
  assign n14349 = ~n14347 & ~n14348 ;
  assign n14350 = n5583 & ~n14349 ;
  assign n14351 = ~n14346 & ~n14350 ;
  assign n14352 = \P1_state_reg[0]/NET0131  & ~n14351 ;
  assign n14353 = ~n14345 & ~n14352 ;
  assign n14356 = \P2_reg1_reg[8]/NET0131  & ~n6380 ;
  assign n14357 = n8913 & n13476 ;
  assign n14358 = ~n14356 & ~n14357 ;
  assign n14359 = n5383 & ~n14358 ;
  assign n14354 = \P2_reg1_reg[8]/NET0131  & ~n8901 ;
  assign n14355 = n8913 & ~n14340 ;
  assign n14360 = ~n14354 & ~n14355 ;
  assign n14361 = ~n14359 & n14360 ;
  assign n14362 = \P1_reg2_reg[3]/NET0131  & ~n6078 ;
  assign n14363 = \P1_reg2_reg[3]/NET0131  & n6095 ;
  assign n14365 = \P1_reg2_reg[3]/NET0131  & ~n6113 ;
  assign n14366 = n6113 & n13507 ;
  assign n14367 = ~n14365 & ~n14366 ;
  assign n14368 = n4011 & ~n14367 ;
  assign n14372 = n6113 & n13519 ;
  assign n14373 = ~n14365 & ~n14372 ;
  assign n14374 = n6282 & ~n14373 ;
  assign n14369 = n6113 & n13513 ;
  assign n14370 = ~n14365 & ~n14369 ;
  assign n14371 = n6207 & ~n14370 ;
  assign n14364 = n6113 & ~n13500 ;
  assign n14375 = ~\P1_reg3_reg[3]/NET0131  & n4112 ;
  assign n14376 = \P1_reg2_reg[3]/NET0131  & ~n11834 ;
  assign n14377 = ~n14375 & ~n14376 ;
  assign n14378 = ~n14364 & n14377 ;
  assign n14379 = ~n14371 & n14378 ;
  assign n14380 = ~n14374 & n14379 ;
  assign n14381 = ~n14368 & n14380 ;
  assign n14382 = n6097 & ~n14381 ;
  assign n14383 = ~n14363 & ~n14382 ;
  assign n14384 = \P1_state_reg[0]/NET0131  & ~n14383 ;
  assign n14385 = ~n14362 & ~n14384 ;
  assign n14386 = \P1_reg2_reg[6]/NET0131  & ~n6078 ;
  assign n14387 = \P1_reg2_reg[6]/NET0131  & n6095 ;
  assign n14389 = \P1_reg2_reg[6]/NET0131  & ~n6113 ;
  assign n14390 = n6113 & n13550 ;
  assign n14391 = ~n14389 & ~n14390 ;
  assign n14392 = n4011 & ~n14391 ;
  assign n14396 = n6113 & ~n13562 ;
  assign n14397 = ~n14389 & ~n14396 ;
  assign n14398 = n6282 & ~n14397 ;
  assign n14393 = n6113 & n13556 ;
  assign n14394 = ~n14389 & ~n14393 ;
  assign n14395 = n6207 & ~n14394 ;
  assign n14388 = n6113 & ~n13542 ;
  assign n14399 = n3739 & n4112 ;
  assign n14400 = \P1_reg2_reg[6]/NET0131  & ~n11834 ;
  assign n14401 = ~n14399 & ~n14400 ;
  assign n14402 = ~n14388 & n14401 ;
  assign n14403 = ~n14395 & n14402 ;
  assign n14404 = ~n14398 & n14403 ;
  assign n14405 = ~n14392 & n14404 ;
  assign n14406 = n6097 & ~n14405 ;
  assign n14407 = ~n14387 & ~n14406 ;
  assign n14408 = \P1_state_reg[0]/NET0131  & ~n14407 ;
  assign n14409 = ~n14386 & ~n14408 ;
  assign n14410 = \P1_reg2_reg[7]/NET0131  & ~n6078 ;
  assign n14411 = \P1_reg2_reg[7]/NET0131  & n6095 ;
  assign n14413 = \P1_reg2_reg[7]/NET0131  & ~n6113 ;
  assign n14414 = n6113 & ~n13592 ;
  assign n14415 = ~n14413 & ~n14414 ;
  assign n14416 = n4011 & ~n14415 ;
  assign n14420 = n6113 & ~n13604 ;
  assign n14421 = ~n14413 & ~n14420 ;
  assign n14422 = n6282 & ~n14421 ;
  assign n14417 = n6113 & n13598 ;
  assign n14418 = ~n14413 & ~n14417 ;
  assign n14419 = n6207 & ~n14418 ;
  assign n14412 = n6113 & ~n13585 ;
  assign n14423 = n3573 & n4112 ;
  assign n14424 = \P1_reg2_reg[7]/NET0131  & ~n11834 ;
  assign n14425 = ~n14423 & ~n14424 ;
  assign n14426 = ~n14412 & n14425 ;
  assign n14427 = ~n14419 & n14426 ;
  assign n14428 = ~n14422 & n14427 ;
  assign n14429 = ~n14416 & n14428 ;
  assign n14430 = n6097 & ~n14429 ;
  assign n14431 = ~n14411 & ~n14430 ;
  assign n14432 = \P1_state_reg[0]/NET0131  & ~n14431 ;
  assign n14433 = ~n14410 & ~n14432 ;
  assign n14434 = \P2_reg2_reg[6]/NET0131  & ~n5589 ;
  assign n14435 = \P2_reg2_reg[6]/NET0131  & n5585 ;
  assign n14437 = \P2_reg2_reg[6]/NET0131  & ~n4219 ;
  assign n14438 = n4219 & n13389 ;
  assign n14439 = ~n14437 & ~n14438 ;
  assign n14440 = n5383 & ~n14439 ;
  assign n14444 = n4219 & ~n13401 ;
  assign n14445 = ~n14437 & ~n14444 ;
  assign n14446 = n5329 & ~n14445 ;
  assign n14441 = n4219 & n13395 ;
  assign n14442 = ~n14437 & ~n14441 ;
  assign n14443 = n5526 & ~n14442 ;
  assign n14448 = ~n5107 & n5565 ;
  assign n14449 = ~n13407 & ~n14448 ;
  assign n14450 = n4219 & ~n14449 ;
  assign n14436 = \P2_reg2_reg[6]/NET0131  & ~n6839 ;
  assign n14447 = n5088 & n5574 ;
  assign n14451 = ~n14436 & ~n14447 ;
  assign n14452 = ~n14450 & n14451 ;
  assign n14453 = ~n14443 & n14452 ;
  assign n14454 = ~n14446 & n14453 ;
  assign n14455 = ~n14440 & n14454 ;
  assign n14456 = n5583 & ~n14455 ;
  assign n14457 = ~n14435 & ~n14456 ;
  assign n14458 = \P1_state_reg[0]/NET0131  & ~n14457 ;
  assign n14459 = ~n14434 & ~n14458 ;
  assign n14461 = ~\P2_reg2_reg[7]/NET0131  & ~n4219 ;
  assign n14462 = n13442 & ~n14334 ;
  assign n14463 = n4219 & ~n14462 ;
  assign n14464 = n5525 & n8830 ;
  assign n14465 = n8899 & ~n14464 ;
  assign n14466 = ~n13428 & n14465 ;
  assign n14467 = ~n14463 & n14466 ;
  assign n14468 = ~n14461 & ~n14467 ;
  assign n14460 = n5063 & n5574 ;
  assign n14469 = \P2_reg2_reg[7]/NET0131  & ~n13137 ;
  assign n14470 = ~n14460 & ~n14469 ;
  assign n14471 = ~n14468 & n14470 ;
  assign n14472 = ~\P2_reg2_reg[7]/NET0131  & ~n8899 ;
  assign n14473 = ~n14471 & ~n14472 ;
  assign n14474 = \P2_reg2_reg[8]/NET0131  & ~n9773 ;
  assign n14475 = n5033 & n5574 ;
  assign n14476 = n4219 & ~n14341 ;
  assign n14477 = ~n14475 & ~n14476 ;
  assign n14478 = n8899 & ~n14477 ;
  assign n14479 = ~n14474 & ~n14478 ;
  assign n14480 = \P1_reg0_reg[3]/NET0131  & ~n6078 ;
  assign n14481 = \P1_reg0_reg[3]/NET0131  & n6095 ;
  assign n14483 = \P1_reg0_reg[3]/NET0131  & ~n6409 ;
  assign n14484 = n6409 & n13507 ;
  assign n14485 = ~n14483 & ~n14484 ;
  assign n14486 = n4011 & ~n14485 ;
  assign n14490 = n6409 & n13513 ;
  assign n14491 = ~n14483 & ~n14490 ;
  assign n14492 = n6207 & ~n14491 ;
  assign n14487 = n6409 & n13519 ;
  assign n14488 = ~n14483 & ~n14487 ;
  assign n14489 = n6282 & ~n14488 ;
  assign n14482 = \P1_reg0_reg[3]/NET0131  & ~n11142 ;
  assign n14493 = n6409 & ~n13500 ;
  assign n14494 = ~n14482 & ~n14493 ;
  assign n14495 = ~n14489 & n14494 ;
  assign n14496 = ~n14492 & n14495 ;
  assign n14497 = ~n14486 & n14496 ;
  assign n14498 = n6097 & ~n14497 ;
  assign n14499 = ~n14481 & ~n14498 ;
  assign n14500 = \P1_state_reg[0]/NET0131  & ~n14499 ;
  assign n14501 = ~n14480 & ~n14500 ;
  assign n14502 = \P1_reg0_reg[7]/NET0131  & ~n6078 ;
  assign n14503 = \P1_reg0_reg[7]/NET0131  & n6095 ;
  assign n14505 = \P1_reg0_reg[7]/NET0131  & ~n6409 ;
  assign n14506 = n6409 & ~n13592 ;
  assign n14507 = ~n14505 & ~n14506 ;
  assign n14508 = n4011 & ~n14507 ;
  assign n14512 = n6409 & n13598 ;
  assign n14513 = ~n14505 & ~n14512 ;
  assign n14514 = n6207 & ~n14513 ;
  assign n14509 = n6409 & ~n13604 ;
  assign n14510 = ~n14505 & ~n14509 ;
  assign n14511 = n6282 & ~n14510 ;
  assign n14515 = n6409 & n13583 ;
  assign n14516 = ~n14505 & ~n14515 ;
  assign n14517 = n6359 & ~n14516 ;
  assign n14504 = \P1_reg0_reg[7]/NET0131  & ~n6424 ;
  assign n14518 = n3568 & n6409 ;
  assign n14519 = ~n14505 & ~n14518 ;
  assign n14520 = n6365 & ~n14519 ;
  assign n14521 = ~n14504 & ~n14520 ;
  assign n14522 = ~n14517 & n14521 ;
  assign n14523 = ~n14511 & n14522 ;
  assign n14524 = ~n14514 & n14523 ;
  assign n14525 = ~n14508 & n14524 ;
  assign n14526 = n6097 & ~n14525 ;
  assign n14527 = ~n14503 & ~n14526 ;
  assign n14528 = \P1_state_reg[0]/NET0131  & ~n14527 ;
  assign n14529 = ~n14502 & ~n14528 ;
  assign n14532 = n5199 & n5585 ;
  assign n14534 = n5199 & ~n7453 ;
  assign n14535 = n4231 & ~n5226 ;
  assign n14536 = n5117 & ~n14229 ;
  assign n14537 = ~n4231 & ~n5351 ;
  assign n14538 = ~n14536 & n14537 ;
  assign n14539 = ~n14535 & ~n14538 ;
  assign n14540 = n7453 & ~n14539 ;
  assign n14541 = ~n14534 & ~n14540 ;
  assign n14542 = n5383 & ~n14541 ;
  assign n14549 = ~n5815 & n5994 ;
  assign n14550 = n5815 & ~n5994 ;
  assign n14551 = ~n14549 & ~n14550 ;
  assign n14552 = n7453 & n14551 ;
  assign n14553 = ~n14534 & ~n14552 ;
  assign n14554 = n5526 & ~n14553 ;
  assign n14543 = n5994 & ~n6735 ;
  assign n14544 = ~n5994 & n6735 ;
  assign n14545 = ~n14543 & ~n14544 ;
  assign n14546 = n7453 & ~n14545 ;
  assign n14547 = ~n14534 & ~n14546 ;
  assign n14548 = n5329 & ~n14547 ;
  assign n14555 = ~n5218 & ~n5531 ;
  assign n14556 = ~n5532 & n5563 ;
  assign n14557 = ~n14555 & n14556 ;
  assign n14558 = n7453 & n14557 ;
  assign n14533 = ~n5218 & ~n7504 ;
  assign n14559 = n5199 & ~n7484 ;
  assign n14560 = ~n14533 & ~n14559 ;
  assign n14561 = ~n14558 & n14560 ;
  assign n14562 = ~n14548 & n14561 ;
  assign n14563 = ~n14554 & n14562 ;
  assign n14564 = ~n14542 & n14563 ;
  assign n14565 = n5583 & ~n14564 ;
  assign n14566 = ~n14532 & ~n14565 ;
  assign n14567 = \P1_state_reg[0]/NET0131  & ~n14566 ;
  assign n14530 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[4]/NET0131  ;
  assign n14531 = n5199 & n5786 ;
  assign n14568 = ~n14530 & ~n14531 ;
  assign n14569 = ~n14567 & n14568 ;
  assign n14570 = \P1_reg3_reg[2]/NET0131  & ~n6078 ;
  assign n14571 = \P1_reg3_reg[2]/NET0131  & n6095 ;
  assign n14573 = \P1_reg3_reg[2]/NET0131  & ~n6568 ;
  assign n14586 = n3756 & ~n6287 ;
  assign n14587 = ~n6288 & ~n14586 ;
  assign n14588 = ~n2713 & ~n14587 ;
  assign n14589 = n2713 & n3704 ;
  assign n14590 = ~n14588 & ~n14589 ;
  assign n14591 = n6568 & n14590 ;
  assign n14592 = ~n14573 & ~n14591 ;
  assign n14593 = n4011 & ~n14592 ;
  assign n14580 = ~n3381 & ~n4042 ;
  assign n14581 = n3381 & n4042 ;
  assign n14582 = ~n14580 & ~n14581 ;
  assign n14583 = n6568 & n14582 ;
  assign n14584 = ~n14573 & ~n14583 ;
  assign n14585 = n6282 & ~n14584 ;
  assign n14574 = n3381 & n6138 ;
  assign n14575 = ~n3381 & ~n6138 ;
  assign n14576 = ~n14574 & ~n14575 ;
  assign n14577 = n6568 & ~n14576 ;
  assign n14578 = ~n14573 & ~n14577 ;
  assign n14579 = n6207 & ~n14578 ;
  assign n14595 = ~n3378 & n6365 ;
  assign n14596 = ~n3378 & ~n6328 ;
  assign n14597 = ~n6329 & n6359 ;
  assign n14598 = ~n14596 & n14597 ;
  assign n14599 = ~n14595 & ~n14598 ;
  assign n14600 = n6568 & ~n14599 ;
  assign n14572 = \P1_reg3_reg[2]/NET0131  & ~n12757 ;
  assign n14594 = ~n3378 & n4112 ;
  assign n14601 = ~n14572 & ~n14594 ;
  assign n14602 = ~n14600 & n14601 ;
  assign n14603 = ~n14579 & n14602 ;
  assign n14604 = ~n14585 & n14603 ;
  assign n14605 = ~n14593 & n14604 ;
  assign n14606 = n6097 & ~n14605 ;
  assign n14607 = ~n14571 & ~n14606 ;
  assign n14608 = \P1_state_reg[0]/NET0131  & ~n14607 ;
  assign n14609 = ~n14570 & ~n14608 ;
  assign n14610 = \P3_reg3_reg[2]/NET0131  & ~n2143 ;
  assign n14611 = \P3_reg3_reg[2]/NET0131  & n2145 ;
  assign n14627 = \P3_reg3_reg[2]/NET0131  & ~n2163 ;
  assign n14628 = n1852 & ~n2245 ;
  assign n14629 = ~n2239 & ~n2246 ;
  assign n14630 = ~n14628 & n14629 ;
  assign n14631 = ~n1877 & n2239 ;
  assign n14632 = ~n14630 & ~n14631 ;
  assign n14633 = n2163 & ~n14632 ;
  assign n14634 = ~n14627 & ~n14633 ;
  assign n14635 = n737 & ~n14634 ;
  assign n14613 = \P3_reg3_reg[2]/NET0131  & ~n2236 ;
  assign n14614 = n2047 & ~n2310 ;
  assign n14615 = ~n2047 & n2310 ;
  assign n14616 = ~n14614 & ~n14615 ;
  assign n14617 = n2236 & ~n14616 ;
  assign n14618 = ~n14613 & ~n14617 ;
  assign n14619 = n2391 & ~n14618 ;
  assign n14612 = ~n1844 & n2580 ;
  assign n14620 = \P3_reg3_reg[2]/NET0131  & ~n2583 ;
  assign n14639 = ~n14612 & ~n14620 ;
  assign n14640 = ~n14619 & n14639 ;
  assign n14621 = ~n1967 & n2047 ;
  assign n14622 = n1967 & ~n2047 ;
  assign n14623 = ~n14621 & ~n14622 ;
  assign n14624 = n2236 & n14623 ;
  assign n14625 = ~n14613 & ~n14624 ;
  assign n14626 = n2234 & ~n14625 ;
  assign n14636 = n2163 & ~n14616 ;
  assign n14637 = ~n14627 & ~n14636 ;
  assign n14638 = n2393 & ~n14637 ;
  assign n14641 = ~n14626 & ~n14638 ;
  assign n14642 = n14640 & n14641 ;
  assign n14643 = ~n14635 & n14642 ;
  assign n14644 = n2147 & ~n14643 ;
  assign n14645 = ~n14611 & ~n14644 ;
  assign n14646 = \P1_state_reg[0]/NET0131  & ~n14645 ;
  assign n14647 = ~n14610 & ~n14646 ;
  assign n14648 = \P2_reg0_reg[4]/NET0131  & ~n5589 ;
  assign n14649 = \P2_reg0_reg[4]/NET0131  & n5585 ;
  assign n14653 = \P2_reg0_reg[4]/NET0131  & ~n6706 ;
  assign n14654 = n6706 & ~n14539 ;
  assign n14655 = ~n14653 & ~n14654 ;
  assign n14656 = n5383 & ~n14655 ;
  assign n14660 = n6706 & n14551 ;
  assign n14661 = ~n14653 & ~n14660 ;
  assign n14662 = n5526 & ~n14661 ;
  assign n14657 = n6706 & ~n14545 ;
  assign n14658 = ~n14653 & ~n14657 ;
  assign n14659 = n5329 & ~n14658 ;
  assign n14650 = ~n5218 & n5565 ;
  assign n14651 = ~n14557 & ~n14650 ;
  assign n14652 = n6706 & ~n14651 ;
  assign n14663 = \P2_reg0_reg[4]/NET0131  & ~n6717 ;
  assign n14664 = ~n14652 & ~n14663 ;
  assign n14665 = ~n14659 & n14664 ;
  assign n14666 = ~n14662 & n14665 ;
  assign n14667 = ~n14656 & n14666 ;
  assign n14668 = n5583 & ~n14667 ;
  assign n14669 = ~n14649 & ~n14668 ;
  assign n14670 = \P1_state_reg[0]/NET0131  & ~n14669 ;
  assign n14671 = ~n14648 & ~n14670 ;
  assign n14672 = \P2_reg1_reg[4]/NET0131  & ~n5589 ;
  assign n14673 = \P2_reg1_reg[4]/NET0131  & n5585 ;
  assign n14675 = \P2_reg1_reg[4]/NET0131  & ~n6380 ;
  assign n14676 = n6380 & ~n14539 ;
  assign n14677 = ~n14675 & ~n14676 ;
  assign n14678 = n5383 & ~n14677 ;
  assign n14682 = n6380 & n14551 ;
  assign n14683 = ~n14675 & ~n14682 ;
  assign n14684 = n5526 & ~n14683 ;
  assign n14679 = n6380 & ~n14545 ;
  assign n14680 = ~n14675 & ~n14679 ;
  assign n14681 = n5329 & ~n14680 ;
  assign n14674 = n6380 & ~n14651 ;
  assign n14685 = \P2_reg1_reg[4]/NET0131  & ~n6397 ;
  assign n14686 = ~n14674 & ~n14685 ;
  assign n14687 = ~n14681 & n14686 ;
  assign n14688 = ~n14684 & n14687 ;
  assign n14689 = ~n14678 & n14688 ;
  assign n14690 = n5583 & ~n14689 ;
  assign n14691 = ~n14673 & ~n14690 ;
  assign n14692 = \P1_state_reg[0]/NET0131  & ~n14691 ;
  assign n14693 = ~n14672 & ~n14692 ;
  assign n14694 = \P1_reg1_reg[6]/NET0131  & ~n6078 ;
  assign n14695 = \P1_reg1_reg[6]/NET0131  & n6095 ;
  assign n14697 = \P1_reg1_reg[6]/NET0131  & ~n6683 ;
  assign n14698 = n6683 & n13550 ;
  assign n14699 = ~n14697 & ~n14698 ;
  assign n14700 = n4011 & ~n14699 ;
  assign n14704 = n6683 & n13556 ;
  assign n14705 = ~n14697 & ~n14704 ;
  assign n14706 = n6207 & ~n14705 ;
  assign n14701 = n6683 & ~n13562 ;
  assign n14702 = ~n14697 & ~n14701 ;
  assign n14703 = n6282 & ~n14702 ;
  assign n14696 = n6683 & ~n13542 ;
  assign n14707 = \P1_reg1_reg[6]/NET0131  & ~n6695 ;
  assign n14708 = ~n14696 & ~n14707 ;
  assign n14709 = ~n14703 & n14708 ;
  assign n14710 = ~n14706 & n14709 ;
  assign n14711 = ~n14700 & n14710 ;
  assign n14712 = n6097 & ~n14711 ;
  assign n14713 = ~n14695 & ~n14712 ;
  assign n14714 = \P1_state_reg[0]/NET0131  & ~n14713 ;
  assign n14715 = ~n14694 & ~n14714 ;
  assign n14716 = \P2_reg0_reg[3]/NET0131  & ~n13732 ;
  assign n14718 = n5383 & n14233 ;
  assign n14717 = ~n5240 & n5565 ;
  assign n14719 = n14225 & ~n14717 ;
  assign n14720 = ~n14718 & n14719 ;
  assign n14721 = n9533 & ~n14720 ;
  assign n14722 = ~n14716 & ~n14721 ;
  assign n14723 = \P2_reg0_reg[6]/NET0131  & ~n5589 ;
  assign n14724 = \P2_reg0_reg[6]/NET0131  & n5585 ;
  assign n14726 = \P2_reg0_reg[6]/NET0131  & ~n6706 ;
  assign n14727 = n6706 & n13389 ;
  assign n14728 = ~n14726 & ~n14727 ;
  assign n14729 = n5383 & ~n14728 ;
  assign n14733 = n6706 & n13395 ;
  assign n14734 = ~n14726 & ~n14733 ;
  assign n14735 = n5526 & ~n14734 ;
  assign n14730 = n6706 & ~n13401 ;
  assign n14731 = ~n14726 & ~n14730 ;
  assign n14732 = n5329 & ~n14731 ;
  assign n14725 = \P2_reg0_reg[6]/NET0131  & ~n6717 ;
  assign n14736 = n6706 & ~n14449 ;
  assign n14737 = ~n14725 & ~n14736 ;
  assign n14738 = ~n14732 & n14737 ;
  assign n14739 = ~n14735 & n14738 ;
  assign n14740 = ~n14729 & n14739 ;
  assign n14741 = n5583 & ~n14740 ;
  assign n14742 = ~n14724 & ~n14741 ;
  assign n14743 = \P1_state_reg[0]/NET0131  & ~n14742 ;
  assign n14744 = ~n14723 & ~n14743 ;
  assign n14745 = \P2_reg1_reg[3]/NET0131  & ~n8902 ;
  assign n14746 = n8913 & ~n14720 ;
  assign n14747 = ~n14745 & ~n14746 ;
  assign n14748 = \P2_reg1_reg[6]/NET0131  & ~n5589 ;
  assign n14749 = \P2_reg1_reg[6]/NET0131  & n5585 ;
  assign n14751 = \P2_reg1_reg[6]/NET0131  & ~n6380 ;
  assign n14752 = n6380 & n13389 ;
  assign n14753 = ~n14751 & ~n14752 ;
  assign n14754 = n5383 & ~n14753 ;
  assign n14758 = n6380 & n13395 ;
  assign n14759 = ~n14751 & ~n14758 ;
  assign n14760 = n5526 & ~n14759 ;
  assign n14755 = n6380 & ~n13401 ;
  assign n14756 = ~n14751 & ~n14755 ;
  assign n14757 = n5329 & ~n14756 ;
  assign n14750 = \P2_reg1_reg[6]/NET0131  & ~n6397 ;
  assign n14761 = n6380 & ~n14449 ;
  assign n14762 = ~n14750 & ~n14761 ;
  assign n14763 = ~n14757 & n14762 ;
  assign n14764 = ~n14760 & n14763 ;
  assign n14765 = ~n14754 & n14764 ;
  assign n14766 = n5583 & ~n14765 ;
  assign n14767 = ~n14749 & ~n14766 ;
  assign n14768 = \P1_state_reg[0]/NET0131  & ~n14767 ;
  assign n14769 = ~n14748 & ~n14768 ;
  assign n14770 = n4219 & ~n14720 ;
  assign n14771 = ~\P2_reg3_reg[3]/NET0131  & n5574 ;
  assign n14772 = ~n14770 & ~n14771 ;
  assign n14773 = n8899 & ~n14772 ;
  assign n14774 = \P2_reg2_reg[3]/NET0131  & ~n9773 ;
  assign n14775 = ~n14773 & ~n14774 ;
  assign n14776 = \P3_reg0_reg[3]/NET0131  & ~n2143 ;
  assign n14777 = \P3_reg0_reg[3]/NET0131  & n2145 ;
  assign n14783 = \P3_reg0_reg[3]/NET0131  & ~n2236 ;
  assign n14786 = n2236 & ~n14267 ;
  assign n14787 = ~n14783 & ~n14786 ;
  assign n14788 = n737 & ~n14787 ;
  assign n14784 = ~n14256 & ~n14783 ;
  assign n14785 = n2393 & ~n14784 ;
  assign n14780 = \P3_reg0_reg[3]/NET0131  & ~n2163 ;
  assign n14781 = ~n14260 & ~n14780 ;
  assign n14782 = n2391 & ~n14781 ;
  assign n14789 = n2163 & n14274 ;
  assign n14790 = ~n14780 & ~n14789 ;
  assign n14791 = n2234 & ~n14790 ;
  assign n14778 = ~n1868 & n2285 ;
  assign n14779 = n2163 & n14778 ;
  assign n14792 = \P3_reg0_reg[3]/NET0131  & ~n2287 ;
  assign n14793 = ~n14779 & ~n14792 ;
  assign n14794 = ~n14791 & n14793 ;
  assign n14795 = ~n14782 & n14794 ;
  assign n14796 = ~n14785 & n14795 ;
  assign n14797 = ~n14788 & n14796 ;
  assign n14798 = n2147 & ~n14797 ;
  assign n14799 = ~n14777 & ~n14798 ;
  assign n14800 = \P1_state_reg[0]/NET0131  & ~n14799 ;
  assign n14801 = ~n14776 & ~n14800 ;
  assign n14802 = \P3_reg0_reg[4]/NET0131  & ~n2143 ;
  assign n14803 = \P3_reg0_reg[4]/NET0131  & n2145 ;
  assign n14805 = \P3_reg0_reg[4]/NET0131  & ~n2236 ;
  assign n14806 = n2236 & ~n13644 ;
  assign n14807 = ~n14805 & ~n14806 ;
  assign n14808 = n737 & ~n14807 ;
  assign n14809 = ~n1820 & n2285 ;
  assign n14810 = n13637 & ~n14809 ;
  assign n14811 = n2163 & ~n14810 ;
  assign n14804 = \P3_reg0_reg[4]/NET0131  & ~n12214 ;
  assign n14812 = n2236 & ~n13628 ;
  assign n14813 = ~n14805 & ~n14812 ;
  assign n14814 = n2393 & ~n14813 ;
  assign n14815 = ~n14804 & ~n14814 ;
  assign n14816 = ~n14811 & n14815 ;
  assign n14817 = ~n14808 & n14816 ;
  assign n14818 = n2147 & ~n14817 ;
  assign n14819 = ~n14803 & ~n14818 ;
  assign n14820 = \P1_state_reg[0]/NET0131  & ~n14819 ;
  assign n14821 = ~n14802 & ~n14820 ;
  assign n14822 = \P1_reg0_reg[6]/NET0131  & ~n6078 ;
  assign n14823 = \P1_reg0_reg[6]/NET0131  & n6095 ;
  assign n14825 = \P1_reg0_reg[6]/NET0131  & ~n6409 ;
  assign n14826 = n6409 & n13550 ;
  assign n14827 = ~n14825 & ~n14826 ;
  assign n14828 = n4011 & ~n14827 ;
  assign n14832 = n6409 & n13556 ;
  assign n14833 = ~n14825 & ~n14832 ;
  assign n14834 = n6207 & ~n14833 ;
  assign n14829 = n6409 & ~n13562 ;
  assign n14830 = ~n14825 & ~n14829 ;
  assign n14831 = n6282 & ~n14830 ;
  assign n14835 = n6409 & n13540 ;
  assign n14836 = ~n14825 & ~n14835 ;
  assign n14837 = n6359 & ~n14836 ;
  assign n14824 = \P1_reg0_reg[6]/NET0131  & ~n6424 ;
  assign n14838 = n3737 & n6409 ;
  assign n14839 = ~n14825 & ~n14838 ;
  assign n14840 = n6365 & ~n14839 ;
  assign n14841 = ~n14824 & ~n14840 ;
  assign n14842 = ~n14837 & n14841 ;
  assign n14843 = ~n14831 & n14842 ;
  assign n14844 = ~n14834 & n14843 ;
  assign n14845 = ~n14828 & n14844 ;
  assign n14846 = n6097 & ~n14845 ;
  assign n14847 = ~n14823 & ~n14846 ;
  assign n14848 = \P1_state_reg[0]/NET0131  & ~n14847 ;
  assign n14849 = ~n14822 & ~n14848 ;
  assign n14850 = \P3_reg1_reg[3]/NET0131  & ~n2143 ;
  assign n14851 = \P3_reg1_reg[3]/NET0131  & n2145 ;
  assign n14858 = \P3_reg1_reg[3]/NET0131  & ~n2427 ;
  assign n14862 = n2427 & ~n14267 ;
  assign n14863 = ~n14858 & ~n14862 ;
  assign n14864 = n737 & ~n14863 ;
  assign n14853 = \P3_reg1_reg[3]/NET0131  & ~n2408 ;
  assign n14854 = n2408 & ~n14255 ;
  assign n14855 = ~n14853 & ~n14854 ;
  assign n14856 = n714 & ~n14855 ;
  assign n14865 = n2408 & n14274 ;
  assign n14866 = ~n14853 & ~n14865 ;
  assign n14867 = ~n2518 & ~n14866 ;
  assign n14859 = n2427 & n14274 ;
  assign n14860 = ~n14858 & ~n14859 ;
  assign n14861 = n2425 & ~n14860 ;
  assign n14852 = n2408 & n14778 ;
  assign n14857 = \P3_reg1_reg[3]/NET0131  & ~n6449 ;
  assign n14868 = ~n14852 & ~n14857 ;
  assign n14869 = ~n14861 & n14868 ;
  assign n14870 = ~n14867 & n14869 ;
  assign n14871 = ~n14856 & n14870 ;
  assign n14872 = ~n14864 & n14871 ;
  assign n14873 = n2147 & ~n14872 ;
  assign n14874 = ~n14851 & ~n14873 ;
  assign n14875 = \P1_state_reg[0]/NET0131  & ~n14874 ;
  assign n14876 = ~n14850 & ~n14875 ;
  assign n14877 = \P3_reg1_reg[4]/NET0131  & ~n2143 ;
  assign n14878 = \P3_reg1_reg[4]/NET0131  & n2145 ;
  assign n14880 = \P3_reg1_reg[4]/NET0131  & ~n2427 ;
  assign n14889 = n2427 & ~n13644 ;
  assign n14890 = ~n14880 & ~n14889 ;
  assign n14891 = n737 & ~n14890 ;
  assign n14881 = n2427 & n13635 ;
  assign n14882 = ~n14880 & ~n14881 ;
  assign n14883 = n2425 & ~n14882 ;
  assign n14879 = n2408 & n14809 ;
  assign n14884 = \P3_reg1_reg[4]/NET0131  & ~n6449 ;
  assign n14895 = ~n14879 & ~n14884 ;
  assign n14896 = ~n14883 & n14895 ;
  assign n14885 = \P3_reg1_reg[4]/NET0131  & ~n2408 ;
  assign n14886 = n2408 & n13635 ;
  assign n14887 = ~n14885 & ~n14886 ;
  assign n14888 = ~n2518 & ~n14887 ;
  assign n14892 = n2408 & ~n13628 ;
  assign n14893 = ~n14885 & ~n14892 ;
  assign n14894 = n714 & ~n14893 ;
  assign n14897 = ~n14888 & ~n14894 ;
  assign n14898 = n14896 & n14897 ;
  assign n14899 = ~n14891 & n14898 ;
  assign n14900 = n2147 & ~n14899 ;
  assign n14901 = ~n14878 & ~n14900 ;
  assign n14902 = \P1_state_reg[0]/NET0131  & ~n14901 ;
  assign n14903 = ~n14877 & ~n14902 ;
  assign n14904 = \P3_reg2_reg[3]/NET0131  & ~n2143 ;
  assign n14905 = \P3_reg2_reg[3]/NET0131  & n2145 ;
  assign n14911 = \P3_reg2_reg[3]/NET0131  & ~n2408 ;
  assign n14914 = n2408 & ~n14267 ;
  assign n14915 = ~n14911 & ~n14914 ;
  assign n14916 = n737 & ~n14915 ;
  assign n14907 = \P3_reg2_reg[3]/NET0131  & ~n2427 ;
  assign n14908 = n2427 & ~n14255 ;
  assign n14909 = ~n14907 & ~n14908 ;
  assign n14910 = n714 & ~n14909 ;
  assign n14917 = ~n14859 & ~n14907 ;
  assign n14918 = ~n2518 & ~n14917 ;
  assign n14912 = ~n14865 & ~n14911 ;
  assign n14913 = n2425 & ~n14912 ;
  assign n14920 = \P3_reg2_reg[3]/NET0131  & ~n2429 ;
  assign n14906 = n2427 & n14778 ;
  assign n14919 = ~\P3_reg3_reg[3]/NET0131  & n2283 ;
  assign n14921 = ~n14906 & ~n14919 ;
  assign n14922 = ~n14920 & n14921 ;
  assign n14923 = ~n14913 & n14922 ;
  assign n14924 = ~n14918 & n14923 ;
  assign n14925 = ~n14910 & n14924 ;
  assign n14926 = ~n14916 & n14925 ;
  assign n14927 = n2147 & ~n14926 ;
  assign n14928 = ~n14905 & ~n14927 ;
  assign n14929 = \P1_state_reg[0]/NET0131  & ~n14928 ;
  assign n14930 = ~n14904 & ~n14929 ;
  assign n14931 = \P3_reg2_reg[4]/NET0131  & ~n2143 ;
  assign n14932 = \P3_reg2_reg[4]/NET0131  & n2145 ;
  assign n14934 = \P3_reg2_reg[4]/NET0131  & ~n2408 ;
  assign n14941 = n2408 & ~n13644 ;
  assign n14942 = ~n14934 & ~n14941 ;
  assign n14943 = n737 & ~n14942 ;
  assign n14935 = ~n14886 & ~n14934 ;
  assign n14936 = n2425 & ~n14935 ;
  assign n14947 = \P3_reg2_reg[4]/NET0131  & ~n2429 ;
  assign n14933 = n2427 & n14809 ;
  assign n14946 = ~n1801 & n2283 ;
  assign n14948 = ~n14933 & ~n14946 ;
  assign n14949 = ~n14947 & n14948 ;
  assign n14950 = ~n14936 & n14949 ;
  assign n14937 = \P3_reg2_reg[4]/NET0131  & ~n2427 ;
  assign n14938 = n2427 & ~n13628 ;
  assign n14939 = ~n14937 & ~n14938 ;
  assign n14940 = n714 & ~n14939 ;
  assign n14944 = ~n14881 & ~n14937 ;
  assign n14945 = ~n2518 & ~n14944 ;
  assign n14951 = ~n14940 & ~n14945 ;
  assign n14952 = n14950 & n14951 ;
  assign n14953 = ~n14943 & n14952 ;
  assign n14954 = n2147 & ~n14953 ;
  assign n14955 = ~n14932 & ~n14954 ;
  assign n14956 = \P1_state_reg[0]/NET0131  & ~n14955 ;
  assign n14957 = ~n14931 & ~n14956 ;
  assign n14958 = n8899 & n12691 ;
  assign n14959 = \P2_reg3_reg[2]/NET0131  & ~n14958 ;
  assign n14960 = n5226 & ~n5348 ;
  assign n14961 = ~n5349 & ~n14960 ;
  assign n14962 = ~n4231 & ~n14961 ;
  assign n14963 = n4231 & n5161 ;
  assign n14964 = ~n14962 & ~n14963 ;
  assign n14965 = n5383 & n14964 ;
  assign n14974 = ~n5193 & n5974 ;
  assign n14973 = n5193 & ~n5974 ;
  assign n14975 = n5329 & ~n14973 ;
  assign n14976 = ~n14974 & n14975 ;
  assign n14967 = n5811 & n5974 ;
  assign n14966 = ~n5811 & ~n5974 ;
  assign n14968 = n5526 & ~n14966 ;
  assign n14969 = ~n14967 & n14968 ;
  assign n14970 = ~n5153 & ~n5529 ;
  assign n14971 = ~n5530 & n5563 ;
  assign n14972 = ~n14970 & n14971 ;
  assign n14977 = ~n14969 & ~n14972 ;
  assign n14978 = ~n14976 & n14977 ;
  assign n14979 = ~n14965 & n14978 ;
  assign n14980 = n7453 & ~n14979 ;
  assign n14981 = ~n5153 & ~n7504 ;
  assign n14982 = ~n14980 & ~n14981 ;
  assign n14983 = n8899 & ~n14982 ;
  assign n14984 = ~n14959 & ~n14983 ;
  assign n14985 = \P3_reg3_reg[1]/NET0131  & ~n2143 ;
  assign n14986 = \P3_reg3_reg[1]/NET0131  & n2145 ;
  assign n14996 = \P3_reg3_reg[1]/NET0131  & ~n2163 ;
  assign n15000 = n1830 & ~n2244 ;
  assign n15001 = ~n2239 & ~n2245 ;
  assign n15002 = ~n15000 & n15001 ;
  assign n15003 = ~n1899 & n2239 ;
  assign n15004 = ~n15002 & ~n15003 ;
  assign n15005 = n2163 & ~n15004 ;
  assign n15006 = ~n14996 & ~n15005 ;
  assign n15007 = n737 & ~n15006 ;
  assign n14988 = \P3_reg3_reg[1]/NET0131  & ~n2236 ;
  assign n14989 = n2054 & ~n2308 ;
  assign n14990 = ~n2054 & n2308 ;
  assign n14991 = ~n14989 & ~n14990 ;
  assign n14992 = n2236 & n14991 ;
  assign n14993 = ~n14988 & ~n14992 ;
  assign n14994 = n2391 & ~n14993 ;
  assign n14987 = ~n1891 & n2580 ;
  assign n14995 = \P3_reg3_reg[1]/NET0131  & ~n2583 ;
  assign n15013 = ~n14987 & ~n14995 ;
  assign n15014 = ~n14994 & n15013 ;
  assign n14997 = n2163 & n14991 ;
  assign n14998 = ~n14996 & ~n14997 ;
  assign n14999 = n2393 & ~n14998 ;
  assign n15008 = n1965 & ~n2054 ;
  assign n15009 = ~n2055 & ~n15008 ;
  assign n15010 = n2236 & n15009 ;
  assign n15011 = ~n14988 & ~n15010 ;
  assign n15012 = n2234 & ~n15011 ;
  assign n15015 = ~n14999 & ~n15012 ;
  assign n15016 = n15014 & n15015 ;
  assign n15017 = ~n15007 & n15016 ;
  assign n15018 = n2147 & ~n15017 ;
  assign n15019 = ~n14986 & ~n15018 ;
  assign n15020 = \P1_state_reg[0]/NET0131  & ~n15019 ;
  assign n15021 = ~n14985 & ~n15020 ;
  assign n15022 = \P1_reg2_reg[2]/NET0131  & ~n6078 ;
  assign n15023 = \P1_reg2_reg[2]/NET0131  & n6095 ;
  assign n15025 = \P1_reg2_reg[2]/NET0131  & ~n6113 ;
  assign n15032 = n6113 & n14590 ;
  assign n15033 = ~n15025 & ~n15032 ;
  assign n15034 = n4011 & ~n15033 ;
  assign n15029 = n6113 & n14582 ;
  assign n15030 = ~n15025 & ~n15029 ;
  assign n15031 = n6282 & ~n15030 ;
  assign n15026 = n6113 & ~n14576 ;
  assign n15027 = ~n15025 & ~n15026 ;
  assign n15028 = n6207 & ~n15027 ;
  assign n15036 = n6113 & ~n14599 ;
  assign n15024 = \P1_reg2_reg[2]/NET0131  & ~n11834 ;
  assign n15035 = \P1_reg3_reg[2]/NET0131  & n4112 ;
  assign n15037 = ~n15024 & ~n15035 ;
  assign n15038 = ~n15036 & n15037 ;
  assign n15039 = ~n15028 & n15038 ;
  assign n15040 = ~n15031 & n15039 ;
  assign n15041 = ~n15034 & n15040 ;
  assign n15042 = n6097 & ~n15041 ;
  assign n15043 = ~n15023 & ~n15042 ;
  assign n15044 = \P1_state_reg[0]/NET0131  & ~n15043 ;
  assign n15045 = ~n15022 & ~n15044 ;
  assign n15051 = \P1_reg1_reg[2]/NET0131  & ~n6683 ;
  assign n15052 = n9045 & n14590 ;
  assign n15053 = ~n15051 & ~n15052 ;
  assign n15054 = n4011 & ~n15053 ;
  assign n15047 = n6207 & ~n14576 ;
  assign n15046 = n6282 & n14582 ;
  assign n15048 = n14599 & ~n15046 ;
  assign n15049 = ~n15047 & n15048 ;
  assign n15050 = n9045 & ~n15049 ;
  assign n15055 = n9044 & ~n11197 ;
  assign n15056 = n6695 & n15055 ;
  assign n15057 = \P1_reg1_reg[2]/NET0131  & ~n15056 ;
  assign n15058 = ~n15050 & ~n15057 ;
  assign n15059 = ~n15054 & n15058 ;
  assign n15060 = \P2_reg0_reg[2]/NET0131  & ~n5589 ;
  assign n15061 = \P2_reg0_reg[2]/NET0131  & n5585 ;
  assign n15063 = ~n5153 & n5565 ;
  assign n15064 = n14978 & ~n15063 ;
  assign n15065 = n6706 & ~n15064 ;
  assign n15062 = \P2_reg0_reg[2]/NET0131  & ~n8886 ;
  assign n15066 = n6706 & ~n14964 ;
  assign n15067 = ~\P2_reg0_reg[2]/NET0131  & ~n6706 ;
  assign n15068 = n5383 & ~n15067 ;
  assign n15069 = ~n15066 & n15068 ;
  assign n15070 = ~n15062 & ~n15069 ;
  assign n15071 = ~n15065 & n15070 ;
  assign n15072 = n5583 & ~n15071 ;
  assign n15073 = ~n15061 & ~n15072 ;
  assign n15074 = \P1_state_reg[0]/NET0131  & ~n15073 ;
  assign n15075 = ~n15060 & ~n15074 ;
  assign n15076 = ~n14965 & n15064 ;
  assign n15077 = n8913 & ~n15076 ;
  assign n15078 = n5525 & n9650 ;
  assign n15079 = n8900 & ~n15078 ;
  assign n15080 = \P2_reg1_reg[2]/NET0131  & ~n15079 ;
  assign n15081 = ~n15077 & ~n15080 ;
  assign n15082 = \P2_reg2_reg[4]/NET0131  & ~n5589 ;
  assign n15083 = \P2_reg2_reg[4]/NET0131  & n5585 ;
  assign n15085 = \P2_reg2_reg[4]/NET0131  & ~n4219 ;
  assign n15086 = n4219 & ~n14539 ;
  assign n15087 = ~n15085 & ~n15086 ;
  assign n15088 = n5383 & ~n15087 ;
  assign n15092 = n4219 & n14551 ;
  assign n15093 = ~n15085 & ~n15092 ;
  assign n15094 = n5526 & ~n15093 ;
  assign n15089 = n4219 & ~n14545 ;
  assign n15090 = ~n15085 & ~n15089 ;
  assign n15091 = n5329 & ~n15090 ;
  assign n15084 = n4219 & ~n14651 ;
  assign n15095 = n5199 & n5574 ;
  assign n15096 = \P2_reg2_reg[4]/NET0131  & ~n6839 ;
  assign n15097 = ~n15095 & ~n15096 ;
  assign n15098 = ~n15084 & n15097 ;
  assign n15099 = ~n15091 & n15098 ;
  assign n15100 = ~n15094 & n15099 ;
  assign n15101 = ~n15088 & n15100 ;
  assign n15102 = n5583 & ~n15101 ;
  assign n15103 = ~n15083 & ~n15102 ;
  assign n15104 = \P1_state_reg[0]/NET0131  & ~n15103 ;
  assign n15105 = ~n15082 & ~n15104 ;
  assign n15106 = \P1_reg0_reg[2]/NET0131  & n6095 ;
  assign n15108 = n6409 & ~n15049 ;
  assign n15107 = \P1_reg0_reg[2]/NET0131  & ~n13177 ;
  assign n15109 = n10016 & n14590 ;
  assign n15110 = ~n15107 & ~n15109 ;
  assign n15111 = ~n15108 & n15110 ;
  assign n15112 = n6097 & ~n15111 ;
  assign n15113 = ~n15106 & ~n15112 ;
  assign n15114 = \P1_state_reg[0]/NET0131  & ~n15113 ;
  assign n15115 = \P1_reg0_reg[2]/NET0131  & ~n6078 ;
  assign n15116 = ~n15114 & ~n15115 ;
  assign n15117 = \P3_reg0_reg[2]/NET0131  & ~n2143 ;
  assign n15118 = \P3_reg0_reg[2]/NET0131  & n2145 ;
  assign n15128 = \P3_reg0_reg[2]/NET0131  & ~n2236 ;
  assign n15129 = n2236 & ~n14632 ;
  assign n15130 = ~n15128 & ~n15129 ;
  assign n15131 = n737 & ~n15130 ;
  assign n15121 = \P3_reg0_reg[2]/NET0131  & ~n2163 ;
  assign n15122 = n2163 & n14623 ;
  assign n15123 = ~n15121 & ~n15122 ;
  assign n15124 = n2234 & ~n15123 ;
  assign n15119 = ~n1844 & n2285 ;
  assign n15120 = n2163 & n15119 ;
  assign n15125 = \P3_reg0_reg[2]/NET0131  & ~n2287 ;
  assign n15134 = ~n15120 & ~n15125 ;
  assign n15135 = ~n15124 & n15134 ;
  assign n15126 = ~n14636 & ~n15121 ;
  assign n15127 = n2391 & ~n15126 ;
  assign n15132 = ~n14617 & ~n15128 ;
  assign n15133 = n2393 & ~n15132 ;
  assign n15136 = ~n15127 & ~n15133 ;
  assign n15137 = n15135 & n15136 ;
  assign n15138 = ~n15131 & n15137 ;
  assign n15139 = n2147 & ~n15138 ;
  assign n15140 = ~n15118 & ~n15139 ;
  assign n15141 = \P1_state_reg[0]/NET0131  & ~n15140 ;
  assign n15142 = ~n15117 & ~n15141 ;
  assign n15143 = \P3_reg1_reg[2]/NET0131  & ~n2143 ;
  assign n15144 = \P3_reg1_reg[2]/NET0131  & n2145 ;
  assign n15154 = \P3_reg1_reg[2]/NET0131  & ~n2427 ;
  assign n15155 = n2427 & ~n14632 ;
  assign n15156 = ~n15154 & ~n15155 ;
  assign n15157 = n737 & ~n15156 ;
  assign n15146 = \P3_reg1_reg[2]/NET0131  & ~n2408 ;
  assign n15147 = n2408 & ~n14616 ;
  assign n15148 = ~n15146 & ~n15147 ;
  assign n15149 = n714 & ~n15148 ;
  assign n15145 = n2408 & n15119 ;
  assign n15150 = \P3_reg1_reg[2]/NET0131  & ~n6449 ;
  assign n15161 = ~n15145 & ~n15150 ;
  assign n15162 = ~n15149 & n15161 ;
  assign n15151 = n2408 & n14623 ;
  assign n15152 = ~n15146 & ~n15151 ;
  assign n15153 = ~n2518 & ~n15152 ;
  assign n15158 = n2427 & n14623 ;
  assign n15159 = ~n15154 & ~n15158 ;
  assign n15160 = n2425 & ~n15159 ;
  assign n15163 = ~n15153 & ~n15160 ;
  assign n15164 = n15162 & n15163 ;
  assign n15165 = ~n15157 & n15164 ;
  assign n15166 = n2147 & ~n15165 ;
  assign n15167 = ~n15144 & ~n15166 ;
  assign n15168 = \P1_state_reg[0]/NET0131  & ~n15167 ;
  assign n15169 = ~n15143 & ~n15168 ;
  assign n15170 = \P3_reg2_reg[2]/NET0131  & ~n2143 ;
  assign n15171 = \P3_reg2_reg[2]/NET0131  & n2145 ;
  assign n15176 = \P3_reg2_reg[2]/NET0131  & ~n2408 ;
  assign n15179 = n2408 & ~n14632 ;
  assign n15180 = ~n15176 & ~n15179 ;
  assign n15181 = n737 & ~n15180 ;
  assign n15173 = \P3_reg2_reg[2]/NET0131  & ~n2427 ;
  assign n15174 = ~n15158 & ~n15173 ;
  assign n15175 = ~n2518 & ~n15174 ;
  assign n15186 = \P3_reg2_reg[2]/NET0131  & ~n2429 ;
  assign n15172 = n2427 & n15119 ;
  assign n15185 = \P3_reg3_reg[2]/NET0131  & n2283 ;
  assign n15187 = ~n15172 & ~n15185 ;
  assign n15188 = ~n15186 & n15187 ;
  assign n15189 = ~n15175 & n15188 ;
  assign n15177 = ~n15151 & ~n15176 ;
  assign n15178 = n2425 & ~n15177 ;
  assign n15182 = n2427 & ~n14616 ;
  assign n15183 = ~n15173 & ~n15182 ;
  assign n15184 = n714 & ~n15183 ;
  assign n15190 = ~n15178 & ~n15184 ;
  assign n15191 = n15189 & n15190 ;
  assign n15192 = ~n15181 & n15191 ;
  assign n15193 = n2147 & ~n15192 ;
  assign n15194 = ~n15171 & ~n15193 ;
  assign n15195 = \P1_state_reg[0]/NET0131  & ~n15194 ;
  assign n15196 = ~n15170 & ~n15195 ;
  assign n15201 = n5139 & ~n5347 ;
  assign n15202 = ~n5348 & ~n15201 ;
  assign n15203 = ~n4231 & ~n15202 ;
  assign n15204 = n4231 & n5184 ;
  assign n15205 = ~n15203 & ~n15204 ;
  assign n15206 = n5383 & n15205 ;
  assign n15208 = n5419 & ~n5972 ;
  assign n15209 = n5526 & ~n5973 ;
  assign n15210 = ~n15208 & n15209 ;
  assign n15198 = ~n5191 & n5972 ;
  assign n15197 = n5191 & ~n5972 ;
  assign n15199 = n5329 & ~n15197 ;
  assign n15200 = ~n15198 & n15199 ;
  assign n15207 = ~n5175 & n5565 ;
  assign n15211 = ~n5175 & ~n5190 ;
  assign n15212 = ~n5529 & n5563 ;
  assign n15213 = ~n15211 & n15212 ;
  assign n15214 = ~n15207 & ~n15213 ;
  assign n15215 = ~n15200 & n15214 ;
  assign n15216 = ~n15210 & n15215 ;
  assign n15217 = ~n15206 & n15216 ;
  assign n15218 = n7453 & ~n15217 ;
  assign n15219 = ~n5175 & n5574 ;
  assign n15220 = ~n15218 & ~n15219 ;
  assign n15221 = n8899 & ~n15220 ;
  assign n15222 = n8899 & n10415 ;
  assign n15223 = ~n15206 & n15222 ;
  assign n15224 = \P2_reg3_reg[1]/NET0131  & ~n15223 ;
  assign n15225 = ~n15221 & ~n15224 ;
  assign n15226 = \P1_reg3_reg[1]/NET0131  & ~n6078 ;
  assign n15227 = \P1_reg3_reg[1]/NET0131  & n6095 ;
  assign n15229 = \P1_reg3_reg[1]/NET0131  & ~n6568 ;
  assign n15239 = n3364 & ~n6286 ;
  assign n15240 = ~n6287 & ~n15239 ;
  assign n15241 = ~n2713 & ~n15240 ;
  assign n15242 = n2713 & n3687 ;
  assign n15243 = ~n15241 & ~n15242 ;
  assign n15244 = n6568 & n15243 ;
  assign n15245 = ~n15229 & ~n15244 ;
  assign n15246 = n4011 & ~n15245 ;
  assign n15230 = n3721 & ~n6136 ;
  assign n15231 = ~n3721 & n6136 ;
  assign n15232 = ~n15230 & ~n15231 ;
  assign n15233 = ~n3694 & ~n15232 ;
  assign n15234 = n3694 & ~n3721 ;
  assign n15235 = ~n15233 & ~n15234 ;
  assign n15236 = n6568 & ~n15235 ;
  assign n15237 = ~n15229 & ~n15236 ;
  assign n15238 = n6282 & ~n15237 ;
  assign n15247 = n6568 & n15232 ;
  assign n15248 = ~n15229 & ~n15247 ;
  assign n15249 = n6207 & ~n15248 ;
  assign n15251 = ~n3718 & n6365 ;
  assign n15252 = ~n3694 & ~n3718 ;
  assign n15253 = ~n6328 & n6359 ;
  assign n15254 = ~n15252 & n15253 ;
  assign n15255 = ~n15251 & ~n15254 ;
  assign n15256 = n6568 & ~n15255 ;
  assign n15228 = \P1_reg3_reg[1]/NET0131  & ~n12757 ;
  assign n15250 = ~n3718 & n4112 ;
  assign n15257 = ~n15228 & ~n15250 ;
  assign n15258 = ~n15256 & n15257 ;
  assign n15259 = ~n15249 & n15258 ;
  assign n15260 = ~n15238 & n15259 ;
  assign n15261 = ~n15246 & n15260 ;
  assign n15262 = n6097 & ~n15261 ;
  assign n15263 = ~n15227 & ~n15262 ;
  assign n15264 = \P1_state_reg[0]/NET0131  & ~n15263 ;
  assign n15265 = ~n15226 & ~n15264 ;
  assign n15266 = n9533 & ~n15217 ;
  assign n15267 = \P2_reg0_reg[1]/NET0131  & ~n13732 ;
  assign n15268 = ~n15266 & ~n15267 ;
  assign n15269 = n8913 & ~n15217 ;
  assign n15270 = n6394 & n8913 ;
  assign n15271 = \P2_reg1_reg[1]/NET0131  & ~n15270 ;
  assign n15272 = ~n15269 & ~n15271 ;
  assign n15273 = \P2_reg2_reg[2]/NET0131  & ~n5589 ;
  assign n15274 = \P2_reg2_reg[2]/NET0131  & n5585 ;
  assign n15277 = n4219 & ~n15076 ;
  assign n15275 = \P2_reg2_reg[2]/NET0131  & ~n9772 ;
  assign n15276 = \P2_reg3_reg[2]/NET0131  & n5574 ;
  assign n15278 = ~n15275 & ~n15276 ;
  assign n15279 = ~n15277 & n15278 ;
  assign n15280 = n5583 & ~n15279 ;
  assign n15281 = ~n15274 & ~n15280 ;
  assign n15282 = \P1_state_reg[0]/NET0131  & ~n15281 ;
  assign n15283 = ~n15273 & ~n15282 ;
  assign n15289 = \P1_reg0_reg[1]/NET0131  & ~n6409 ;
  assign n15290 = n9829 & n15243 ;
  assign n15291 = ~n15289 & ~n15290 ;
  assign n15292 = n4011 & ~n15291 ;
  assign n15284 = n6282 & ~n15235 ;
  assign n15285 = n6207 & n15232 ;
  assign n15286 = n15255 & ~n15285 ;
  assign n15287 = ~n15284 & n15286 ;
  assign n15288 = n9829 & ~n15287 ;
  assign n15293 = ~n6409 & ~n8656 ;
  assign n15294 = n11119 & ~n15293 ;
  assign n15295 = \P1_reg0_reg[1]/NET0131  & ~n15294 ;
  assign n15296 = ~n15288 & ~n15295 ;
  assign n15297 = ~n15292 & n15296 ;
  assign n15298 = \P3_reg0_reg[1]/NET0131  & ~n2143 ;
  assign n15299 = \P3_reg0_reg[1]/NET0131  & n2145 ;
  assign n15307 = \P3_reg0_reg[1]/NET0131  & ~n2236 ;
  assign n15310 = n2236 & ~n15004 ;
  assign n15311 = ~n15307 & ~n15310 ;
  assign n15312 = n737 & ~n15311 ;
  assign n15302 = \P3_reg0_reg[1]/NET0131  & ~n2163 ;
  assign n15303 = n2163 & n15009 ;
  assign n15304 = ~n15302 & ~n15303 ;
  assign n15305 = n2234 & ~n15304 ;
  assign n15300 = ~n1891 & n2285 ;
  assign n15301 = n2163 & n15300 ;
  assign n15306 = \P3_reg0_reg[1]/NET0131  & ~n2287 ;
  assign n15315 = ~n15301 & ~n15306 ;
  assign n15316 = ~n15305 & n15315 ;
  assign n15308 = ~n14992 & ~n15307 ;
  assign n15309 = n2393 & ~n15308 ;
  assign n15313 = ~n14997 & ~n15302 ;
  assign n15314 = n2391 & ~n15313 ;
  assign n15317 = ~n15309 & ~n15314 ;
  assign n15318 = n15316 & n15317 ;
  assign n15319 = ~n15312 & n15318 ;
  assign n15320 = n2147 & ~n15319 ;
  assign n15321 = ~n15299 & ~n15320 ;
  assign n15322 = \P1_state_reg[0]/NET0131  & ~n15321 ;
  assign n15323 = ~n15298 & ~n15322 ;
  assign n15324 = \P3_reg1_reg[1]/NET0131  & ~n2143 ;
  assign n15325 = \P3_reg1_reg[1]/NET0131  & n2145 ;
  assign n15326 = \P3_reg1_reg[1]/NET0131  & ~n2427 ;
  assign n15339 = n2427 & ~n15004 ;
  assign n15340 = ~n15326 & ~n15339 ;
  assign n15341 = n737 & ~n15340 ;
  assign n15331 = ~n2518 & n15009 ;
  assign n15330 = n714 & n14991 ;
  assign n15332 = ~n15300 & ~n15330 ;
  assign n15333 = ~n15331 & n15332 ;
  assign n15334 = n2408 & ~n15333 ;
  assign n15327 = n2427 & n15009 ;
  assign n15328 = ~n15326 & ~n15327 ;
  assign n15329 = n2425 & ~n15328 ;
  assign n15335 = ~n714 & n2518 ;
  assign n15336 = ~n2408 & ~n15335 ;
  assign n15337 = n6449 & ~n15336 ;
  assign n15338 = \P3_reg1_reg[1]/NET0131  & ~n15337 ;
  assign n15342 = ~n15329 & ~n15338 ;
  assign n15343 = ~n15334 & n15342 ;
  assign n15344 = ~n15341 & n15343 ;
  assign n15345 = n2147 & ~n15344 ;
  assign n15346 = ~n15325 & ~n15345 ;
  assign n15347 = \P1_state_reg[0]/NET0131  & ~n15346 ;
  assign n15348 = ~n15324 & ~n15347 ;
  assign n15349 = \P3_reg2_reg[1]/NET0131  & ~n2143 ;
  assign n15350 = \P3_reg2_reg[1]/NET0131  & n2145 ;
  assign n15355 = \P3_reg2_reg[1]/NET0131  & ~n2408 ;
  assign n15359 = n2408 & ~n15004 ;
  assign n15360 = ~n15355 & ~n15359 ;
  assign n15361 = n737 & ~n15360 ;
  assign n15352 = \P3_reg2_reg[1]/NET0131  & ~n2427 ;
  assign n15353 = ~n15327 & ~n15352 ;
  assign n15354 = ~n2518 & ~n15353 ;
  assign n15366 = \P3_reg2_reg[1]/NET0131  & ~n2429 ;
  assign n15351 = n2427 & n15300 ;
  assign n15365 = \P3_reg3_reg[1]/NET0131  & n2283 ;
  assign n15367 = ~n15351 & ~n15365 ;
  assign n15368 = ~n15366 & n15367 ;
  assign n15369 = ~n15354 & n15368 ;
  assign n15356 = n2408 & n15009 ;
  assign n15357 = ~n15355 & ~n15356 ;
  assign n15358 = n2425 & ~n15357 ;
  assign n15362 = n2427 & n14991 ;
  assign n15363 = ~n15352 & ~n15362 ;
  assign n15364 = n714 & ~n15363 ;
  assign n15370 = ~n15358 & ~n15364 ;
  assign n15371 = n15369 & n15370 ;
  assign n15372 = ~n15361 & n15371 ;
  assign n15373 = n2147 & ~n15372 ;
  assign n15374 = ~n15350 & ~n15373 ;
  assign n15375 = \P1_state_reg[0]/NET0131  & ~n15374 ;
  assign n15376 = ~n15349 & ~n15375 ;
  assign n15378 = \P1_reg1_reg[1]/NET0131  & ~n6683 ;
  assign n15379 = n9045 & n15243 ;
  assign n15380 = ~n15378 & ~n15379 ;
  assign n15381 = n4011 & ~n15380 ;
  assign n15377 = n9045 & ~n15287 ;
  assign n15382 = \P1_reg1_reg[1]/NET0131  & ~n15056 ;
  assign n15383 = ~n15377 & ~n15382 ;
  assign n15384 = ~n15381 & n15383 ;
  assign n15385 = \P3_reg3_reg[0]/NET0131  & ~n2143 ;
  assign n15386 = \P3_reg3_reg[0]/NET0131  & n2145 ;
  assign n15393 = \P3_reg3_reg[0]/NET0131  & ~n2163 ;
  assign n15394 = n1877 & ~n2243 ;
  assign n15395 = ~n2239 & ~n2244 ;
  assign n15396 = ~n15394 & n15395 ;
  assign n15397 = n2163 & n15396 ;
  assign n15398 = ~n15393 & ~n15397 ;
  assign n15399 = n737 & ~n15398 ;
  assign n15389 = ~n1908 & ~n1965 ;
  assign n15400 = n2163 & ~n15389 ;
  assign n15401 = ~n15393 & ~n15400 ;
  assign n15402 = n2393 & ~n15401 ;
  assign n15388 = \P3_reg3_reg[0]/NET0131  & ~n2236 ;
  assign n15390 = n2236 & ~n15389 ;
  assign n15391 = ~n15388 & ~n15390 ;
  assign n15392 = ~n12212 & ~n15391 ;
  assign n15403 = n1907 & n2236 ;
  assign n15404 = ~n15388 & ~n15403 ;
  assign n15405 = n2285 & ~n15404 ;
  assign n15387 = \P3_reg3_reg[0]/NET0131  & n710 ;
  assign n15406 = n1907 & n2283 ;
  assign n15407 = ~n15387 & ~n15406 ;
  assign n15408 = ~n15405 & n15407 ;
  assign n15409 = ~n15392 & n15408 ;
  assign n15410 = ~n15402 & n15409 ;
  assign n15411 = ~n15399 & n15410 ;
  assign n15412 = n2147 & ~n15411 ;
  assign n15413 = ~n15386 & ~n15412 ;
  assign n15414 = \P1_state_reg[0]/NET0131  & ~n15413 ;
  assign n15415 = ~n15385 & ~n15414 ;
  assign n15416 = \P1_reg2_reg[1]/NET0131  & ~n6078 ;
  assign n15417 = \P1_reg2_reg[1]/NET0131  & n6095 ;
  assign n15419 = \P1_reg2_reg[1]/NET0131  & ~n6113 ;
  assign n15423 = n6113 & n15243 ;
  assign n15424 = ~n15419 & ~n15423 ;
  assign n15425 = n4011 & ~n15424 ;
  assign n15420 = n6113 & ~n15235 ;
  assign n15421 = ~n15419 & ~n15420 ;
  assign n15422 = n6282 & ~n15421 ;
  assign n15426 = n6113 & n15232 ;
  assign n15427 = ~n15419 & ~n15426 ;
  assign n15428 = n6207 & ~n15427 ;
  assign n15430 = \P1_reg2_reg[1]/NET0131  & ~n11834 ;
  assign n15418 = n6113 & ~n15255 ;
  assign n15429 = \P1_reg3_reg[1]/NET0131  & n4112 ;
  assign n15431 = ~n15418 & ~n15429 ;
  assign n15432 = ~n15430 & n15431 ;
  assign n15433 = ~n15428 & n15432 ;
  assign n15434 = ~n15422 & n15433 ;
  assign n15435 = ~n15425 & n15434 ;
  assign n15436 = n6097 & ~n15435 ;
  assign n15437 = ~n15417 & ~n15436 ;
  assign n15438 = \P1_state_reg[0]/NET0131  & ~n15437 ;
  assign n15439 = ~n15416 & ~n15438 ;
  assign n15440 = n4219 & ~n15217 ;
  assign n15441 = \P2_reg3_reg[1]/NET0131  & n5574 ;
  assign n15442 = ~n15440 & ~n15441 ;
  assign n15443 = n8899 & ~n15442 ;
  assign n15444 = n4219 & ~n15205 ;
  assign n15445 = n5383 & ~n15444 ;
  assign n15446 = n13807 & ~n15445 ;
  assign n15447 = \P2_reg2_reg[1]/NET0131  & ~n15446 ;
  assign n15448 = ~n15443 & ~n15447 ;
  assign n15449 = \P3_reg0_reg[0]/NET0131  & ~n2143 ;
  assign n15450 = \P3_reg0_reg[0]/NET0131  & n2145 ;
  assign n15456 = \P3_reg0_reg[0]/NET0131  & ~n2236 ;
  assign n15459 = n2236 & n15396 ;
  assign n15460 = ~n15456 & ~n15459 ;
  assign n15461 = n737 & ~n15460 ;
  assign n15452 = \P3_reg0_reg[0]/NET0131  & ~n2163 ;
  assign n15462 = ~n15400 & ~n15452 ;
  assign n15463 = ~n12212 & ~n15462 ;
  assign n15457 = ~n15390 & ~n15456 ;
  assign n15458 = n2393 & ~n15457 ;
  assign n15451 = \P3_reg0_reg[0]/NET0131  & ~n2284 ;
  assign n15453 = n1907 & n2163 ;
  assign n15454 = ~n15452 & ~n15453 ;
  assign n15455 = n2285 & ~n15454 ;
  assign n15464 = ~n15451 & ~n15455 ;
  assign n15465 = ~n15458 & n15464 ;
  assign n15466 = ~n15463 & n15465 ;
  assign n15467 = ~n15461 & n15466 ;
  assign n15468 = n2147 & ~n15467 ;
  assign n15469 = ~n15450 & ~n15468 ;
  assign n15470 = \P1_state_reg[0]/NET0131  & ~n15469 ;
  assign n15471 = ~n15449 & ~n15470 ;
  assign n15472 = \P3_reg1_reg[0]/NET0131  & ~n2143 ;
  assign n15473 = \P3_reg1_reg[0]/NET0131  & n2145 ;
  assign n15482 = \P3_reg1_reg[0]/NET0131  & ~n2427 ;
  assign n15483 = n2427 & n15396 ;
  assign n15484 = ~n15482 & ~n15483 ;
  assign n15485 = n737 & ~n15484 ;
  assign n15486 = n2427 & ~n15389 ;
  assign n15487 = ~n15482 & ~n15486 ;
  assign n15488 = n2425 & ~n15487 ;
  assign n15475 = \P3_reg1_reg[0]/NET0131  & ~n2408 ;
  assign n15479 = n2408 & ~n15389 ;
  assign n15480 = ~n15475 & ~n15479 ;
  assign n15481 = ~n15335 & ~n15480 ;
  assign n15474 = \P3_reg1_reg[0]/NET0131  & ~n2284 ;
  assign n15476 = n1907 & n2408 ;
  assign n15477 = ~n15475 & ~n15476 ;
  assign n15478 = n2285 & ~n15477 ;
  assign n15489 = ~n15474 & ~n15478 ;
  assign n15490 = ~n15481 & n15489 ;
  assign n15491 = ~n15488 & n15490 ;
  assign n15492 = ~n15485 & n15491 ;
  assign n15493 = n2147 & ~n15492 ;
  assign n15494 = ~n15473 & ~n15493 ;
  assign n15495 = \P1_state_reg[0]/NET0131  & ~n15494 ;
  assign n15496 = ~n15472 & ~n15495 ;
  assign n15497 = \P3_reg2_reg[0]/NET0131  & ~n2143 ;
  assign n15498 = \P3_reg2_reg[0]/NET0131  & n2145 ;
  assign n15503 = \P3_reg2_reg[0]/NET0131  & ~n2408 ;
  assign n15504 = n2408 & n15396 ;
  assign n15505 = ~n15503 & ~n15504 ;
  assign n15506 = n737 & ~n15505 ;
  assign n15507 = ~n15479 & ~n15503 ;
  assign n15508 = n2425 & ~n15507 ;
  assign n15500 = \P3_reg2_reg[0]/NET0131  & ~n2427 ;
  assign n15501 = ~n15486 & ~n15500 ;
  assign n15502 = ~n15335 & ~n15501 ;
  assign n15509 = n1907 & n2427 ;
  assign n15510 = ~n15500 & ~n15509 ;
  assign n15511 = n2285 & ~n15510 ;
  assign n15499 = \P3_reg3_reg[0]/NET0131  & n2283 ;
  assign n15512 = \P3_reg2_reg[0]/NET0131  & n710 ;
  assign n15513 = ~n15499 & ~n15512 ;
  assign n15514 = ~n15511 & n15513 ;
  assign n15515 = ~n15502 & n15514 ;
  assign n15516 = ~n15508 & n15515 ;
  assign n15517 = ~n15506 & n15516 ;
  assign n15518 = n2147 & ~n15517 ;
  assign n15519 = ~n15498 & ~n15518 ;
  assign n15520 = \P1_state_reg[0]/NET0131  & ~n15519 ;
  assign n15521 = ~n15497 & ~n15520 ;
  assign n15522 = ~n3694 & n4112 ;
  assign n15525 = n3704 & ~n6285 ;
  assign n15526 = ~n2713 & ~n6286 ;
  assign n15527 = ~n15525 & n15526 ;
  assign n15528 = n4011 & n15527 ;
  assign n15523 = ~n3694 & n6693 ;
  assign n15524 = ~n3697 & ~n8656 ;
  assign n15529 = ~n15523 & ~n15524 ;
  assign n15530 = ~n15528 & n15529 ;
  assign n15531 = n6568 & ~n15530 ;
  assign n15532 = ~n15522 & ~n15531 ;
  assign n15533 = n9044 & ~n15532 ;
  assign n15534 = ~n4011 & ~n6693 ;
  assign n15535 = n8656 & n15534 ;
  assign n15536 = ~n6568 & ~n15535 ;
  assign n15537 = n10960 & ~n15536 ;
  assign n15538 = \P1_reg3_reg[0]/NET0131  & ~n15537 ;
  assign n15539 = ~n15533 & ~n15538 ;
  assign n15540 = \P2_reg3_reg[0]/NET0131  & ~n5589 ;
  assign n15541 = \P2_reg3_reg[0]/NET0131  & n5585 ;
  assign n15543 = \P2_reg3_reg[0]/NET0131  & ~n7453 ;
  assign n15551 = n5161 & ~n5346 ;
  assign n15552 = ~n4231 & ~n5347 ;
  assign n15553 = ~n15551 & n15552 ;
  assign n15554 = n7453 & n15553 ;
  assign n15555 = ~n15543 & ~n15554 ;
  assign n15556 = n5383 & ~n15555 ;
  assign n15547 = ~n5419 & ~n5919 ;
  assign n15548 = n7453 & ~n15547 ;
  assign n15549 = ~n15543 & ~n15548 ;
  assign n15550 = ~n8884 & ~n15549 ;
  assign n15544 = ~n5190 & n7453 ;
  assign n15545 = ~n15543 & ~n15544 ;
  assign n15546 = ~n6395 & ~n15545 ;
  assign n15542 = \P2_reg3_reg[0]/NET0131  & n5568 ;
  assign n15557 = ~n5190 & n5574 ;
  assign n15558 = ~n15542 & ~n15557 ;
  assign n15559 = ~n15546 & n15558 ;
  assign n15560 = ~n15550 & n15559 ;
  assign n15561 = ~n15556 & n15560 ;
  assign n15562 = n5583 & ~n15561 ;
  assign n15563 = ~n15541 & ~n15562 ;
  assign n15564 = \P1_state_reg[0]/NET0131  & ~n15563 ;
  assign n15565 = ~n15540 & ~n15564 ;
  assign n15566 = \P1_reg2_reg[0]/NET0131  & ~n6078 ;
  assign n15567 = \P1_reg2_reg[0]/NET0131  & n6095 ;
  assign n15568 = n6113 & ~n15530 ;
  assign n15569 = \P1_reg3_reg[0]/NET0131  & n4112 ;
  assign n15570 = ~n6113 & ~n15535 ;
  assign n15571 = ~n6361 & ~n15570 ;
  assign n15572 = \P1_reg2_reg[0]/NET0131  & ~n15571 ;
  assign n15573 = ~n15569 & ~n15572 ;
  assign n15574 = ~n15568 & n15573 ;
  assign n15575 = n6097 & ~n15574 ;
  assign n15576 = ~n15567 & ~n15575 ;
  assign n15577 = \P1_state_reg[0]/NET0131  & ~n15576 ;
  assign n15578 = ~n15566 & ~n15577 ;
  assign n15579 = \P2_reg1_reg[0]/NET0131  & ~n8902 ;
  assign n15581 = n5383 & n15553 ;
  assign n15580 = ~n8884 & ~n15547 ;
  assign n15582 = ~n5190 & ~n6395 ;
  assign n15583 = ~n15580 & ~n15582 ;
  assign n15584 = ~n15581 & n15583 ;
  assign n15585 = n8913 & ~n15584 ;
  assign n15586 = ~n15579 & ~n15585 ;
  assign n15588 = \P1_reg0_reg[0]/NET0131  & ~n6409 ;
  assign n15589 = n6409 & n15527 ;
  assign n15590 = ~n15588 & ~n15589 ;
  assign n15591 = n4011 & ~n15590 ;
  assign n15592 = ~n3697 & n6409 ;
  assign n15593 = ~n15588 & ~n15592 ;
  assign n15594 = ~n8656 & ~n15593 ;
  assign n15587 = n6409 & n15523 ;
  assign n15595 = \P1_reg0_reg[0]/NET0131  & ~n11118 ;
  assign n15596 = ~n15587 & ~n15595 ;
  assign n15597 = ~n15594 & n15596 ;
  assign n15598 = ~n15591 & n15597 ;
  assign n15599 = n6097 & ~n15598 ;
  assign n15600 = \P1_reg0_reg[0]/NET0131  & n6095 ;
  assign n15601 = ~n15599 & ~n15600 ;
  assign n15602 = \P1_state_reg[0]/NET0131  & ~n15601 ;
  assign n15603 = \P1_reg0_reg[0]/NET0131  & ~n6078 ;
  assign n15604 = ~n15602 & ~n15603 ;
  assign n15605 = \P2_reg3_reg[0]/NET0131  & n5574 ;
  assign n15606 = n4219 & ~n15584 ;
  assign n15607 = ~n15605 & ~n15606 ;
  assign n15608 = n8899 & ~n15607 ;
  assign n15609 = \P2_reg2_reg[0]/NET0131  & ~n9773 ;
  assign n15610 = ~n15608 & ~n15609 ;
  assign n15612 = \P1_reg1_reg[0]/NET0131  & ~n6683 ;
  assign n15613 = n6683 & n15527 ;
  assign n15614 = ~n15612 & ~n15613 ;
  assign n15615 = n4011 & ~n15614 ;
  assign n15616 = ~n3697 & n6683 ;
  assign n15617 = ~n15612 & ~n15616 ;
  assign n15618 = ~n8656 & ~n15617 ;
  assign n15611 = n6683 & n15523 ;
  assign n15619 = \P1_reg1_reg[0]/NET0131  & ~n6695 ;
  assign n15620 = ~n15611 & ~n15619 ;
  assign n15621 = ~n15618 & n15620 ;
  assign n15622 = ~n15615 & n15621 ;
  assign n15623 = n6097 & ~n15622 ;
  assign n15624 = \P1_reg1_reg[0]/NET0131  & n6095 ;
  assign n15625 = ~n15623 & ~n15624 ;
  assign n15626 = \P1_state_reg[0]/NET0131  & ~n15625 ;
  assign n15627 = \P1_reg1_reg[0]/NET0131  & ~n6078 ;
  assign n15628 = ~n15626 & ~n15627 ;
  assign n15629 = \P2_reg0_reg[0]/NET0131  & ~n13732 ;
  assign n15630 = n9533 & ~n15584 ;
  assign n15631 = ~n15629 & ~n15630 ;
  assign n15632 = n1318 & n2289 ;
  assign n15634 = n1336 & ~n2273 ;
  assign n15633 = n1944 & n2272 ;
  assign n15635 = n2242 & ~n15633 ;
  assign n15636 = ~n15634 & n15635 ;
  assign n15637 = n737 & n2236 ;
  assign n15638 = n15636 & n15637 ;
  assign n15639 = ~n15632 & ~n15638 ;
  assign n15640 = ~n757 & n2143 ;
  assign n15641 = ~n15639 & n15640 ;
  assign n15642 = ~n737 & ~n2393 ;
  assign n15643 = ~n2236 & ~n15642 ;
  assign n15644 = n15640 & ~n15643 ;
  assign n15645 = n12214 & n15644 ;
  assign n15646 = \P3_reg0_reg[30]/NET0131  & ~n15645 ;
  assign n15647 = ~n15641 & ~n15646 ;
  assign n15648 = n1367 & n2285 ;
  assign n15649 = n2163 & n15648 ;
  assign n15650 = ~n15638 & ~n15649 ;
  assign n15651 = n15640 & ~n15650 ;
  assign n15652 = n15645 & ~n15648 ;
  assign n15653 = \P3_reg0_reg[31]/NET0131  & ~n15652 ;
  assign n15654 = ~n15651 & ~n15653 ;
  assign n15655 = n1318 & n6451 ;
  assign n15656 = n737 & n2427 ;
  assign n15657 = n15636 & n15656 ;
  assign n15658 = ~n15655 & ~n15657 ;
  assign n15659 = n15640 & ~n15658 ;
  assign n15660 = ~n737 & ~n2425 ;
  assign n15661 = ~n2427 & ~n15660 ;
  assign n15662 = n15640 & ~n15661 ;
  assign n15663 = n15337 & n15662 ;
  assign n15664 = \P3_reg1_reg[30]/NET0131  & ~n15663 ;
  assign n15665 = ~n15659 & ~n15664 ;
  assign n15666 = n1367 & n6451 ;
  assign n15667 = ~n15657 & ~n15666 ;
  assign n15668 = n15640 & ~n15667 ;
  assign n15669 = \P3_reg1_reg[31]/NET0131  & ~n15663 ;
  assign n15670 = ~n15668 & ~n15669 ;
  assign n15677 = n737 & n2408 ;
  assign n15678 = n15636 & n15677 ;
  assign n15679 = ~n6513 & ~n15678 ;
  assign n15680 = n15640 & ~n15679 ;
  assign n15671 = ~n2408 & ~n15660 ;
  assign n15672 = n15640 & ~n15671 ;
  assign n15673 = ~n2427 & ~n15335 ;
  assign n15674 = ~n710 & ~n15673 ;
  assign n15675 = n15672 & n15674 ;
  assign n15676 = \P3_reg2_reg[30]/NET0131  & ~n15675 ;
  assign n15681 = \P3_reg2_reg[30]/NET0131  & ~n2427 ;
  assign n15682 = n2427 & n15640 ;
  assign n15683 = n1318 & n15682 ;
  assign n15684 = ~n15681 & ~n15683 ;
  assign n15685 = n2285 & ~n15684 ;
  assign n15686 = ~n15676 & ~n15685 ;
  assign n15687 = ~n15680 & n15686 ;
  assign n15688 = ~n688 & ~n2424 ;
  assign n15689 = ~n2282 & n15688 ;
  assign n15690 = ~n2427 & n15689 ;
  assign n15691 = ~n710 & ~n15690 ;
  assign n15692 = n15672 & n15691 ;
  assign n15693 = \P3_reg2_reg[31]/NET0131  & ~n15692 ;
  assign n15694 = \P3_reg2_reg[31]/NET0131  & ~n2427 ;
  assign n15695 = n1367 & n15682 ;
  assign n15696 = ~n15694 & ~n15695 ;
  assign n15697 = n2285 & ~n15696 ;
  assign n15698 = ~n15693 & ~n15697 ;
  assign n15699 = ~n15680 & n15698 ;
  assign n15700 = ~\P1_state_reg[0]/NET0131  & ~n4612 ;
  assign n15701 = \P1_state_reg[0]/NET0131  & ~n4197 ;
  assign n15702 = ~n15700 & ~n15701 ;
  assign n15703 = ~\P1_state_reg[0]/NET0131  & ~n4591 ;
  assign n15704 = \P1_state_reg[0]/NET0131  & ~n4205 ;
  assign n15705 = ~n15703 & ~n15704 ;
  assign n15706 = ~\P1_state_reg[0]/NET0131  & ~n4542 ;
  assign n15707 = \P1_state_reg[0]/NET0131  & n4225 ;
  assign n15708 = ~n15706 & ~n15707 ;
  assign n15709 = \P1_state_reg[0]/NET0131  & ~n745 ;
  assign n15710 = ~\P1_state_reg[0]/NET0131  & n1261 ;
  assign n15711 = ~n15709 & ~n15710 ;
  assign n15712 = \P1_state_reg[0]/NET0131  & n752 ;
  assign n15713 = ~\P1_state_reg[0]/NET0131  & n1464 ;
  assign n15714 = ~n15712 & ~n15713 ;
  assign n15715 = \P1_state_reg[0]/NET0131  & n724 ;
  assign n15716 = ~\P1_state_reg[0]/NET0131  & n1435 ;
  assign n15717 = ~n15715 & ~n15716 ;
  assign n15718 = \P1_state_reg[0]/NET0131  & ~n6087 ;
  assign n15719 = ~\P1_state_reg[0]/NET0131  & n3164 ;
  assign n15720 = ~n15718 & ~n15719 ;
  assign n15721 = ~\P1_state_reg[0]/NET0131  & ~n3426 ;
  assign n15722 = \P1_state_reg[0]/NET0131  & n2725 ;
  assign n15723 = ~n15721 & ~n15722 ;
  assign n15724 = ~\P1_state_reg[0]/NET0131  & ~n3517 ;
  assign n15725 = \P1_state_reg[0]/NET0131  & ~n6082 ;
  assign n15726 = ~n15724 & ~n15725 ;
  assign n15727 = ~\P1_state_reg[0]/NET0131  & ~n5894 ;
  assign n15728 = \P1_state_reg[0]/NET0131  & n4378 ;
  assign n15729 = ~n15727 & ~n15728 ;
  assign n15730 = \P1_state_reg[0]/NET0131  & ~n4735 ;
  assign n15731 = ~\P1_state_reg[0]/NET0131  & n4743 ;
  assign n15732 = ~n15730 & ~n15731 ;
  assign n15733 = \P1_state_reg[0]/NET0131  & ~n5012 ;
  assign n15734 = ~\P1_state_reg[0]/NET0131  & n5020 ;
  assign n15735 = ~n15733 & ~n15734 ;
  assign n15736 = ~\P1_state_reg[0]/NET0131  & ~n5048 ;
  assign n15737 = \P1_state_reg[0]/NET0131  & n5056 ;
  assign n15738 = ~n15736 & ~n15737 ;
  assign n15739 = \P1_state_reg[0]/NET0131  & ~n4963 ;
  assign n15740 = ~\P1_state_reg[0]/NET0131  & n4971 ;
  assign n15741 = ~n15739 & ~n15740 ;
  assign n15742 = \P1_state_reg[0]/NET0131  & ~n4938 ;
  assign n15743 = ~\P1_state_reg[0]/NET0131  & n4946 ;
  assign n15744 = ~n15742 & ~n15743 ;
  assign n15745 = \P1_state_reg[0]/NET0131  & ~n4779 ;
  assign n15746 = ~\P1_state_reg[0]/NET0131  & n4787 ;
  assign n15747 = ~n15745 & ~n15746 ;
  assign n15748 = ~\P1_state_reg[0]/NET0131  & ~n4890 ;
  assign n15749 = \P1_state_reg[0]/NET0131  & ~n4882 ;
  assign n15750 = ~n15748 & ~n15749 ;
  assign n15751 = \P1_state_reg[0]/NET0131  & n5326 ;
  assign n15752 = ~\P1_state_reg[0]/NET0131  & n4693 ;
  assign n15753 = ~n15751 & ~n15752 ;
  assign n15754 = ~\P1_state_reg[0]/NET0131  & ~n4865 ;
  assign n15755 = \P1_state_reg[0]/NET0131  & ~n4857 ;
  assign n15756 = ~n15754 & ~n15755 ;
  assign n15757 = \P1_state_reg[0]/NET0131  & ~n4385 ;
  assign n15758 = ~\P1_state_reg[0]/NET0131  & n4370 ;
  assign n15759 = ~n15757 & ~n15758 ;
  assign n15760 = ~\P1_state_reg[0]/NET0131  & ~n4991 ;
  assign n15761 = \P1_state_reg[0]/NET0131  & ~n4995 ;
  assign n15762 = ~n15760 & ~n15761 ;
  assign n15763 = \P1_state_reg[0]/NET0131  & ~n4833 ;
  assign n15764 = ~\P1_state_reg[0]/NET0131  & n4841 ;
  assign n15765 = ~n15763 & ~n15764 ;
  assign n15766 = \P1_state_reg[0]/NET0131  & ~n4907 ;
  assign n15767 = ~\P1_state_reg[0]/NET0131  & n4916 ;
  assign n15768 = ~n15766 & ~n15767 ;
  assign n15769 = \P1_state_reg[0]/NET0131  & ~n4804 ;
  assign n15770 = ~\P1_state_reg[0]/NET0131  & n4812 ;
  assign n15771 = ~n15769 & ~n15770 ;
  assign n15772 = \P1_state_reg[0]/NET0131  & ~n5322 ;
  assign n15773 = ~\P1_state_reg[0]/NET0131  & n4753 ;
  assign n15774 = ~n15772 & ~n15773 ;
  assign n15775 = \P1_state_reg[0]/NET0131  & ~n5311 ;
  assign n15776 = ~\P1_state_reg[0]/NET0131  & n4674 ;
  assign n15777 = ~n15775 & ~n15776 ;
  assign n15778 = ~\P1_state_reg[0]/NET0131  & n4655 ;
  assign n15779 = ~n5589 & ~n15778 ;
  assign n15780 = ~\P1_state_reg[0]/NET0131  & ~n4634 ;
  assign n15781 = \P1_state_reg[0]/NET0131  & n4190 ;
  assign n15782 = ~n15780 & ~n15781 ;
  assign n15783 = ~\P1_state_reg[0]/NET0131  & ~n4486 ;
  assign n15784 = \P1_state_reg[0]/NET0131  & n4231 ;
  assign n15785 = ~n15783 & ~n15784 ;
  assign n15786 = ~\P1_state_reg[0]/NET0131  & ~n5146 ;
  assign n15787 = \P1_state_reg[0]/NET0131  & n5151 ;
  assign n15788 = ~n15786 & ~n15787 ;
  assign n15789 = ~\P1_state_reg[0]/NET0131  & ~n5233 ;
  assign n15790 = \P1_state_reg[0]/NET0131  & n5238 ;
  assign n15791 = ~n15789 & ~n15790 ;
  assign n15792 = \P1_state_reg[0]/NET0131  & ~n5207 ;
  assign n15793 = ~\P1_state_reg[0]/NET0131  & n5216 ;
  assign n15794 = ~n15792 & ~n15793 ;
  assign n15795 = ~\P1_state_reg[0]/NET0131  & ~n5129 ;
  assign n15796 = \P1_state_reg[0]/NET0131  & n5121 ;
  assign n15797 = ~n15795 & ~n15796 ;
  assign n15798 = \P1_state_reg[0]/NET0131  & ~n5096 ;
  assign n15799 = ~\P1_state_reg[0]/NET0131  & n5105 ;
  assign n15800 = ~n15798 & ~n15799 ;
  assign n15801 = ~\P1_state_reg[0]/NET0131  & ~n5075 ;
  assign n15802 = \P1_state_reg[0]/NET0131  & n5079 ;
  assign n15803 = ~n15801 & ~n15802 ;
  assign n15804 = \P1_state_reg[0]/NET0131  & ~n5165 ;
  assign n15805 = ~\P1_state_reg[0]/NET0131  & n5173 ;
  assign n15806 = ~n15804 & ~n15805 ;
  assign n15807 = ~\P1_state_reg[0]/NET0131  & ~n5878 ;
  assign n15808 = \P1_state_reg[0]/NET0131  & ~\P2_IR_reg[27]/NET0131  ;
  assign n15809 = ~\P2_IR_reg[30]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n15810 = n15808 & n15809 ;
  assign n15811 = n4372 & n15810 ;
  assign n15812 = n4221 & n15811 ;
  assign n15813 = ~n15807 & ~n15812 ;
  assign n15814 = ~\P1_state_reg[0]/NET0131  & ~n885 ;
  assign n15815 = ~n765 & ~n15814 ;
  assign n15816 = ~\P1_state_reg[0]/NET0131  & ~n1644 ;
  assign n15817 = \P1_state_reg[0]/NET0131  & n1649 ;
  assign n15818 = ~n15816 & ~n15817 ;
  assign n15819 = ~\P1_state_reg[0]/NET0131  & ~n1620 ;
  assign n15820 = \P1_state_reg[0]/NET0131  & n1625 ;
  assign n15821 = ~n15819 & ~n15820 ;
  assign n15822 = \P1_state_reg[0]/NET0131  & ~n1574 ;
  assign n15823 = ~\P1_state_reg[0]/NET0131  & n1582 ;
  assign n15824 = ~n15822 & ~n15823 ;
  assign n15825 = ~\P1_state_reg[0]/NET0131  & ~n1553 ;
  assign n15826 = \P1_state_reg[0]/NET0131  & n1558 ;
  assign n15827 = ~n15825 & ~n15826 ;
  assign n15828 = ~\P1_state_reg[0]/NET0131  & ~n1538 ;
  assign n15829 = \P1_state_reg[0]/NET0131  & n1542 ;
  assign n15830 = ~n15828 & ~n15829 ;
  assign n15831 = \P1_state_reg[0]/NET0131  & ~n1502 ;
  assign n15832 = ~\P1_state_reg[0]/NET0131  & ~n1510 ;
  assign n15833 = ~n15831 & ~n15832 ;
  assign n15834 = ~\P1_state_reg[0]/NET0131  & ~n1177 ;
  assign n15835 = \P1_state_reg[0]/NET0131  & n1183 ;
  assign n15836 = ~n15834 & ~n15835 ;
  assign n15837 = ~\P1_state_reg[0]/NET0131  & ~n1159 ;
  assign n15838 = \P1_state_reg[0]/NET0131  & ~n1164 ;
  assign n15839 = ~n15837 & ~n15838 ;
  assign n15840 = ~\P1_state_reg[0]/NET0131  & ~n1128 ;
  assign n15841 = \P1_state_reg[0]/NET0131  & n1135 ;
  assign n15842 = ~n15840 & ~n15841 ;
  assign n15843 = ~\P1_state_reg[0]/NET0131  & ~n1104 ;
  assign n15844 = \P1_state_reg[0]/NET0131  & n1108 ;
  assign n15845 = ~n15843 & ~n15844 ;
  assign n15846 = \P1_state_reg[0]/NET0131  & ~n1881 ;
  assign n15847 = ~\P1_state_reg[0]/NET0131  & ~n1889 ;
  assign n15848 = ~n15846 & ~n15847 ;
  assign n15849 = ~\P1_state_reg[0]/NET0131  & ~n1062 ;
  assign n15850 = \P1_state_reg[0]/NET0131  & n708 ;
  assign n15851 = ~n15849 & ~n15850 ;
  assign n15852 = ~\P1_state_reg[0]/NET0131  & ~n1028 ;
  assign n15853 = \P1_state_reg[0]/NET0131  & n701 ;
  assign n15854 = ~n15852 & ~n15853 ;
  assign n15855 = ~\P1_state_reg[0]/NET0131  & ~n990 ;
  assign n15856 = \P1_state_reg[0]/NET0131  & n687 ;
  assign n15857 = ~n15855 & ~n15856 ;
  assign n15858 = ~\P1_state_reg[0]/NET0131  & ~n1222 ;
  assign n15859 = \P1_state_reg[0]/NET0131  & n755 ;
  assign n15860 = ~n15858 & ~n15859 ;
  assign n15861 = ~\P1_state_reg[0]/NET0131  & ~n1407 ;
  assign n15862 = \P1_state_reg[0]/NET0131  & n733 ;
  assign n15863 = ~n15861 & ~n15862 ;
  assign n15864 = \P1_state_reg[0]/NET0131  & ~n894 ;
  assign n15865 = ~\P1_state_reg[0]/NET0131  & n1384 ;
  assign n15866 = ~n15864 & ~n15865 ;
  assign n15867 = ~\P1_state_reg[0]/NET0131  & ~n1837 ;
  assign n15868 = \P1_state_reg[0]/NET0131  & n1842 ;
  assign n15869 = ~n15867 & ~n15868 ;
  assign n15870 = \P1_state_reg[0]/NET0131  & ~n900 ;
  assign n15871 = ~\P1_state_reg[0]/NET0131  & n1317 ;
  assign n15872 = ~n15870 & ~n15871 ;
  assign n15873 = ~\P1_state_reg[0]/NET0131  & ~n1366 ;
  assign n15874 = \P1_state_reg[0]/NET0131  & ~\P3_IR_reg[29]/NET0131  ;
  assign n15875 = ~\P3_IR_reg[30]/NET0131  & \P3_IR_reg[31]/NET0131  ;
  assign n15876 = n15874 & n15875 ;
  assign n15877 = n887 & n15876 ;
  assign n15878 = n720 & n15877 ;
  assign n15879 = ~n15873 & ~n15878 ;
  assign n15880 = \P1_state_reg[0]/NET0131  & n1857 ;
  assign n15881 = ~\P1_state_reg[0]/NET0131  & n1866 ;
  assign n15882 = ~n15880 & ~n15881 ;
  assign n15883 = ~\P1_state_reg[0]/NET0131  & ~n1813 ;
  assign n15884 = \P1_state_reg[0]/NET0131  & ~n1818 ;
  assign n15885 = ~n15883 & ~n15884 ;
  assign n15886 = ~\P1_state_reg[0]/NET0131  & ~n1787 ;
  assign n15887 = \P1_state_reg[0]/NET0131  & ~n1792 ;
  assign n15888 = ~n15886 & ~n15887 ;
  assign n15889 = ~\P1_state_reg[0]/NET0131  & ~n1762 ;
  assign n15890 = \P1_state_reg[0]/NET0131  & ~n1766 ;
  assign n15891 = ~n15889 & ~n15890 ;
  assign n15892 = ~\P1_state_reg[0]/NET0131  & ~n1736 ;
  assign n15893 = \P1_state_reg[0]/NET0131  & n1742 ;
  assign n15894 = ~n15892 & ~n15893 ;
  assign n15895 = ~\P1_state_reg[0]/NET0131  & ~n1695 ;
  assign n15896 = \P1_state_reg[0]/NET0131  & n1702 ;
  assign n15897 = ~n15895 & ~n15896 ;
  assign n15898 = ~\P1_state_reg[0]/NET0131  & ~n1670 ;
  assign n15899 = \P1_state_reg[0]/NET0131  & n1675 ;
  assign n15900 = ~n15898 & ~n15899 ;
  assign n15901 = \P1_state_reg[0]/NET0131  & ~n3658 ;
  assign n15902 = ~\P1_state_reg[0]/NET0131  & n3666 ;
  assign n15903 = ~n15901 & ~n15902 ;
  assign n15904 = ~\P1_state_reg[0]/NET0131  & ~n3244 ;
  assign n15905 = \P1_state_reg[0]/NET0131  & ~n3236 ;
  assign n15906 = ~n15904 & ~n15905 ;
  assign n15907 = \P1_state_reg[0]/NET0131  & ~n3631 ;
  assign n15908 = ~\P1_state_reg[0]/NET0131  & n3639 ;
  assign n15909 = ~n15907 & ~n15908 ;
  assign n15910 = \P1_state_reg[0]/NET0131  & ~n3335 ;
  assign n15911 = ~\P1_state_reg[0]/NET0131  & n3343 ;
  assign n15912 = ~n15910 & ~n15911 ;
  assign n15913 = ~\P1_state_reg[0]/NET0131  & ~n3217 ;
  assign n15914 = \P1_state_reg[0]/NET0131  & ~n3209 ;
  assign n15915 = ~n15913 & ~n15914 ;
  assign n15916 = \P1_state_reg[0]/NET0131  & ~n3184 ;
  assign n15917 = ~\P1_state_reg[0]/NET0131  & n3192 ;
  assign n15918 = ~n15916 & ~n15917 ;
  assign n15919 = \P1_state_reg[0]/NET0131  & ~n3044 ;
  assign n15920 = ~\P1_state_reg[0]/NET0131  & n3070 ;
  assign n15921 = ~n15919 & ~n15920 ;
  assign n15922 = ~\P1_state_reg[0]/NET0131  & ~n3612 ;
  assign n15923 = \P1_state_reg[0]/NET0131  & n3604 ;
  assign n15924 = ~n15922 & ~n15923 ;
  assign n15925 = \P1_state_reg[0]/NET0131  & ~n3090 ;
  assign n15926 = ~\P1_state_reg[0]/NET0131  & n3098 ;
  assign n15927 = ~n15925 & ~n15926 ;
  assign n15928 = ~\P1_state_reg[0]/NET0131  & ~n2940 ;
  assign n15929 = \P1_state_reg[0]/NET0131  & n2893 ;
  assign n15930 = ~n15928 & ~n15929 ;
  assign n15931 = \P1_state_reg[0]/NET0131  & ~n3708 ;
  assign n15932 = ~\P1_state_reg[0]/NET0131  & n3716 ;
  assign n15933 = ~n15931 & ~n15932 ;
  assign n15934 = ~\P1_state_reg[0]/NET0131  & ~n3587 ;
  assign n15935 = \P1_state_reg[0]/NET0131  & n2702 ;
  assign n15936 = ~n15934 & ~n15935 ;
  assign n15937 = ~\P1_state_reg[0]/NET0131  & ~n3293 ;
  assign n15938 = \P1_state_reg[0]/NET0131  & n2699 ;
  assign n15939 = ~n15937 & ~n15938 ;
  assign n15940 = ~\P1_state_reg[0]/NET0131  & n3272 ;
  assign n15941 = ~n6078 & ~n15940 ;
  assign n15942 = \P1_state_reg[0]/NET0131  & ~n2690 ;
  assign n15943 = ~\P1_state_reg[0]/NET0131  & n2829 ;
  assign n15944 = ~n15942 & ~n15943 ;
  assign n15945 = \P1_state_reg[0]/NET0131  & ~n6092 ;
  assign n15946 = ~\P1_state_reg[0]/NET0131  & n3538 ;
  assign n15947 = ~n15945 & ~n15946 ;
  assign n15948 = ~\P1_state_reg[0]/NET0131  & ~n3018 ;
  assign n15949 = \P1_state_reg[0]/NET0131  & n2713 ;
  assign n15950 = ~n15948 & ~n15949 ;
  assign n15951 = ~\P1_state_reg[0]/NET0131  & ~n3402 ;
  assign n15952 = \P1_state_reg[0]/NET0131  & n2850 ;
  assign n15953 = ~n15951 & ~n15952 ;
  assign n15954 = ~\P1_state_reg[0]/NET0131  & ~n3371 ;
  assign n15955 = \P1_state_reg[0]/NET0131  & ~n3376 ;
  assign n15956 = ~n15954 & ~n15955 ;
  assign n15957 = ~\P1_state_reg[0]/NET0131  & ~n3499 ;
  assign n15958 = \P1_state_reg[0]/NET0131  & n2840 ;
  assign n15959 = ~n15957 & ~n15958 ;
  assign n15960 = ~\P1_state_reg[0]/NET0131  & n3466 ;
  assign n15961 = ~\P1_IR_reg[29]/NET0131  & ~\P1_IR_reg[30]/NET0131  ;
  assign n15962 = \P1_IR_reg[31]/NET0131  & \P1_state_reg[0]/NET0131  ;
  assign n15963 = n15961 & n15962 ;
  assign n15964 = n2833 & n15963 ;
  assign n15965 = n2720 & n15964 ;
  assign n15966 = n2718 & n15965 ;
  assign n15967 = ~n15960 & ~n15966 ;
  assign n15968 = ~\P1_state_reg[0]/NET0131  & ~n3763 ;
  assign n15969 = \P1_state_reg[0]/NET0131  & ~n3768 ;
  assign n15970 = ~n15968 & ~n15969 ;
  assign n15971 = ~\P1_state_reg[0]/NET0131  & ~n3780 ;
  assign n15972 = \P1_state_reg[0]/NET0131  & ~n3784 ;
  assign n15973 = ~n15971 & ~n15972 ;
  assign n15974 = ~\P1_state_reg[0]/NET0131  & ~n3119 ;
  assign n15975 = \P1_state_reg[0]/NET0131  & n3126 ;
  assign n15976 = ~n15974 & ~n15975 ;
  assign n15977 = ~\P1_state_reg[0]/NET0131  & ~n3729 ;
  assign n15978 = \P1_state_reg[0]/NET0131  & ~n3735 ;
  assign n15979 = ~n15977 & ~n15978 ;
  assign n15980 = ~\P1_state_reg[0]/NET0131  & ~n3566 ;
  assign n15981 = \P1_state_reg[0]/NET0131  & ~n3558 ;
  assign n15982 = ~n15980 & ~n15981 ;
  assign n15983 = \P1_state_reg[0]/NET0131  & ~n3803 ;
  assign n15984 = ~\P1_state_reg[0]/NET0131  & n3811 ;
  assign n15985 = ~n15983 & ~n15984 ;
  assign n15986 = ~\P1_state_reg[0]/NET0131  & ~n3318 ;
  assign n15987 = \P1_state_reg[0]/NET0131  & ~n3310 ;
  assign n15988 = ~n15986 & ~n15987 ;
  assign n16064 = \P2_reg1_reg[16]/NET0131  & ~n4882 ;
  assign n16065 = ~\P2_reg1_reg[16]/NET0131  & n4882 ;
  assign n16066 = ~n16064 & ~n16065 ;
  assign n16067 = ~\P2_reg1_reg[15]/NET0131  & ~n4907 ;
  assign n16068 = ~\P2_reg1_reg[14]/NET0131  & ~n4833 ;
  assign n16069 = ~\P2_reg1_reg[13]/NET0131  & n4857 ;
  assign n16072 = ~\P2_reg1_reg[12]/NET0131  & ~n4963 ;
  assign n16073 = ~\P2_reg1_reg[11]/NET0131  & ~n4938 ;
  assign n16075 = ~\P2_reg1_reg[10]/NET0131  & n4995 ;
  assign n16076 = \P2_reg1_reg[9]/NET0131  & n5012 ;
  assign n16077 = ~\P2_reg1_reg[9]/NET0131  & ~n5012 ;
  assign n16078 = \P2_reg1_reg[8]/NET0131  & n5056 ;
  assign n16079 = ~\P2_reg1_reg[8]/NET0131  & ~n5056 ;
  assign n16080 = \P2_reg1_reg[7]/NET0131  & n5079 ;
  assign n16081 = ~\P2_reg1_reg[7]/NET0131  & ~n5079 ;
  assign n16082 = \P2_reg1_reg[6]/NET0131  & ~n5096 ;
  assign n16083 = ~\P2_reg1_reg[6]/NET0131  & n5096 ;
  assign n16084 = \P2_reg1_reg[5]/NET0131  & n5121 ;
  assign n16085 = ~\P2_reg1_reg[5]/NET0131  & ~n5121 ;
  assign n16086 = \P2_reg1_reg[4]/NET0131  & ~n5207 ;
  assign n16087 = ~\P2_reg1_reg[4]/NET0131  & n5207 ;
  assign n16088 = \P2_reg1_reg[3]/NET0131  & n5238 ;
  assign n16089 = ~\P2_reg1_reg[3]/NET0131  & ~n5238 ;
  assign n16090 = \P2_reg1_reg[2]/NET0131  & n5151 ;
  assign n16091 = ~\P2_reg1_reg[2]/NET0131  & ~n5151 ;
  assign n16092 = \P2_reg1_reg[1]/NET0131  & ~n5165 ;
  assign n16093 = ~\P2_reg1_reg[1]/NET0131  & n5165 ;
  assign n16094 = \P2_IR_reg[0]/NET0131  & \P2_reg1_reg[0]/NET0131  ;
  assign n16095 = ~n16093 & n16094 ;
  assign n16096 = ~n16092 & ~n16095 ;
  assign n16097 = ~n16091 & ~n16096 ;
  assign n16098 = ~n16090 & ~n16097 ;
  assign n16099 = ~n16089 & ~n16098 ;
  assign n16100 = ~n16088 & ~n16099 ;
  assign n16101 = ~n16087 & ~n16100 ;
  assign n16102 = ~n16086 & ~n16101 ;
  assign n16103 = ~n16085 & ~n16102 ;
  assign n16104 = ~n16084 & ~n16103 ;
  assign n16105 = ~n16083 & ~n16104 ;
  assign n16106 = ~n16082 & ~n16105 ;
  assign n16107 = ~n16081 & ~n16106 ;
  assign n16108 = ~n16080 & ~n16107 ;
  assign n16109 = ~n16079 & ~n16108 ;
  assign n16110 = ~n16078 & ~n16109 ;
  assign n16111 = ~n16077 & ~n16110 ;
  assign n16112 = ~n16076 & ~n16111 ;
  assign n16113 = ~n16075 & ~n16112 ;
  assign n16074 = \P2_reg1_reg[11]/NET0131  & n4938 ;
  assign n16114 = \P2_reg1_reg[10]/NET0131  & ~n4995 ;
  assign n16115 = ~n16074 & ~n16114 ;
  assign n16116 = ~n16113 & n16115 ;
  assign n16117 = ~n16073 & ~n16116 ;
  assign n16118 = ~n16072 & n16117 ;
  assign n16070 = \P2_reg1_reg[12]/NET0131  & n4963 ;
  assign n16071 = \P2_reg1_reg[13]/NET0131  & ~n4857 ;
  assign n16119 = ~n16070 & ~n16071 ;
  assign n16120 = ~n16118 & n16119 ;
  assign n16121 = ~n16069 & ~n16120 ;
  assign n16122 = ~n16068 & n16121 ;
  assign n16123 = \P2_reg1_reg[14]/NET0131  & n4833 ;
  assign n16124 = \P2_reg1_reg[15]/NET0131  & n4907 ;
  assign n16125 = ~n16123 & ~n16124 ;
  assign n16126 = ~n16122 & n16125 ;
  assign n16127 = ~n16067 & ~n16126 ;
  assign n16129 = n16066 & n16127 ;
  assign n16063 = ~n4225 & n4231 ;
  assign n16128 = ~n16066 & ~n16127 ;
  assign n16130 = n16063 & ~n16128 ;
  assign n16131 = ~n16129 & n16130 ;
  assign n15989 = ~n4225 & ~n5585 ;
  assign n15991 = n4882 & ~n15989 ;
  assign n15990 = ~\P2_addr_reg[16]/NET0131  & n15989 ;
  assign n15992 = ~n4231 & ~n15990 ;
  assign n15993 = ~n15991 & n15992 ;
  assign n15995 = \P2_reg2_reg[16]/NET0131  & ~n4882 ;
  assign n15996 = ~\P2_reg2_reg[16]/NET0131  & n4882 ;
  assign n15997 = ~n15995 & ~n15996 ;
  assign n15998 = ~\P2_reg2_reg[15]/NET0131  & ~n4907 ;
  assign n15999 = ~\P2_reg2_reg[14]/NET0131  & ~n4833 ;
  assign n16000 = ~\P2_reg2_reg[13]/NET0131  & n4857 ;
  assign n16003 = ~\P2_reg2_reg[12]/NET0131  & ~n4963 ;
  assign n16004 = ~\P2_reg2_reg[11]/NET0131  & ~n4938 ;
  assign n16006 = ~\P2_reg2_reg[10]/NET0131  & n4995 ;
  assign n16007 = ~\P2_reg2_reg[9]/NET0131  & ~n5012 ;
  assign n16009 = ~\P2_reg2_reg[8]/NET0131  & ~n5056 ;
  assign n16010 = \P2_reg2_reg[7]/NET0131  & n5079 ;
  assign n16011 = ~\P2_reg2_reg[7]/NET0131  & ~n5079 ;
  assign n16012 = \P2_reg2_reg[6]/NET0131  & ~n5096 ;
  assign n16013 = ~\P2_reg2_reg[6]/NET0131  & n5096 ;
  assign n16014 = \P2_reg2_reg[5]/NET0131  & n5121 ;
  assign n16015 = ~\P2_reg2_reg[5]/NET0131  & ~n5121 ;
  assign n16016 = \P2_reg2_reg[4]/NET0131  & ~n5207 ;
  assign n16017 = ~\P2_reg2_reg[4]/NET0131  & n5207 ;
  assign n16018 = \P2_reg2_reg[3]/NET0131  & n5238 ;
  assign n16019 = ~\P2_reg2_reg[3]/NET0131  & ~n5238 ;
  assign n16020 = \P2_reg2_reg[2]/NET0131  & n5151 ;
  assign n16021 = ~\P2_reg2_reg[2]/NET0131  & ~n5151 ;
  assign n16022 = \P2_reg2_reg[1]/NET0131  & ~n5165 ;
  assign n16023 = ~\P2_reg2_reg[1]/NET0131  & n5165 ;
  assign n16024 = \P2_IR_reg[0]/NET0131  & \P2_reg2_reg[0]/NET0131  ;
  assign n16025 = ~n16023 & n16024 ;
  assign n16026 = ~n16022 & ~n16025 ;
  assign n16027 = ~n16021 & ~n16026 ;
  assign n16028 = ~n16020 & ~n16027 ;
  assign n16029 = ~n16019 & ~n16028 ;
  assign n16030 = ~n16018 & ~n16029 ;
  assign n16031 = ~n16017 & ~n16030 ;
  assign n16032 = ~n16016 & ~n16031 ;
  assign n16033 = ~n16015 & ~n16032 ;
  assign n16034 = ~n16014 & ~n16033 ;
  assign n16035 = ~n16013 & ~n16034 ;
  assign n16036 = ~n16012 & ~n16035 ;
  assign n16037 = ~n16011 & ~n16036 ;
  assign n16038 = ~n16010 & ~n16037 ;
  assign n16039 = ~n16009 & ~n16038 ;
  assign n16008 = \P2_reg2_reg[8]/NET0131  & n5056 ;
  assign n16040 = \P2_reg2_reg[9]/NET0131  & n5012 ;
  assign n16041 = ~n16008 & ~n16040 ;
  assign n16042 = ~n16039 & n16041 ;
  assign n16043 = ~n16007 & ~n16042 ;
  assign n16044 = ~n16006 & n16043 ;
  assign n16005 = \P2_reg2_reg[11]/NET0131  & n4938 ;
  assign n16045 = \P2_reg2_reg[10]/NET0131  & ~n4995 ;
  assign n16046 = ~n16005 & ~n16045 ;
  assign n16047 = ~n16044 & n16046 ;
  assign n16048 = ~n16004 & ~n16047 ;
  assign n16049 = ~n16003 & n16048 ;
  assign n16001 = \P2_reg2_reg[12]/NET0131  & n4963 ;
  assign n16002 = \P2_reg2_reg[13]/NET0131  & ~n4857 ;
  assign n16050 = ~n16001 & ~n16002 ;
  assign n16051 = ~n16049 & n16050 ;
  assign n16052 = ~n16000 & ~n16051 ;
  assign n16053 = ~n15999 & n16052 ;
  assign n16054 = \P2_reg2_reg[14]/NET0131  & n4833 ;
  assign n16055 = \P2_reg2_reg[15]/NET0131  & n4907 ;
  assign n16056 = ~n16054 & ~n16055 ;
  assign n16057 = ~n16053 & n16056 ;
  assign n16058 = ~n15998 & ~n16057 ;
  assign n16060 = n15997 & n16058 ;
  assign n15994 = n4225 & n4231 ;
  assign n16059 = ~n15997 & ~n16058 ;
  assign n16061 = n15994 & ~n16059 ;
  assign n16062 = ~n16060 & n16061 ;
  assign n16132 = ~n15993 & ~n16062 ;
  assign n16133 = ~n16131 & n16132 ;
  assign n16134 = \P1_state_reg[0]/NET0131  & ~n16133 ;
  assign n16135 = ~n11529 & ~n16134 ;
  assign n16136 = \P1_reg3_reg[1]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n16140 = n3708 & n6095 ;
  assign n16139 = ~\P1_addr_reg[1]/NET0131  & ~n6095 ;
  assign n16141 = n2726 & ~n16139 ;
  assign n16142 = ~n16140 & n16141 ;
  assign n16152 = n2713 & n2725 ;
  assign n16153 = \P1_IR_reg[0]/NET0131  & \P1_reg2_reg[0]/NET0131  ;
  assign n16154 = ~\P1_reg2_reg[1]/NET0131  & n3708 ;
  assign n16155 = \P1_reg2_reg[1]/NET0131  & ~n3708 ;
  assign n16156 = ~n16154 & ~n16155 ;
  assign n16157 = ~n16153 & ~n16156 ;
  assign n16158 = n16153 & n16156 ;
  assign n16159 = ~n16157 & ~n16158 ;
  assign n16160 = n16152 & n16159 ;
  assign n16137 = ~n2713 & n2725 ;
  assign n16138 = ~n3708 & n16137 ;
  assign n16148 = n2713 & ~n2725 ;
  assign n16143 = \P1_IR_reg[0]/NET0131  & \P1_reg1_reg[0]/NET0131  ;
  assign n16144 = ~\P1_reg1_reg[1]/NET0131  & n3708 ;
  assign n16145 = \P1_reg1_reg[1]/NET0131  & ~n3708 ;
  assign n16146 = ~n16144 & ~n16145 ;
  assign n16147 = n16143 & n16146 ;
  assign n16149 = ~n16143 & ~n16146 ;
  assign n16150 = ~n16147 & ~n16149 ;
  assign n16151 = n16148 & n16150 ;
  assign n16161 = ~n16138 & ~n16151 ;
  assign n16162 = ~n16160 & n16161 ;
  assign n16163 = ~n16142 & n16162 ;
  assign n16164 = \P1_state_reg[0]/NET0131  & ~n16163 ;
  assign n16165 = ~n16136 & ~n16164 ;
  assign n16166 = \P1_reg3_reg[2]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n16169 = n3376 & n6095 ;
  assign n16168 = ~\P1_addr_reg[2]/NET0131  & ~n6095 ;
  assign n16170 = n2726 & ~n16168 ;
  assign n16171 = ~n16169 & n16170 ;
  assign n16181 = \P1_reg1_reg[2]/NET0131  & ~n3376 ;
  assign n16182 = ~\P1_reg1_reg[2]/NET0131  & n3376 ;
  assign n16183 = ~n16181 & ~n16182 ;
  assign n16184 = ~n16143 & ~n16145 ;
  assign n16185 = ~n16144 & ~n16184 ;
  assign n16186 = ~n16183 & ~n16185 ;
  assign n16187 = n16183 & n16185 ;
  assign n16188 = ~n16186 & ~n16187 ;
  assign n16189 = n16148 & n16188 ;
  assign n16167 = ~n3376 & n16137 ;
  assign n16172 = \P1_reg2_reg[2]/NET0131  & ~n3376 ;
  assign n16173 = ~\P1_reg2_reg[2]/NET0131  & n3376 ;
  assign n16174 = ~n16172 & ~n16173 ;
  assign n16175 = ~n16153 & ~n16155 ;
  assign n16176 = ~n16154 & ~n16175 ;
  assign n16177 = ~n16174 & ~n16176 ;
  assign n16178 = n16174 & n16176 ;
  assign n16179 = ~n16177 & ~n16178 ;
  assign n16180 = n16152 & n16179 ;
  assign n16190 = ~n16167 & ~n16180 ;
  assign n16191 = ~n16189 & n16190 ;
  assign n16192 = ~n16171 & n16191 ;
  assign n16193 = \P1_state_reg[0]/NET0131  & ~n16192 ;
  assign n16194 = ~n16166 & ~n16193 ;
  assign n16200 = ~n16008 & ~n16009 ;
  assign n16201 = n16038 & ~n16200 ;
  assign n16202 = ~n16038 & n16200 ;
  assign n16203 = ~n16201 & ~n16202 ;
  assign n16204 = n4225 & ~n16203 ;
  assign n16195 = ~n16078 & ~n16079 ;
  assign n16197 = ~n16108 & ~n16195 ;
  assign n16196 = n16108 & n16195 ;
  assign n16198 = ~n4225 & ~n16196 ;
  assign n16199 = ~n16197 & n16198 ;
  assign n16205 = n4231 & ~n16199 ;
  assign n16206 = ~n16204 & n16205 ;
  assign n16208 = ~n5056 & ~n15989 ;
  assign n16207 = ~\P2_addr_reg[8]/NET0131  & n15989 ;
  assign n16209 = ~n4231 & ~n16207 ;
  assign n16210 = ~n16208 & n16209 ;
  assign n16211 = ~n16206 & ~n16210 ;
  assign n16212 = \P1_state_reg[0]/NET0131  & ~n16211 ;
  assign n16213 = ~n13457 & ~n16212 ;
  assign n16216 = n3768 & n6095 ;
  assign n16215 = ~\P1_addr_reg[3]/NET0131  & ~n6095 ;
  assign n16217 = n2726 & ~n16215 ;
  assign n16218 = ~n16216 & n16217 ;
  assign n16228 = \P1_reg2_reg[3]/NET0131  & ~n3768 ;
  assign n16229 = ~\P1_reg2_reg[3]/NET0131  & n3768 ;
  assign n16230 = ~n16228 & ~n16229 ;
  assign n16231 = ~n16172 & ~n16176 ;
  assign n16232 = ~n16173 & ~n16231 ;
  assign n16233 = ~n16230 & ~n16232 ;
  assign n16234 = n16230 & n16232 ;
  assign n16235 = ~n16233 & ~n16234 ;
  assign n16236 = n16152 & n16235 ;
  assign n16214 = ~n3768 & n16137 ;
  assign n16219 = \P1_reg1_reg[3]/NET0131  & ~n3768 ;
  assign n16220 = ~\P1_reg1_reg[3]/NET0131  & n3768 ;
  assign n16221 = ~n16219 & ~n16220 ;
  assign n16222 = ~n16181 & ~n16185 ;
  assign n16223 = ~n16182 & ~n16222 ;
  assign n16224 = ~n16221 & ~n16223 ;
  assign n16225 = n16221 & n16223 ;
  assign n16226 = ~n16224 & ~n16225 ;
  assign n16227 = n16148 & n16226 ;
  assign n16237 = ~n16214 & ~n16227 ;
  assign n16238 = ~n16236 & n16237 ;
  assign n16239 = ~n16218 & n16238 ;
  assign n16240 = \P1_state_reg[0]/NET0131  & ~n16239 ;
  assign n16241 = ~n13493 & ~n16240 ;
  assign n16244 = ~n3784 & n6095 ;
  assign n16243 = ~\P1_addr_reg[4]/NET0131  & ~n6095 ;
  assign n16245 = n2726 & ~n16243 ;
  assign n16246 = ~n16244 & n16245 ;
  assign n16256 = \P1_reg1_reg[4]/NET0131  & n3784 ;
  assign n16257 = ~\P1_reg1_reg[4]/NET0131  & ~n3784 ;
  assign n16258 = ~n16256 & ~n16257 ;
  assign n16259 = ~n16219 & ~n16223 ;
  assign n16260 = ~n16220 & ~n16259 ;
  assign n16261 = ~n16258 & ~n16260 ;
  assign n16262 = n16258 & n16260 ;
  assign n16263 = ~n16261 & ~n16262 ;
  assign n16264 = n16148 & n16263 ;
  assign n16242 = n3784 & n16137 ;
  assign n16247 = \P1_reg2_reg[4]/NET0131  & n3784 ;
  assign n16248 = ~\P1_reg2_reg[4]/NET0131  & ~n3784 ;
  assign n16249 = ~n16247 & ~n16248 ;
  assign n16250 = ~n16228 & ~n16232 ;
  assign n16251 = ~n16229 & ~n16250 ;
  assign n16252 = ~n16249 & ~n16251 ;
  assign n16253 = n16249 & n16251 ;
  assign n16254 = ~n16252 & ~n16253 ;
  assign n16255 = n16152 & n16254 ;
  assign n16265 = ~n16242 & ~n16255 ;
  assign n16266 = ~n16264 & n16265 ;
  assign n16267 = ~n16246 & n16266 ;
  assign n16268 = \P1_state_reg[0]/NET0131  & ~n16267 ;
  assign n16269 = ~n12724 & ~n16268 ;
  assign n16272 = ~n3126 & n6095 ;
  assign n16271 = ~\P1_addr_reg[5]/NET0131  & ~n6095 ;
  assign n16273 = n2726 & ~n16271 ;
  assign n16274 = ~n16272 & n16273 ;
  assign n16284 = \P1_reg1_reg[5]/NET0131  & n3126 ;
  assign n16285 = ~\P1_reg1_reg[5]/NET0131  & ~n3126 ;
  assign n16286 = ~n16284 & ~n16285 ;
  assign n16287 = ~n16256 & ~n16260 ;
  assign n16288 = ~n16257 & ~n16287 ;
  assign n16290 = n16286 & n16288 ;
  assign n16289 = ~n16286 & ~n16288 ;
  assign n16291 = n16148 & ~n16289 ;
  assign n16292 = ~n16290 & n16291 ;
  assign n16270 = n3126 & n16137 ;
  assign n16275 = \P1_reg2_reg[5]/NET0131  & n3126 ;
  assign n16276 = ~\P1_reg2_reg[5]/NET0131  & ~n3126 ;
  assign n16277 = ~n16275 & ~n16276 ;
  assign n16278 = ~n16247 & ~n16251 ;
  assign n16279 = ~n16248 & ~n16278 ;
  assign n16281 = n16277 & n16279 ;
  assign n16280 = ~n16277 & ~n16279 ;
  assign n16282 = n16152 & ~n16280 ;
  assign n16283 = ~n16281 & n16282 ;
  assign n16293 = ~n16270 & ~n16283 ;
  assign n16294 = ~n16292 & n16293 ;
  assign n16295 = ~n16274 & n16294 ;
  assign n16296 = \P1_state_reg[0]/NET0131  & ~n16295 ;
  assign n16297 = ~n12769 & ~n16296 ;
  assign n16316 = ~n2725 & ~n6095 ;
  assign n16318 = ~n3735 & ~n16316 ;
  assign n16317 = ~\P1_addr_reg[6]/NET0131  & n16316 ;
  assign n16319 = ~n2713 & ~n16317 ;
  assign n16320 = ~n16318 & n16319 ;
  assign n16298 = \P1_reg1_reg[6]/NET0131  & n3735 ;
  assign n16299 = ~\P1_reg1_reg[6]/NET0131  & ~n3735 ;
  assign n16300 = ~n16298 & ~n16299 ;
  assign n16301 = ~n16284 & ~n16288 ;
  assign n16302 = ~n16285 & ~n16301 ;
  assign n16304 = n16300 & n16302 ;
  assign n16303 = ~n16300 & ~n16302 ;
  assign n16305 = n16148 & ~n16303 ;
  assign n16306 = ~n16304 & n16305 ;
  assign n16307 = \P1_reg2_reg[6]/NET0131  & n3735 ;
  assign n16308 = ~\P1_reg2_reg[6]/NET0131  & ~n3735 ;
  assign n16309 = ~n16307 & ~n16308 ;
  assign n16310 = ~n16275 & ~n16279 ;
  assign n16311 = ~n16276 & ~n16310 ;
  assign n16313 = n16309 & n16311 ;
  assign n16312 = ~n16309 & ~n16311 ;
  assign n16314 = n16152 & ~n16312 ;
  assign n16315 = ~n16313 & n16314 ;
  assign n16321 = ~n16306 & ~n16315 ;
  assign n16322 = ~n16320 & n16321 ;
  assign n16323 = \P1_state_reg[0]/NET0131  & ~n16322 ;
  assign n16324 = ~n13535 & ~n16323 ;
  assign n16350 = \P1_reg1_reg[10]/NET0131  & n3658 ;
  assign n16351 = ~\P1_reg1_reg[10]/NET0131  & ~n3658 ;
  assign n16352 = ~n16350 & ~n16351 ;
  assign n16353 = \P1_reg1_reg[9]/NET0131  & ~n3310 ;
  assign n16354 = ~\P1_reg1_reg[9]/NET0131  & n3310 ;
  assign n16355 = ~\P1_reg1_reg[8]/NET0131  & ~n3803 ;
  assign n16356 = \P1_reg1_reg[8]/NET0131  & n3803 ;
  assign n16357 = ~\P1_reg1_reg[7]/NET0131  & n3558 ;
  assign n16358 = \P1_reg1_reg[7]/NET0131  & ~n3558 ;
  assign n16359 = ~n16298 & ~n16302 ;
  assign n16360 = ~n16299 & ~n16359 ;
  assign n16361 = ~n16358 & ~n16360 ;
  assign n16362 = ~n16357 & ~n16361 ;
  assign n16363 = ~n16356 & ~n16362 ;
  assign n16364 = ~n16355 & ~n16363 ;
  assign n16365 = ~n16354 & n16364 ;
  assign n16366 = ~n16353 & ~n16365 ;
  assign n16368 = n16352 & ~n16366 ;
  assign n16367 = ~n16352 & n16366 ;
  assign n16369 = n16148 & ~n16367 ;
  assign n16370 = ~n16368 & n16369 ;
  assign n16326 = ~n3658 & ~n16316 ;
  assign n16325 = ~\P1_addr_reg[10]/NET0131  & n16316 ;
  assign n16327 = ~n2713 & ~n16325 ;
  assign n16328 = ~n16326 & n16327 ;
  assign n16329 = \P1_reg2_reg[10]/NET0131  & n3658 ;
  assign n16330 = ~\P1_reg2_reg[10]/NET0131  & ~n3658 ;
  assign n16331 = ~n16329 & ~n16330 ;
  assign n16332 = \P1_reg2_reg[9]/NET0131  & ~n3310 ;
  assign n16333 = ~\P1_reg2_reg[7]/NET0131  & n3558 ;
  assign n16334 = ~n16307 & ~n16311 ;
  assign n16335 = ~n16308 & ~n16334 ;
  assign n16336 = ~n16333 & n16335 ;
  assign n16337 = \P1_reg2_reg[8]/NET0131  & n3803 ;
  assign n16338 = \P1_reg2_reg[7]/NET0131  & ~n3558 ;
  assign n16339 = ~n16337 & ~n16338 ;
  assign n16340 = ~n16336 & n16339 ;
  assign n16341 = ~\P1_reg2_reg[9]/NET0131  & n3310 ;
  assign n16342 = ~\P1_reg2_reg[8]/NET0131  & ~n3803 ;
  assign n16343 = ~n16341 & ~n16342 ;
  assign n16344 = ~n16340 & n16343 ;
  assign n16345 = ~n16332 & ~n16344 ;
  assign n16347 = n16331 & ~n16345 ;
  assign n16346 = ~n16331 & n16345 ;
  assign n16348 = n16152 & ~n16346 ;
  assign n16349 = ~n16347 & n16348 ;
  assign n16371 = ~n16328 & ~n16349 ;
  assign n16372 = ~n16370 & n16371 ;
  assign n16373 = \P1_state_reg[0]/NET0131  & ~n16372 ;
  assign n16374 = ~n11653 & ~n16373 ;
  assign n16384 = ~n16333 & ~n16338 ;
  assign n16386 = n16335 & n16384 ;
  assign n16385 = ~n16335 & ~n16384 ;
  assign n16387 = n16152 & ~n16385 ;
  assign n16388 = ~n16386 & n16387 ;
  assign n16375 = ~n16357 & ~n16358 ;
  assign n16377 = n16360 & n16375 ;
  assign n16376 = ~n16360 & ~n16375 ;
  assign n16378 = n16148 & ~n16376 ;
  assign n16379 = ~n16377 & n16378 ;
  assign n16381 = n3558 & ~n16316 ;
  assign n16380 = ~\P1_addr_reg[7]/NET0131  & n16316 ;
  assign n16382 = ~n2713 & ~n16380 ;
  assign n16383 = ~n16381 & n16382 ;
  assign n16389 = ~n16379 & ~n16383 ;
  assign n16390 = ~n16388 & n16389 ;
  assign n16391 = \P1_state_reg[0]/NET0131  & ~n16390 ;
  assign n16392 = ~n13578 & ~n16391 ;
  assign n16403 = ~n16355 & ~n16356 ;
  assign n16405 = ~n16362 & ~n16403 ;
  assign n16404 = n16362 & n16403 ;
  assign n16406 = n16148 & ~n16404 ;
  assign n16407 = ~n16405 & n16406 ;
  assign n16393 = ~n16337 & ~n16342 ;
  assign n16394 = ~n16336 & ~n16338 ;
  assign n16396 = ~n16393 & n16394 ;
  assign n16395 = n16393 & ~n16394 ;
  assign n16397 = n16152 & ~n16395 ;
  assign n16398 = ~n16396 & n16397 ;
  assign n16400 = ~n3803 & ~n16316 ;
  assign n16399 = ~\P1_addr_reg[8]/NET0131  & n16316 ;
  assign n16401 = ~n2713 & ~n16399 ;
  assign n16402 = ~n16400 & n16401 ;
  assign n16408 = ~n16398 & ~n16402 ;
  assign n16409 = ~n16407 & n16408 ;
  assign n16410 = \P1_state_reg[0]/NET0131  & ~n16409 ;
  assign n16411 = ~n11532 & ~n16410 ;
  assign n16422 = ~n16353 & ~n16354 ;
  assign n16424 = ~n16364 & ~n16422 ;
  assign n16423 = n16364 & n16422 ;
  assign n16425 = n16148 & ~n16423 ;
  assign n16426 = ~n16424 & n16425 ;
  assign n16413 = n3310 & ~n16316 ;
  assign n16412 = ~\P1_addr_reg[9]/NET0131  & n16316 ;
  assign n16414 = ~n2713 & ~n16412 ;
  assign n16415 = ~n16413 & n16414 ;
  assign n16416 = ~n16332 & ~n16341 ;
  assign n16417 = ~n16340 & ~n16342 ;
  assign n16419 = n16416 & n16417 ;
  assign n16418 = ~n16416 & ~n16417 ;
  assign n16420 = n16152 & ~n16418 ;
  assign n16421 = ~n16419 & n16420 ;
  assign n16427 = ~n16415 & ~n16421 ;
  assign n16428 = ~n16426 & n16427 ;
  assign n16429 = \P1_state_reg[0]/NET0131  & ~n16428 ;
  assign n16430 = ~n11725 & ~n16429 ;
  assign n16431 = \P1_reg3_reg[17]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n16472 = ~\P1_reg1_reg[16]/NET0131  & ~n3184 ;
  assign n16473 = ~\P1_reg1_reg[15]/NET0131  & ~n3604 ;
  assign n16474 = ~\P1_reg1_reg[14]/NET0131  & n3209 ;
  assign n16475 = ~\P1_reg1_reg[13]/NET0131  & ~n3335 ;
  assign n16476 = \P1_reg1_reg[12]/NET0131  & n3631 ;
  assign n16477 = \P1_reg1_reg[11]/NET0131  & ~n3236 ;
  assign n16478 = ~n16354 & ~n16355 ;
  assign n16479 = ~n16351 & n16478 ;
  assign n16480 = ~n16363 & n16479 ;
  assign n16481 = ~n16350 & ~n16353 ;
  assign n16482 = ~n16351 & ~n16481 ;
  assign n16483 = ~n16480 & ~n16482 ;
  assign n16484 = ~n16477 & n16483 ;
  assign n16485 = ~\P1_reg1_reg[11]/NET0131  & n3236 ;
  assign n16486 = ~\P1_reg1_reg[12]/NET0131  & ~n3631 ;
  assign n16487 = ~n16485 & ~n16486 ;
  assign n16488 = ~n16484 & n16487 ;
  assign n16489 = ~n16476 & ~n16488 ;
  assign n16490 = ~n16475 & ~n16489 ;
  assign n16491 = \P1_reg1_reg[13]/NET0131  & n3335 ;
  assign n16492 = \P1_reg1_reg[14]/NET0131  & ~n3209 ;
  assign n16493 = ~n16491 & ~n16492 ;
  assign n16494 = ~n16490 & n16493 ;
  assign n16495 = ~n16474 & ~n16494 ;
  assign n16496 = ~n16473 & n16495 ;
  assign n16497 = \P1_reg1_reg[15]/NET0131  & n3604 ;
  assign n16498 = \P1_reg1_reg[16]/NET0131  & n3184 ;
  assign n16499 = ~n16497 & ~n16498 ;
  assign n16500 = ~n16496 & n16499 ;
  assign n16501 = ~n16472 & ~n16500 ;
  assign n16502 = \P1_reg1_reg[17]/NET0131  & n3044 ;
  assign n16503 = ~\P1_reg1_reg[17]/NET0131  & ~n3044 ;
  assign n16504 = ~n16502 & ~n16503 ;
  assign n16506 = n16501 & n16504 ;
  assign n16505 = ~n16501 & ~n16504 ;
  assign n16507 = n16148 & ~n16505 ;
  assign n16508 = ~n16506 & n16507 ;
  assign n16432 = \P1_reg2_reg[17]/NET0131  & n3044 ;
  assign n16435 = ~\P1_reg2_reg[15]/NET0131  & ~n3604 ;
  assign n16436 = ~\P1_reg2_reg[14]/NET0131  & n3209 ;
  assign n16437 = ~\P1_reg2_reg[13]/NET0131  & ~n3335 ;
  assign n16438 = \P1_reg2_reg[12]/NET0131  & n3631 ;
  assign n16439 = \P1_reg2_reg[11]/NET0131  & ~n3236 ;
  assign n16440 = ~n16329 & ~n16332 ;
  assign n16441 = ~n16344 & n16440 ;
  assign n16442 = ~n16330 & ~n16441 ;
  assign n16443 = ~n16439 & ~n16442 ;
  assign n16444 = ~\P1_reg2_reg[11]/NET0131  & n3236 ;
  assign n16445 = ~\P1_reg2_reg[12]/NET0131  & ~n3631 ;
  assign n16446 = ~n16444 & ~n16445 ;
  assign n16447 = ~n16443 & n16446 ;
  assign n16448 = ~n16438 & ~n16447 ;
  assign n16449 = ~n16437 & ~n16448 ;
  assign n16450 = \P1_reg2_reg[13]/NET0131  & n3335 ;
  assign n16451 = \P1_reg2_reg[14]/NET0131  & ~n3209 ;
  assign n16452 = ~n16450 & ~n16451 ;
  assign n16453 = ~n16449 & n16452 ;
  assign n16454 = ~n16436 & ~n16453 ;
  assign n16455 = ~n16435 & n16454 ;
  assign n16456 = \P1_reg2_reg[15]/NET0131  & n3604 ;
  assign n16457 = \P1_reg2_reg[16]/NET0131  & n3184 ;
  assign n16458 = ~n16456 & ~n16457 ;
  assign n16459 = ~n16455 & n16458 ;
  assign n16433 = ~\P1_reg2_reg[17]/NET0131  & ~n3044 ;
  assign n16460 = ~\P1_reg2_reg[16]/NET0131  & ~n3184 ;
  assign n16463 = ~n16433 & ~n16460 ;
  assign n16464 = ~n16459 & n16463 ;
  assign n16465 = ~n16432 & n16464 ;
  assign n16434 = ~n16432 & ~n16433 ;
  assign n16461 = ~n16459 & ~n16460 ;
  assign n16462 = ~n16434 & ~n16461 ;
  assign n16466 = n16152 & ~n16462 ;
  assign n16467 = ~n16465 & n16466 ;
  assign n16469 = ~n3044 & ~n16316 ;
  assign n16468 = ~\P1_addr_reg[17]/NET0131  & n16316 ;
  assign n16470 = ~n2713 & ~n16468 ;
  assign n16471 = ~n16469 & n16470 ;
  assign n16509 = ~n16467 & ~n16471 ;
  assign n16510 = ~n16508 & n16509 ;
  assign n16511 = \P1_state_reg[0]/NET0131  & ~n16510 ;
  assign n16512 = ~n16431 & ~n16511 ;
  assign n16516 = ~n5238 & n5585 ;
  assign n16515 = ~\P2_addr_reg[3]/NET0131  & ~n5585 ;
  assign n16517 = n4232 & ~n16515 ;
  assign n16518 = ~n16516 & n16517 ;
  assign n16524 = ~n16018 & ~n16019 ;
  assign n16525 = n16028 & ~n16524 ;
  assign n16526 = ~n16028 & n16524 ;
  assign n16527 = ~n16525 & ~n16526 ;
  assign n16528 = n15994 & n16527 ;
  assign n16513 = n4225 & ~n4231 ;
  assign n16514 = n5238 & n16513 ;
  assign n16519 = ~n16088 & ~n16089 ;
  assign n16520 = ~n16098 & n16519 ;
  assign n16521 = n16098 & ~n16519 ;
  assign n16522 = ~n16520 & ~n16521 ;
  assign n16523 = n16063 & n16522 ;
  assign n16529 = ~n16514 & ~n16523 ;
  assign n16530 = ~n16528 & n16529 ;
  assign n16531 = ~n16518 & n16530 ;
  assign n16532 = \P1_state_reg[0]/NET0131  & ~n16531 ;
  assign n16533 = ~n14208 & ~n16532 ;
  assign n16534 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[2]/NET0131  ;
  assign n16537 = ~n5151 & n5585 ;
  assign n16536 = ~\P2_addr_reg[2]/NET0131  & ~n5585 ;
  assign n16538 = n4232 & ~n16536 ;
  assign n16539 = ~n16537 & n16538 ;
  assign n16545 = ~n16090 & ~n16091 ;
  assign n16546 = n16096 & ~n16545 ;
  assign n16547 = ~n16096 & n16545 ;
  assign n16548 = ~n16546 & ~n16547 ;
  assign n16549 = n16063 & n16548 ;
  assign n16535 = n5151 & n16513 ;
  assign n16540 = ~n16020 & ~n16021 ;
  assign n16541 = ~n16026 & n16540 ;
  assign n16542 = n16026 & ~n16540 ;
  assign n16543 = ~n16541 & ~n16542 ;
  assign n16544 = n15994 & n16543 ;
  assign n16550 = ~n16535 & ~n16544 ;
  assign n16551 = ~n16549 & n16550 ;
  assign n16552 = ~n16539 & n16551 ;
  assign n16553 = \P1_state_reg[0]/NET0131  & ~n16552 ;
  assign n16554 = ~n16534 & ~n16553 ;
  assign n16555 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[0]/NET0131  ;
  assign n16558 = ~\P2_IR_reg[0]/NET0131  & n5585 ;
  assign n16557 = ~\P2_addr_reg[0]/NET0131  & ~n5585 ;
  assign n16559 = n4232 & ~n16557 ;
  assign n16560 = ~n16558 & n16559 ;
  assign n16564 = ~\P2_IR_reg[0]/NET0131  & ~\P2_reg1_reg[0]/NET0131  ;
  assign n16565 = ~n16094 & ~n16564 ;
  assign n16566 = n16063 & n16565 ;
  assign n16556 = \P2_IR_reg[0]/NET0131  & n16513 ;
  assign n16561 = ~\P2_IR_reg[0]/NET0131  & ~\P2_reg2_reg[0]/NET0131  ;
  assign n16562 = ~n16024 & ~n16561 ;
  assign n16563 = n15994 & n16562 ;
  assign n16567 = ~n16556 & ~n16563 ;
  assign n16568 = ~n16566 & n16567 ;
  assign n16569 = ~n16560 & n16568 ;
  assign n16570 = \P1_state_reg[0]/NET0131  & ~n16569 ;
  assign n16571 = ~n16555 & ~n16570 ;
  assign n16572 = \P1_reg3_reg[0]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n16575 = ~\P1_IR_reg[0]/NET0131  & n6095 ;
  assign n16574 = ~\P1_addr_reg[0]/NET0131  & ~n6095 ;
  assign n16576 = n2726 & ~n16574 ;
  assign n16577 = ~n16575 & n16576 ;
  assign n16581 = ~\P1_IR_reg[0]/NET0131  & ~\P1_reg2_reg[0]/NET0131  ;
  assign n16582 = ~n16153 & ~n16581 ;
  assign n16583 = n16152 & n16582 ;
  assign n16573 = \P1_IR_reg[0]/NET0131  & n16137 ;
  assign n16578 = ~\P1_IR_reg[0]/NET0131  & ~\P1_reg1_reg[0]/NET0131  ;
  assign n16579 = ~n16143 & ~n16578 ;
  assign n16580 = n16148 & n16579 ;
  assign n16584 = ~n16573 & ~n16580 ;
  assign n16585 = ~n16583 & n16584 ;
  assign n16586 = ~n16577 & n16585 ;
  assign n16587 = \P1_state_reg[0]/NET0131  & ~n16586 ;
  assign n16588 = ~n16572 & ~n16587 ;
  assign n16598 = ~n16010 & ~n16011 ;
  assign n16600 = ~n16036 & n16598 ;
  assign n16599 = n16036 & ~n16598 ;
  assign n16601 = n15994 & ~n16599 ;
  assign n16602 = ~n16600 & n16601 ;
  assign n16590 = ~n5079 & ~n15989 ;
  assign n16589 = ~\P2_addr_reg[7]/NET0131  & n15989 ;
  assign n16591 = ~n4231 & ~n16589 ;
  assign n16592 = ~n16590 & n16591 ;
  assign n16593 = ~n16080 & ~n16081 ;
  assign n16595 = ~n16106 & n16593 ;
  assign n16594 = n16106 & ~n16593 ;
  assign n16596 = n16063 & ~n16594 ;
  assign n16597 = ~n16595 & n16596 ;
  assign n16603 = ~n16592 & ~n16597 ;
  assign n16604 = ~n16602 & n16603 ;
  assign n16605 = \P1_state_reg[0]/NET0131  & ~n16604 ;
  assign n16606 = ~n13420 & ~n16605 ;
  assign n16623 = ~n16073 & ~n16074 ;
  assign n16624 = ~n16076 & ~n16114 ;
  assign n16625 = ~n16111 & n16624 ;
  assign n16626 = ~n16075 & ~n16625 ;
  assign n16628 = ~n16623 & ~n16626 ;
  assign n16627 = n16623 & n16626 ;
  assign n16629 = n16063 & ~n16627 ;
  assign n16630 = ~n16628 & n16629 ;
  assign n16607 = ~n16004 & ~n16005 ;
  assign n16608 = ~n16008 & ~n16010 ;
  assign n16609 = ~n16037 & n16608 ;
  assign n16610 = ~n16009 & ~n16609 ;
  assign n16611 = ~n16007 & n16610 ;
  assign n16612 = ~n16040 & ~n16045 ;
  assign n16613 = ~n16611 & n16612 ;
  assign n16614 = ~n16006 & ~n16613 ;
  assign n16616 = ~n16607 & ~n16614 ;
  assign n16615 = n16607 & n16614 ;
  assign n16617 = n15994 & ~n16615 ;
  assign n16618 = ~n16616 & n16617 ;
  assign n16620 = ~n4938 & ~n15989 ;
  assign n16619 = ~\P2_addr_reg[11]/NET0131  & n15989 ;
  assign n16621 = ~n4231 & ~n16619 ;
  assign n16622 = ~n16620 & n16621 ;
  assign n16631 = ~n16618 & ~n16622 ;
  assign n16632 = ~n16630 & n16631 ;
  assign n16633 = \P1_state_reg[0]/NET0131  & ~n16632 ;
  assign n16634 = ~n11325 & ~n16633 ;
  assign n16644 = ~n16439 & ~n16444 ;
  assign n16646 = n16442 & n16644 ;
  assign n16645 = ~n16442 & ~n16644 ;
  assign n16647 = n16152 & ~n16645 ;
  assign n16648 = ~n16646 & n16647 ;
  assign n16635 = ~n16477 & ~n16485 ;
  assign n16637 = ~n16483 & n16635 ;
  assign n16636 = n16483 & ~n16635 ;
  assign n16638 = n16148 & ~n16636 ;
  assign n16639 = ~n16637 & n16638 ;
  assign n16641 = n3236 & ~n16316 ;
  assign n16640 = ~\P1_addr_reg[11]/NET0131  & n16316 ;
  assign n16642 = ~n2713 & ~n16640 ;
  assign n16643 = ~n16641 & n16642 ;
  assign n16649 = ~n16639 & ~n16643 ;
  assign n16650 = ~n16648 & n16649 ;
  assign n16651 = \P1_state_reg[0]/NET0131  & ~n16650 ;
  assign n16652 = ~n11322 & ~n16651 ;
  assign n16662 = ~n16075 & ~n16114 ;
  assign n16664 = ~n16112 & n16662 ;
  assign n16663 = n16112 & ~n16662 ;
  assign n16665 = n16063 & ~n16663 ;
  assign n16666 = ~n16664 & n16665 ;
  assign n16654 = n4995 & ~n15989 ;
  assign n16653 = ~\P2_addr_reg[10]/NET0131  & n15989 ;
  assign n16655 = ~n4231 & ~n16653 ;
  assign n16656 = ~n16654 & n16655 ;
  assign n16657 = ~n16006 & ~n16045 ;
  assign n16659 = n16043 & n16657 ;
  assign n16658 = ~n16043 & ~n16657 ;
  assign n16660 = n15994 & ~n16658 ;
  assign n16661 = ~n16659 & n16660 ;
  assign n16667 = ~n16656 & ~n16661 ;
  assign n16668 = ~n16666 & n16667 ;
  assign n16669 = \P1_state_reg[0]/NET0131  & ~n16668 ;
  assign n16670 = ~n10325 & ~n16669 ;
  assign n16682 = ~n5121 & ~n15989 ;
  assign n16681 = ~\P2_addr_reg[5]/NET0131  & n15989 ;
  assign n16683 = ~n4231 & ~n16681 ;
  assign n16684 = ~n16682 & n16683 ;
  assign n16671 = ~n16014 & ~n16015 ;
  assign n16672 = ~n16032 & n16671 ;
  assign n16673 = n16032 & ~n16671 ;
  assign n16674 = ~n16672 & ~n16673 ;
  assign n16675 = n15994 & n16674 ;
  assign n16676 = ~n16084 & ~n16085 ;
  assign n16677 = n16102 & ~n16676 ;
  assign n16678 = ~n16102 & n16676 ;
  assign n16679 = ~n16677 & ~n16678 ;
  assign n16680 = n16063 & n16679 ;
  assign n16685 = ~n16675 & ~n16680 ;
  assign n16686 = ~n16684 & n16685 ;
  assign n16687 = \P1_state_reg[0]/NET0131  & ~n16686 ;
  assign n16688 = ~n12688 & ~n16687 ;
  assign n16698 = ~n16068 & ~n16123 ;
  assign n16700 = n16121 & n16698 ;
  assign n16699 = ~n16121 & ~n16698 ;
  assign n16701 = n16063 & ~n16699 ;
  assign n16702 = ~n16700 & n16701 ;
  assign n16690 = ~n4833 & ~n15989 ;
  assign n16689 = ~\P2_addr_reg[14]/NET0131  & n15989 ;
  assign n16691 = ~n4231 & ~n16689 ;
  assign n16692 = ~n16690 & n16691 ;
  assign n16693 = ~n15999 & ~n16054 ;
  assign n16695 = n16052 & n16693 ;
  assign n16694 = ~n16052 & ~n16693 ;
  assign n16696 = n15994 & ~n16694 ;
  assign n16697 = ~n16695 & n16696 ;
  assign n16703 = ~n16692 & ~n16697 ;
  assign n16704 = ~n16702 & n16703 ;
  assign n16705 = \P1_state_reg[0]/NET0131  & ~n16704 ;
  assign n16706 = ~n11405 & ~n16705 ;
  assign n16720 = ~n16476 & ~n16486 ;
  assign n16721 = ~n16351 & ~n16366 ;
  assign n16722 = ~n16350 & ~n16477 ;
  assign n16723 = ~n16721 & n16722 ;
  assign n16724 = ~n16485 & ~n16723 ;
  assign n16726 = n16720 & n16724 ;
  assign n16725 = ~n16720 & ~n16724 ;
  assign n16727 = n16148 & ~n16725 ;
  assign n16728 = ~n16726 & n16727 ;
  assign n16708 = ~n3631 & ~n16316 ;
  assign n16707 = ~\P1_addr_reg[12]/NET0131  & n16316 ;
  assign n16709 = ~n2713 & ~n16707 ;
  assign n16710 = ~n16708 & n16709 ;
  assign n16711 = ~n16438 & ~n16445 ;
  assign n16712 = ~n16330 & ~n16345 ;
  assign n16713 = ~n16329 & ~n16439 ;
  assign n16714 = ~n16712 & n16713 ;
  assign n16715 = ~n16444 & ~n16714 ;
  assign n16717 = n16711 & n16715 ;
  assign n16716 = ~n16711 & ~n16715 ;
  assign n16718 = n16152 & ~n16716 ;
  assign n16719 = ~n16717 & n16718 ;
  assign n16729 = ~n16710 & ~n16719 ;
  assign n16730 = ~n16728 & n16729 ;
  assign n16731 = \P1_state_reg[0]/NET0131  & ~n16730 ;
  assign n16732 = ~n9093 & ~n16731 ;
  assign n16756 = ~\P2_reg1_reg[17]/NET0131  & ~n4779 ;
  assign n16757 = \P2_reg1_reg[17]/NET0131  & n4779 ;
  assign n16758 = ~n16756 & ~n16757 ;
  assign n16759 = ~n16074 & ~n16626 ;
  assign n16760 = ~n16072 & ~n16073 ;
  assign n16761 = ~n16759 & n16760 ;
  assign n16762 = ~n16070 & ~n16761 ;
  assign n16763 = ~n16069 & ~n16762 ;
  assign n16764 = ~n16071 & ~n16123 ;
  assign n16765 = ~n16763 & n16764 ;
  assign n16766 = ~n16068 & ~n16765 ;
  assign n16767 = ~n16067 & n16766 ;
  assign n16768 = ~n16064 & ~n16124 ;
  assign n16769 = ~n16767 & n16768 ;
  assign n16770 = ~n16065 & ~n16769 ;
  assign n16772 = n16758 & n16770 ;
  assign n16771 = ~n16758 & ~n16770 ;
  assign n16773 = n16063 & ~n16771 ;
  assign n16774 = ~n16772 & n16773 ;
  assign n16733 = ~\P2_reg2_reg[17]/NET0131  & ~n4779 ;
  assign n16734 = \P2_reg2_reg[17]/NET0131  & n4779 ;
  assign n16735 = ~n16733 & ~n16734 ;
  assign n16736 = ~n16005 & ~n16614 ;
  assign n16737 = ~n16003 & ~n16004 ;
  assign n16738 = ~n16736 & n16737 ;
  assign n16739 = ~n16001 & ~n16738 ;
  assign n16740 = ~n16000 & ~n16739 ;
  assign n16741 = ~n16002 & ~n16054 ;
  assign n16742 = ~n16740 & n16741 ;
  assign n16743 = ~n15999 & ~n16742 ;
  assign n16744 = ~n15998 & n16743 ;
  assign n16745 = ~n15995 & ~n16055 ;
  assign n16746 = ~n16744 & n16745 ;
  assign n16747 = ~n15996 & ~n16746 ;
  assign n16749 = n16735 & n16747 ;
  assign n16748 = ~n16735 & ~n16747 ;
  assign n16750 = n15994 & ~n16748 ;
  assign n16751 = ~n16749 & n16750 ;
  assign n16753 = ~n4779 & ~n15989 ;
  assign n16752 = ~\P2_addr_reg[17]/NET0131  & n15989 ;
  assign n16754 = ~n4231 & ~n16752 ;
  assign n16755 = ~n16753 & n16754 ;
  assign n16775 = ~n16751 & ~n16755 ;
  assign n16776 = ~n16774 & n16775 ;
  assign n16777 = \P1_state_reg[0]/NET0131  & ~n16776 ;
  assign n16778 = ~n8466 & ~n16777 ;
  assign n16788 = ~n16437 & ~n16450 ;
  assign n16790 = ~n16448 & n16788 ;
  assign n16789 = n16448 & ~n16788 ;
  assign n16791 = n16152 & ~n16789 ;
  assign n16792 = ~n16790 & n16791 ;
  assign n16780 = ~n3335 & ~n16316 ;
  assign n16779 = ~\P1_addr_reg[13]/NET0131  & n16316 ;
  assign n16781 = ~n2713 & ~n16779 ;
  assign n16782 = ~n16780 & n16781 ;
  assign n16783 = ~n16475 & ~n16491 ;
  assign n16785 = ~n16489 & n16783 ;
  assign n16784 = n16489 & ~n16783 ;
  assign n16786 = n16148 & ~n16784 ;
  assign n16787 = ~n16785 & n16786 ;
  assign n16793 = ~n16782 & ~n16787 ;
  assign n16794 = ~n16792 & n16793 ;
  assign n16795 = \P1_state_reg[0]/NET0131  & ~n16794 ;
  assign n16796 = ~n11692 & ~n16795 ;
  assign n16797 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[1]/NET0131  ;
  assign n16800 = n5165 & n5585 ;
  assign n16799 = ~\P2_addr_reg[1]/NET0131  & ~n5585 ;
  assign n16801 = n4232 & ~n16799 ;
  assign n16802 = ~n16800 & n16801 ;
  assign n16808 = ~n16092 & ~n16093 ;
  assign n16809 = ~n16094 & ~n16808 ;
  assign n16810 = n16094 & n16808 ;
  assign n16811 = ~n16809 & ~n16810 ;
  assign n16812 = n16063 & n16811 ;
  assign n16798 = ~n5165 & n16513 ;
  assign n16803 = ~n16022 & ~n16023 ;
  assign n16804 = n16024 & n16803 ;
  assign n16805 = ~n16024 & ~n16803 ;
  assign n16806 = ~n16804 & ~n16805 ;
  assign n16807 = n15994 & n16806 ;
  assign n16813 = ~n16798 & ~n16807 ;
  assign n16814 = ~n16812 & n16813 ;
  assign n16815 = ~n16802 & n16814 ;
  assign n16816 = \P1_state_reg[0]/NET0131  & ~n16815 ;
  assign n16817 = ~n16797 & ~n16816 ;
  assign n16831 = ~n16474 & ~n16492 ;
  assign n16832 = ~n16486 & n16724 ;
  assign n16833 = ~n16476 & ~n16491 ;
  assign n16834 = ~n16832 & n16833 ;
  assign n16835 = ~n16475 & ~n16834 ;
  assign n16837 = n16831 & n16835 ;
  assign n16836 = ~n16831 & ~n16835 ;
  assign n16838 = n16148 & ~n16836 ;
  assign n16839 = ~n16837 & n16838 ;
  assign n16819 = n3209 & ~n16316 ;
  assign n16818 = ~\P1_addr_reg[14]/NET0131  & n16316 ;
  assign n16820 = ~n2713 & ~n16818 ;
  assign n16821 = ~n16819 & n16820 ;
  assign n16822 = ~n16436 & ~n16451 ;
  assign n16823 = ~n16445 & n16715 ;
  assign n16824 = ~n16438 & ~n16450 ;
  assign n16825 = ~n16823 & n16824 ;
  assign n16826 = ~n16437 & ~n16825 ;
  assign n16828 = n16822 & n16826 ;
  assign n16827 = ~n16822 & ~n16826 ;
  assign n16829 = n16152 & ~n16827 ;
  assign n16830 = ~n16828 & n16829 ;
  assign n16840 = ~n16821 & ~n16830 ;
  assign n16841 = ~n16839 & n16840 ;
  assign n16842 = \P1_state_reg[0]/NET0131  & ~n16841 ;
  assign n16843 = ~n12652 & ~n16842 ;
  assign n16853 = ~n16070 & ~n16072 ;
  assign n16855 = n16117 & n16853 ;
  assign n16854 = ~n16117 & ~n16853 ;
  assign n16856 = n16063 & ~n16854 ;
  assign n16857 = ~n16855 & n16856 ;
  assign n16845 = ~n4963 & ~n15989 ;
  assign n16844 = ~\P2_addr_reg[12]/NET0131  & n15989 ;
  assign n16846 = ~n4231 & ~n16844 ;
  assign n16847 = ~n16845 & n16846 ;
  assign n16848 = ~n16001 & ~n16003 ;
  assign n16850 = n16048 & n16848 ;
  assign n16849 = ~n16048 & ~n16848 ;
  assign n16851 = n15994 & ~n16849 ;
  assign n16852 = ~n16850 & n16851 ;
  assign n16858 = ~n16847 & ~n16852 ;
  assign n16859 = ~n16857 & n16858 ;
  assign n16860 = \P1_state_reg[0]/NET0131  & ~n16859 ;
  assign n16861 = ~n10368 & ~n16860 ;
  assign n16864 = ~n16076 & n16111 ;
  assign n16862 = ~n16076 & ~n16077 ;
  assign n16863 = n16110 & ~n16862 ;
  assign n16865 = n16063 & ~n16863 ;
  assign n16866 = ~n16864 & n16865 ;
  assign n16868 = ~n5012 & ~n15989 ;
  assign n16867 = ~\P2_addr_reg[9]/NET0131  & n15989 ;
  assign n16869 = ~n4231 & ~n16867 ;
  assign n16870 = ~n16868 & n16869 ;
  assign n16871 = ~n16007 & ~n16040 ;
  assign n16873 = n16610 & n16871 ;
  assign n16872 = ~n16610 & ~n16871 ;
  assign n16874 = n15994 & ~n16872 ;
  assign n16875 = ~n16873 & n16874 ;
  assign n16876 = ~n16870 & ~n16875 ;
  assign n16877 = ~n16866 & n16876 ;
  assign n16878 = \P1_state_reg[0]/NET0131  & ~n16877 ;
  assign n16879 = ~n10449 & ~n16878 ;
  assign n16889 = ~n16435 & ~n16456 ;
  assign n16891 = n16454 & n16889 ;
  assign n16890 = ~n16454 & ~n16889 ;
  assign n16892 = n16152 & ~n16890 ;
  assign n16893 = ~n16891 & n16892 ;
  assign n16881 = ~n3604 & ~n16316 ;
  assign n16880 = ~\P1_addr_reg[15]/NET0131  & n16316 ;
  assign n16882 = ~n2713 & ~n16880 ;
  assign n16883 = ~n16881 & n16882 ;
  assign n16884 = ~n16473 & ~n16497 ;
  assign n16886 = n16495 & n16884 ;
  assign n16885 = ~n16495 & ~n16884 ;
  assign n16887 = n16148 & ~n16885 ;
  assign n16888 = ~n16886 & n16887 ;
  assign n16894 = ~n16883 & ~n16888 ;
  assign n16895 = ~n16893 & n16894 ;
  assign n16896 = \P1_state_reg[0]/NET0131  & ~n16895 ;
  assign n16897 = ~n11366 & ~n16896 ;
  assign n16911 = ~n16472 & ~n16498 ;
  assign n16912 = ~n16474 & n16835 ;
  assign n16913 = ~n16492 & ~n16497 ;
  assign n16914 = ~n16912 & n16913 ;
  assign n16915 = ~n16473 & ~n16914 ;
  assign n16917 = n16911 & n16915 ;
  assign n16916 = ~n16911 & ~n16915 ;
  assign n16918 = n16148 & ~n16916 ;
  assign n16919 = ~n16917 & n16918 ;
  assign n16898 = ~n16457 & ~n16460 ;
  assign n16899 = ~n16436 & n16826 ;
  assign n16900 = ~n16451 & ~n16456 ;
  assign n16901 = ~n16899 & n16900 ;
  assign n16902 = ~n16435 & ~n16901 ;
  assign n16904 = n16898 & n16902 ;
  assign n16903 = ~n16898 & ~n16902 ;
  assign n16905 = n16152 & ~n16903 ;
  assign n16906 = ~n16904 & n16905 ;
  assign n16908 = ~n3184 & ~n16316 ;
  assign n16907 = ~\P1_addr_reg[16]/NET0131  & n16316 ;
  assign n16909 = ~n2713 & ~n16907 ;
  assign n16910 = ~n16908 & n16909 ;
  assign n16920 = ~n16906 & ~n16910 ;
  assign n16921 = ~n16919 & n16920 ;
  assign n16922 = \P1_state_reg[0]/NET0131  & ~n16921 ;
  assign n16923 = ~n9096 & ~n16922 ;
  assign n16933 = ~n16069 & ~n16071 ;
  assign n16935 = ~n16762 & n16933 ;
  assign n16934 = n16762 & ~n16933 ;
  assign n16936 = n16063 & ~n16934 ;
  assign n16937 = ~n16935 & n16936 ;
  assign n16925 = n4857 & ~n15989 ;
  assign n16924 = ~\P2_addr_reg[13]/NET0131  & n15989 ;
  assign n16926 = ~n4231 & ~n16924 ;
  assign n16927 = ~n16925 & n16926 ;
  assign n16928 = ~n16000 & ~n16002 ;
  assign n16930 = ~n16739 & n16928 ;
  assign n16929 = n16739 & ~n16928 ;
  assign n16931 = n15994 & ~n16929 ;
  assign n16932 = ~n16930 & n16931 ;
  assign n16938 = ~n16927 & ~n16932 ;
  assign n16939 = ~n16937 & n16938 ;
  assign n16940 = \P1_state_reg[0]/NET0131  & ~n16939 ;
  assign n16941 = ~n10412 & ~n16940 ;
  assign n16953 = n5096 & ~n15989 ;
  assign n16952 = ~\P2_addr_reg[6]/NET0131  & n15989 ;
  assign n16954 = ~n4231 & ~n16952 ;
  assign n16955 = ~n16953 & n16954 ;
  assign n16942 = ~n16082 & ~n16083 ;
  assign n16944 = ~n16104 & n16942 ;
  assign n16943 = n16104 & ~n16942 ;
  assign n16945 = n16063 & ~n16943 ;
  assign n16946 = ~n16944 & n16945 ;
  assign n16947 = ~n16012 & ~n16013 ;
  assign n16949 = ~n16034 & n16947 ;
  assign n16948 = n16034 & ~n16947 ;
  assign n16950 = n15994 & ~n16948 ;
  assign n16951 = ~n16949 & n16950 ;
  assign n16956 = ~n16946 & ~n16951 ;
  assign n16957 = ~n16955 & n16956 ;
  assign n16958 = \P1_state_reg[0]/NET0131  & ~n16957 ;
  assign n16959 = ~n13380 & ~n16958 ;
  assign n16962 = n5207 & n5585 ;
  assign n16961 = ~\P2_addr_reg[4]/NET0131  & ~n5585 ;
  assign n16963 = n4232 & ~n16961 ;
  assign n16964 = ~n16962 & n16963 ;
  assign n16970 = ~n16016 & ~n16017 ;
  assign n16971 = n16030 & ~n16970 ;
  assign n16972 = ~n16030 & n16970 ;
  assign n16973 = ~n16971 & ~n16972 ;
  assign n16974 = n15994 & n16973 ;
  assign n16960 = ~n5207 & n16513 ;
  assign n16965 = ~n16086 & ~n16087 ;
  assign n16966 = ~n16100 & n16965 ;
  assign n16967 = n16100 & ~n16965 ;
  assign n16968 = ~n16966 & ~n16967 ;
  assign n16969 = n16063 & n16968 ;
  assign n16975 = ~n16960 & ~n16969 ;
  assign n16976 = ~n16974 & n16975 ;
  assign n16977 = ~n16964 & n16976 ;
  assign n16978 = \P1_state_reg[0]/NET0131  & ~n16977 ;
  assign n16979 = ~n14530 & ~n16978 ;
  assign n16989 = ~n16067 & ~n16124 ;
  assign n16991 = n16766 & n16989 ;
  assign n16990 = ~n16766 & ~n16989 ;
  assign n16992 = n16063 & ~n16990 ;
  assign n16993 = ~n16991 & n16992 ;
  assign n16981 = ~n4907 & ~n15989 ;
  assign n16980 = ~\P2_addr_reg[15]/NET0131  & n15989 ;
  assign n16982 = ~n4231 & ~n16980 ;
  assign n16983 = ~n16981 & n16982 ;
  assign n16984 = ~n15998 & ~n16055 ;
  assign n16986 = n16743 & n16984 ;
  assign n16985 = ~n16743 & ~n16984 ;
  assign n16987 = n15994 & ~n16985 ;
  assign n16988 = ~n16986 & n16987 ;
  assign n16994 = ~n16983 & ~n16988 ;
  assign n16995 = ~n16993 & n16994 ;
  assign n16996 = \P1_state_reg[0]/NET0131  & ~n16995 ;
  assign n16997 = ~n11447 & ~n16996 ;
  assign n17014 = ~\P1_reg1_reg[18]/NET0131  & ~n3090 ;
  assign n17016 = n16501 & ~n16503 ;
  assign n17015 = \P1_reg1_reg[18]/NET0131  & n3090 ;
  assign n17017 = ~n16502 & ~n17015 ;
  assign n17018 = ~n17016 & n17017 ;
  assign n17019 = ~n17014 & ~n17018 ;
  assign n17020 = \P1_reg1_reg[19]/NET0131  & n17019 ;
  assign n17021 = ~\P1_reg1_reg[19]/NET0131  & ~n17019 ;
  assign n17022 = ~n17020 & ~n17021 ;
  assign n17024 = ~n2893 & ~n17022 ;
  assign n17023 = n2893 & n17022 ;
  assign n17025 = n16148 & ~n17023 ;
  assign n17026 = ~n17024 & n17025 ;
  assign n16998 = ~\P1_reg2_reg[18]/NET0131  & ~n3090 ;
  assign n16999 = \P1_reg2_reg[18]/NET0131  & n3090 ;
  assign n17000 = ~n16432 & ~n16999 ;
  assign n17001 = ~n16464 & n17000 ;
  assign n17002 = ~n16998 & ~n17001 ;
  assign n17003 = \P1_reg2_reg[19]/NET0131  & n17002 ;
  assign n17004 = ~\P1_reg2_reg[19]/NET0131  & ~n17002 ;
  assign n17005 = ~n17003 & ~n17004 ;
  assign n17007 = ~n2893 & ~n17005 ;
  assign n17006 = n2893 & n17005 ;
  assign n17008 = n16152 & ~n17006 ;
  assign n17009 = ~n17007 & n17008 ;
  assign n17011 = ~n2893 & ~n16316 ;
  assign n17010 = ~\P1_addr_reg[19]/NET0131  & n16316 ;
  assign n17012 = ~n2713 & ~n17010 ;
  assign n17013 = ~n17011 & n17012 ;
  assign n17027 = ~n17009 & ~n17013 ;
  assign n17028 = ~n17026 & n17027 ;
  assign n17029 = \P1_state_reg[0]/NET0131  & ~n17028 ;
  assign n17030 = ~n9228 & ~n17029 ;
  assign n17043 = ~n17014 & ~n17015 ;
  assign n17044 = ~n16498 & ~n16915 ;
  assign n17045 = ~n16472 & ~n16503 ;
  assign n17046 = ~n17044 & n17045 ;
  assign n17047 = ~n16502 & ~n17046 ;
  assign n17049 = n17043 & ~n17047 ;
  assign n17048 = ~n17043 & n17047 ;
  assign n17050 = n16148 & ~n17048 ;
  assign n17051 = ~n17049 & n17050 ;
  assign n17031 = ~n16998 & ~n16999 ;
  assign n17032 = ~n16457 & ~n16902 ;
  assign n17033 = n16463 & ~n17032 ;
  assign n17034 = ~n16432 & ~n17033 ;
  assign n17036 = n17031 & ~n17034 ;
  assign n17035 = ~n17031 & n17034 ;
  assign n17037 = n16152 & ~n17035 ;
  assign n17038 = ~n17036 & n17037 ;
  assign n17040 = ~n3090 & ~n16316 ;
  assign n17039 = ~\P1_addr_reg[18]/NET0131  & n16316 ;
  assign n17041 = ~n2713 & ~n17039 ;
  assign n17042 = ~n17040 & n17041 ;
  assign n17052 = ~n17038 & ~n17042 ;
  assign n17053 = ~n17051 & n17052 ;
  assign n17054 = \P1_state_reg[0]/NET0131  & ~n17053 ;
  assign n17055 = ~n9187 & ~n17054 ;
  assign n17071 = \P2_reg1_reg[18]/NET0131  & n4804 ;
  assign n17072 = ~\P2_reg1_reg[18]/NET0131  & ~n4804 ;
  assign n17073 = ~n17071 & ~n17072 ;
  assign n17074 = ~n16065 & n16127 ;
  assign n17075 = ~n16064 & ~n16757 ;
  assign n17076 = ~n17074 & n17075 ;
  assign n17077 = ~n16756 & ~n17076 ;
  assign n17079 = n17073 & n17077 ;
  assign n17078 = ~n17073 & ~n17077 ;
  assign n17080 = n16063 & ~n17078 ;
  assign n17081 = ~n17079 & n17080 ;
  assign n17056 = \P2_reg2_reg[18]/NET0131  & n4804 ;
  assign n17057 = ~\P2_reg2_reg[18]/NET0131  & ~n4804 ;
  assign n17058 = ~n17056 & ~n17057 ;
  assign n17059 = ~n15996 & n16058 ;
  assign n17060 = ~n15995 & ~n16734 ;
  assign n17061 = ~n17059 & n17060 ;
  assign n17062 = ~n16733 & ~n17061 ;
  assign n17064 = n17058 & n17062 ;
  assign n17063 = ~n17058 & ~n17062 ;
  assign n17065 = n15994 & ~n17063 ;
  assign n17066 = ~n17064 & n17065 ;
  assign n17068 = ~n4804 & ~n15989 ;
  assign n17067 = ~\P2_addr_reg[18]/NET0131  & n15989 ;
  assign n17069 = ~n4231 & ~n17067 ;
  assign n17070 = ~n17068 & n17069 ;
  assign n17082 = ~n17066 & ~n17070 ;
  assign n17083 = ~n17081 & n17082 ;
  assign n17084 = \P1_state_reg[0]/NET0131  & ~n17083 ;
  assign n17085 = ~n8423 & ~n17084 ;
  assign n17101 = ~n16734 & ~n16747 ;
  assign n17102 = ~n16733 & ~n17057 ;
  assign n17103 = ~n17101 & n17102 ;
  assign n17104 = ~n17056 & ~n17103 ;
  assign n17105 = \P2_reg2_reg[19]/NET0131  & ~n17104 ;
  assign n17106 = ~\P2_reg2_reg[19]/NET0131  & n17104 ;
  assign n17107 = ~n17105 & ~n17106 ;
  assign n17109 = ~n4735 & ~n17107 ;
  assign n17108 = n4735 & n17107 ;
  assign n17110 = n15994 & ~n17108 ;
  assign n17111 = ~n17109 & n17110 ;
  assign n17086 = ~n16757 & ~n16770 ;
  assign n17087 = ~n16756 & ~n17072 ;
  assign n17088 = ~n17086 & n17087 ;
  assign n17089 = ~n17071 & ~n17088 ;
  assign n17090 = \P2_reg1_reg[19]/NET0131  & n4735 ;
  assign n17091 = ~\P2_reg1_reg[19]/NET0131  & ~n4735 ;
  assign n17092 = ~n17090 & ~n17091 ;
  assign n17094 = ~n17089 & n17092 ;
  assign n17093 = n17089 & ~n17092 ;
  assign n17095 = n16063 & ~n17093 ;
  assign n17096 = ~n17094 & n17095 ;
  assign n17098 = ~n4735 & ~n15989 ;
  assign n17097 = ~\P2_addr_reg[19]/NET0131  & n15989 ;
  assign n17099 = ~n4231 & ~n17097 ;
  assign n17100 = ~n17098 & n17099 ;
  assign n17112 = ~n17096 & ~n17100 ;
  assign n17113 = ~n17111 & n17112 ;
  assign n17114 = \P1_state_reg[0]/NET0131  & ~n17113 ;
  assign n17115 = ~n8550 & ~n17114 ;
  assign n17116 = ~n4232 & ~n5585 ;
  assign n17117 = \P1_state_reg[0]/NET0131  & ~n17116 ;
  assign n17119 = ~\P3_reg2_reg[12]/NET0131  & n1574 ;
  assign n17120 = \P3_reg2_reg[12]/NET0131  & ~n1574 ;
  assign n17121 = ~n17119 & ~n17120 ;
  assign n17122 = \P3_reg2_reg[11]/NET0131  & ~n1625 ;
  assign n17123 = ~\P3_reg2_reg[11]/NET0131  & n1625 ;
  assign n17124 = \P3_reg2_reg[10]/NET0131  & ~n1649 ;
  assign n17163 = ~\P3_reg2_reg[10]/NET0131  & n1649 ;
  assign n17126 = \P3_reg2_reg[9]/NET0131  & ~n1675 ;
  assign n17125 = ~\P3_reg2_reg[9]/NET0131  & n1675 ;
  assign n17127 = \P3_reg2_reg[8]/NET0131  & ~n1702 ;
  assign n17128 = ~\P3_reg2_reg[8]/NET0131  & n1702 ;
  assign n17129 = \P3_reg2_reg[7]/NET0131  & ~n1742 ;
  assign n17130 = ~\P3_reg2_reg[7]/NET0131  & n1742 ;
  assign n17131 = \P3_reg2_reg[6]/NET0131  & n1766 ;
  assign n17132 = ~\P3_reg2_reg[6]/NET0131  & ~n1766 ;
  assign n17133 = \P3_reg2_reg[5]/NET0131  & n1792 ;
  assign n17134 = ~\P3_reg2_reg[5]/NET0131  & ~n1792 ;
  assign n17135 = \P3_reg2_reg[4]/NET0131  & n1818 ;
  assign n17136 = ~\P3_reg2_reg[4]/NET0131  & ~n1818 ;
  assign n17137 = \P3_reg2_reg[3]/NET0131  & ~n1857 ;
  assign n17138 = ~\P3_reg2_reg[3]/NET0131  & n1857 ;
  assign n17139 = \P3_reg2_reg[2]/NET0131  & ~n1842 ;
  assign n17140 = ~\P3_reg2_reg[2]/NET0131  & n1842 ;
  assign n17142 = \P3_reg2_reg[1]/NET0131  & n1881 ;
  assign n17141 = ~\P3_reg2_reg[1]/NET0131  & ~n1881 ;
  assign n17257 = \P3_IR_reg[0]/NET0131  & ~\P3_reg2_reg[0]/NET0131  ;
  assign n17258 = ~n17141 & ~n17257 ;
  assign n17259 = ~n17142 & ~n17258 ;
  assign n17260 = ~n17140 & ~n17259 ;
  assign n17261 = ~n17139 & ~n17260 ;
  assign n17262 = ~n17138 & ~n17261 ;
  assign n17263 = ~n17137 & ~n17262 ;
  assign n17264 = ~n17136 & ~n17263 ;
  assign n17265 = ~n17135 & ~n17264 ;
  assign n17266 = ~n17134 & ~n17265 ;
  assign n17267 = ~n17133 & ~n17266 ;
  assign n17268 = ~n17132 & ~n17267 ;
  assign n17269 = ~n17131 & ~n17268 ;
  assign n17270 = ~n17130 & ~n17269 ;
  assign n17271 = ~n17129 & ~n17270 ;
  assign n17272 = ~n17128 & ~n17271 ;
  assign n17273 = ~n17127 & ~n17272 ;
  assign n17274 = ~n17125 & ~n17273 ;
  assign n17275 = ~n17126 & ~n17274 ;
  assign n17276 = ~n17163 & ~n17275 ;
  assign n17277 = ~n17124 & ~n17276 ;
  assign n17278 = ~n17123 & ~n17277 ;
  assign n17279 = ~n17122 & ~n17278 ;
  assign n17281 = ~n17121 & n17279 ;
  assign n17223 = n724 & ~n733 ;
  assign n17280 = n17121 & ~n17279 ;
  assign n17282 = n17223 & ~n17280 ;
  assign n17283 = ~n17281 & n17282 ;
  assign n17171 = ~\P3_reg1_reg[12]/NET0131  & n1574 ;
  assign n17172 = \P3_reg1_reg[12]/NET0131  & ~n1574 ;
  assign n17173 = ~n17171 & ~n17172 ;
  assign n17174 = \P3_reg1_reg[11]/NET0131  & ~n1625 ;
  assign n17214 = ~\P3_reg1_reg[11]/NET0131  & n1625 ;
  assign n17175 = \P3_reg1_reg[10]/NET0131  & ~n1649 ;
  assign n17215 = ~\P3_reg1_reg[10]/NET0131  & n1649 ;
  assign n17176 = \P3_reg1_reg[9]/NET0131  & ~n1675 ;
  assign n17208 = ~\P3_reg1_reg[9]/NET0131  & n1675 ;
  assign n17177 = \P3_reg1_reg[8]/NET0131  & ~n1702 ;
  assign n17209 = ~\P3_reg1_reg[8]/NET0131  & n1702 ;
  assign n17179 = \P3_reg1_reg[7]/NET0131  & ~n1742 ;
  assign n17178 = ~\P3_reg1_reg[7]/NET0131  & n1742 ;
  assign n17180 = \P3_reg1_reg[6]/NET0131  & n1766 ;
  assign n17181 = ~\P3_reg1_reg[6]/NET0131  & ~n1766 ;
  assign n17182 = \P3_reg1_reg[5]/NET0131  & n1792 ;
  assign n17183 = ~\P3_reg1_reg[5]/NET0131  & ~n1792 ;
  assign n17184 = \P3_reg1_reg[4]/NET0131  & n1818 ;
  assign n17185 = ~\P3_reg1_reg[4]/NET0131  & ~n1818 ;
  assign n17186 = \P3_reg1_reg[3]/NET0131  & ~n1857 ;
  assign n17187 = ~\P3_reg1_reg[3]/NET0131  & n1857 ;
  assign n17188 = \P3_reg1_reg[2]/NET0131  & ~n1842 ;
  assign n17189 = ~\P3_reg1_reg[2]/NET0131  & n1842 ;
  assign n17191 = \P3_reg1_reg[1]/NET0131  & n1881 ;
  assign n17190 = ~\P3_reg1_reg[1]/NET0131  & ~n1881 ;
  assign n17230 = \P3_IR_reg[0]/NET0131  & ~\P3_reg1_reg[0]/NET0131  ;
  assign n17231 = ~n17190 & ~n17230 ;
  assign n17232 = ~n17191 & ~n17231 ;
  assign n17233 = ~n17189 & ~n17232 ;
  assign n17234 = ~n17188 & ~n17233 ;
  assign n17235 = ~n17187 & ~n17234 ;
  assign n17236 = ~n17186 & ~n17235 ;
  assign n17237 = ~n17185 & ~n17236 ;
  assign n17238 = ~n17184 & ~n17237 ;
  assign n17239 = ~n17183 & ~n17238 ;
  assign n17240 = ~n17182 & ~n17239 ;
  assign n17241 = ~n17181 & ~n17240 ;
  assign n17242 = ~n17180 & ~n17241 ;
  assign n17243 = ~n17178 & ~n17242 ;
  assign n17244 = ~n17179 & ~n17243 ;
  assign n17245 = ~n17209 & ~n17244 ;
  assign n17246 = ~n17177 & ~n17245 ;
  assign n17247 = ~n17208 & ~n17246 ;
  assign n17248 = ~n17176 & ~n17247 ;
  assign n17249 = ~n17215 & ~n17248 ;
  assign n17250 = ~n17175 & ~n17249 ;
  assign n17251 = ~n17214 & ~n17250 ;
  assign n17252 = ~n17174 & ~n17251 ;
  assign n17254 = n17173 & ~n17252 ;
  assign n17253 = ~n17173 & n17252 ;
  assign n17255 = n767 & ~n17253 ;
  assign n17256 = ~n17254 & n17255 ;
  assign n17229 = n733 & n1574 ;
  assign n17284 = n2145 & ~n17229 ;
  assign n17285 = ~n17256 & n17284 ;
  assign n17286 = ~n17283 & n17285 ;
  assign n17143 = ~\P3_IR_reg[0]/NET0131  & \P3_reg2_reg[0]/NET0131  ;
  assign n17144 = ~n17142 & ~n17143 ;
  assign n17145 = ~n17141 & ~n17144 ;
  assign n17146 = ~n17140 & n17145 ;
  assign n17147 = ~n17139 & ~n17146 ;
  assign n17148 = ~n17138 & ~n17147 ;
  assign n17149 = ~n17137 & ~n17148 ;
  assign n17150 = ~n17136 & ~n17149 ;
  assign n17151 = ~n17135 & ~n17150 ;
  assign n17152 = ~n17134 & ~n17151 ;
  assign n17153 = ~n17133 & ~n17152 ;
  assign n17154 = ~n17132 & ~n17153 ;
  assign n17155 = ~n17131 & ~n17154 ;
  assign n17156 = ~n17130 & ~n17155 ;
  assign n17157 = ~n17129 & ~n17156 ;
  assign n17158 = ~n17128 & ~n17157 ;
  assign n17159 = ~n17127 & ~n17158 ;
  assign n17160 = ~n17126 & n17159 ;
  assign n17161 = ~n17125 & ~n17160 ;
  assign n17162 = ~n17124 & ~n17161 ;
  assign n17164 = ~n17123 & ~n17163 ;
  assign n17165 = ~n17162 & n17164 ;
  assign n17166 = ~n17122 & ~n17165 ;
  assign n17168 = n17121 & n17166 ;
  assign n17167 = ~n17121 & ~n17166 ;
  assign n17169 = n2238 & ~n17167 ;
  assign n17170 = ~n17168 & n17169 ;
  assign n17192 = ~\P3_IR_reg[0]/NET0131  & \P3_reg1_reg[0]/NET0131  ;
  assign n17193 = ~n17191 & ~n17192 ;
  assign n17194 = ~n17190 & ~n17193 ;
  assign n17195 = ~n17189 & n17194 ;
  assign n17196 = ~n17188 & ~n17195 ;
  assign n17197 = ~n17187 & ~n17196 ;
  assign n17198 = ~n17186 & ~n17197 ;
  assign n17199 = ~n17185 & ~n17198 ;
  assign n17200 = ~n17184 & ~n17199 ;
  assign n17201 = ~n17183 & ~n17200 ;
  assign n17202 = ~n17182 & ~n17201 ;
  assign n17203 = ~n17181 & ~n17202 ;
  assign n17204 = ~n17180 & ~n17203 ;
  assign n17205 = ~n17179 & n17204 ;
  assign n17206 = ~n17178 & ~n17205 ;
  assign n17207 = ~n17177 & ~n17206 ;
  assign n17210 = ~n17208 & ~n17209 ;
  assign n17211 = ~n17207 & n17210 ;
  assign n17212 = ~n17176 & ~n17211 ;
  assign n17213 = ~n17175 & n17212 ;
  assign n17216 = ~n17214 & ~n17215 ;
  assign n17217 = ~n17213 & n17216 ;
  assign n17218 = ~n17174 & ~n17217 ;
  assign n17220 = n17173 & n17218 ;
  assign n17219 = ~n17173 & ~n17218 ;
  assign n17221 = n734 & ~n17219 ;
  assign n17222 = ~n17220 & n17221 ;
  assign n17224 = n1574 & n17223 ;
  assign n17118 = \P3_addr_reg[12]/NET0131  & n767 ;
  assign n17225 = ~n2145 & ~n17118 ;
  assign n17226 = ~n17224 & n17225 ;
  assign n17227 = ~n17222 & n17226 ;
  assign n17228 = ~n17170 & n17227 ;
  assign n17287 = \P1_state_reg[0]/NET0131  & ~n17228 ;
  assign n17288 = ~n17286 & n17287 ;
  assign n17289 = ~n10568 & ~n17288 ;
  assign n17290 = ~\P1_state_reg[0]/NET0131  & ~\P3_reg3_reg[0]/NET0131  ;
  assign n17291 = \P3_addr_reg[0]/NET0131  & n767 ;
  assign n17297 = ~n2145 & ~n17291 ;
  assign n17295 = ~n17192 & ~n17230 ;
  assign n17296 = n734 & ~n17295 ;
  assign n17292 = \P3_IR_reg[0]/NET0131  & n17223 ;
  assign n17293 = ~n17143 & ~n17257 ;
  assign n17294 = n2238 & ~n17293 ;
  assign n17298 = ~n17292 & ~n17294 ;
  assign n17299 = ~n17296 & n17298 ;
  assign n17300 = n17297 & n17299 ;
  assign n17303 = n767 & ~n17295 ;
  assign n17301 = n17223 & ~n17293 ;
  assign n17302 = \P3_IR_reg[0]/NET0131  & n733 ;
  assign n17304 = n2145 & ~n17302 ;
  assign n17305 = ~n17301 & n17304 ;
  assign n17306 = ~n17303 & n17305 ;
  assign n17307 = ~n17300 & ~n17306 ;
  assign n17308 = \P1_state_reg[0]/NET0131  & ~n17307 ;
  assign n17309 = ~n17290 & ~n17308 ;
  assign n17316 = ~n17124 & ~n17163 ;
  assign n17318 = n17275 & ~n17316 ;
  assign n17317 = ~n17275 & n17316 ;
  assign n17319 = n17223 & ~n17317 ;
  assign n17320 = ~n17318 & n17319 ;
  assign n17311 = ~n17175 & ~n17215 ;
  assign n17313 = ~n17248 & n17311 ;
  assign n17312 = n17248 & ~n17311 ;
  assign n17314 = n767 & ~n17312 ;
  assign n17315 = ~n17313 & n17314 ;
  assign n17310 = n733 & n1649 ;
  assign n17321 = n2145 & ~n17310 ;
  assign n17322 = ~n17315 & n17321 ;
  assign n17323 = ~n17320 & n17322 ;
  assign n17330 = n17161 & ~n17316 ;
  assign n17329 = ~n17161 & n17316 ;
  assign n17331 = n2238 & ~n17329 ;
  assign n17332 = ~n17330 & n17331 ;
  assign n17326 = n17212 & n17311 ;
  assign n17325 = ~n17212 & ~n17311 ;
  assign n17327 = n734 & ~n17325 ;
  assign n17328 = ~n17326 & n17327 ;
  assign n17333 = n1649 & n17223 ;
  assign n17324 = \P3_addr_reg[10]/NET0131  & n767 ;
  assign n17334 = ~n2145 & ~n17324 ;
  assign n17335 = ~n17333 & n17334 ;
  assign n17336 = ~n17328 & n17335 ;
  assign n17337 = ~n17332 & n17336 ;
  assign n17338 = \P1_state_reg[0]/NET0131  & ~n17337 ;
  assign n17339 = ~n17323 & n17338 ;
  assign n17340 = ~n10487 & ~n17339 ;
  assign n17350 = ~n17174 & ~n17214 ;
  assign n17373 = n17250 & ~n17350 ;
  assign n17372 = ~n17250 & n17350 ;
  assign n17374 = n767 & ~n17372 ;
  assign n17375 = ~n17373 & n17374 ;
  assign n17342 = ~n17122 & ~n17123 ;
  assign n17369 = ~n17277 & n17342 ;
  assign n17368 = n17277 & ~n17342 ;
  assign n17370 = n17223 & ~n17368 ;
  assign n17371 = ~n17369 & n17370 ;
  assign n17367 = n733 & n1625 ;
  assign n17376 = n2145 & ~n17367 ;
  assign n17377 = ~n17371 & n17376 ;
  assign n17378 = ~n17375 & n17377 ;
  assign n17343 = ~n17125 & ~n17163 ;
  assign n17344 = ~n17160 & n17343 ;
  assign n17345 = ~n17124 & ~n17344 ;
  assign n17347 = n17342 & n17345 ;
  assign n17346 = ~n17342 & ~n17345 ;
  assign n17348 = n2238 & ~n17346 ;
  assign n17349 = ~n17347 & n17348 ;
  assign n17351 = ~n17178 & ~n17209 ;
  assign n17352 = ~n17205 & n17351 ;
  assign n17353 = ~n17177 & ~n17352 ;
  assign n17354 = ~n17176 & n17353 ;
  assign n17355 = ~n17208 & ~n17215 ;
  assign n17356 = ~n17354 & n17355 ;
  assign n17357 = ~n17175 & ~n17356 ;
  assign n17359 = n17350 & n17357 ;
  assign n17358 = ~n17350 & ~n17357 ;
  assign n17360 = n734 & ~n17358 ;
  assign n17361 = ~n17359 & n17360 ;
  assign n17362 = n1625 & n17223 ;
  assign n17341 = \P3_addr_reg[11]/NET0131  & n767 ;
  assign n17363 = ~n2145 & ~n17341 ;
  assign n17364 = ~n17362 & n17363 ;
  assign n17365 = ~n17361 & n17364 ;
  assign n17366 = ~n17349 & n17365 ;
  assign n17379 = \P1_state_reg[0]/NET0131  & ~n17366 ;
  assign n17380 = ~n17378 & n17379 ;
  assign n17381 = ~n10528 & ~n17380 ;
  assign n17394 = ~\P3_reg1_reg[13]/NET0131  & n1558 ;
  assign n17395 = \P3_reg1_reg[13]/NET0131  & ~n1558 ;
  assign n17396 = ~n17394 & ~n17395 ;
  assign n17418 = ~n17172 & ~n17174 ;
  assign n17419 = ~n17251 & n17418 ;
  assign n17420 = ~n17171 & ~n17419 ;
  assign n17422 = ~n17396 & ~n17420 ;
  assign n17421 = n17396 & n17420 ;
  assign n17423 = n767 & ~n17421 ;
  assign n17424 = ~n17422 & n17423 ;
  assign n17383 = ~\P3_reg2_reg[13]/NET0131  & n1558 ;
  assign n17384 = \P3_reg2_reg[13]/NET0131  & ~n1558 ;
  assign n17385 = ~n17383 & ~n17384 ;
  assign n17411 = ~n17120 & ~n17122 ;
  assign n17412 = ~n17278 & n17411 ;
  assign n17413 = ~n17119 & ~n17412 ;
  assign n17415 = n17385 & n17413 ;
  assign n17414 = ~n17385 & ~n17413 ;
  assign n17416 = n17223 & ~n17414 ;
  assign n17417 = ~n17415 & n17416 ;
  assign n17410 = n733 & n1558 ;
  assign n17425 = n2145 & ~n17410 ;
  assign n17426 = ~n17417 & n17425 ;
  assign n17427 = ~n17424 & n17426 ;
  assign n17386 = ~n17122 & n17345 ;
  assign n17387 = ~n17119 & ~n17123 ;
  assign n17388 = ~n17386 & n17387 ;
  assign n17389 = ~n17120 & ~n17388 ;
  assign n17391 = n17385 & n17389 ;
  assign n17390 = ~n17385 & ~n17389 ;
  assign n17392 = n2238 & ~n17390 ;
  assign n17393 = ~n17391 & n17392 ;
  assign n17397 = ~n17174 & n17357 ;
  assign n17398 = ~n17171 & ~n17214 ;
  assign n17399 = ~n17397 & n17398 ;
  assign n17400 = ~n17172 & ~n17399 ;
  assign n17402 = n17396 & n17400 ;
  assign n17401 = ~n17396 & ~n17400 ;
  assign n17403 = n734 & ~n17401 ;
  assign n17404 = ~n17402 & n17403 ;
  assign n17405 = n1558 & n17223 ;
  assign n17382 = \P3_addr_reg[13]/NET0131  & n767 ;
  assign n17406 = ~n2145 & ~n17382 ;
  assign n17407 = ~n17405 & n17406 ;
  assign n17408 = ~n17404 & n17407 ;
  assign n17409 = ~n17393 & n17408 ;
  assign n17428 = \P1_state_reg[0]/NET0131  & ~n17409 ;
  assign n17429 = ~n17427 & n17428 ;
  assign n17430 = ~n10608 & ~n17429 ;
  assign n17446 = ~\P3_reg2_reg[15]/NET0131  & ~n1502 ;
  assign n17447 = \P3_reg2_reg[15]/NET0131  & n1502 ;
  assign n17448 = ~n17446 & ~n17447 ;
  assign n17449 = ~\P3_reg2_reg[14]/NET0131  & n1542 ;
  assign n17450 = ~n17383 & ~n17449 ;
  assign n17451 = n17413 & n17450 ;
  assign n17452 = \P3_reg2_reg[14]/NET0131  & ~n1542 ;
  assign n17453 = n17384 & ~n17449 ;
  assign n17454 = ~n17452 & ~n17453 ;
  assign n17455 = ~n17451 & n17454 ;
  assign n17457 = ~n17448 & n17455 ;
  assign n17456 = n17448 & ~n17455 ;
  assign n17458 = n17223 & ~n17456 ;
  assign n17459 = ~n17457 & n17458 ;
  assign n17432 = ~\P3_reg1_reg[15]/NET0131  & ~n1502 ;
  assign n17433 = \P3_reg1_reg[15]/NET0131  & n1502 ;
  assign n17434 = ~n17432 & ~n17433 ;
  assign n17435 = ~\P3_reg1_reg[14]/NET0131  & n1542 ;
  assign n17436 = ~n17394 & ~n17435 ;
  assign n17437 = n17420 & n17436 ;
  assign n17438 = \P3_reg1_reg[14]/NET0131  & ~n1542 ;
  assign n17439 = n17395 & ~n17435 ;
  assign n17440 = ~n17438 & ~n17439 ;
  assign n17441 = ~n17437 & n17440 ;
  assign n17443 = n17434 & ~n17441 ;
  assign n17442 = ~n17434 & n17441 ;
  assign n17444 = n767 & ~n17442 ;
  assign n17445 = ~n17443 & n17444 ;
  assign n17431 = n733 & ~n1502 ;
  assign n17460 = n2145 & ~n17431 ;
  assign n17461 = ~n17445 & n17460 ;
  assign n17462 = ~n17459 & n17461 ;
  assign n17471 = ~n17384 & n17389 ;
  assign n17472 = n17450 & ~n17471 ;
  assign n17473 = ~n17452 & ~n17472 ;
  assign n17475 = n17448 & n17473 ;
  assign n17474 = ~n17448 & ~n17473 ;
  assign n17476 = n2238 & ~n17474 ;
  assign n17477 = ~n17475 & n17476 ;
  assign n17464 = ~n17395 & n17400 ;
  assign n17465 = n17436 & ~n17464 ;
  assign n17466 = ~n17438 & ~n17465 ;
  assign n17468 = n17434 & n17466 ;
  assign n17467 = ~n17434 & ~n17466 ;
  assign n17469 = n734 & ~n17467 ;
  assign n17470 = ~n17468 & n17469 ;
  assign n17478 = ~n1502 & n17223 ;
  assign n17463 = \P3_addr_reg[15]/NET0131  & n767 ;
  assign n17479 = ~n2145 & ~n17463 ;
  assign n17480 = ~n17478 & n17479 ;
  assign n17481 = ~n17470 & n17480 ;
  assign n17482 = ~n17477 & n17481 ;
  assign n17483 = \P1_state_reg[0]/NET0131  & ~n17482 ;
  assign n17484 = ~n17462 & n17483 ;
  assign n17485 = ~n11574 & ~n17484 ;
  assign n17504 = ~\P3_reg2_reg[16]/NET0131  & n1183 ;
  assign n17505 = \P3_reg2_reg[16]/NET0131  & ~n1183 ;
  assign n17506 = ~n17504 & ~n17505 ;
  assign n17507 = ~n17447 & ~n17452 ;
  assign n17508 = ~n17119 & ~n17279 ;
  assign n17509 = ~n17120 & ~n17384 ;
  assign n17510 = ~n17508 & n17509 ;
  assign n17511 = ~n17383 & ~n17510 ;
  assign n17512 = ~n17449 & n17511 ;
  assign n17513 = n17507 & ~n17512 ;
  assign n17514 = ~n17446 & ~n17513 ;
  assign n17516 = ~n17506 & ~n17514 ;
  assign n17515 = n17506 & n17514 ;
  assign n17517 = n17223 & ~n17515 ;
  assign n17518 = ~n17516 & n17517 ;
  assign n17487 = ~\P3_reg1_reg[16]/NET0131  & n1183 ;
  assign n17488 = \P3_reg1_reg[16]/NET0131  & ~n1183 ;
  assign n17489 = ~n17487 & ~n17488 ;
  assign n17490 = ~n17433 & ~n17438 ;
  assign n17491 = ~n17432 & ~n17490 ;
  assign n17492 = ~n17432 & ~n17435 ;
  assign n17494 = ~n17171 & ~n17394 ;
  assign n17495 = ~n17252 & n17494 ;
  assign n17493 = n17172 & ~n17394 ;
  assign n17496 = ~n17395 & ~n17493 ;
  assign n17497 = ~n17495 & n17496 ;
  assign n17498 = n17492 & ~n17497 ;
  assign n17499 = ~n17491 & ~n17498 ;
  assign n17501 = n17489 & ~n17499 ;
  assign n17500 = ~n17489 & n17499 ;
  assign n17502 = n767 & ~n17500 ;
  assign n17503 = ~n17501 & n17502 ;
  assign n17486 = n733 & n1183 ;
  assign n17519 = n2145 & ~n17486 ;
  assign n17520 = ~n17503 & n17519 ;
  assign n17521 = ~n17518 & n17520 ;
  assign n17533 = ~n17120 & n17166 ;
  assign n17534 = ~n17119 & ~n17383 ;
  assign n17535 = ~n17533 & n17534 ;
  assign n17536 = ~n17384 & ~n17535 ;
  assign n17537 = n17507 & n17536 ;
  assign n17538 = ~n17447 & n17449 ;
  assign n17539 = ~n17446 & ~n17538 ;
  assign n17540 = ~n17537 & n17539 ;
  assign n17542 = n17506 & ~n17540 ;
  assign n17541 = ~n17506 & n17540 ;
  assign n17543 = n2238 & ~n17541 ;
  assign n17544 = ~n17542 & n17543 ;
  assign n17523 = ~n17172 & n17218 ;
  assign n17524 = n17494 & ~n17523 ;
  assign n17525 = ~n17395 & ~n17524 ;
  assign n17526 = ~n17438 & n17525 ;
  assign n17527 = n17492 & ~n17526 ;
  assign n17528 = ~n17433 & ~n17527 ;
  assign n17530 = n17489 & n17528 ;
  assign n17529 = ~n17489 & ~n17528 ;
  assign n17531 = n734 & ~n17529 ;
  assign n17532 = ~n17530 & n17531 ;
  assign n17545 = \P3_addr_reg[16]/NET0131  & n767 ;
  assign n17522 = n1183 & n17223 ;
  assign n17546 = ~n2145 & ~n17522 ;
  assign n17547 = ~n17545 & n17546 ;
  assign n17548 = ~n17532 & n17547 ;
  assign n17549 = ~n17544 & n17548 ;
  assign n17550 = \P1_state_reg[0]/NET0131  & ~n17549 ;
  assign n17551 = ~n17521 & n17550 ;
  assign n17552 = ~n9142 & ~n17551 ;
  assign n17567 = ~\P3_reg2_reg[18]/NET0131  & n1135 ;
  assign n17568 = \P3_reg2_reg[18]/NET0131  & ~n1135 ;
  assign n17569 = ~n17567 & ~n17568 ;
  assign n17570 = ~\P3_reg2_reg[17]/NET0131  & ~n1164 ;
  assign n17572 = ~n17504 & n17514 ;
  assign n17571 = \P3_reg2_reg[17]/NET0131  & n1164 ;
  assign n17573 = ~n17505 & ~n17571 ;
  assign n17574 = ~n17572 & n17573 ;
  assign n17575 = ~n17570 & ~n17574 ;
  assign n17577 = n17569 & n17575 ;
  assign n17576 = ~n17569 & ~n17575 ;
  assign n17578 = n17223 & ~n17576 ;
  assign n17579 = ~n17577 & n17578 ;
  assign n17554 = ~\P3_reg1_reg[18]/NET0131  & n1135 ;
  assign n17555 = \P3_reg1_reg[18]/NET0131  & ~n1135 ;
  assign n17556 = ~n17554 & ~n17555 ;
  assign n17557 = ~\P3_reg1_reg[17]/NET0131  & ~n1164 ;
  assign n17558 = ~n17487 & ~n17499 ;
  assign n17559 = \P3_reg1_reg[17]/NET0131  & n1164 ;
  assign n17560 = ~n17488 & ~n17559 ;
  assign n17561 = ~n17558 & n17560 ;
  assign n17562 = ~n17557 & ~n17561 ;
  assign n17564 = ~n17556 & ~n17562 ;
  assign n17563 = n17556 & n17562 ;
  assign n17565 = n767 & ~n17563 ;
  assign n17566 = ~n17564 & n17565 ;
  assign n17553 = n733 & n1135 ;
  assign n17580 = n2145 & ~n17553 ;
  assign n17581 = ~n17566 & n17580 ;
  assign n17582 = ~n17579 & n17581 ;
  assign n17593 = ~n17505 & ~n17540 ;
  assign n17594 = ~n17504 & ~n17570 ;
  assign n17595 = ~n17593 & n17594 ;
  assign n17596 = ~n17571 & ~n17595 ;
  assign n17598 = ~n17569 & ~n17596 ;
  assign n17597 = n17569 & n17596 ;
  assign n17599 = n2238 & ~n17597 ;
  assign n17600 = ~n17598 & n17599 ;
  assign n17583 = ~n17488 & n17528 ;
  assign n17584 = ~n17487 & ~n17557 ;
  assign n17585 = ~n17583 & n17584 ;
  assign n17586 = ~n17559 & ~n17585 ;
  assign n17588 = ~n17556 & ~n17586 ;
  assign n17587 = n17556 & n17586 ;
  assign n17589 = n734 & ~n17587 ;
  assign n17590 = ~n17588 & n17589 ;
  assign n17592 = \P3_addr_reg[18]/NET0131  & n767 ;
  assign n17591 = n1135 & n17223 ;
  assign n17601 = ~n2145 & ~n17591 ;
  assign n17602 = ~n17592 & n17601 ;
  assign n17603 = ~n17590 & n17602 ;
  assign n17604 = ~n17600 & n17603 ;
  assign n17605 = \P1_state_reg[0]/NET0131  & ~n17604 ;
  assign n17606 = ~n17582 & n17605 ;
  assign n17607 = ~n8553 & ~n17606 ;
  assign n17614 = ~n17133 & ~n17134 ;
  assign n17629 = n17151 & n17614 ;
  assign n17628 = ~n17151 & ~n17614 ;
  assign n17630 = n2238 & ~n17628 ;
  assign n17631 = ~n17629 & n17630 ;
  assign n17609 = ~n17182 & ~n17183 ;
  assign n17623 = n17200 & n17609 ;
  assign n17622 = ~n17200 & ~n17609 ;
  assign n17624 = n734 & ~n17622 ;
  assign n17625 = ~n17623 & n17624 ;
  assign n17627 = \P3_addr_reg[5]/NET0131  & n767 ;
  assign n17626 = ~n1792 & n17223 ;
  assign n17632 = ~n2145 & ~n17626 ;
  assign n17633 = ~n17627 & n17632 ;
  assign n17634 = ~n17625 & n17633 ;
  assign n17635 = ~n17631 & n17634 ;
  assign n17616 = n17265 & ~n17614 ;
  assign n17615 = ~n17265 & n17614 ;
  assign n17617 = n17223 & ~n17615 ;
  assign n17618 = ~n17616 & n17617 ;
  assign n17611 = n17238 & ~n17609 ;
  assign n17610 = ~n17238 & n17609 ;
  assign n17612 = n767 & ~n17610 ;
  assign n17613 = ~n17611 & n17612 ;
  assign n17608 = n733 & ~n1792 ;
  assign n17619 = n2145 & ~n17608 ;
  assign n17620 = ~n17613 & n17619 ;
  assign n17621 = ~n17618 & n17620 ;
  assign n17636 = \P1_state_reg[0]/NET0131  & ~n17621 ;
  assign n17637 = ~n17635 & n17636 ;
  assign n17638 = ~n12811 & ~n17637 ;
  assign n17640 = ~n17180 & ~n17181 ;
  assign n17661 = n17240 & ~n17640 ;
  assign n17660 = ~n17240 & n17640 ;
  assign n17662 = n767 & ~n17660 ;
  assign n17663 = ~n17661 & n17662 ;
  assign n17645 = ~n17131 & ~n17132 ;
  assign n17657 = ~n17267 & n17645 ;
  assign n17656 = n17267 & ~n17645 ;
  assign n17658 = n17223 & ~n17656 ;
  assign n17659 = ~n17657 & n17658 ;
  assign n17655 = n733 & ~n1766 ;
  assign n17664 = n2145 & ~n17655 ;
  assign n17665 = ~n17659 & n17664 ;
  assign n17666 = ~n17663 & n17665 ;
  assign n17647 = n17153 & n17645 ;
  assign n17646 = ~n17153 & ~n17645 ;
  assign n17648 = n2238 & ~n17646 ;
  assign n17649 = ~n17647 & n17648 ;
  assign n17642 = n17202 & n17640 ;
  assign n17641 = ~n17202 & ~n17640 ;
  assign n17643 = n734 & ~n17641 ;
  assign n17644 = ~n17642 & n17643 ;
  assign n17650 = ~n1766 & n17223 ;
  assign n17639 = \P3_addr_reg[6]/NET0131  & n767 ;
  assign n17651 = ~n2145 & ~n17639 ;
  assign n17652 = ~n17650 & n17651 ;
  assign n17653 = ~n17644 & n17652 ;
  assign n17654 = ~n17649 & n17653 ;
  assign n17667 = \P1_state_reg[0]/NET0131  & ~n17654 ;
  assign n17668 = ~n17666 & n17667 ;
  assign n17669 = ~n12853 & ~n17668 ;
  assign n17676 = ~n17127 & ~n17128 ;
  assign n17692 = n17271 & ~n17676 ;
  assign n17691 = ~n17271 & n17676 ;
  assign n17693 = n17223 & ~n17691 ;
  assign n17694 = ~n17692 & n17693 ;
  assign n17671 = ~n17177 & ~n17209 ;
  assign n17688 = ~n17244 & n17671 ;
  assign n17687 = n17244 & ~n17671 ;
  assign n17689 = n767 & ~n17687 ;
  assign n17690 = ~n17688 & n17689 ;
  assign n17686 = n733 & n1702 ;
  assign n17695 = n2145 & ~n17686 ;
  assign n17696 = ~n17690 & n17695 ;
  assign n17697 = ~n17694 & n17696 ;
  assign n17678 = n17157 & n17676 ;
  assign n17677 = ~n17157 & ~n17676 ;
  assign n17679 = n2238 & ~n17677 ;
  assign n17680 = ~n17678 & n17679 ;
  assign n17673 = n17206 & ~n17671 ;
  assign n17672 = ~n17206 & n17671 ;
  assign n17674 = n734 & ~n17672 ;
  assign n17675 = ~n17673 & n17674 ;
  assign n17681 = n1702 & n17223 ;
  assign n17670 = \P3_addr_reg[8]/NET0131  & n767 ;
  assign n17682 = ~n2145 & ~n17670 ;
  assign n17683 = ~n17681 & n17682 ;
  assign n17684 = ~n17675 & n17683 ;
  assign n17685 = ~n17680 & n17684 ;
  assign n17698 = \P1_state_reg[0]/NET0131  & ~n17685 ;
  assign n17699 = ~n17697 & n17698 ;
  assign n17700 = ~n11613 & ~n17699 ;
  assign n17718 = ~n17567 & ~n17570 ;
  assign n17719 = ~n17446 & ~n17504 ;
  assign n17720 = ~n17447 & n17473 ;
  assign n17721 = n17719 & ~n17720 ;
  assign n17722 = ~n17505 & ~n17721 ;
  assign n17723 = ~n17571 & n17722 ;
  assign n17724 = n17718 & ~n17723 ;
  assign n17725 = ~n17568 & ~n17724 ;
  assign n17726 = ~\P3_reg2_reg[19]/NET0131  & ~n1108 ;
  assign n17727 = \P3_reg2_reg[19]/NET0131  & n1108 ;
  assign n17728 = ~n17726 & ~n17727 ;
  assign n17730 = n17725 & ~n17728 ;
  assign n17729 = ~n17725 & n17728 ;
  assign n17731 = n2238 & ~n17729 ;
  assign n17732 = ~n17730 & n17731 ;
  assign n17701 = ~n17554 & ~n17557 ;
  assign n17702 = ~n17432 & ~n17487 ;
  assign n17703 = ~n17433 & n17466 ;
  assign n17704 = n17702 & ~n17703 ;
  assign n17705 = ~n17488 & ~n17704 ;
  assign n17706 = ~n17559 & n17705 ;
  assign n17707 = n17701 & ~n17706 ;
  assign n17708 = ~n17555 & ~n17707 ;
  assign n17709 = ~\P3_reg1_reg[19]/NET0131  & ~n1108 ;
  assign n17710 = \P3_reg1_reg[19]/NET0131  & n1108 ;
  assign n17711 = ~n17709 & ~n17710 ;
  assign n17713 = n17708 & ~n17711 ;
  assign n17712 = ~n17708 & n17711 ;
  assign n17714 = n734 & ~n17712 ;
  assign n17715 = ~n17713 & n17714 ;
  assign n17717 = \P3_addr_reg[19]/NET0131  & n767 ;
  assign n17716 = n1108 & n17223 ;
  assign n17733 = ~n2145 & ~n17716 ;
  assign n17734 = ~n17717 & n17733 ;
  assign n17735 = ~n17715 & n17734 ;
  assign n17736 = ~n17732 & n17735 ;
  assign n17749 = ~n17441 & n17702 ;
  assign n17750 = n17433 & ~n17487 ;
  assign n17751 = ~n17488 & ~n17750 ;
  assign n17752 = ~n17749 & n17751 ;
  assign n17753 = ~n17559 & n17752 ;
  assign n17754 = n17701 & ~n17753 ;
  assign n17755 = ~n17555 & ~n17754 ;
  assign n17757 = ~n17711 & ~n17755 ;
  assign n17756 = n17711 & n17755 ;
  assign n17758 = n767 & ~n17756 ;
  assign n17759 = ~n17757 & n17758 ;
  assign n17738 = ~n17455 & n17719 ;
  assign n17739 = n17447 & ~n17504 ;
  assign n17740 = ~n17505 & ~n17739 ;
  assign n17741 = ~n17571 & n17740 ;
  assign n17742 = ~n17738 & n17741 ;
  assign n17743 = n17718 & ~n17742 ;
  assign n17744 = ~n17568 & ~n17743 ;
  assign n17746 = n17728 & n17744 ;
  assign n17745 = ~n17728 & ~n17744 ;
  assign n17747 = n17223 & ~n17745 ;
  assign n17748 = ~n17746 & n17747 ;
  assign n17737 = n733 & n1108 ;
  assign n17760 = n2145 & ~n17737 ;
  assign n17761 = ~n17748 & n17760 ;
  assign n17762 = ~n17759 & n17761 ;
  assign n17763 = \P1_state_reg[0]/NET0131  & ~n17762 ;
  assign n17764 = ~n17736 & n17763 ;
  assign n17765 = ~n6525 & ~n17764 ;
  assign n17767 = ~n17449 & ~n17452 ;
  assign n17784 = n17511 & n17767 ;
  assign n17783 = ~n17511 & ~n17767 ;
  assign n17785 = n17223 & ~n17783 ;
  assign n17786 = ~n17784 & n17785 ;
  assign n17772 = ~n17435 & ~n17438 ;
  assign n17788 = n17497 & ~n17772 ;
  assign n17787 = ~n17497 & n17772 ;
  assign n17789 = n767 & ~n17787 ;
  assign n17790 = ~n17788 & n17789 ;
  assign n17782 = n733 & n1542 ;
  assign n17791 = n2145 & ~n17782 ;
  assign n17792 = ~n17790 & n17791 ;
  assign n17793 = ~n17786 & n17792 ;
  assign n17769 = n17536 & n17767 ;
  assign n17768 = ~n17536 & ~n17767 ;
  assign n17770 = n2238 & ~n17768 ;
  assign n17771 = ~n17769 & n17770 ;
  assign n17774 = n17525 & n17772 ;
  assign n17773 = ~n17525 & ~n17772 ;
  assign n17775 = n734 & ~n17773 ;
  assign n17776 = ~n17774 & n17775 ;
  assign n17777 = n1542 & n17223 ;
  assign n17766 = \P3_addr_reg[14]/NET0131  & n767 ;
  assign n17778 = ~n2145 & ~n17766 ;
  assign n17779 = ~n17777 & n17778 ;
  assign n17780 = ~n17776 & n17779 ;
  assign n17781 = ~n17771 & n17780 ;
  assign n17794 = \P1_state_reg[0]/NET0131  & ~n17781 ;
  assign n17795 = ~n17793 & n17794 ;
  assign n17796 = ~n10650 & ~n17795 ;
  assign n17803 = ~n17570 & ~n17571 ;
  assign n17814 = ~n17384 & ~n17413 ;
  assign n17815 = n17450 & ~n17814 ;
  assign n17816 = ~n17452 & ~n17815 ;
  assign n17817 = n17719 & ~n17816 ;
  assign n17818 = n17740 & ~n17817 ;
  assign n17820 = ~n17803 & n17818 ;
  assign n17819 = n17803 & ~n17818 ;
  assign n17821 = n17223 & ~n17819 ;
  assign n17822 = ~n17820 & n17821 ;
  assign n17798 = ~n17557 & ~n17559 ;
  assign n17824 = n17752 & ~n17798 ;
  assign n17823 = ~n17752 & n17798 ;
  assign n17825 = n767 & ~n17823 ;
  assign n17826 = ~n17824 & n17825 ;
  assign n17813 = n733 & ~n1164 ;
  assign n17827 = n2145 & ~n17813 ;
  assign n17828 = ~n17826 & n17827 ;
  assign n17829 = ~n17822 & n17828 ;
  assign n17805 = n17722 & n17803 ;
  assign n17804 = ~n17722 & ~n17803 ;
  assign n17806 = n2238 & ~n17804 ;
  assign n17807 = ~n17805 & n17806 ;
  assign n17800 = n17705 & n17798 ;
  assign n17799 = ~n17705 & ~n17798 ;
  assign n17801 = n734 & ~n17799 ;
  assign n17802 = ~n17800 & n17801 ;
  assign n17808 = ~n1164 & n17223 ;
  assign n17797 = \P3_addr_reg[17]/NET0131  & n767 ;
  assign n17809 = ~n2145 & ~n17797 ;
  assign n17810 = ~n17808 & n17809 ;
  assign n17811 = ~n17802 & n17810 ;
  assign n17812 = ~n17807 & n17811 ;
  assign n17830 = \P1_state_reg[0]/NET0131  & ~n17812 ;
  assign n17831 = ~n17829 & n17830 ;
  assign n17832 = ~n8593 & ~n17831 ;
  assign n17839 = ~n17125 & ~n17126 ;
  assign n17841 = n17273 & ~n17839 ;
  assign n17840 = ~n17273 & n17839 ;
  assign n17842 = n17223 & ~n17840 ;
  assign n17843 = ~n17841 & n17842 ;
  assign n17834 = ~n17176 & ~n17208 ;
  assign n17836 = ~n17246 & n17834 ;
  assign n17835 = n17246 & ~n17834 ;
  assign n17837 = n767 & ~n17835 ;
  assign n17838 = ~n17836 & n17837 ;
  assign n17833 = n733 & n1675 ;
  assign n17844 = n2145 & ~n17833 ;
  assign n17845 = ~n17838 & n17844 ;
  assign n17846 = ~n17843 & n17845 ;
  assign n17853 = n17159 & n17839 ;
  assign n17852 = ~n17159 & ~n17839 ;
  assign n17854 = n2238 & ~n17852 ;
  assign n17855 = ~n17853 & n17854 ;
  assign n17849 = n17353 & n17834 ;
  assign n17848 = ~n17353 & ~n17834 ;
  assign n17850 = n734 & ~n17848 ;
  assign n17851 = ~n17849 & n17850 ;
  assign n17856 = n1675 & n17223 ;
  assign n17847 = \P3_addr_reg[9]/NET0131  & n767 ;
  assign n17857 = ~n2145 & ~n17847 ;
  assign n17858 = ~n17856 & n17857 ;
  assign n17859 = ~n17851 & n17858 ;
  assign n17860 = ~n17855 & n17859 ;
  assign n17861 = \P1_state_reg[0]/NET0131  & ~n17860 ;
  assign n17862 = ~n17846 & n17861 ;
  assign n17863 = ~n10284 & ~n17862 ;
  assign n17870 = ~n17178 & ~n17179 ;
  assign n17886 = n17242 & ~n17870 ;
  assign n17885 = ~n17242 & n17870 ;
  assign n17887 = n767 & ~n17885 ;
  assign n17888 = ~n17886 & n17887 ;
  assign n17865 = ~n17129 & ~n17130 ;
  assign n17882 = ~n17269 & n17865 ;
  assign n17881 = n17269 & ~n17865 ;
  assign n17883 = n17223 & ~n17881 ;
  assign n17884 = ~n17882 & n17883 ;
  assign n17880 = n733 & n1742 ;
  assign n17889 = n2145 & ~n17880 ;
  assign n17890 = ~n17884 & n17889 ;
  assign n17891 = ~n17888 & n17890 ;
  assign n17872 = n17204 & n17870 ;
  assign n17871 = ~n17204 & ~n17870 ;
  assign n17873 = n734 & ~n17871 ;
  assign n17874 = ~n17872 & n17873 ;
  assign n17867 = n17155 & n17865 ;
  assign n17866 = ~n17155 & ~n17865 ;
  assign n17868 = n2238 & ~n17866 ;
  assign n17869 = ~n17867 & n17868 ;
  assign n17875 = n1742 & n17223 ;
  assign n17864 = \P3_addr_reg[7]/NET0131  & n767 ;
  assign n17876 = ~n2145 & ~n17864 ;
  assign n17877 = ~n17875 & n17876 ;
  assign n17878 = ~n17869 & n17877 ;
  assign n17879 = ~n17874 & n17878 ;
  assign n17892 = \P1_state_reg[0]/NET0131  & ~n17879 ;
  assign n17893 = ~n17891 & n17892 ;
  assign n17894 = ~n12894 & ~n17893 ;
  assign n17895 = ~\P1_state_reg[0]/NET0131  & ~\P3_reg3_reg[2]/NET0131  ;
  assign n17896 = \P3_addr_reg[2]/NET0131  & n767 ;
  assign n17908 = ~n2145 & ~n17896 ;
  assign n17903 = ~n17188 & ~n17189 ;
  assign n17904 = n17194 & ~n17903 ;
  assign n17905 = ~n17194 & n17903 ;
  assign n17906 = ~n17904 & ~n17905 ;
  assign n17907 = n734 & n17906 ;
  assign n17897 = n1842 & n17223 ;
  assign n17898 = ~n17139 & ~n17140 ;
  assign n17899 = n17145 & ~n17898 ;
  assign n17900 = ~n17145 & n17898 ;
  assign n17901 = ~n17899 & ~n17900 ;
  assign n17902 = n2238 & n17901 ;
  assign n17909 = ~n17897 & ~n17902 ;
  assign n17910 = ~n17907 & n17909 ;
  assign n17911 = n17908 & n17910 ;
  assign n17917 = ~n17232 & n17903 ;
  assign n17918 = n17232 & ~n17903 ;
  assign n17919 = ~n17917 & ~n17918 ;
  assign n17920 = n767 & n17919 ;
  assign n17912 = ~n17259 & n17898 ;
  assign n17913 = n17259 & ~n17898 ;
  assign n17914 = ~n17912 & ~n17913 ;
  assign n17915 = n17223 & n17914 ;
  assign n17916 = n733 & n1842 ;
  assign n17921 = n2145 & ~n17916 ;
  assign n17922 = ~n17915 & n17921 ;
  assign n17923 = ~n17920 & n17922 ;
  assign n17924 = ~n17911 & ~n17923 ;
  assign n17925 = \P1_state_reg[0]/NET0131  & ~n17924 ;
  assign n17926 = ~n17895 & ~n17925 ;
  assign n17927 = \P3_addr_reg[3]/NET0131  & n767 ;
  assign n17939 = ~n2145 & ~n17927 ;
  assign n17934 = ~n17137 & ~n17138 ;
  assign n17935 = ~n17147 & ~n17934 ;
  assign n17936 = n17147 & n17934 ;
  assign n17937 = ~n17935 & ~n17936 ;
  assign n17938 = n2238 & n17937 ;
  assign n17928 = n1857 & n17223 ;
  assign n17929 = ~n17186 & ~n17187 ;
  assign n17930 = ~n17196 & ~n17929 ;
  assign n17931 = n17196 & n17929 ;
  assign n17932 = ~n17930 & ~n17931 ;
  assign n17933 = n734 & n17932 ;
  assign n17940 = ~n17928 & ~n17933 ;
  assign n17941 = ~n17938 & n17940 ;
  assign n17942 = n17939 & n17941 ;
  assign n17948 = ~n17234 & n17929 ;
  assign n17949 = n17234 & ~n17929 ;
  assign n17950 = ~n17948 & ~n17949 ;
  assign n17951 = n767 & n17950 ;
  assign n17944 = n17261 & ~n17934 ;
  assign n17945 = ~n17261 & n17934 ;
  assign n17946 = ~n17944 & ~n17945 ;
  assign n17947 = n17223 & n17946 ;
  assign n17943 = n733 & n1857 ;
  assign n17952 = n2145 & ~n17943 ;
  assign n17953 = ~n17947 & n17952 ;
  assign n17954 = ~n17951 & n17953 ;
  assign n17955 = \P1_state_reg[0]/NET0131  & ~n17954 ;
  assign n17956 = ~n17942 & n17955 ;
  assign n17957 = ~n14247 & ~n17956 ;
  assign n17958 = \P3_addr_reg[4]/NET0131  & n767 ;
  assign n17970 = ~n2145 & ~n17958 ;
  assign n17965 = ~n17135 & ~n17136 ;
  assign n17966 = ~n17149 & ~n17965 ;
  assign n17967 = n17149 & n17965 ;
  assign n17968 = ~n17966 & ~n17967 ;
  assign n17969 = n2238 & n17968 ;
  assign n17959 = ~n1818 & n17223 ;
  assign n17960 = ~n17184 & ~n17185 ;
  assign n17961 = ~n17198 & ~n17960 ;
  assign n17962 = n17198 & n17960 ;
  assign n17963 = ~n17961 & ~n17962 ;
  assign n17964 = n734 & n17963 ;
  assign n17971 = ~n17959 & ~n17964 ;
  assign n17972 = ~n17969 & n17971 ;
  assign n17973 = n17970 & n17972 ;
  assign n17979 = ~n17236 & n17960 ;
  assign n17980 = n17236 & ~n17960 ;
  assign n17981 = ~n17979 & ~n17980 ;
  assign n17982 = n767 & n17981 ;
  assign n17975 = n17263 & ~n17965 ;
  assign n17976 = ~n17263 & n17965 ;
  assign n17977 = ~n17975 & ~n17976 ;
  assign n17978 = n17223 & n17977 ;
  assign n17974 = n733 & ~n1818 ;
  assign n17983 = n2145 & ~n17974 ;
  assign n17984 = ~n17978 & n17983 ;
  assign n17985 = ~n17982 & n17984 ;
  assign n17986 = \P1_state_reg[0]/NET0131  & ~n17985 ;
  assign n17987 = ~n17973 & n17986 ;
  assign n17988 = ~n13620 & ~n17987 ;
  assign n17989 = ~\P1_state_reg[0]/NET0131  & ~\P3_reg3_reg[1]/NET0131  ;
  assign n17996 = ~n17141 & ~n17142 ;
  assign n17997 = ~n17257 & n17996 ;
  assign n17998 = n17257 & ~n17996 ;
  assign n17999 = ~n17997 & ~n17998 ;
  assign n18000 = n17223 & n17999 ;
  assign n17991 = ~n17190 & ~n17191 ;
  assign n17992 = n17230 & ~n17991 ;
  assign n17993 = ~n17230 & n17991 ;
  assign n17994 = ~n17992 & ~n17993 ;
  assign n17995 = n767 & n17994 ;
  assign n17990 = n733 & ~n1881 ;
  assign n18001 = n2145 & ~n17990 ;
  assign n18002 = ~n17995 & n18001 ;
  assign n18003 = ~n18000 & n18002 ;
  assign n18004 = ~n1881 & n17223 ;
  assign n18014 = ~n2145 & ~n18004 ;
  assign n18013 = \P3_addr_reg[1]/NET0131  & n767 ;
  assign n18005 = n17143 & ~n17996 ;
  assign n18006 = ~n17143 & n17996 ;
  assign n18007 = ~n18005 & ~n18006 ;
  assign n18008 = n2238 & n18007 ;
  assign n18009 = ~n17192 & n17991 ;
  assign n18010 = n17192 & ~n17991 ;
  assign n18011 = ~n18009 & ~n18010 ;
  assign n18012 = n734 & n18011 ;
  assign n18015 = ~n18008 & ~n18012 ;
  assign n18016 = ~n18013 & n18015 ;
  assign n18017 = n18014 & n18016 ;
  assign n18018 = ~n18003 & ~n18017 ;
  assign n18019 = \P1_state_reg[0]/NET0131  & ~n18018 ;
  assign n18020 = ~n17989 & ~n18019 ;
  assign n18021 = ~n2726 & ~n6095 ;
  assign n18022 = \P1_state_reg[0]/NET0131  & ~n18021 ;
  assign n18023 = ~n767 & ~n2145 ;
  assign n18024 = \P1_state_reg[0]/NET0131  & ~n18023 ;
  assign n18025 = \P1_state_reg[0]/NET0131  & n6095 ;
  assign n18026 = \P1_state_reg[0]/NET0131  & n5585 ;
  assign n18027 = \P1_state_reg[0]/NET0131  & n2145 ;
  assign n18028 = \P1_reg2_reg[27]/NET0131  & ~n10960 ;
  assign n18029 = \P1_reg2_reg[27]/NET0131  & ~n6113 ;
  assign n18031 = n6113 & ~n6603 ;
  assign n18032 = ~n18029 & ~n18031 ;
  assign n18033 = n6282 & ~n18032 ;
  assign n18034 = n6113 & ~n6644 ;
  assign n18035 = ~n18029 & ~n18034 ;
  assign n18036 = n6207 & ~n18035 ;
  assign n18037 = n6113 & ~n8133 ;
  assign n18030 = ~n15534 & n18029 ;
  assign n18038 = n3433 & n4112 ;
  assign n18039 = ~n18030 & ~n18038 ;
  assign n18040 = ~n18037 & n18039 ;
  assign n18041 = ~n18036 & n18040 ;
  assign n18042 = ~n18033 & n18041 ;
  assign n18043 = n9044 & ~n18042 ;
  assign n18044 = ~n18028 & ~n18043 ;
  assign n18046 = \P1_reg1_reg[27]/NET0131  & ~n6683 ;
  assign n18047 = ~n6603 & n9045 ;
  assign n18048 = ~n18046 & ~n18047 ;
  assign n18049 = n6282 & ~n18048 ;
  assign n18050 = ~n6644 & n9045 ;
  assign n18051 = ~n18046 & ~n18050 ;
  assign n18052 = n6207 & ~n18051 ;
  assign n18045 = \P1_reg1_reg[27]/NET0131  & ~n11258 ;
  assign n18053 = ~n8133 & n9045 ;
  assign n18054 = ~n18045 & ~n18053 ;
  assign n18055 = ~n18052 & n18054 ;
  assign n18056 = ~n18049 & n18055 ;
  assign n18058 = n3077 & n6095 ;
  assign n18060 = n3077 & ~n6568 ;
  assign n18061 = n6568 & ~n9420 ;
  assign n18062 = ~n18060 & ~n18061 ;
  assign n18063 = n6207 & ~n18062 ;
  assign n18067 = n6568 & n9433 ;
  assign n18068 = ~n18060 & ~n18067 ;
  assign n18069 = n6282 & ~n18068 ;
  assign n18070 = n6568 & n9441 ;
  assign n18071 = ~n18060 & ~n18070 ;
  assign n18072 = n4011 & ~n18071 ;
  assign n18064 = n6568 & n9425 ;
  assign n18065 = ~n18060 & ~n18064 ;
  assign n18066 = n6359 & ~n18065 ;
  assign n18059 = n3072 & ~n6649 ;
  assign n18073 = n3077 & ~n6666 ;
  assign n18074 = ~n18059 & ~n18073 ;
  assign n18075 = ~n18066 & n18074 ;
  assign n18076 = ~n18072 & n18075 ;
  assign n18077 = ~n18069 & n18076 ;
  assign n18078 = ~n18063 & n18077 ;
  assign n18079 = n6097 & ~n18078 ;
  assign n18080 = ~n18058 & ~n18079 ;
  assign n18081 = \P1_state_reg[0]/NET0131  & ~n18080 ;
  assign n18057 = n3077 & n4130 ;
  assign n18082 = ~n16431 & ~n18057 ;
  assign n18083 = ~n18081 & n18082 ;
  assign n18084 = \P1_reg1_reg[21]/NET0131  & ~n6078 ;
  assign n18085 = \P1_reg1_reg[21]/NET0131  & n6095 ;
  assign n18087 = \P1_reg1_reg[21]/NET0131  & ~n6683 ;
  assign n18097 = n6683 & n9329 ;
  assign n18098 = ~n18087 & ~n18097 ;
  assign n18099 = n6359 & ~n18098 ;
  assign n18091 = n6683 & ~n9318 ;
  assign n18092 = ~n18087 & ~n18091 ;
  assign n18093 = n6282 & ~n18092 ;
  assign n18086 = \P1_reg1_reg[21]/NET0131  & ~n7806 ;
  assign n18100 = n6683 & n9346 ;
  assign n18101 = ~n18086 & ~n18100 ;
  assign n18102 = ~n18093 & n18101 ;
  assign n18103 = ~n18099 & n18102 ;
  assign n18088 = n6683 & n9312 ;
  assign n18089 = ~n18087 & ~n18088 ;
  assign n18090 = n4011 & ~n18089 ;
  assign n18094 = n6683 & ~n9324 ;
  assign n18095 = ~n18087 & ~n18094 ;
  assign n18096 = n6207 & ~n18095 ;
  assign n18104 = ~n18090 & ~n18096 ;
  assign n18105 = n18103 & n18104 ;
  assign n18106 = n6097 & ~n18105 ;
  assign n18107 = ~n18085 & ~n18106 ;
  assign n18108 = \P1_state_reg[0]/NET0131  & ~n18107 ;
  assign n18109 = ~n18084 & ~n18108 ;
  assign n18110 = \P2_reg0_reg[28]/NET0131  & ~n6706 ;
  assign n18111 = ~n6801 & n9533 ;
  assign n18112 = ~n18110 & ~n18111 ;
  assign n18113 = n5329 & ~n18112 ;
  assign n18114 = n5526 & ~n6818 ;
  assign n18115 = n6835 & ~n18114 ;
  assign n18116 = n9533 & ~n18115 ;
  assign n18117 = ~n7984 & n9530 ;
  assign n18118 = \P2_reg0_reg[28]/NET0131  & ~n18117 ;
  assign n18119 = ~n18116 & ~n18118 ;
  assign n18120 = ~n18113 & n18119 ;
  assign n18121 = \P2_reg2_reg[24]/NET0131  & ~n5589 ;
  assign n18122 = \P2_reg2_reg[24]/NET0131  & n5585 ;
  assign n18123 = n4219 & ~n8921 ;
  assign n18124 = \P2_reg2_reg[24]/NET0131  & ~n9772 ;
  assign n18125 = n4643 & n5574 ;
  assign n18126 = ~n18124 & ~n18125 ;
  assign n18127 = ~n18123 & n18126 ;
  assign n18128 = n5583 & ~n18127 ;
  assign n18129 = ~n18122 & ~n18128 ;
  assign n18130 = \P1_state_reg[0]/NET0131  & ~n18129 ;
  assign n18131 = ~n18121 & ~n18130 ;
  assign n18132 = \P1_reg2_reg[26]/NET0131  & ~n10960 ;
  assign n18134 = \P1_reg2_reg[26]/NET0131  & ~n6113 ;
  assign n18135 = n6113 & ~n7156 ;
  assign n18136 = ~n18134 & ~n18135 ;
  assign n18137 = n6282 & ~n18136 ;
  assign n18138 = n6113 & ~n7192 ;
  assign n18139 = ~n18134 & ~n18138 ;
  assign n18140 = n6207 & ~n18139 ;
  assign n18141 = n6113 & n7203 ;
  assign n18142 = ~n18134 & ~n18141 ;
  assign n18143 = n6359 & ~n18142 ;
  assign n18144 = n6113 & ~n7200 ;
  assign n18145 = ~n18134 & ~n18144 ;
  assign n18146 = n4011 & ~n18145 ;
  assign n18133 = n3523 & n4112 ;
  assign n18147 = n3518 & n6113 ;
  assign n18148 = ~n18134 & ~n18147 ;
  assign n18149 = n6365 & ~n18148 ;
  assign n18150 = ~n18133 & ~n18149 ;
  assign n18151 = ~n18146 & n18150 ;
  assign n18152 = ~n18143 & n18151 ;
  assign n18153 = ~n18140 & n18152 ;
  assign n18154 = ~n18137 & n18153 ;
  assign n18155 = n9044 & ~n18154 ;
  assign n18156 = ~n18132 & ~n18155 ;
  assign n18157 = \P1_reg2_reg[24]/NET0131  & ~n10960 ;
  assign n18159 = \P1_reg2_reg[24]/NET0131  & ~n6113 ;
  assign n18163 = n6113 & ~n7031 ;
  assign n18164 = ~n18159 & ~n18163 ;
  assign n18165 = n6207 & ~n18164 ;
  assign n18160 = n6113 & ~n6964 ;
  assign n18161 = ~n18159 & ~n18160 ;
  assign n18162 = n6282 & ~n18161 ;
  assign n18166 = n6113 & n7044 ;
  assign n18167 = ~n18159 & ~n18166 ;
  assign n18168 = n4011 & ~n18167 ;
  assign n18169 = n6113 & n7049 ;
  assign n18170 = ~n18159 & ~n18169 ;
  assign n18171 = n6359 & ~n18170 ;
  assign n18158 = n3544 & n4112 ;
  assign n18172 = n3539 & n6113 ;
  assign n18173 = ~n18159 & ~n18172 ;
  assign n18174 = n6365 & ~n18173 ;
  assign n18175 = ~n18158 & ~n18174 ;
  assign n18176 = ~n18171 & n18175 ;
  assign n18177 = ~n18168 & n18176 ;
  assign n18178 = ~n18162 & n18177 ;
  assign n18179 = ~n18165 & n18178 ;
  assign n18180 = n9044 & ~n18179 ;
  assign n18181 = ~n18157 & ~n18180 ;
  assign n18182 = \P1_rd_reg/NET0131  & ~\P2_rd_reg/NET0131  ;
  assign n18183 = ~\P1_rd_reg/NET0131  & \P2_rd_reg/NET0131  ;
  assign n18184 = ~n18182 & ~n18183 ;
  assign n18185 = ~\P3_rd_reg/NET0131  & ~n18184 ;
  assign n18186 = \P1_addr_reg[0]/NET0131  & \P2_addr_reg[0]/NET0131  ;
  assign n18187 = ~\P1_addr_reg[0]/NET0131  & ~\P2_addr_reg[0]/NET0131  ;
  assign n18188 = ~n18186 & ~n18187 ;
  assign n18189 = ~\P3_addr_reg[0]/NET0131  & n18188 ;
  assign n18190 = \P3_addr_reg[0]/NET0131  & ~n18188 ;
  assign n18191 = ~n18189 & ~n18190 ;
  assign n18192 = \P1_addr_reg[10]/NET0131  & \P2_addr_reg[10]/NET0131  ;
  assign n18193 = ~\P1_addr_reg[10]/NET0131  & ~\P2_addr_reg[10]/NET0131  ;
  assign n18194 = ~n18192 & ~n18193 ;
  assign n18195 = ~\P1_addr_reg[9]/NET0131  & ~\P2_addr_reg[9]/NET0131  ;
  assign n18196 = \P1_addr_reg[9]/NET0131  & \P2_addr_reg[9]/NET0131  ;
  assign n18197 = ~\P1_addr_reg[8]/NET0131  & ~\P2_addr_reg[8]/NET0131  ;
  assign n18198 = \P1_addr_reg[8]/NET0131  & \P2_addr_reg[8]/NET0131  ;
  assign n18199 = ~\P1_addr_reg[7]/NET0131  & ~\P2_addr_reg[7]/NET0131  ;
  assign n18200 = \P1_addr_reg[7]/NET0131  & \P2_addr_reg[7]/NET0131  ;
  assign n18201 = ~\P1_addr_reg[6]/NET0131  & ~\P2_addr_reg[6]/NET0131  ;
  assign n18202 = \P1_addr_reg[6]/NET0131  & \P2_addr_reg[6]/NET0131  ;
  assign n18203 = ~\P1_addr_reg[5]/NET0131  & ~\P2_addr_reg[5]/NET0131  ;
  assign n18204 = \P1_addr_reg[5]/NET0131  & \P2_addr_reg[5]/NET0131  ;
  assign n18205 = ~\P1_addr_reg[4]/NET0131  & ~\P2_addr_reg[4]/NET0131  ;
  assign n18206 = \P1_addr_reg[4]/NET0131  & \P2_addr_reg[4]/NET0131  ;
  assign n18207 = ~\P1_addr_reg[3]/NET0131  & ~\P2_addr_reg[3]/NET0131  ;
  assign n18208 = \P1_addr_reg[3]/NET0131  & \P2_addr_reg[3]/NET0131  ;
  assign n18209 = ~\P1_addr_reg[2]/NET0131  & ~\P2_addr_reg[2]/NET0131  ;
  assign n18210 = \P1_addr_reg[2]/NET0131  & \P2_addr_reg[2]/NET0131  ;
  assign n18211 = ~\P1_addr_reg[1]/NET0131  & ~\P2_addr_reg[1]/NET0131  ;
  assign n18212 = \P1_addr_reg[1]/NET0131  & \P2_addr_reg[1]/NET0131  ;
  assign n18213 = ~n18186 & ~n18212 ;
  assign n18214 = ~n18211 & ~n18213 ;
  assign n18215 = ~n18210 & ~n18214 ;
  assign n18216 = ~n18209 & ~n18215 ;
  assign n18217 = ~n18208 & ~n18216 ;
  assign n18218 = ~n18207 & ~n18217 ;
  assign n18219 = ~n18206 & ~n18218 ;
  assign n18220 = ~n18205 & ~n18219 ;
  assign n18221 = ~n18204 & ~n18220 ;
  assign n18222 = ~n18203 & ~n18221 ;
  assign n18223 = ~n18202 & ~n18222 ;
  assign n18224 = ~n18201 & ~n18223 ;
  assign n18225 = ~n18200 & ~n18224 ;
  assign n18226 = ~n18199 & ~n18225 ;
  assign n18227 = ~n18198 & ~n18226 ;
  assign n18228 = ~n18197 & ~n18227 ;
  assign n18229 = ~n18196 & ~n18228 ;
  assign n18230 = ~n18195 & ~n18229 ;
  assign n18231 = ~n18194 & n18230 ;
  assign n18232 = n18194 & ~n18230 ;
  assign n18233 = ~n18231 & ~n18232 ;
  assign n18234 = ~\P3_addr_reg[10]/NET0131  & ~n18233 ;
  assign n18235 = \P3_addr_reg[10]/NET0131  & n18233 ;
  assign n18236 = ~n18234 & ~n18235 ;
  assign n18237 = ~n18195 & ~n18196 ;
  assign n18238 = n18228 & ~n18237 ;
  assign n18239 = ~n18228 & n18237 ;
  assign n18240 = ~n18238 & ~n18239 ;
  assign n18241 = ~\P3_addr_reg[9]/NET0131  & ~n18240 ;
  assign n18242 = \P3_addr_reg[9]/NET0131  & n18240 ;
  assign n18243 = ~n18197 & ~n18198 ;
  assign n18244 = n18226 & ~n18243 ;
  assign n18245 = ~n18226 & n18243 ;
  assign n18246 = ~n18244 & ~n18245 ;
  assign n18247 = ~\P3_addr_reg[8]/NET0131  & ~n18246 ;
  assign n18248 = \P3_addr_reg[8]/NET0131  & n18246 ;
  assign n18249 = ~n18199 & ~n18200 ;
  assign n18250 = n18224 & ~n18249 ;
  assign n18251 = ~n18224 & n18249 ;
  assign n18252 = ~n18250 & ~n18251 ;
  assign n18253 = ~\P3_addr_reg[7]/NET0131  & ~n18252 ;
  assign n18254 = \P3_addr_reg[7]/NET0131  & n18252 ;
  assign n18255 = ~n18201 & ~n18202 ;
  assign n18256 = n18222 & ~n18255 ;
  assign n18257 = ~n18222 & n18255 ;
  assign n18258 = ~n18256 & ~n18257 ;
  assign n18259 = ~\P3_addr_reg[6]/NET0131  & ~n18258 ;
  assign n18260 = \P3_addr_reg[6]/NET0131  & n18258 ;
  assign n18261 = ~n18203 & ~n18204 ;
  assign n18262 = n18220 & ~n18261 ;
  assign n18263 = ~n18220 & n18261 ;
  assign n18264 = ~n18262 & ~n18263 ;
  assign n18265 = ~\P3_addr_reg[5]/NET0131  & ~n18264 ;
  assign n18266 = \P3_addr_reg[5]/NET0131  & n18264 ;
  assign n18267 = ~n18205 & ~n18206 ;
  assign n18268 = n18218 & ~n18267 ;
  assign n18269 = ~n18218 & n18267 ;
  assign n18270 = ~n18268 & ~n18269 ;
  assign n18271 = \P3_addr_reg[4]/NET0131  & n18270 ;
  assign n18272 = ~n18207 & ~n18208 ;
  assign n18273 = n18216 & ~n18272 ;
  assign n18274 = ~n18216 & n18272 ;
  assign n18275 = ~n18273 & ~n18274 ;
  assign n18276 = ~\P3_addr_reg[3]/NET0131  & ~n18275 ;
  assign n18277 = \P3_addr_reg[3]/NET0131  & n18275 ;
  assign n18278 = ~n18209 & ~n18210 ;
  assign n18279 = n18214 & ~n18278 ;
  assign n18280 = ~n18214 & n18278 ;
  assign n18281 = ~n18279 & ~n18280 ;
  assign n18282 = ~\P3_addr_reg[2]/NET0131  & ~n18281 ;
  assign n18283 = \P3_addr_reg[2]/NET0131  & n18281 ;
  assign n18284 = ~n18211 & ~n18212 ;
  assign n18285 = n18186 & ~n18284 ;
  assign n18286 = ~n18186 & n18284 ;
  assign n18287 = ~n18285 & ~n18286 ;
  assign n18288 = \P3_addr_reg[1]/NET0131  & n18287 ;
  assign n18289 = ~n18190 & ~n18288 ;
  assign n18290 = ~\P3_addr_reg[1]/NET0131  & ~n18287 ;
  assign n18291 = ~n18289 & ~n18290 ;
  assign n18292 = ~n18283 & ~n18291 ;
  assign n18293 = ~n18282 & ~n18292 ;
  assign n18294 = ~n18277 & ~n18293 ;
  assign n18295 = ~n18276 & ~n18294 ;
  assign n18296 = ~n18271 & ~n18295 ;
  assign n18297 = ~\P3_addr_reg[4]/NET0131  & ~n18270 ;
  assign n18298 = ~n18296 & ~n18297 ;
  assign n18299 = ~n18266 & ~n18298 ;
  assign n18300 = ~n18265 & ~n18299 ;
  assign n18301 = ~n18260 & ~n18300 ;
  assign n18302 = ~n18259 & ~n18301 ;
  assign n18303 = ~n18254 & ~n18302 ;
  assign n18304 = ~n18253 & ~n18303 ;
  assign n18305 = ~n18248 & ~n18304 ;
  assign n18306 = ~n18247 & ~n18305 ;
  assign n18307 = ~n18242 & ~n18306 ;
  assign n18308 = ~n18241 & ~n18307 ;
  assign n18309 = ~n18236 & n18308 ;
  assign n18310 = n18236 & ~n18308 ;
  assign n18311 = ~n18309 & ~n18310 ;
  assign n18312 = \P1_addr_reg[11]/NET0131  & \P2_addr_reg[11]/NET0131  ;
  assign n18313 = ~\P1_addr_reg[11]/NET0131  & ~\P2_addr_reg[11]/NET0131  ;
  assign n18314 = ~n18312 & ~n18313 ;
  assign n18315 = ~n18192 & ~n18230 ;
  assign n18316 = ~n18193 & ~n18315 ;
  assign n18317 = ~n18314 & n18316 ;
  assign n18318 = n18314 & ~n18316 ;
  assign n18319 = ~n18317 & ~n18318 ;
  assign n18320 = ~\P3_addr_reg[11]/NET0131  & ~n18319 ;
  assign n18321 = \P3_addr_reg[11]/NET0131  & n18319 ;
  assign n18322 = ~n18320 & ~n18321 ;
  assign n18323 = ~n18235 & ~n18308 ;
  assign n18324 = ~n18234 & ~n18323 ;
  assign n18325 = n18322 & n18324 ;
  assign n18326 = ~n18322 & ~n18324 ;
  assign n18327 = ~n18325 & ~n18326 ;
  assign n18328 = \P1_addr_reg[12]/NET0131  & \P2_addr_reg[12]/NET0131  ;
  assign n18329 = ~\P1_addr_reg[12]/NET0131  & ~\P2_addr_reg[12]/NET0131  ;
  assign n18330 = ~n18328 & ~n18329 ;
  assign n18331 = ~n18312 & ~n18316 ;
  assign n18332 = ~n18313 & ~n18331 ;
  assign n18333 = ~n18330 & n18332 ;
  assign n18334 = n18330 & ~n18332 ;
  assign n18335 = ~n18333 & ~n18334 ;
  assign n18336 = ~\P3_addr_reg[12]/NET0131  & ~n18335 ;
  assign n18337 = \P3_addr_reg[12]/NET0131  & n18335 ;
  assign n18338 = ~n18336 & ~n18337 ;
  assign n18339 = ~n18321 & ~n18324 ;
  assign n18340 = ~n18320 & ~n18339 ;
  assign n18341 = n18338 & n18340 ;
  assign n18342 = ~n18338 & ~n18340 ;
  assign n18343 = ~n18341 & ~n18342 ;
  assign n18344 = \P1_addr_reg[13]/NET0131  & \P2_addr_reg[13]/NET0131  ;
  assign n18345 = ~\P1_addr_reg[13]/NET0131  & ~\P2_addr_reg[13]/NET0131  ;
  assign n18346 = ~n18344 & ~n18345 ;
  assign n18347 = ~n18328 & ~n18332 ;
  assign n18348 = ~n18329 & ~n18347 ;
  assign n18349 = ~n18346 & n18348 ;
  assign n18350 = n18346 & ~n18348 ;
  assign n18351 = ~n18349 & ~n18350 ;
  assign n18352 = ~\P3_addr_reg[13]/NET0131  & ~n18351 ;
  assign n18353 = \P3_addr_reg[13]/NET0131  & n18351 ;
  assign n18354 = ~n18352 & ~n18353 ;
  assign n18355 = ~n18337 & ~n18340 ;
  assign n18356 = ~n18336 & ~n18355 ;
  assign n18357 = n18354 & n18356 ;
  assign n18358 = ~n18354 & ~n18356 ;
  assign n18359 = ~n18357 & ~n18358 ;
  assign n18360 = \P1_addr_reg[14]/NET0131  & \P2_addr_reg[14]/NET0131  ;
  assign n18361 = ~\P1_addr_reg[14]/NET0131  & ~\P2_addr_reg[14]/NET0131  ;
  assign n18362 = ~n18360 & ~n18361 ;
  assign n18363 = ~n18344 & ~n18348 ;
  assign n18364 = ~n18345 & ~n18363 ;
  assign n18365 = ~n18362 & n18364 ;
  assign n18366 = n18362 & ~n18364 ;
  assign n18367 = ~n18365 & ~n18366 ;
  assign n18368 = ~\P3_addr_reg[14]/NET0131  & ~n18367 ;
  assign n18369 = \P3_addr_reg[14]/NET0131  & n18367 ;
  assign n18370 = ~n18368 & ~n18369 ;
  assign n18371 = ~n18353 & ~n18356 ;
  assign n18372 = ~n18352 & ~n18371 ;
  assign n18373 = n18370 & n18372 ;
  assign n18374 = ~n18370 & ~n18372 ;
  assign n18375 = ~n18373 & ~n18374 ;
  assign n18376 = \P1_addr_reg[15]/NET0131  & \P2_addr_reg[15]/NET0131  ;
  assign n18377 = ~\P1_addr_reg[15]/NET0131  & ~\P2_addr_reg[15]/NET0131  ;
  assign n18378 = ~n18376 & ~n18377 ;
  assign n18379 = ~n18360 & ~n18364 ;
  assign n18380 = ~n18361 & ~n18379 ;
  assign n18381 = ~n18378 & n18380 ;
  assign n18382 = n18378 & ~n18380 ;
  assign n18383 = ~n18381 & ~n18382 ;
  assign n18384 = ~\P3_addr_reg[15]/NET0131  & ~n18383 ;
  assign n18385 = \P3_addr_reg[15]/NET0131  & n18383 ;
  assign n18386 = ~n18384 & ~n18385 ;
  assign n18387 = ~n18369 & ~n18372 ;
  assign n18388 = ~n18368 & ~n18387 ;
  assign n18389 = n18386 & n18388 ;
  assign n18390 = ~n18386 & ~n18388 ;
  assign n18391 = ~n18389 & ~n18390 ;
  assign n18392 = \P1_addr_reg[16]/NET0131  & \P2_addr_reg[16]/NET0131  ;
  assign n18393 = ~\P1_addr_reg[16]/NET0131  & ~\P2_addr_reg[16]/NET0131  ;
  assign n18394 = ~n18392 & ~n18393 ;
  assign n18395 = ~n18376 & ~n18380 ;
  assign n18396 = ~n18377 & ~n18395 ;
  assign n18397 = n18394 & ~n18396 ;
  assign n18398 = ~n18394 & n18396 ;
  assign n18399 = ~n18397 & ~n18398 ;
  assign n18400 = ~\P3_addr_reg[16]/NET0131  & ~n18399 ;
  assign n18401 = \P3_addr_reg[16]/NET0131  & n18399 ;
  assign n18402 = ~n18400 & ~n18401 ;
  assign n18403 = ~n18385 & ~n18388 ;
  assign n18404 = ~n18384 & ~n18403 ;
  assign n18405 = n18402 & n18404 ;
  assign n18406 = ~n18402 & ~n18404 ;
  assign n18407 = ~n18405 & ~n18406 ;
  assign n18408 = \P1_addr_reg[17]/NET0131  & \P2_addr_reg[17]/NET0131  ;
  assign n18409 = ~\P1_addr_reg[17]/NET0131  & ~\P2_addr_reg[17]/NET0131  ;
  assign n18410 = ~n18408 & ~n18409 ;
  assign n18411 = ~n18393 & n18396 ;
  assign n18412 = ~n18392 & ~n18411 ;
  assign n18413 = ~n18410 & n18412 ;
  assign n18414 = n18410 & ~n18412 ;
  assign n18415 = ~n18413 & ~n18414 ;
  assign n18416 = ~\P3_addr_reg[17]/NET0131  & n18415 ;
  assign n18417 = \P3_addr_reg[17]/NET0131  & ~n18415 ;
  assign n18418 = ~n18416 & ~n18417 ;
  assign n18419 = ~n18401 & ~n18404 ;
  assign n18420 = ~n18400 & ~n18419 ;
  assign n18421 = n18418 & ~n18420 ;
  assign n18422 = ~n18418 & n18420 ;
  assign n18423 = ~n18421 & ~n18422 ;
  assign n18424 = \P1_addr_reg[18]/NET0131  & \P2_addr_reg[18]/NET0131  ;
  assign n18425 = ~\P1_addr_reg[18]/NET0131  & ~\P2_addr_reg[18]/NET0131  ;
  assign n18426 = ~n18424 & ~n18425 ;
  assign n18427 = ~n18392 & ~n18408 ;
  assign n18428 = ~n18411 & n18427 ;
  assign n18429 = ~n18409 & ~n18428 ;
  assign n18430 = n18426 & ~n18429 ;
  assign n18431 = ~n18426 & n18429 ;
  assign n18432 = ~n18430 & ~n18431 ;
  assign n18433 = ~\P3_addr_reg[18]/NET0131  & ~n18432 ;
  assign n18434 = \P3_addr_reg[18]/NET0131  & n18432 ;
  assign n18435 = ~n18433 & ~n18434 ;
  assign n18436 = ~n18416 & n18420 ;
  assign n18437 = ~n18417 & ~n18436 ;
  assign n18438 = n18435 & n18437 ;
  assign n18439 = ~n18435 & ~n18437 ;
  assign n18440 = ~n18438 & ~n18439 ;
  assign n18441 = ~n18417 & ~n18434 ;
  assign n18442 = ~n18436 & n18441 ;
  assign n18443 = ~n18433 & ~n18442 ;
  assign n18444 = ~n768 & ~n771 ;
  assign n18445 = \P3_addr_reg[19]/NET0131  & ~n18444 ;
  assign n18446 = ~\P3_addr_reg[19]/NET0131  & n18444 ;
  assign n18447 = ~n18445 & ~n18446 ;
  assign n18448 = ~n18424 & ~n18429 ;
  assign n18449 = ~n18425 & ~n18448 ;
  assign n18450 = n18447 & ~n18449 ;
  assign n18451 = ~n18447 & n18449 ;
  assign n18452 = ~n18450 & ~n18451 ;
  assign n18453 = n18443 & n18452 ;
  assign n18454 = ~n18443 & ~n18452 ;
  assign n18455 = ~n18453 & ~n18454 ;
  assign n18456 = ~n18288 & ~n18290 ;
  assign n18457 = n18190 & n18456 ;
  assign n18458 = ~n18190 & ~n18456 ;
  assign n18459 = ~n18457 & ~n18458 ;
  assign n18460 = ~n18282 & ~n18283 ;
  assign n18461 = ~n18291 & n18460 ;
  assign n18462 = n18291 & ~n18460 ;
  assign n18463 = ~n18461 & ~n18462 ;
  assign n18464 = ~n18276 & ~n18277 ;
  assign n18465 = ~n18293 & n18464 ;
  assign n18466 = n18293 & ~n18464 ;
  assign n18467 = ~n18465 & ~n18466 ;
  assign n18468 = ~n18271 & ~n18297 ;
  assign n18469 = n18295 & ~n18468 ;
  assign n18470 = ~n18295 & n18468 ;
  assign n18471 = ~n18469 & ~n18470 ;
  assign n18472 = ~n18265 & ~n18266 ;
  assign n18473 = n18298 & n18472 ;
  assign n18474 = ~n18298 & ~n18472 ;
  assign n18475 = ~n18473 & ~n18474 ;
  assign n18476 = ~n18259 & ~n18260 ;
  assign n18477 = n18300 & n18476 ;
  assign n18478 = ~n18300 & ~n18476 ;
  assign n18479 = ~n18477 & ~n18478 ;
  assign n18480 = ~n18253 & ~n18254 ;
  assign n18481 = n18302 & n18480 ;
  assign n18482 = ~n18302 & ~n18480 ;
  assign n18483 = ~n18481 & ~n18482 ;
  assign n18484 = ~n18247 & ~n18248 ;
  assign n18485 = n18304 & n18484 ;
  assign n18486 = ~n18304 & ~n18484 ;
  assign n18487 = ~n18485 & ~n18486 ;
  assign n18488 = ~n18241 & ~n18242 ;
  assign n18489 = n18306 & n18488 ;
  assign n18490 = ~n18306 & ~n18488 ;
  assign n18491 = ~n18489 & ~n18490 ;
  assign n18492 = \P1_wr_reg/NET0131  & ~\P2_wr_reg/NET0131  ;
  assign n18493 = ~\P1_wr_reg/NET0131  & \P2_wr_reg/NET0131  ;
  assign n18494 = ~n18492 & ~n18493 ;
  assign n18495 = ~\P3_wr_reg/NET0131  & ~n18494 ;
  assign \P1_state_reg[0]/NET0131_syn_2  = ~\P1_state_reg[0]/NET0131  ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g106254/_0_  = ~n2142 ;
  assign \g106255/_0_  = ~n2405 ;
  assign \g106267/_0_  = ~n2529 ;
  assign \g106268/_0_  = ~n2635 ;
  assign \g106269/_0_  = ~n2664 ;
  assign \g106270/_0_  = ~n4133 ;
  assign \g106271/_0_  = ~n4162 ;
  assign \g106272/_0_  = ~n5591 ;
  assign \g106288/_0_  = ~n5649 ;
  assign \g106289/_0_  = ~n5694 ;
  assign \g106290/_0_  = ~n5785 ;
  assign \g106291/_0_  = ~n6077 ;
  assign \g106292/_0_  = ~n6377 ;
  assign \g106293/_0_  = ~n6406 ;
  assign \g106294/_0_  = ~n6437 ;
  assign \g106295/_0_  = ~n6467 ;
  assign \g106296/_0_  = ~n6496 ;
  assign \g106297/_0_  = ~n6523 ;
  assign \g106352/_0_  = ~n6566 ;
  assign \g106356/_0_  = ~n6680 ;
  assign \g106359/_0_  = ~n6704 ;
  assign \g106360/_0_  = ~n6727 ;
  assign \g106361/_0_  = ~n6850 ;
  assign \g106362/_0_  = ~n6875 ;
  assign \g106363/_0_  = ~n6900 ;
  assign \g106364/_0_  = ~n6925 ;
  assign \g106365/_0_  = ~n6950 ;
  assign \g106406/_0_  = ~n7062 ;
  assign \g106407/_0_  = ~n7123 ;
  assign \g106408/_0_  = ~n7219 ;
  assign \g106410/_0_  = ~n7248 ;
  assign \g106411/_0_  = ~n7289 ;
  assign \g106412/_0_  = ~n7329 ;
  assign \g106413/_0_  = ~n7377 ;
  assign \g106414/_0_  = ~n7420 ;
  assign \g106417/_0_  = ~n7449 ;
  assign \g106418/_0_  = ~n7515 ;
  assign \g106419/_0_  = ~n7624 ;
  assign \g106420/_0_  = ~n7654 ;
  assign \g106421/_0_  = ~n7712 ;
  assign \g106422/_0_  = ~n7741 ;
  assign \g106423/_0_  = ~n7770 ;
  assign \g106424/_0_  = ~n7793 ;
  assign \g106425/_0_  = ~n7818 ;
  assign \g106426/_0_  = ~n7875 ;
  assign \g106427/_0_  = ~n7970 ;
  assign \g106428/_0_  = ~n7994 ;
  assign \g106430/_0_  = ~n8016 ;
  assign \g106431/_0_  = ~n8035 ;
  assign \g106432/_0_  = ~n8053 ;
  assign \g106433/_0_  = ~n8075 ;
  assign \g106434/_0_  = ~n8103 ;
  assign \g106436/_0_  = ~n8124 ;
  assign \g106437/_0_  = ~n8144 ;
  assign \g106438/_0_  = ~n8166 ;
  assign \g106439/_0_  = ~n8191 ;
  assign \g106440/_0_  = ~n8216 ;
  assign \g106441/_0_  = ~n8234 ;
  assign \g106442/_0_  = ~n8259 ;
  assign \g106443/_0_  = ~n8284 ;
  assign \g106444/_0_  = ~n8309 ;
  assign \g106445/_0_  = ~n8334 ;
  assign \g106446/_0_  = ~n8363 ;
  assign \g106447/_0_  = ~n8392 ;
  assign \g106448/_0_  = ~n8421 ;
  assign \g106530/_0_  = ~n8464 ;
  assign \g106531/_0_  = ~n8510 ;
  assign \g106532/_0_  = ~n8552 ;
  assign \g106533/_0_  = ~n8592 ;
  assign \g106534/_0_  = ~n8632 ;
  assign \g106554/_0_  = ~n8654 ;
  assign \g106556/_0_  = ~n8705 ;
  assign \g106557/_0_  = ~n8731 ;
  assign \g106559/_0_  = ~n8784 ;
  assign \g106560/_0_  = ~n8810 ;
  assign \g106561/_0_  = ~n8840 ;
  assign \g106562/_0_  = ~n8858 ;
  assign \g106563/_0_  = ~n8881 ;
  assign \g106564/_0_  = ~n8897 ;
  assign \g106565/_0_  = ~n8915 ;
  assign \g106566/_0_  = ~n8927 ;
  assign \g106567/_0_  = ~n8949 ;
  assign \g106568/_0_  = ~n8973 ;
  assign \g106569/_0_  = ~n9001 ;
  assign \g106570/_0_  = ~n9025 ;
  assign \g106571/_0_  = ~n9043 ;
  assign \g106572/_0_  = ~n9055 ;
  assign \g106633/_0_  = ~n9095 ;
  assign \g106634/_0_  = ~n9141 ;
  assign \g106640/_0_  = ~n9186 ;
  assign \g106654/_0_  = ~n9227 ;
  assign \g106655/_0_  = ~n9259 ;
  assign \g106679/_0_  = ~n9301 ;
  assign \g106682/_0_  = ~n9343 ;
  assign \g106684/_0_  = ~n9372 ;
  assign \g106687/_0_  = ~n9411 ;
  assign \g106690/_0_  = ~n9457 ;
  assign \g106691/_0_  = ~n9480 ;
  assign \g106692/_0_  = ~n9505 ;
  assign \g106693/_0_  = ~n9527 ;
  assign \g106694/_0_  = ~n9535 ;
  assign \g106695/_0_  = ~n9557 ;
  assign \g106696/_0_  = ~n9577 ;
  assign \g106697/_0_  = ~n9595 ;
  assign \g106698/_0_  = ~n9617 ;
  assign \g106699/_0_  = ~n9635 ;
  assign \g106700/_0_  = ~n9642 ;
  assign \g106701/_0_  = ~n9649 ;
  assign \g106702/_0_  = ~n9666 ;
  assign \g106703/_0_  = ~n9690 ;
  assign \g106704/_0_  = ~n9714 ;
  assign \g106705/_0_  = ~n9742 ;
  assign \g106706/_0_  = ~n9769 ;
  assign \g106707/_0_  = ~n9779 ;
  assign \g106708/_0_  = ~n9797 ;
  assign \g106710/_0_  = ~n9823 ;
  assign \g106711/_0_  = ~n9831 ;
  assign \g106712/_0_  = ~n9856 ;
  assign \g106713/_0_  = ~n9882 ;
  assign \g106714/_0_  = ~n9907 ;
  assign \g106715/_0_  = ~n9932 ;
  assign \g106716/_0_  = ~n9957 ;
  assign \g106717/_0_  = ~n9982 ;
  assign \g106718/_0_  = ~n10007 ;
  assign \g106719/_0_  = ~n10024 ;
  assign \g106720/_0_  = ~n10051 ;
  assign \g106721/_0_  = ~n10076 ;
  assign \g106722/_0_  = ~n10103 ;
  assign \g106723/_0_  = ~n10128 ;
  assign \g106724/_0_  = ~n10153 ;
  assign \g106725/_0_  = ~n10178 ;
  assign \g106726/_0_  = ~n10203 ;
  assign \g106727/_0_  = ~n10230 ;
  assign \g106728/_0_  = ~n10257 ;
  assign \g106729/_0_  = ~n10283 ;
  assign \g106830/_0_  = ~n10324 ;
  assign \g106836/_0_  = ~n10367 ;
  assign \g106837/_0_  = ~n10411 ;
  assign \g106838/_0_  = ~n10448 ;
  assign \g106843/_0_  = ~n10486 ;
  assign \g106850/_0_  = ~n10527 ;
  assign \g106851/_0_  = ~n10567 ;
  assign \g106852/_0_  = ~n10607 ;
  assign \g106853/_0_  = ~n10648 ;
  assign \g106854/_0_  = ~n10688 ;
  assign \g106899/_0_  = ~n10728 ;
  assign \g106901/_0_  = ~n10776 ;
  assign \g106902/_0_  = ~n10798 ;
  assign \g106903/_0_  = ~n10801 ;
  assign \g106904/_0_  = ~n10820 ;
  assign \g106905/_0_  = ~n10844 ;
  assign \g106906/_0_  = ~n10873 ;
  assign \g106907/_0_  = ~n10902 ;
  assign \g106908/_0_  = ~n10931 ;
  assign \g106909/_0_  = ~n10953 ;
  assign \g106910/_0_  = ~n10966 ;
  assign \g106911/_0_  = ~n11012 ;
  assign \g106912/_0_  = ~n11031 ;
  assign \g106913/_0_  = ~n11053 ;
  assign \g106914/_0_  = ~n11063 ;
  assign \g106915/_0_  = ~n11089 ;
  assign \g106916/_0_  = ~n11115 ;
  assign \g106917/_0_  = ~n11126 ;
  assign \g106918/_0_  = ~n11151 ;
  assign \g106919/_0_  = ~n11177 ;
  assign \g106920/_0_  = ~n11194 ;
  assign \g106921/_0_  = ~n11205 ;
  assign \g106922/_0_  = ~n11231 ;
  assign \g106923/_0_  = ~n11257 ;
  assign \g106924/_0_  = ~n11262 ;
  assign \g106925/_0_  = ~n11284 ;
  assign \g106994/_0_  = ~n11324 ;
  assign \g106995/_0_  = ~n11365 ;
  assign \g106996/_0_  = ~n11404 ;
  assign \g106997/_0_  = ~n11445 ;
  assign \g106998/_0_  = ~n11488 ;
  assign \g106999/_0_  = ~n11531 ;
  assign \g107002/_0_  = ~n11572 ;
  assign \g107007/_0_  = ~n11612 ;
  assign \g107008/_0_  = ~n11652 ;
  assign \g107038/_0_  = ~n11691 ;
  assign \g107041/_0_  = ~n11724 ;
  assign \g107048/_0_  = ~n11767 ;
  assign \g107091/_0_  = ~n11787 ;
  assign \g107093/_0_  = ~n11816 ;
  assign \g107094/_0_  = ~n11844 ;
  assign \g107096/_0_  = ~n11849 ;
  assign \g107097/_0_  = ~n11867 ;
  assign \g107098/_0_  = ~n11882 ;
  assign \g107099/_0_  = ~n11904 ;
  assign \g107100/_0_  = ~n11913 ;
  assign \g107101/_0_  = ~n11920 ;
  assign \g107102/_0_  = ~n11925 ;
  assign \g107103/_0_  = ~n11943 ;
  assign \g107104/_0_  = ~n11955 ;
  assign \g107105/_0_  = ~n11958 ;
  assign \g107106/_0_  = ~n11964 ;
  assign \g107107/_0_  = ~n11991 ;
  assign \g107108/_0_  = ~n11997 ;
  assign \g107109/_0_  = ~n12015 ;
  assign \g107110/_0_  = ~n12021 ;
  assign \g107111/_0_  = ~n12047 ;
  assign \g107112/_0_  = ~n12052 ;
  assign \g107113/_0_  = ~n12056 ;
  assign \g107114/_0_  = ~n12082 ;
  assign \g107115/_0_  = ~n12107 ;
  assign \g107116/_0_  = ~n12132 ;
  assign \g107117/_0_  = ~n12158 ;
  assign \g107118/_0_  = ~n12184 ;
  assign \g107119/_0_  = ~n12209 ;
  assign \g107120/_0_  = ~n12234 ;
  assign \g107121/_0_  = ~n12261 ;
  assign \g107122/_0_  = ~n12288 ;
  assign \g107123/_0_  = ~n12315 ;
  assign \g107124/_0_  = ~n12342 ;
  assign \g107125/_0_  = ~n12369 ;
  assign \g107126/_0_  = ~n12396 ;
  assign \g107127/_0_  = ~n12423 ;
  assign \g107128/_0_  = ~n12450 ;
  assign \g107129/_0_  = ~n12477 ;
  assign \g107130/_0_  = ~n12504 ;
  assign \g107131/_0_  = ~n12531 ;
  assign \g107132/_0_  = ~n12558 ;
  assign \g107133/_0_  = ~n12585 ;
  assign \g107134/_0_  = ~n12610 ;
  assign \g107135/_0_  = ~n12615 ;
  assign \g107136/_0_  = ~n12618 ;
  assign \g107137/_0_  = ~n12645 ;
  assign \g107138/_0_  = ~n12651 ;
  assign \g107248/_0_  = ~n12687 ;
  assign \g107252/_0_  = ~n12723 ;
  assign \g107254/_0_  = ~n12768 ;
  assign \g107255/_0_  = ~n12810 ;
  assign \g107280/_0_  = ~n12852 ;
  assign \g107281/_0_  = ~n12893 ;
  assign \g107282/_0_  = ~n12933 ;
  assign \g107370/_0_  = ~n12953 ;
  assign \g107371/_0_  = ~n12964 ;
  assign \g107372/_0_  = ~n12970 ;
  assign \g107373/_0_  = ~n12992 ;
  assign \g107374/_0_  = ~n13014 ;
  assign \g107375/_0_  = ~n13043 ;
  assign \g107376/_0_  = ~n13066 ;
  assign \g107377/_0_  = ~n13093 ;
  assign \g107378/_0_  = ~n13105 ;
  assign \g107379/_0_  = ~n13133 ;
  assign \g107380/_0_  = ~n13154 ;
  assign \g107381/_0_  = ~n13176 ;
  assign \g107382/_0_  = ~n13182 ;
  assign \g107383/_0_  = ~n13207 ;
  assign \g107384/_0_  = ~n13234 ;
  assign \g107385/_0_  = ~n13256 ;
  assign \g107386/_0_  = ~n13283 ;
  assign \g107387/_0_  = ~n13309 ;
  assign \g107388/_0_  = ~n13313 ;
  assign \g107389/_0_  = ~n13335 ;
  assign \g107390/_0_  = ~n13361 ;
  assign \g107391/_0_  = ~n13379 ;
  assign \g107488/_0_  = ~n13419 ;
  assign \g107489/_0_  = ~n13456 ;
  assign \g107490/_0_  = ~n13492 ;
  assign \g107491/_0_  = ~n13534 ;
  assign \g107492/_0_  = ~n13577 ;
  assign \g107493/_0_  = ~n13619 ;
  assign \g107500/_0_  = ~n13659 ;
  assign \g107615/_0_  = ~n13683 ;
  assign \g107623/_0_  = ~n13705 ;
  assign \g107624/_0_  = ~n13727 ;
  assign \g107625/_0_  = ~n13734 ;
  assign \g107626/_0_  = ~n13744 ;
  assign \g107627/_0_  = ~n13766 ;
  assign \g107628/_0_  = ~n13769 ;
  assign \g107629/_0_  = ~n13777 ;
  assign \g107630/_0_  = ~n13801 ;
  assign \g107631/_0_  = n13812 ;
  assign \g107632/_0_  = ~n13815 ;
  assign \g107634/_0_  = ~n13818 ;
  assign \g107637/_0_  = ~n13840 ;
  assign \g107638/_0_  = ~n13862 ;
  assign \g107639/_0_  = ~n13888 ;
  assign \g107640/_0_  = ~n13910 ;
  assign \g107641/_0_  = ~n13932 ;
  assign \g107642/_0_  = ~n13960 ;
  assign \g107643/_0_  = ~n13987 ;
  assign \g107644/_0_  = ~n14014 ;
  assign \g107645/_0_  = ~n14041 ;
  assign \g107646/_0_  = ~n14068 ;
  assign \g107647/_0_  = ~n14071 ;
  assign \g107650/_0_  = ~n14098 ;
  assign \g107651/_0_  = ~n14125 ;
  assign \g107652/_0_  = ~n14128 ;
  assign \g107653/_0_  = ~n14155 ;
  assign \g107654/_0_  = ~n14182 ;
  assign \g107655/_0_  = ~n14204 ;
  assign \g107656/_0_  = ~n14207 ;
  assign \g107743/_0_  = ~n14246 ;
  assign \g107787/_0_  = ~n14288 ;
  assign \g107954/_0_  = ~n14310 ;
  assign \g107955/_0_  = ~n14332 ;
  assign \g107956/_0_  = ~n14337 ;
  assign \g107957/_0_  = ~n14344 ;
  assign \g107958/_0_  = ~n14353 ;
  assign \g107959/_0_  = ~n14361 ;
  assign \g107960/_0_  = ~n14385 ;
  assign \g107961/_0_  = ~n14409 ;
  assign \g107962/_0_  = ~n14433 ;
  assign \g107963/_0_  = ~n14459 ;
  assign \g107964/_0_  = n14473 ;
  assign \g107965/_0_  = ~n14479 ;
  assign \g107966/_0_  = ~n14501 ;
  assign \g107967/_0_  = ~n14529 ;
  assign \g108118/_0_  = ~n14569 ;
  assign \g108125/_0_  = ~n14609 ;
  assign \g108169/_0_  = ~n14647 ;
  assign \g108269/_0_  = ~n14671 ;
  assign \g108270/_0_  = ~n14693 ;
  assign \g108319/_0_  = ~n14715 ;
  assign \g108320/_0_  = ~n14722 ;
  assign \g108321/_0_  = ~n14744 ;
  assign \g108322/_0_  = ~n14747 ;
  assign \g108323/_0_  = ~n14769 ;
  assign \g108324/_0_  = ~n14775 ;
  assign \g108326/_0_  = ~n14801 ;
  assign \g108327/_0_  = ~n14821 ;
  assign \g108328/_0_  = ~n14849 ;
  assign \g108329/_0_  = ~n14876 ;
  assign \g108330/_0_  = ~n14903 ;
  assign \g108334/_0_  = ~n14930 ;
  assign \g108335/_0_  = ~n14957 ;
  assign \g108468/_0_  = ~n14984 ;
  assign \g108538/_0_  = ~n15021 ;
  assign \g108801/_0_  = ~n15045 ;
  assign \g108812/_0_  = ~n15059 ;
  assign \g108813/_0_  = ~n15075 ;
  assign \g108814/_0_  = ~n15081 ;
  assign \g108815/_0_  = ~n15105 ;
  assign \g108817/_0_  = ~n15116 ;
  assign \g108818/_0_  = ~n15142 ;
  assign \g108819/_0_  = ~n15169 ;
  assign \g108822/_0_  = ~n15196 ;
  assign \g109052/_0_  = ~n15225 ;
  assign \g109053/_0_  = ~n15265 ;
  assign \g109401/_0_  = ~n15268 ;
  assign \g109402/_0_  = ~n15272 ;
  assign \g109403/_0_  = ~n15283 ;
  assign \g109410/_0_  = ~n15297 ;
  assign \g109411/_0_  = ~n15323 ;
  assign \g109415/_0_  = ~n15348 ;
  assign \g109420/_0_  = ~n15376 ;
  assign \g109425/_0_  = ~n15384 ;
  assign \g109693/_0_  = ~n15415 ;
  assign \g110116/_0_  = ~n15439 ;
  assign \g110117/_0_  = ~n15448 ;
  assign \g110905/_0_  = ~n15471 ;
  assign \g110906/_0_  = ~n15496 ;
  assign \g110907/_0_  = ~n15521 ;
  assign \g111086/_0_  = ~n15539 ;
  assign \g111094/_0_  = ~n15565 ;
  assign \g112422/_0_  = ~n15578 ;
  assign \g112423/_0_  = ~n15586 ;
  assign \g112424/_0_  = ~n15604 ;
  assign \g112425/_0_  = ~n15610 ;
  assign \g112426/_0_  = ~n15628 ;
  assign \g112427/_0_  = ~n15631 ;
  assign \g113647/_0_  = ~n15647 ;
  assign \g113648/_0_  = ~n15654 ;
  assign \g113649/_0_  = ~n15665 ;
  assign \g113650/_0_  = ~n15670 ;
  assign \g113651/_0_  = ~n15687 ;
  assign \g114133/_0_  = ~n15699 ;
  assign \g117884/_0_  = ~n15702 ;
  assign \g117885/_0_  = ~n15705 ;
  assign \g117886/_0_  = ~n15708 ;
  assign \g117895/_3_  = ~n15711 ;
  assign \g117896/_3_  = ~n15714 ;
  assign \g117897/_0_  = ~n15717 ;
  assign \g117898/_0_  = n15720 ;
  assign \g117899/_0_  = ~n15723 ;
  assign \g117900/_3_  = ~n15726 ;
  assign \g120982/_0_  = ~n15729 ;
  assign \g120983/_0_  = n15732 ;
  assign \g120984/_0_  = n15735 ;
  assign \g120985/_0_  = ~n15738 ;
  assign \g120986/_0_  = n15741 ;
  assign \g120987/_0_  = n15744 ;
  assign \g120988/_3_  = n15747 ;
  assign \g120989/_0_  = ~n15750 ;
  assign \g120990/_0_  = n15753 ;
  assign \g120991/_0_  = ~n15756 ;
  assign \g120992/_0_  = n15759 ;
  assign \g120993/_0_  = ~n15762 ;
  assign \g120994/_0_  = n15765 ;
  assign \g120995/_0_  = n15768 ;
  assign \g120996/_3_  = n15771 ;
  assign \g120997/_0_  = n15774 ;
  assign \g120998/_0_  = n15777 ;
  assign \g120999/_0_  = n15779 ;
  assign \g121000/_0_  = ~n15782 ;
  assign \g121001/_0_  = ~n15785 ;
  assign \g121002/_3_  = ~n15788 ;
  assign \g121003/_0_  = ~n15791 ;
  assign \g121004/_0_  = ~n15794 ;
  assign \g121005/_3_  = ~n15797 ;
  assign \g121006/_0_  = ~n15800 ;
  assign \g121007/_0_  = ~n15803 ;
  assign \g121008/_0_  = ~n15806 ;
  assign \g121029/_0_  = ~n15813 ;
  assign \g121030/_3_  = ~n15815 ;
  assign \g121032/_3_  = ~n15818 ;
  assign \g121033/_3_  = ~n15821 ;
  assign \g121034/_3_  = n15824 ;
  assign \g121035/_3_  = ~n15827 ;
  assign \g121036/_3_  = ~n15830 ;
  assign \g121037/_3_  = ~n15833 ;
  assign \g121038/_3_  = ~n15836 ;
  assign \g121039/_3_  = ~n15839 ;
  assign \g121040/_3_  = ~n15842 ;
  assign \g121041/_3_  = ~n15845 ;
  assign \g121042/_3_  = ~n15848 ;
  assign \g121043/_3_  = ~n15851 ;
  assign \g121044/_3_  = ~n15854 ;
  assign \g121045/_3_  = ~n15857 ;
  assign \g121046/_3_  = ~n15860 ;
  assign \g121047/_3_  = ~n15863 ;
  assign \g121048/_3_  = n15866 ;
  assign \g121049/_3_  = ~n15869 ;
  assign \g121050/_3_  = n15872 ;
  assign \g121051/_0_  = ~n15879 ;
  assign \g121052/_3_  = ~n15882 ;
  assign \g121053/_3_  = ~n15885 ;
  assign \g121054/_3_  = ~n15888 ;
  assign \g121055/_3_  = ~n15891 ;
  assign \g121056/_3_  = ~n15894 ;
  assign \g121057/_3_  = ~n15897 ;
  assign \g121058/_3_  = ~n15900 ;
  assign \g121060/_3_  = n15903 ;
  assign \g121061/_3_  = ~n15906 ;
  assign \g121062/_3_  = n15909 ;
  assign \g121063/_3_  = n15912 ;
  assign \g121064/_3_  = ~n15915 ;
  assign \g121065/_3_  = n15918 ;
  assign \g121066/_3_  = n15921 ;
  assign \g121067/_3_  = ~n15924 ;
  assign \g121068/_3_  = n15927 ;
  assign \g121069/_3_  = ~n15930 ;
  assign \g121070/_3_  = ~n15933 ;
  assign \g121071/_3_  = ~n15936 ;
  assign \g121072/_3_  = ~n15939 ;
  assign \g121073/_3_  = n15941 ;
  assign \g121074/_3_  = n15944 ;
  assign \g121075/_3_  = n15947 ;
  assign \g121076/_3_  = ~n15950 ;
  assign \g121077/_3_  = ~n15953 ;
  assign \g121078/_3_  = ~n15956 ;
  assign \g121079/_3_  = ~n15959 ;
  assign \g121080/_0_  = ~n15967 ;
  assign \g121081/_3_  = ~n15970 ;
  assign \g121082/_0_  = n15973 ;
  assign \g121083/_3_  = ~n15976 ;
  assign \g121084/_3_  = n15979 ;
  assign \g121085/_3_  = ~n15982 ;
  assign \g121086/_3_  = n15985 ;
  assign \g121087/_3_  = ~n15988 ;
  assign \g121626/_0_  = n3691 ;
  assign \g121633/_0_  = ~n1904 ;
  assign \g121669/_0_  = n5187 ;
  assign \g122948/_0_  = ~n16135 ;
  assign \g122949/_0_  = ~n16165 ;
  assign \g122951/_0_  = ~n16194 ;
  assign \g122952/_0_  = ~n16213 ;
  assign \g122953/_0_  = ~n16241 ;
  assign \g122954/_0_  = ~n16269 ;
  assign \g122955/_0_  = ~n16297 ;
  assign \g122956/_0_  = ~n16324 ;
  assign \g122957/_0_  = ~n16374 ;
  assign \g122958/_0_  = ~n16392 ;
  assign \g122959/_0_  = ~n16411 ;
  assign \g122960/_0_  = ~n16430 ;
  assign \g122963/_0_  = ~n16512 ;
  assign \g122965/_0_  = ~n16533 ;
  assign \g122967/_0_  = ~n16554 ;
  assign \g122968/_0_  = ~n16571 ;
  assign \g122972/_0_  = ~n16588 ;
  assign \g122973/_0_  = ~n16606 ;
  assign \g122974/_0_  = ~n16634 ;
  assign \g122975/_0_  = ~n16652 ;
  assign \g122976/_0_  = ~n16670 ;
  assign \g122977/_0_  = ~n16688 ;
  assign \g122978/_0_  = ~n16706 ;
  assign \g122979/_0_  = ~n16732 ;
  assign \g122980/_0_  = ~n16778 ;
  assign \g122981/_0_  = ~n16796 ;
  assign \g122982/_0_  = ~n16817 ;
  assign \g122983/_0_  = ~n16843 ;
  assign \g122984/_0_  = ~n16861 ;
  assign \g122985/_0_  = ~n16879 ;
  assign \g122986/_0_  = ~n16897 ;
  assign \g122987/_0_  = ~n16923 ;
  assign \g122988/_0_  = ~n16941 ;
  assign \g122989/_0_  = ~n16959 ;
  assign \g122990/_0_  = ~n16979 ;
  assign \g122991/_0_  = ~n16997 ;
  assign \g122997/_0_  = ~n17030 ;
  assign \g122998/_0_  = ~n17055 ;
  assign \g122999/_0_  = ~n17085 ;
  assign \g123000/_0_  = ~n17115 ;
  assign \g123740/_0_  = ~n17117 ;
  assign \g123811/_0_  = ~n17289 ;
  assign \g123812/_0_  = n17309 ;
  assign \g123813/_0_  = ~n17340 ;
  assign \g123814/_0_  = ~n17381 ;
  assign \g123815/_0_  = ~n17430 ;
  assign \g123816/_0_  = ~n17485 ;
  assign \g123817/_0_  = ~n17552 ;
  assign \g123818/_0_  = ~n17607 ;
  assign \g123819/_0_  = ~n17638 ;
  assign \g123820/_0_  = ~n17669 ;
  assign \g123821/_0_  = ~n17700 ;
  assign \g123822/_0_  = ~n17765 ;
  assign \g123823/_0_  = ~n17796 ;
  assign \g123824/_0_  = ~n17832 ;
  assign \g123825/_0_  = ~n17863 ;
  assign \g123826/_0_  = ~n17894 ;
  assign \g123827/_0_  = n17926 ;
  assign \g123828/_0_  = ~n17957 ;
  assign \g123829/_0_  = ~n17988 ;
  assign \g123830/_0_  = n18020 ;
  assign \g123853/u3_syn_4  = n8899 ;
  assign \g123854/u3_syn_4  = n15640 ;
  assign \g123871/_0_  = ~n18022 ;
  assign \g124519/_0_  = ~n18024 ;
  assign \g124554/_0_  = ~n6107 ;
  assign \g124798/_0_  = ~n2157 ;
  assign \g124897/_0_  = ~n6112 ;
  assign \g125133/_0_  = n4218 ;
  assign \g125231/_0_  = ~n2162 ;
  assign \g125318/u3_syn_4  = n18025 ;
  assign \g125495/u3_syn_4  = n18026 ;
  assign \g126480/_0_  = ~n3473 ;
  assign \g126501/_0_  = ~n3410 ;
  assign \g127137/_0_  = ~n3795 ;
  assign \g127147/_0_  = ~n3650 ;
  assign \g127163/_0_  = ~n3229 ;
  assign \g127173/_0_  = ~n3255 ;
  assign \g127202/_0_  = ~n2887 ;
  assign \g127211/_0_  = ~n3329 ;
  assign \g127223/_0_  = ~n3746 ;
  assign \g127234/_0_  = ~n3137 ;
  assign \g127241/_0_  = ~n3756 ;
  assign \g127251/_0_  = ~n3364 ;
  assign \g127257/_0_  = ~n3687 ;
  assign \g127262/_0_  = ~n3704 ;
  assign \g127271/_0_  = ~n3203 ;
  assign \g127285/_0_  = ~n2952 ;
  assign \g127292/_0_  = ~n3109 ;
  assign \g127302/_0_  = ~n3623 ;
  assign \g127313/_0_  = ~n3677 ;
  assign \g127324/_0_  = ~n3597 ;
  assign \g127334/_0_  = ~n3527 ;
  assign \g127348/_0_  = ~n3437 ;
  assign \g127366/_0_  = ~n3577 ;
  assign \g127396/_0_  = ~n3176 ;
  assign \g127405/_0_  = ~n5345 ;
  assign \g127411/_0_  = ~n4421 ;
  assign \g127427/_0_  = ~n3034 ;
  assign \g127439/_0_  = ~n3283 ;
  assign \g127464/_0_  = ~n5339 ;
  assign \g127893/_0_  = n18027 ;
  assign \g128290/_0_  = ~n5117 ;
  assign \g128431/_0_  = ~n5092 ;
  assign \g128477/_0_  = ~n4958 ;
  assign \g128501/_0_  = ~n5008 ;
  assign \g128540/_0_  = ~n5161 ;
  assign \g128566/_0_  = ~n4799 ;
  assign \g128575/_0_  = ~n4728 ;
  assign \g128586/_0_  = ~n4774 ;
  assign \g128594/_1_  = ~n4500 ;
  assign \g128631/_0_  = ~n4552 ;
  assign \g128648/_0_  = ~n4622 ;
  assign \g128698/_0_  = ~n5184 ;
  assign \g131281/_1_  = n6078 ;
  assign \g140384/_0_  = ~n3303 ;
  assign \g140411/_0_  = ~n3081 ;
  assign \g140627/_0_  = ~n18044 ;
  assign \g140741/_0_  = ~n18056 ;
  assign \g140774/_0_  = ~n3548 ;
  assign \g140804/_0_  = ~n3822 ;
  assign \g140955/_0_  = ~n4984 ;
  assign \g140986/_0_  = ~n5068 ;
  assign \g141163/_0_  = ~n3354 ;
  assign \g141237/_0_  = ~n4647 ;
  assign \g141301/_0_  = ~n18083 ;
  assign \g141328/_0_  = ~n4211 ;
  assign \g141367/_0_  = ~n18109 ;
  assign \g141441/_0_  = ~n4703 ;
  assign \g141474/_0_  = ~n18120 ;
  assign \g141548/_0_  = ~n18131 ;
  assign \g141640/_0_  = ~n4684 ;
  assign \g141838/_0_  = ~n5203 ;
  assign \g141844/_0_  = ~n5226 ;
  assign \g141853/_0_  = ~n4879 ;
  assign \g141855/_0_  = ~n4902 ;
  assign \g141860/_0_  = ~n4827 ;
  assign \g141896/_0_  = ~n5040 ;
  assign \g141915/_0_  = ~n4931 ;
  assign \g141952/_0_  = ~n4601 ;
  assign \g142033/_0_  = ~n4665 ;
  assign \g142046/_0_  = ~n5139 ;
  assign \g29/_0_  = ~n18156 ;
  assign \g33/_0_  = ~n18181 ;
  assign \g53/_0_  = ~n3506 ;
  assign \g71/_0_  = ~n4763 ;
  assign \g90/_0_  = ~n4854 ;
  assign rd_pad = ~n18185 ;
  assign \so[0]_pad  = ~n18191 ;
  assign \so[10]_pad  = n18311 ;
  assign \so[11]_pad  = ~n18327 ;
  assign \so[12]_pad  = ~n18343 ;
  assign \so[13]_pad  = ~n18359 ;
  assign \so[14]_pad  = ~n18375 ;
  assign \so[15]_pad  = ~n18391 ;
  assign \so[16]_pad  = ~n18407 ;
  assign \so[17]_pad  = n18423 ;
  assign \so[18]_pad  = n18440 ;
  assign \so[19]_pad  = n18455 ;
  assign \so[1]_pad  = ~n18459 ;
  assign \so[2]_pad  = n18463 ;
  assign \so[3]_pad  = n18467 ;
  assign \so[4]_pad  = n18471 ;
  assign \so[5]_pad  = ~n18475 ;
  assign \so[6]_pad  = ~n18479 ;
  assign \so[7]_pad  = ~n18483 ;
  assign \so[8]_pad  = ~n18487 ;
  assign \so[9]_pad  = ~n18491 ;
  assign wr_pad = ~n18495 ;
endmodule
