module top (CLR_pad, \v0_pad , \v10_reg/NET0131 , \v11_reg/NET0131 , \v12_reg/NET0131 , \v1_pad , \v2_pad , \v3_pad , \v4_pad , \v5_pad , \v6_pad , \v7_reg/NET0131 , \v8_reg/NET0131 , \v9_reg/NET0131 , \_al_n0 , \_al_n1 , \g1757/_0_ , \g1763/_1_ , \g1787/_3_ , \g1800/_3_ , \g1821/_2_ , \g1940/_1_ , \g25/_0_ , \g2783/_3_ , \g2823/_0_ , \g38/_1_ , \g40/_1_ , \v13_D_11_pad , \v13_D_12_pad , \v13_D_13_pad , \v13_D_14_pad , \v13_D_16_pad , \v13_D_18_pad , \v13_D_19_pad , \v13_D_21_pad , \v13_D_22_pad , \v13_D_23_pad , \v13_D_24_pad , \v13_D_7_pad , \v13_D_8_pad , \v13_D_9_pad );
	input CLR_pad ;
	input \v0_pad  ;
	input \v10_reg/NET0131  ;
	input \v11_reg/NET0131  ;
	input \v12_reg/NET0131  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input \v4_pad  ;
	input \v5_pad  ;
	input \v6_pad  ;
	input \v7_reg/NET0131  ;
	input \v8_reg/NET0131  ;
	input \v9_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1757/_0_  ;
	output \g1763/_1_  ;
	output \g1787/_3_  ;
	output \g1800/_3_  ;
	output \g1821/_2_  ;
	output \g1940/_1_  ;
	output \g25/_0_  ;
	output \g2783/_3_  ;
	output \g2823/_0_  ;
	output \g38/_1_  ;
	output \g40/_1_  ;
	output \v13_D_11_pad  ;
	output \v13_D_12_pad  ;
	output \v13_D_13_pad  ;
	output \v13_D_14_pad  ;
	output \v13_D_16_pad  ;
	output \v13_D_18_pad  ;
	output \v13_D_19_pad  ;
	output \v13_D_21_pad  ;
	output \v13_D_22_pad  ;
	output \v13_D_23_pad  ;
	output \v13_D_24_pad  ;
	output \v13_D_7_pad  ;
	output \v13_D_8_pad  ;
	output \v13_D_9_pad  ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w16_ ;
	wire _w17_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	LUT4 #(
		.INIT('h9998)
	) name0 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v3_pad ,
		\v6_pad ,
		_w16_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\v12_reg/NET0131 ,
		_w16_,
		_w17_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w18_
	);
	LUT3 #(
		.INIT('hbc)
	) name3 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w19_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\v4_pad ,
		\v5_pad ,
		_w20_
	);
	LUT3 #(
		.INIT('h40)
	) name5 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w21_
	);
	LUT3 #(
		.INIT('h45)
	) name6 (
		_w18_,
		_w19_,
		_w21_,
		_w22_
	);
	LUT3 #(
		.INIT('h45)
	) name7 (
		\v8_reg/NET0131 ,
		_w17_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\v10_reg/NET0131 ,
		\v1_pad ,
		_w24_
	);
	LUT4 #(
		.INIT('h0040)
	) name9 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w25_
	);
	LUT4 #(
		.INIT('h0008)
	) name10 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v8_reg/NET0131 ,
		_w26_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w27_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12 (
		\v2_pad ,
		_w26_,
		_w27_,
		_w25_,
		_w28_
	);
	LUT3 #(
		.INIT('h80)
	) name13 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w29_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w31_
	);
	LUT4 #(
		.INIT('h0010)
	) name16 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w32_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w29_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		_w28_,
		_w33_,
		_w34_
	);
	LUT3 #(
		.INIT('h45)
	) name19 (
		\v7_reg/NET0131 ,
		_w23_,
		_w34_,
		_w35_
	);
	LUT3 #(
		.INIT('h8c)
	) name20 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w36_
	);
	LUT4 #(
		.INIT('h0804)
	) name21 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w38_
	);
	LUT4 #(
		.INIT('h0800)
	) name23 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w40_
	);
	LUT3 #(
		.INIT('ha2)
	) name25 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w41_
	);
	LUT4 #(
		.INIT('h0031)
	) name26 (
		_w30_,
		_w39_,
		_w41_,
		_w37_,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\v7_reg/NET0131 ,
		_w42_,
		_w43_
	);
	LUT3 #(
		.INIT('h40)
	) name28 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w44_
	);
	LUT4 #(
		.INIT('h4000)
	) name29 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v8_reg/NET0131 ,
		_w45_
	);
	LUT3 #(
		.INIT('h02)
	) name30 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v7_reg/NET0131 ,
		_w46_
	);
	LUT3 #(
		.INIT('he0)
	) name31 (
		_w44_,
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w48_
	);
	LUT3 #(
		.INIT('h08)
	) name33 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w49_
	);
	LUT3 #(
		.INIT('h08)
	) name34 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w50_
	);
	LUT3 #(
		.INIT('ha8)
	) name35 (
		_w48_,
		_w49_,
		_w50_,
		_w51_
	);
	LUT4 #(
		.INIT('hef23)
	) name36 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT3 #(
		.INIT('h01)
	) name39 (
		_w51_,
		_w54_,
		_w47_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		_w43_,
		_w55_,
		_w56_
	);
	LUT3 #(
		.INIT('h8a)
	) name41 (
		CLR_pad,
		_w35_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w58_
	);
	LUT3 #(
		.INIT('h40)
	) name43 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w59_
	);
	LUT4 #(
		.INIT('hcf73)
	) name44 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w60_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		_w58_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\v10_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w62_
	);
	LUT3 #(
		.INIT('h40)
	) name47 (
		\v11_reg/NET0131 ,
		_w21_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w64_
	);
	LUT4 #(
		.INIT('h0100)
	) name49 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w65_
	);
	LUT4 #(
		.INIT('h0800)
	) name50 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w66_
	);
	LUT3 #(
		.INIT('ha8)
	) name51 (
		_w24_,
		_w65_,
		_w66_,
		_w67_
	);
	LUT3 #(
		.INIT('h01)
	) name52 (
		_w63_,
		_w67_,
		_w61_,
		_w68_
	);
	LUT3 #(
		.INIT('h07)
	) name53 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w69_
	);
	LUT3 #(
		.INIT('h40)
	) name54 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w70_
	);
	LUT4 #(
		.INIT('h8acf)
	) name55 (
		\v10_reg/NET0131 ,
		_w69_,
		_w70_,
		_w65_,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\v2_pad ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w73_
	);
	LUT3 #(
		.INIT('h70)
	) name58 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\v11_reg/NET0131 ,
		\v6_pad ,
		_w76_
	);
	LUT4 #(
		.INIT('h0100)
	) name61 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w77_
	);
	LUT3 #(
		.INIT('h70)
	) name62 (
		\v4_pad ,
		\v5_pad ,
		\v9_reg/NET0131 ,
		_w78_
	);
	LUT4 #(
		.INIT('h153f)
	) name63 (
		_w70_,
		_w76_,
		_w77_,
		_w78_,
		_w79_
	);
	LUT3 #(
		.INIT('h20)
	) name64 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v2_pad ,
		_w80_
	);
	LUT4 #(
		.INIT('h002a)
	) name65 (
		\v10_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v8_reg/NET0131 ,
		_w81_
	);
	LUT3 #(
		.INIT('ha8)
	) name66 (
		_w31_,
		_w80_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		_w83_
	);
	LUT3 #(
		.INIT('h10)
	) name68 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w84_
	);
	LUT4 #(
		.INIT('h2000)
	) name69 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w85_
	);
	LUT4 #(
		.INIT('h0111)
	) name70 (
		\v7_reg/NET0131 ,
		_w85_,
		_w83_,
		_w84_,
		_w86_
	);
	LUT4 #(
		.INIT('h1000)
	) name71 (
		_w82_,
		_w75_,
		_w86_,
		_w79_,
		_w87_
	);
	LUT3 #(
		.INIT('h0e)
	) name72 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w88_
	);
	LUT4 #(
		.INIT('hf100)
	) name73 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w89_
	);
	LUT3 #(
		.INIT('hc4)
	) name74 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w90_
	);
	LUT4 #(
		.INIT('h9010)
	) name75 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w91_
	);
	LUT3 #(
		.INIT('h02)
	) name76 (
		\v8_reg/NET0131 ,
		_w91_,
		_w89_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w93_
	);
	LUT4 #(
		.INIT('h0c04)
	) name78 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\v7_reg/NET0131 ,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w92_,
		_w95_,
		_w96_
	);
	LUT4 #(
		.INIT('h00bf)
	) name81 (
		_w72_,
		_w68_,
		_w87_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		_w98_
	);
	LUT3 #(
		.INIT('h01)
	) name83 (
		\v10_reg/NET0131 ,
		\v6_pad ,
		\v8_reg/NET0131 ,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w100_
	);
	LUT4 #(
		.INIT('h0002)
	) name85 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w101_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name86 (
		_w32_,
		_w98_,
		_w99_,
		_w101_,
		_w102_
	);
	LUT3 #(
		.INIT('h8a)
	) name87 (
		CLR_pad,
		_w97_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w104_
	);
	LUT4 #(
		.INIT('h4000)
	) name89 (
		\v11_reg/NET0131 ,
		_w21_,
		_w62_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w106_
	);
	LUT4 #(
		.INIT('h33f8)
	) name91 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w107_
	);
	LUT3 #(
		.INIT('hc8)
	) name92 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w108_
	);
	LUT4 #(
		.INIT('hc080)
	) name93 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w109_
	);
	LUT4 #(
		.INIT('h3302)
	) name94 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w107_,
		_w109_,
		_w110_
	);
	LUT4 #(
		.INIT('h0f04)
	) name95 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w111_
	);
	LUT4 #(
		.INIT('h0080)
	) name96 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w112_
	);
	LUT3 #(
		.INIT('ha8)
	) name97 (
		\v7_reg/NET0131 ,
		_w111_,
		_w112_,
		_w113_
	);
	LUT4 #(
		.INIT('heeec)
	) name98 (
		\v2_pad ,
		_w105_,
		_w110_,
		_w113_,
		_w114_
	);
	LUT4 #(
		.INIT('hd3df)
	) name99 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v9_reg/NET0131 ,
		_w115_
	);
	LUT3 #(
		.INIT('hc8)
	) name100 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w115_,
		_w116_
	);
	LUT3 #(
		.INIT('hc8)
	) name101 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\v4_pad ,
		\v5_pad ,
		_w118_
	);
	LUT4 #(
		.INIT('h00ba)
	) name103 (
		\v10_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v9_reg/NET0131 ,
		_w119_
	);
	LUT3 #(
		.INIT('h04)
	) name104 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w120_
	);
	LUT4 #(
		.INIT('h00ab)
	) name105 (
		\v12_reg/NET0131 ,
		_w117_,
		_w119_,
		_w120_,
		_w121_
	);
	LUT4 #(
		.INIT('h3323)
	) name106 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w122_
	);
	LUT4 #(
		.INIT('h0010)
	) name107 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w123_
	);
	LUT4 #(
		.INIT('h10f0)
	) name108 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w124_
	);
	LUT3 #(
		.INIT('h04)
	) name109 (
		_w123_,
		_w124_,
		_w122_,
		_w125_
	);
	LUT4 #(
		.INIT('hff54)
	) name110 (
		\v7_reg/NET0131 ,
		_w116_,
		_w121_,
		_w125_,
		_w126_
	);
	LUT4 #(
		.INIT('h2000)
	) name111 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w128_
	);
	LUT4 #(
		.INIT('h0004)
	) name113 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v7_reg/NET0131 ,
		_w129_
	);
	LUT4 #(
		.INIT('hf400)
	) name114 (
		_w19_,
		_w58_,
		_w127_,
		_w129_,
		_w130_
	);
	LUT3 #(
		.INIT('hb0)
	) name115 (
		\v1_pad ,
		\v6_pad ,
		\v8_reg/NET0131 ,
		_w131_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w132_
	);
	LUT4 #(
		.INIT('h8000)
	) name117 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w133_
	);
	LUT3 #(
		.INIT('h80)
	) name118 (
		_w131_,
		_w132_,
		_w133_,
		_w134_
	);
	LUT4 #(
		.INIT('h0222)
	) name119 (
		\v10_reg/NET0131 ,
		\v2_pad ,
		\v4_pad ,
		\v5_pad ,
		_w135_
	);
	LUT4 #(
		.INIT('h50d0)
	) name120 (
		\v9_reg/NET0131 ,
		_w93_,
		_w108_,
		_w135_,
		_w136_
	);
	LUT3 #(
		.INIT('h10)
	) name121 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v6_pad ,
		_w137_
	);
	LUT4 #(
		.INIT('h1000)
	) name122 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v6_pad ,
		_w138_
	);
	LUT4 #(
		.INIT('h2000)
	) name123 (
		\v11_reg/NET0131 ,
		\v1_pad ,
		\v6_pad ,
		\v8_reg/NET0131 ,
		_w139_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		_w140_
	);
	LUT4 #(
		.INIT('h4000)
	) name125 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		_w141_
	);
	LUT4 #(
		.INIT('h0777)
	) name126 (
		_w58_,
		_w138_,
		_w139_,
		_w141_,
		_w142_
	);
	LUT4 #(
		.INIT('h0001)
	) name127 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w143_
	);
	LUT3 #(
		.INIT('h80)
	) name128 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w144_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name129 (
		_w131_,
		_w140_,
		_w143_,
		_w144_,
		_w145_
	);
	LUT3 #(
		.INIT('h54)
	) name130 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w146_
	);
	LUT4 #(
		.INIT('h0a11)
	) name131 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w147_
	);
	LUT3 #(
		.INIT('h08)
	) name132 (
		\v4_pad ,
		\v5_pad ,
		\v9_reg/NET0131 ,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\v0_pad ,
		\v12_reg/NET0131 ,
		_w149_
	);
	LUT4 #(
		.INIT('ha888)
	) name134 (
		\v10_reg/NET0131 ,
		_w147_,
		_w148_,
		_w149_,
		_w150_
	);
	LUT4 #(
		.INIT('h0100)
	) name135 (
		_w136_,
		_w145_,
		_w150_,
		_w142_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w152_
	);
	LUT4 #(
		.INIT('ha8b8)
	) name137 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w153_
	);
	LUT3 #(
		.INIT('h54)
	) name138 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w154_
	);
	LUT4 #(
		.INIT('h8a88)
	) name139 (
		\v7_reg/NET0131 ,
		_w39_,
		_w153_,
		_w154_,
		_w155_
	);
	LUT3 #(
		.INIT('h08)
	) name140 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		_w90_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w158_
	);
	LUT4 #(
		.INIT('h0200)
	) name143 (
		\v1_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w159_
	);
	LUT3 #(
		.INIT('h80)
	) name144 (
		_w137_,
		_w158_,
		_w159_,
		_w160_
	);
	LUT3 #(
		.INIT('h01)
	) name145 (
		_w157_,
		_w155_,
		_w160_,
		_w161_
	);
	LUT4 #(
		.INIT('h02aa)
	) name146 (
		CLR_pad,
		\v7_reg/NET0131 ,
		_w151_,
		_w161_,
		_w162_
	);
	LUT3 #(
		.INIT('h08)
	) name147 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w163_
	);
	LUT4 #(
		.INIT('h2022)
	) name148 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w164_
	);
	LUT3 #(
		.INIT('ha8)
	) name149 (
		_w100_,
		_w163_,
		_w164_,
		_w165_
	);
	LUT4 #(
		.INIT('h0804)
	) name150 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w166_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name151 (
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w167_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w168_
	);
	LUT4 #(
		.INIT('h8808)
	) name153 (
		\v4_pad ,
		\v5_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w169_
	);
	LUT3 #(
		.INIT('h45)
	) name154 (
		_w166_,
		_w167_,
		_w169_,
		_w170_
	);
	LUT3 #(
		.INIT('ha8)
	) name155 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w171_
	);
	LUT4 #(
		.INIT('h0057)
	) name156 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v7_reg/NET0131 ,
		_w172_
	);
	LUT4 #(
		.INIT('h2220)
	) name157 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w173_
	);
	LUT3 #(
		.INIT('h4c)
	) name158 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w174_
	);
	LUT4 #(
		.INIT('h0100)
	) name159 (
		_w120_,
		_w172_,
		_w173_,
		_w174_,
		_w175_
	);
	LUT4 #(
		.INIT('hff45)
	) name160 (
		\v12_reg/NET0131 ,
		_w165_,
		_w170_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w177_
	);
	LUT4 #(
		.INIT('h8088)
	) name162 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v1_pad ,
		\v6_pad ,
		_w178_
	);
	LUT3 #(
		.INIT('ha8)
	) name163 (
		\v3_pad ,
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w180_
	);
	LUT4 #(
		.INIT('h0020)
	) name165 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w181_
	);
	LUT4 #(
		.INIT('hcd00)
	) name166 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		_w181_,
		_w182_,
		_w183_
	);
	LUT4 #(
		.INIT('h0200)
	) name168 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w184_
	);
	LUT4 #(
		.INIT('h0100)
	) name169 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v6_pad ,
		\v9_reg/NET0131 ,
		_w185_
	);
	LUT4 #(
		.INIT('hc400)
	) name170 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w186_
	);
	LUT4 #(
		.INIT('h5554)
	) name171 (
		\v8_reg/NET0131 ,
		_w185_,
		_w186_,
		_w184_,
		_w187_
	);
	LUT4 #(
		.INIT('h0004)
	) name172 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w188_
	);
	LUT4 #(
		.INIT('h2000)
	) name173 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w188_,
		_w189_,
		_w190_
	);
	LUT4 #(
		.INIT('h0045)
	) name175 (
		_w187_,
		_w179_,
		_w183_,
		_w190_,
		_w191_
	);
	LUT4 #(
		.INIT('h7faa)
	) name176 (
		\v11_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v8_reg/NET0131 ,
		_w192_
	);
	LUT3 #(
		.INIT('h10)
	) name177 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w194_
	);
	LUT4 #(
		.INIT('h0080)
	) name179 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w195_
	);
	LUT4 #(
		.INIT('h5510)
	) name180 (
		\v2_pad ,
		_w192_,
		_w193_,
		_w195_,
		_w196_
	);
	LUT3 #(
		.INIT('h70)
	) name181 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w197_
	);
	LUT3 #(
		.INIT('h40)
	) name182 (
		_w31_,
		_w124_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w196_,
		_w198_,
		_w199_
	);
	LUT4 #(
		.INIT('h02aa)
	) name184 (
		CLR_pad,
		\v7_reg/NET0131 ,
		_w191_,
		_w199_,
		_w200_
	);
	LUT3 #(
		.INIT('h32)
	) name185 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w201_
	);
	LUT4 #(
		.INIT('h4055)
	) name186 (
		\v2_pad ,
		\v4_pad ,
		\v5_pad ,
		\v9_reg/NET0131 ,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w201_,
		_w202_,
		_w203_
	);
	LUT4 #(
		.INIT('h2220)
	) name188 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\v10_reg/NET0131 ,
		_w204_,
		_w205_
	);
	LUT3 #(
		.INIT('h20)
	) name190 (
		\v0_pad ,
		\v1_pad ,
		\v6_pad ,
		_w206_
	);
	LUT3 #(
		.INIT('h80)
	) name191 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w207_
	);
	LUT3 #(
		.INIT('h45)
	) name192 (
		_w146_,
		_w206_,
		_w207_,
		_w208_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name193 (
		\v8_reg/NET0131 ,
		_w205_,
		_w203_,
		_w208_,
		_w209_
	);
	LUT4 #(
		.INIT('hfa77)
	) name194 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name195 (
		_w152_,
		_w210_,
		_w211_
	);
	LUT3 #(
		.INIT('h04)
	) name196 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w212_
	);
	LUT4 #(
		.INIT('h9ddf)
	) name197 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w213_
	);
	LUT4 #(
		.INIT('hab00)
	) name198 (
		\v6_pad ,
		_w77_,
		_w212_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w211_,
		_w214_,
		_w215_
	);
	LUT3 #(
		.INIT('h23)
	) name200 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w216_
	);
	LUT4 #(
		.INIT('h1054)
	) name201 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name202 (
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w218_
	);
	LUT3 #(
		.INIT('h10)
	) name203 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w219_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name204 (
		_w216_,
		_w217_,
		_w218_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		_w222_
	);
	LUT3 #(
		.INIT('h80)
	) name207 (
		_w49_,
		_w221_,
		_w222_,
		_w223_
	);
	LUT4 #(
		.INIT('h3313)
	) name208 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w225_
	);
	LUT3 #(
		.INIT('h10)
	) name210 (
		_w117_,
		_w224_,
		_w225_,
		_w226_
	);
	LUT3 #(
		.INIT('h10)
	) name211 (
		_w223_,
		_w226_,
		_w220_,
		_w227_
	);
	LUT4 #(
		.INIT('hba00)
	) name212 (
		\v7_reg/NET0131 ,
		_w209_,
		_w215_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		CLR_pad,
		_w228_,
		_w229_
	);
	LUT3 #(
		.INIT('h20)
	) name214 (
		\v11_reg/NET0131 ,
		_w206_,
		_w207_,
		_w230_
	);
	LUT4 #(
		.INIT('h0111)
	) name215 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w231_
	);
	LUT3 #(
		.INIT('h01)
	) name216 (
		_w59_,
		_w185_,
		_w231_,
		_w232_
	);
	LUT3 #(
		.INIT('h8a)
	) name217 (
		\v8_reg/NET0131 ,
		_w230_,
		_w232_,
		_w233_
	);
	LUT4 #(
		.INIT('haa67)
	) name218 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v6_pad ,
		\v9_reg/NET0131 ,
		_w234_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		_w180_,
		_w234_,
		_w235_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name220 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w236_
	);
	LUT3 #(
		.INIT('h32)
	) name221 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v8_reg/NET0131 ,
		_w237_
	);
	LUT4 #(
		.INIT('h7077)
	) name222 (
		_w21_,
		_w62_,
		_w236_,
		_w237_,
		_w238_
	);
	LUT4 #(
		.INIT('hcac8)
	) name223 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w239_
	);
	LUT3 #(
		.INIT('h8a)
	) name224 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w240_
	);
	LUT4 #(
		.INIT('h3020)
	) name225 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w241_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name226 (
		_w168_,
		_w239_,
		_w240_,
		_w241_,
		_w242_
	);
	LUT4 #(
		.INIT('h0e00)
	) name227 (
		\v11_reg/NET0131 ,
		_w238_,
		_w235_,
		_w242_,
		_w243_
	);
	LUT3 #(
		.INIT('h90)
	) name228 (
		\v10_reg/NET0131 ,
		_w40_,
		_w53_,
		_w244_
	);
	LUT3 #(
		.INIT('h23)
	) name229 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w245_
	);
	LUT3 #(
		.INIT('h40)
	) name230 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w246_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		_w245_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w244_,
		_w247_,
		_w248_
	);
	LUT4 #(
		.INIT('hba00)
	) name233 (
		\v7_reg/NET0131 ,
		_w233_,
		_w243_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		CLR_pad,
		_w249_,
		_w250_
	);
	LUT4 #(
		.INIT('h0053)
	) name235 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		\v8_reg/NET0131 ,
		_w251_,
		_w252_
	);
	LUT3 #(
		.INIT('hd0)
	) name237 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w253_
	);
	LUT3 #(
		.INIT('h40)
	) name238 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		\v6_pad ,
		_w254_
	);
	LUT4 #(
		.INIT('h80c0)
	) name239 (
		\v11_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v8_reg/NET0131 ,
		_w255_
	);
	LUT4 #(
		.INIT('h1101)
	) name240 (
		\v12_reg/NET0131 ,
		_w255_,
		_w253_,
		_w254_,
		_w256_
	);
	LUT4 #(
		.INIT('h0004)
	) name241 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w124_,
		_w257_,
		_w258_
	);
	LUT4 #(
		.INIT('h45ff)
	) name243 (
		\v7_reg/NET0131 ,
		_w252_,
		_w256_,
		_w258_,
		_w259_
	);
	LUT3 #(
		.INIT('h40)
	) name244 (
		\v10_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w260_
	);
	LUT3 #(
		.INIT('h07)
	) name245 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w261_
	);
	LUT4 #(
		.INIT('h002f)
	) name246 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w262_
	);
	LUT4 #(
		.INIT('h1055)
	) name247 (
		_w39_,
		_w260_,
		_w261_,
		_w262_,
		_w263_
	);
	LUT4 #(
		.INIT('h0004)
	) name248 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w264_
	);
	LUT4 #(
		.INIT('h3301)
	) name249 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w263_,
		_w264_,
		_w265_
	);
	LUT3 #(
		.INIT('h3a)
	) name250 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w266_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name251 (
		\v8_reg/NET0131 ,
		_w171_,
		_w225_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('he)
	) name252 (
		_w265_,
		_w267_,
		_w268_
	);
	LUT4 #(
		.INIT('h004f)
	) name253 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w269_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name254 (
		\v8_reg/NET0131 ,
		_w20_,
		_w127_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w108_,
		_w222_,
		_w271_
	);
	LUT3 #(
		.INIT('hd1)
	) name256 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w272_
	);
	LUT3 #(
		.INIT('h06)
	) name257 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT4 #(
		.INIT('h00ab)
	) name259 (
		\v12_reg/NET0131 ,
		_w270_,
		_w271_,
		_w274_,
		_w275_
	);
	LUT4 #(
		.INIT('hfdea)
	) name260 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w276_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name261 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w257_,
		_w276_,
		_w277_
	);
	LUT4 #(
		.INIT('h54fc)
	) name262 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w278_
	);
	LUT3 #(
		.INIT('h32)
	) name263 (
		\v9_reg/NET0131 ,
		_w177_,
		_w278_,
		_w279_
	);
	LUT4 #(
		.INIT('h1030)
	) name264 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w280_
	);
	LUT2 #(
		.INIT('h2)
	) name265 (
		\v10_reg/NET0131 ,
		_w280_,
		_w281_
	);
	LUT3 #(
		.INIT('h45)
	) name266 (
		_w277_,
		_w279_,
		_w281_,
		_w282_
	);
	LUT3 #(
		.INIT('h1f)
	) name267 (
		\v7_reg/NET0131 ,
		_w275_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		\v8_reg/NET0131 ,
		_w269_,
		_w284_
	);
	LUT3 #(
		.INIT('h15)
	) name269 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w285_
	);
	LUT4 #(
		.INIT('hddd0)
	) name270 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w286_
	);
	LUT3 #(
		.INIT('h40)
	) name271 (
		_w253_,
		_w285_,
		_w286_,
		_w287_
	);
	LUT4 #(
		.INIT('h030b)
	) name272 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w288_
	);
	LUT3 #(
		.INIT('h51)
	) name273 (
		_w124_,
		_w225_,
		_w288_,
		_w289_
	);
	LUT4 #(
		.INIT('h45ff)
	) name274 (
		\v7_reg/NET0131 ,
		_w284_,
		_w287_,
		_w289_,
		_w290_
	);
	LUT4 #(
		.INIT('h135f)
	) name275 (
		_w49_,
		_w193_,
		_w222_,
		_w254_,
		_w291_
	);
	LUT2 #(
		.INIT('h2)
	) name276 (
		_w221_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w20_,
		_w143_,
		_w293_
	);
	LUT3 #(
		.INIT('h40)
	) name278 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w294_
	);
	LUT3 #(
		.INIT('ha8)
	) name279 (
		\v11_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w295_
	);
	LUT3 #(
		.INIT('he0)
	) name280 (
		_w188_,
		_w294_,
		_w295_,
		_w296_
	);
	LUT3 #(
		.INIT('ha8)
	) name281 (
		_w128_,
		_w293_,
		_w296_,
		_w297_
	);
	LUT3 #(
		.INIT('h20)
	) name282 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v6_pad ,
		_w298_
	);
	LUT4 #(
		.INIT('h135f)
	) name283 (
		_w40_,
		_w73_,
		_w99_,
		_w298_,
		_w299_
	);
	LUT3 #(
		.INIT('h04)
	) name284 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		\v7_reg/NET0131 ,
		_w300_
	);
	LUT3 #(
		.INIT('hba)
	) name285 (
		_w223_,
		_w299_,
		_w300_,
		_w301_
	);
	LUT3 #(
		.INIT('h80)
	) name286 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w302_
	);
	LUT3 #(
		.INIT('h01)
	) name287 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w303_
	);
	LUT4 #(
		.INIT('hf800)
	) name288 (
		_w64_,
		_w148_,
		_w302_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		_w184_,
		_w194_,
		_w305_
	);
	LUT4 #(
		.INIT('h0100)
	) name290 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w306_
	);
	LUT3 #(
		.INIT('h20)
	) name291 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w308_
	);
	LUT3 #(
		.INIT('he0)
	) name293 (
		_w306_,
		_w307_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('he)
	) name294 (
		_w305_,
		_w309_,
		_w310_
	);
	LUT4 #(
		.INIT('h0080)
	) name295 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w311_
	);
	LUT4 #(
		.INIT('h8000)
	) name296 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w312_
	);
	LUT4 #(
		.INIT('h00ab)
	) name297 (
		\v9_reg/NET0131 ,
		_w138_,
		_w311_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		_w104_,
		_w313_,
		_w314_
	);
	LUT3 #(
		.INIT('h90)
	) name299 (
		\v10_reg/NET0131 ,
		_w73_,
		_w225_,
		_w315_
	);
	LUT4 #(
		.INIT('hee5f)
	) name300 (
		\v12_reg/NET0131 ,
		\v5_pad ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w316_
	);
	LUT4 #(
		.INIT('h2300)
	) name301 (
		\v10_reg/NET0131 ,
		\v2_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w316_,
		_w317_,
		_w318_
	);
	LUT3 #(
		.INIT('ha8)
	) name303 (
		\v11_reg/NET0131 ,
		_w315_,
		_w318_,
		_w319_
	);
	LUT3 #(
		.INIT('h80)
	) name304 (
		_w83_,
		_w73_,
		_w298_,
		_w320_
	);
	LUT4 #(
		.INIT('h9990)
	) name305 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v5_pad ,
		_w321_
	);
	LUT3 #(
		.INIT('h02)
	) name306 (
		_w58_,
		_w88_,
		_w321_,
		_w322_
	);
	LUT4 #(
		.INIT('h1000)
	) name307 (
		\v10_reg/NET0131 ,
		\v2_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w323_
	);
	LUT3 #(
		.INIT('h08)
	) name308 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v5_pad ,
		_w324_
	);
	LUT3 #(
		.INIT('h01)
	) name309 (
		\v0_pad ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w325_
	);
	LUT4 #(
		.INIT('hec00)
	) name310 (
		_w104_,
		_w323_,
		_w324_,
		_w325_,
		_w326_
	);
	LUT4 #(
		.INIT('h00ab)
	) name311 (
		\v7_reg/NET0131 ,
		_w320_,
		_w322_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('hb)
	) name312 (
		_w319_,
		_w327_,
		_w328_
	);
	LUT3 #(
		.INIT('hc9)
	) name313 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w329_
	);
	LUT4 #(
		.INIT('h3f15)
	) name314 (
		_w53_,
		_w38_,
		_w36_,
		_w329_,
		_w330_
	);
	LUT4 #(
		.INIT('h0042)
	) name315 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w331_
	);
	LUT4 #(
		.INIT('h0200)
	) name316 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w332_
	);
	LUT3 #(
		.INIT('h54)
	) name317 (
		\v9_reg/NET0131 ,
		_w331_,
		_w332_,
		_w333_
	);
	LUT3 #(
		.INIT('h45)
	) name318 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w334_
	);
	LUT3 #(
		.INIT('he0)
	) name319 (
		_w127_,
		_w188_,
		_w334_,
		_w335_
	);
	LUT4 #(
		.INIT('h7772)
	) name320 (
		\v7_reg/NET0131 ,
		_w330_,
		_w333_,
		_w335_,
		_w336_
	);
	LUT3 #(
		.INIT('hc8)
	) name321 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w337_
	);
	LUT4 #(
		.INIT('h00fd)
	) name322 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w338_
	);
	LUT3 #(
		.INIT('h45)
	) name323 (
		\v8_reg/NET0131 ,
		_w337_,
		_w338_,
		_w339_
	);
	LUT4 #(
		.INIT('hfd20)
	) name324 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w340_
	);
	LUT3 #(
		.INIT('h54)
	) name325 (
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w340_,
		_w341_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name326 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w342_
	);
	LUT4 #(
		.INIT('h0054)
	) name327 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w343_
	);
	LUT3 #(
		.INIT('h13)
	) name328 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w344_
	);
	LUT4 #(
		.INIT('h0e00)
	) name329 (
		_w118_,
		_w342_,
		_w343_,
		_w344_,
		_w345_
	);
	LUT3 #(
		.INIT('he0)
	) name330 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w346_
	);
	LUT4 #(
		.INIT('h2a00)
	) name331 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w347_
	);
	LUT4 #(
		.INIT('h2022)
	) name332 (
		\v7_reg/NET0131 ,
		_w257_,
		_w346_,
		_w347_,
		_w348_
	);
	LUT4 #(
		.INIT('h00ef)
	) name333 (
		_w341_,
		_w339_,
		_w345_,
		_w348_,
		_w349_
	);
	LUT4 #(
		.INIT('h5040)
	) name334 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w106_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('he)
	) name336 (
		_w349_,
		_w351_,
		_w352_
	);
	LUT3 #(
		.INIT('h04)
	) name337 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w353_
	);
	LUT3 #(
		.INIT('ha8)
	) name338 (
		_w132_,
		_w163_,
		_w353_,
		_w354_
	);
	LUT3 #(
		.INIT('h35)
	) name339 (
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w355_
	);
	LUT4 #(
		.INIT('hea00)
	) name340 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w356_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w355_,
		_w356_,
		_w357_
	);
	LUT3 #(
		.INIT('h54)
	) name342 (
		\v12_reg/NET0131 ,
		_w354_,
		_w357_,
		_w358_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1757/_0_  = _w57_ ;
	assign \g1763/_1_  = _w103_ ;
	assign \g1787/_3_  = _w114_ ;
	assign \g1800/_3_  = _w126_ ;
	assign \g1821/_2_  = _w130_ ;
	assign \g1940/_1_  = _w134_ ;
	assign \g25/_0_  = _w162_ ;
	assign \g2783/_3_  = _w176_ ;
	assign \g2823/_0_  = _w200_ ;
	assign \g38/_1_  = _w229_ ;
	assign \g40/_1_  = _w250_ ;
	assign \v13_D_11_pad  = _w259_ ;
	assign \v13_D_12_pad  = _w268_ ;
	assign \v13_D_13_pad  = _w283_ ;
	assign \v13_D_14_pad  = _w290_ ;
	assign \v13_D_16_pad  = _w292_ ;
	assign \v13_D_18_pad  = _w297_ ;
	assign \v13_D_19_pad  = _w301_ ;
	assign \v13_D_21_pad  = _w304_ ;
	assign \v13_D_22_pad  = _w310_ ;
	assign \v13_D_23_pad  = _w314_ ;
	assign \v13_D_24_pad  = _w328_ ;
	assign \v13_D_7_pad  = _w336_ ;
	assign \v13_D_8_pad  = _w352_ ;
	assign \v13_D_9_pad  = _w358_ ;
endmodule;