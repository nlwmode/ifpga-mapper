module top( \DataOut_pad_o[0]_pad  , \DataOut_pad_o[1]_pad  , \DataOut_pad_o[2]_pad  , \DataOut_pad_o[3]_pad  , \DataOut_pad_o[4]_pad  , \DataOut_pad_o[5]_pad  , \DataOut_pad_o[6]_pad  , \DataOut_pad_o[7]_pad  , \LineState_pad_i[0]_pad  , \LineState_pad_i[1]_pad  , \LineState_r_reg[0]/P0001  , \LineState_r_reg[1]/P0001  , \OpMode_pad_o[1]_pad  , RxActive_pad_i_pad , RxError_pad_i_pad , RxValid_pad_i_pad , TermSel_pad_o_pad , TxReady_pad_i_pad , TxValid_pad_o_pad , VControl_Load_pad_o_pad , XcvSelect_pad_o_pad , \dma_ack_i[0]_pad  , \dma_ack_i[1]_pad  , \dma_ack_i[2]_pad  , \dma_ack_i[3]_pad  , \dma_req_o[0]_pad  , \dma_req_o[1]_pad  , \dma_req_o[2]_pad  , \dma_req_o[3]_pad  , resume_req_i_pad , \resume_req_r_reg/P0001  , rst_i_pad , \sram_data_i[0]_pad  , \sram_data_i[10]_pad  , \sram_data_i[11]_pad  , \sram_data_i[12]_pad  , \sram_data_i[13]_pad  , \sram_data_i[14]_pad  , \sram_data_i[15]_pad  , \sram_data_i[16]_pad  , \sram_data_i[17]_pad  , \sram_data_i[18]_pad  , \sram_data_i[19]_pad  , \sram_data_i[1]_pad  , \sram_data_i[20]_pad  , \sram_data_i[21]_pad  , \sram_data_i[22]_pad  , \sram_data_i[23]_pad  , \sram_data_i[24]_pad  , \sram_data_i[25]_pad  , \sram_data_i[26]_pad  , \sram_data_i[27]_pad  , \sram_data_i[28]_pad  , \sram_data_i[29]_pad  , \sram_data_i[2]_pad  , \sram_data_i[30]_pad  , \sram_data_i[31]_pad  , \sram_data_i[3]_pad  , \sram_data_i[4]_pad  , \sram_data_i[5]_pad  , \sram_data_i[6]_pad  , \sram_data_i[7]_pad  , \sram_data_i[8]_pad  , \sram_data_i[9]_pad  , susp_o_pad , \suspend_clr_wr_reg/P0001  , \u0_drive_k_r_reg/P0001  , \u0_rx_active_reg/P0001  , \u0_rx_data_reg[0]/P0001  , \u0_rx_data_reg[1]/P0001  , \u0_rx_data_reg[2]/P0001  , \u0_rx_data_reg[3]/P0001  , \u0_rx_data_reg[4]/P0001  , \u0_rx_data_reg[5]/P0001  , \u0_rx_data_reg[6]/P0001  , \u0_rx_data_reg[7]/P0001  , \u0_rx_err_reg/P0001  , \u0_rx_valid_reg/P0001  , \u0_tx_ready_reg/NET0131  , \u0_u0_T1_gt_2_5_uS_reg/P0001  , \u0_u0_T1_gt_3_0_mS_reg/P0001  , \u0_u0_T1_gt_5_0_mS_reg/P0001  , \u0_u0_T1_st_3_0_mS_reg/P0001  , \u0_u0_T2_gt_100_uS_reg/P0001  , \u0_u0_T2_gt_1_0_mS_reg/P0001  , \u0_u0_T2_wakeup_reg/P0001  , \u0_u0_chirp_cnt_is_6_reg/P0001  , \u0_u0_chirp_cnt_reg[0]/P0001  , \u0_u0_chirp_cnt_reg[1]/P0001  , \u0_u0_chirp_cnt_reg[2]/P0001  , \u0_u0_drive_k_reg/P0001  , \u0_u0_idle_cnt1_clr_reg/P0001  , \u0_u0_idle_cnt1_next_reg[0]/P0001  , \u0_u0_idle_cnt1_next_reg[1]/P0001  , \u0_u0_idle_cnt1_next_reg[2]/P0001  , \u0_u0_idle_cnt1_next_reg[3]/P0001  , \u0_u0_idle_cnt1_next_reg[4]/P0001  , \u0_u0_idle_cnt1_next_reg[5]/P0001  , \u0_u0_idle_cnt1_next_reg[6]/P0001  , \u0_u0_idle_cnt1_next_reg[7]/P0001  , \u0_u0_idle_cnt1_reg[0]/P0001  , \u0_u0_idle_cnt1_reg[1]/P0001  , \u0_u0_idle_cnt1_reg[2]/P0001  , \u0_u0_idle_cnt1_reg[3]/P0001  , \u0_u0_idle_cnt1_reg[4]/P0001  , \u0_u0_idle_cnt1_reg[5]/P0001  , \u0_u0_idle_cnt1_reg[6]/P0001  , \u0_u0_idle_cnt1_reg[7]/P0001  , \u0_u0_idle_long_reg/P0001  , \u0_u0_ls_idle_r_reg/P0001  , \u0_u0_ls_j_r_reg/P0001  , \u0_u0_ls_k_r_reg/P0001  , \u0_u0_ls_se0_r_reg/P0001  , \u0_u0_me_cnt_100_ms_reg/P0001  , \u0_u0_me_cnt_reg[0]/P0001  , \u0_u0_me_cnt_reg[1]/P0001  , \u0_u0_me_cnt_reg[2]/P0001  , \u0_u0_me_cnt_reg[3]/P0001  , \u0_u0_me_cnt_reg[4]/P0001  , \u0_u0_me_cnt_reg[5]/P0001  , \u0_u0_me_cnt_reg[6]/P0001  , \u0_u0_me_cnt_reg[7]/P0001  , \u0_u0_me_ps2_0_5_ms_reg/P0001  , \u0_u0_me_ps2_reg[0]/P0001  , \u0_u0_me_ps2_reg[1]/P0001  , \u0_u0_me_ps2_reg[2]/P0001  , \u0_u0_me_ps2_reg[3]/P0001  , \u0_u0_me_ps2_reg[4]/P0001  , \u0_u0_me_ps2_reg[5]/P0001  , \u0_u0_me_ps2_reg[6]/P0001  , \u0_u0_me_ps2_reg[7]/P0001  , \u0_u0_me_ps_2_5_us_reg/P0001  , \u0_u0_me_ps_reg[0]/P0001  , \u0_u0_me_ps_reg[1]/P0001  , \u0_u0_me_ps_reg[2]/P0001  , \u0_u0_me_ps_reg[3]/P0001  , \u0_u0_me_ps_reg[4]/P0001  , \u0_u0_me_ps_reg[5]/P0001  , \u0_u0_me_ps_reg[6]/P0001  , \u0_u0_me_ps_reg[7]/P0001  , \u0_u0_mode_hs_reg/P0001  , \u0_u0_ps_cnt_clr_reg/P0001  , \u0_u0_ps_cnt_reg[0]/P0001  , \u0_u0_ps_cnt_reg[1]/P0001  , \u0_u0_ps_cnt_reg[2]/P0001  , \u0_u0_ps_cnt_reg[3]/P0001  , \u0_u0_resume_req_s_reg/P0001  , \u0_u0_state_reg[0]/NET0131  , \u0_u0_state_reg[10]/P0001  , \u0_u0_state_reg[11]/NET0131  , \u0_u0_state_reg[12]/NET0131  , \u0_u0_state_reg[13]/NET0131  , \u0_u0_state_reg[14]/P0001  , \u0_u0_state_reg[1]/P0001  , \u0_u0_state_reg[2]/NET0131  , \u0_u0_state_reg[3]/P0001  , \u0_u0_state_reg[4]/NET0131  , \u0_u0_state_reg[5]/P0001  , \u0_u0_state_reg[6]/NET0131  , \u0_u0_state_reg[7]/NET0131  , \u0_u0_state_reg[8]/NET0131  , \u0_u0_state_reg[9]/P0001  , \u0_u0_usb_attached_reg/P0001  , \u0_u0_usb_suspend_reg/P0001  , \u1_clr_sof_time_reg/P0001  , \u1_frame_no_r_reg[0]/P0001  , \u1_frame_no_r_reg[10]/P0001  , \u1_frame_no_r_reg[1]/P0001  , \u1_frame_no_r_reg[2]/P0001  , \u1_frame_no_r_reg[3]/P0001  , \u1_frame_no_r_reg[4]/P0001  , \u1_frame_no_r_reg[5]/P0001  , \u1_frame_no_r_reg[6]/P0001  , \u1_frame_no_r_reg[7]/P0001  , \u1_frame_no_r_reg[8]/P0001  , \u1_frame_no_r_reg[9]/P0001  , \u1_frame_no_same_reg/P0001  , \u1_hms_clk_reg/P0001  , \u1_hms_cnt_reg[0]/P0001  , \u1_hms_cnt_reg[1]/P0001  , \u1_hms_cnt_reg[2]/P0001  , \u1_hms_cnt_reg[3]/P0001  , \u1_hms_cnt_reg[4]/P0001  , \u1_mfm_cnt_reg[0]/P0001  , \u1_mfm_cnt_reg[1]/P0001  , \u1_mfm_cnt_reg[2]/P0001  , \u1_mfm_cnt_reg[3]/P0001  , \u1_sof_time_reg[0]/P0001  , \u1_sof_time_reg[10]/P0001  , \u1_sof_time_reg[11]/P0001  , \u1_sof_time_reg[1]/P0001  , \u1_sof_time_reg[2]/P0001  , \u1_sof_time_reg[3]/P0001  , \u1_sof_time_reg[4]/P0001  , \u1_sof_time_reg[5]/P0001  , \u1_sof_time_reg[6]/P0001  , \u1_sof_time_reg[7]/P0001  , \u1_sof_time_reg[8]/P0001  , \u1_sof_time_reg[9]/P0001  , \u1_u0_crc16_sum_reg[0]/P0001  , \u1_u0_crc16_sum_reg[10]/P0001  , \u1_u0_crc16_sum_reg[11]/P0001  , \u1_u0_crc16_sum_reg[12]/P0001  , \u1_u0_crc16_sum_reg[13]/P0001  , \u1_u0_crc16_sum_reg[14]/P0001  , \u1_u0_crc16_sum_reg[15]/P0001  , \u1_u0_crc16_sum_reg[1]/P0001  , \u1_u0_crc16_sum_reg[2]/P0001  , \u1_u0_crc16_sum_reg[3]/P0001  , \u1_u0_crc16_sum_reg[4]/P0001  , \u1_u0_crc16_sum_reg[5]/P0001  , \u1_u0_crc16_sum_reg[6]/P0001  , \u1_u0_crc16_sum_reg[7]/P0001  , \u1_u0_crc16_sum_reg[8]/P0001  , \u1_u0_crc16_sum_reg[9]/P0001  , \u1_u0_data_valid0_reg/P0001  , \u1_u0_pid_reg[0]/NET0131  , \u1_u0_pid_reg[1]/NET0131  , \u1_u0_pid_reg[2]/NET0131  , \u1_u0_pid_reg[3]/NET0131  , \u1_u0_pid_reg[4]/P0001  , \u1_u0_pid_reg[5]/P0001  , \u1_u0_pid_reg[6]/P0001  , \u1_u0_pid_reg[7]/P0001  , \u1_u0_rx_active_r_reg/P0001  , \u1_u0_rxv1_reg/P0001  , \u1_u0_rxv2_reg/P0001  , \u1_u0_state_reg[0]/P0001  , \u1_u0_state_reg[1]/P0001  , \u1_u0_state_reg[2]/P0001  , \u1_u0_state_reg[3]/P0001  , \u1_u0_token0_reg[0]/NET0131  , \u1_u0_token0_reg[1]/P0001  , \u1_u0_token0_reg[2]/NET0131  , \u1_u0_token0_reg[3]/NET0131  , \u1_u0_token0_reg[4]/P0001  , \u1_u0_token0_reg[5]/NET0131  , \u1_u0_token0_reg[6]/P0001  , \u1_u0_token0_reg[7]/P0001  , \u1_u0_token1_reg[0]/P0001  , \u1_u0_token1_reg[1]/P0001  , \u1_u0_token1_reg[2]/P0001  , \u1_u0_token1_reg[3]/P0001  , \u1_u0_token1_reg[4]/P0001  , \u1_u0_token1_reg[5]/P0001  , \u1_u0_token1_reg[6]/P0001  , \u1_u0_token1_reg[7]/P0001  , \u1_u0_token_valid_r1_reg/P0001  , \u1_u0_token_valid_str1_reg/P0001  , \u1_u1_crc16_reg[0]/P0001  , \u1_u1_crc16_reg[10]/P0001  , \u1_u1_crc16_reg[11]/P0001  , \u1_u1_crc16_reg[12]/P0001  , \u1_u1_crc16_reg[13]/P0001  , \u1_u1_crc16_reg[14]/P0001  , \u1_u1_crc16_reg[15]/P0001  , \u1_u1_crc16_reg[1]/P0001  , \u1_u1_crc16_reg[2]/P0001  , \u1_u1_crc16_reg[3]/P0001  , \u1_u1_crc16_reg[4]/P0001  , \u1_u1_crc16_reg[5]/P0001  , \u1_u1_crc16_reg[6]/P0001  , \u1_u1_crc16_reg[7]/P0001  , \u1_u1_crc16_reg[8]/P0001  , \u1_u1_crc16_reg[9]/P0001  , \u1_u1_send_data_r2_reg/P0001  , \u1_u1_send_data_r_reg/P0001  , \u1_u1_send_token_r_reg/P0001  , \u1_u1_send_zero_length_r_reg/P0001  , \u1_u1_state_reg[0]/NET0131  , \u1_u1_state_reg[1]/NET0131  , \u1_u1_state_reg[2]/NET0131  , \u1_u1_state_reg[3]/NET0131  , \u1_u1_state_reg[4]/NET0131  , \u1_u1_tx_first_r_reg/P0001  , \u1_u1_tx_valid_r_reg/NET0131  , \u1_u1_zero_length_r_reg/P0001  , \u1_u2_adr_cb_reg[0]/NET0131  , \u1_u2_adr_cb_reg[1]/NET0131  , \u1_u2_adr_cb_reg[2]/NET0131  , \u1_u2_adr_cw_reg[0]/NET0131  , \u1_u2_adr_cw_reg[10]/P0001  , \u1_u2_adr_cw_reg[11]/P0001  , \u1_u2_adr_cw_reg[12]/P0001  , \u1_u2_adr_cw_reg[13]/P0001  , \u1_u2_adr_cw_reg[14]/P0001  , \u1_u2_adr_cw_reg[1]/P0001  , \u1_u2_adr_cw_reg[2]/P0001  , \u1_u2_adr_cw_reg[3]/NET0131  , \u1_u2_adr_cw_reg[4]/P0001  , \u1_u2_adr_cw_reg[5]/NET0131  , \u1_u2_adr_cw_reg[6]/NET0131  , \u1_u2_adr_cw_reg[7]/NET0131  , \u1_u2_adr_cw_reg[8]/P0001  , \u1_u2_adr_cw_reg[9]/NET0131  , \u1_u2_dout_r_reg[0]/P0001  , \u1_u2_dout_r_reg[10]/P0001  , \u1_u2_dout_r_reg[11]/P0001  , \u1_u2_dout_r_reg[12]/P0001  , \u1_u2_dout_r_reg[13]/P0001  , \u1_u2_dout_r_reg[14]/P0001  , \u1_u2_dout_r_reg[15]/P0001  , \u1_u2_dout_r_reg[16]/P0001  , \u1_u2_dout_r_reg[17]/P0001  , \u1_u2_dout_r_reg[18]/P0001  , \u1_u2_dout_r_reg[19]/P0001  , \u1_u2_dout_r_reg[1]/P0001  , \u1_u2_dout_r_reg[20]/P0001  , \u1_u2_dout_r_reg[21]/P0001  , \u1_u2_dout_r_reg[22]/P0001  , \u1_u2_dout_r_reg[23]/P0001  , \u1_u2_dout_r_reg[24]/P0001  , \u1_u2_dout_r_reg[25]/P0001  , \u1_u2_dout_r_reg[26]/P0001  , \u1_u2_dout_r_reg[27]/P0001  , \u1_u2_dout_r_reg[28]/P0001  , \u1_u2_dout_r_reg[29]/P0001  , \u1_u2_dout_r_reg[2]/P0001  , \u1_u2_dout_r_reg[30]/P0001  , \u1_u2_dout_r_reg[31]/P0001  , \u1_u2_dout_r_reg[3]/P0001  , \u1_u2_dout_r_reg[4]/P0001  , \u1_u2_dout_r_reg[5]/P0001  , \u1_u2_dout_r_reg[6]/P0001  , \u1_u2_dout_r_reg[7]/P0001  , \u1_u2_dout_r_reg[8]/P0001  , \u1_u2_dout_r_reg[9]/P0001  , \u1_u2_dtmp_r_reg[0]/P0001  , \u1_u2_dtmp_r_reg[10]/P0001  , \u1_u2_dtmp_r_reg[11]/P0001  , \u1_u2_dtmp_r_reg[12]/P0001  , \u1_u2_dtmp_r_reg[13]/P0001  , \u1_u2_dtmp_r_reg[14]/P0001  , \u1_u2_dtmp_r_reg[15]/P0001  , \u1_u2_dtmp_r_reg[16]/P0001  , \u1_u2_dtmp_r_reg[17]/P0001  , \u1_u2_dtmp_r_reg[18]/P0001  , \u1_u2_dtmp_r_reg[19]/P0001  , \u1_u2_dtmp_r_reg[1]/P0001  , \u1_u2_dtmp_r_reg[20]/P0001  , \u1_u2_dtmp_r_reg[21]/P0001  , \u1_u2_dtmp_r_reg[22]/P0001  , \u1_u2_dtmp_r_reg[23]/P0001  , \u1_u2_dtmp_r_reg[24]/P0001  , \u1_u2_dtmp_r_reg[25]/P0001  , \u1_u2_dtmp_r_reg[26]/P0001  , \u1_u2_dtmp_r_reg[27]/P0001  , \u1_u2_dtmp_r_reg[28]/P0001  , \u1_u2_dtmp_r_reg[29]/P0001  , \u1_u2_dtmp_r_reg[2]/P0001  , \u1_u2_dtmp_r_reg[30]/P0001  , \u1_u2_dtmp_r_reg[31]/P0001  , \u1_u2_dtmp_r_reg[3]/P0001  , \u1_u2_dtmp_r_reg[4]/P0001  , \u1_u2_dtmp_r_reg[5]/P0001  , \u1_u2_dtmp_r_reg[6]/P0001  , \u1_u2_dtmp_r_reg[7]/P0001  , \u1_u2_dtmp_r_reg[8]/P0001  , \u1_u2_dtmp_r_reg[9]/P0001  , \u1_u2_dtmp_sel_r_reg/P0001  , \u1_u2_idma_done_reg/P0001  , \u1_u2_last_buf_adr_reg[0]/P0001  , \u1_u2_last_buf_adr_reg[10]/P0001  , \u1_u2_last_buf_adr_reg[11]/P0001  , \u1_u2_last_buf_adr_reg[12]/P0001  , \u1_u2_last_buf_adr_reg[13]/P0001  , \u1_u2_last_buf_adr_reg[14]/P0001  , \u1_u2_last_buf_adr_reg[1]/P0001  , \u1_u2_last_buf_adr_reg[2]/P0001  , \u1_u2_last_buf_adr_reg[3]/P0001  , \u1_u2_last_buf_adr_reg[4]/P0001  , \u1_u2_last_buf_adr_reg[5]/P0001  , \u1_u2_last_buf_adr_reg[6]/P0001  , \u1_u2_last_buf_adr_reg[7]/P0001  , \u1_u2_last_buf_adr_reg[8]/P0001  , \u1_u2_last_buf_adr_reg[9]/P0001  , \u1_u2_mack_r_reg/P0001  , \u1_u2_mwe_reg/P0001  , \u1_u2_rd_buf0_reg[0]/NET0131  , \u1_u2_rd_buf0_reg[10]/NET0131  , \u1_u2_rd_buf0_reg[11]/NET0131  , \u1_u2_rd_buf0_reg[12]/P0001  , \u1_u2_rd_buf0_reg[13]/P0001  , \u1_u2_rd_buf0_reg[14]/P0001  , \u1_u2_rd_buf0_reg[15]/P0001  , \u1_u2_rd_buf0_reg[16]/NET0131  , \u1_u2_rd_buf0_reg[17]/NET0131  , \u1_u2_rd_buf0_reg[18]/NET0131  , \u1_u2_rd_buf0_reg[19]/NET0131  , \u1_u2_rd_buf0_reg[1]/NET0131  , \u1_u2_rd_buf0_reg[20]/P0001  , \u1_u2_rd_buf0_reg[21]/P0001  , \u1_u2_rd_buf0_reg[22]/P0001  , \u1_u2_rd_buf0_reg[23]/P0001  , \u1_u2_rd_buf0_reg[24]/NET0131  , \u1_u2_rd_buf0_reg[25]/NET0131  , \u1_u2_rd_buf0_reg[26]/NET0131  , \u1_u2_rd_buf0_reg[27]/NET0131  , \u1_u2_rd_buf0_reg[28]/P0001  , \u1_u2_rd_buf0_reg[29]/P0001  , \u1_u2_rd_buf0_reg[2]/NET0131  , \u1_u2_rd_buf0_reg[30]/P0001  , \u1_u2_rd_buf0_reg[31]/P0001  , \u1_u2_rd_buf0_reg[3]/NET0131  , \u1_u2_rd_buf0_reg[4]/P0001  , \u1_u2_rd_buf0_reg[5]/P0001  , \u1_u2_rd_buf0_reg[6]/P0001  , \u1_u2_rd_buf0_reg[7]/P0001  , \u1_u2_rd_buf0_reg[8]/NET0131  , \u1_u2_rd_buf0_reg[9]/NET0131  , \u1_u2_rd_buf1_reg[0]/NET0131  , \u1_u2_rd_buf1_reg[10]/NET0131  , \u1_u2_rd_buf1_reg[11]/NET0131  , \u1_u2_rd_buf1_reg[12]/P0001  , \u1_u2_rd_buf1_reg[13]/P0001  , \u1_u2_rd_buf1_reg[14]/P0001  , \u1_u2_rd_buf1_reg[15]/P0001  , \u1_u2_rd_buf1_reg[16]/NET0131  , \u1_u2_rd_buf1_reg[17]/NET0131  , \u1_u2_rd_buf1_reg[18]/NET0131  , \u1_u2_rd_buf1_reg[19]/NET0131  , \u1_u2_rd_buf1_reg[1]/NET0131  , \u1_u2_rd_buf1_reg[20]/P0001  , \u1_u2_rd_buf1_reg[21]/P0001  , \u1_u2_rd_buf1_reg[22]/P0001  , \u1_u2_rd_buf1_reg[23]/P0001  , \u1_u2_rd_buf1_reg[24]/NET0131  , \u1_u2_rd_buf1_reg[25]/NET0131  , \u1_u2_rd_buf1_reg[26]/NET0131  , \u1_u2_rd_buf1_reg[27]/NET0131  , \u1_u2_rd_buf1_reg[28]/P0001  , \u1_u2_rd_buf1_reg[29]/P0001  , \u1_u2_rd_buf1_reg[2]/NET0131  , \u1_u2_rd_buf1_reg[30]/P0001  , \u1_u2_rd_buf1_reg[31]/P0001  , \u1_u2_rd_buf1_reg[3]/NET0131  , \u1_u2_rd_buf1_reg[4]/P0001  , \u1_u2_rd_buf1_reg[5]/P0001  , \u1_u2_rd_buf1_reg[6]/P0001  , \u1_u2_rd_buf1_reg[7]/P0001  , \u1_u2_rd_buf1_reg[8]/NET0131  , \u1_u2_rd_buf1_reg[9]/NET0131  , \u1_u2_rx_data_done_r2_reg/P0001  , \u1_u2_rx_data_done_r_reg/P0001  , \u1_u2_rx_data_st_r_reg[0]/P0001  , \u1_u2_rx_data_st_r_reg[1]/P0001  , \u1_u2_rx_data_st_r_reg[2]/P0001  , \u1_u2_rx_data_st_r_reg[3]/P0001  , \u1_u2_rx_data_st_r_reg[4]/P0001  , \u1_u2_rx_data_st_r_reg[5]/P0001  , \u1_u2_rx_data_st_r_reg[6]/P0001  , \u1_u2_rx_data_st_r_reg[7]/P0001  , \u1_u2_rx_data_valid_r_reg/NET0131  , \u1_u2_rx_dma_en_r_reg/P0001  , \u1_u2_send_data_r_reg/NET0131  , \u1_u2_sizd_c_reg[0]/P0001  , \u1_u2_sizd_c_reg[10]/P0001  , \u1_u2_sizd_c_reg[11]/P0001  , \u1_u2_sizd_c_reg[12]/P0001  , \u1_u2_sizd_c_reg[13]/P0001  , \u1_u2_sizd_c_reg[1]/P0001  , \u1_u2_sizd_c_reg[2]/P0001  , \u1_u2_sizd_c_reg[3]/P0001  , \u1_u2_sizd_c_reg[4]/P0001  , \u1_u2_sizd_c_reg[5]/P0001  , \u1_u2_sizd_c_reg[6]/P0001  , \u1_u2_sizd_c_reg[7]/P0001  , \u1_u2_sizd_c_reg[8]/P0001  , \u1_u2_sizd_c_reg[9]/P0001  , \u1_u2_sizd_is_zero_reg/P0001  , \u1_u2_sizu_c_reg[0]/P0001  , \u1_u2_sizu_c_reg[10]/P0001  , \u1_u2_sizu_c_reg[1]/P0001  , \u1_u2_sizu_c_reg[2]/P0001  , \u1_u2_sizu_c_reg[3]/P0001  , \u1_u2_sizu_c_reg[4]/P0001  , \u1_u2_sizu_c_reg[5]/P0001  , \u1_u2_sizu_c_reg[6]/P0001  , \u1_u2_sizu_c_reg[7]/P0001  , \u1_u2_sizu_c_reg[8]/NET0131  , \u1_u2_sizu_c_reg[9]/P0001  , \u1_u2_state_reg[0]/P0001  , \u1_u2_state_reg[1]/NET0131  , \u1_u2_state_reg[2]/NET0131  , \u1_u2_state_reg[3]/NET0131  , \u1_u2_state_reg[4]/NET0131  , \u1_u2_state_reg[5]/NET0131  , \u1_u2_state_reg[6]/NET0131  , \u1_u2_state_reg[7]/NET0131  , \u1_u2_tx_dma_en_r_reg/P0001  , \u1_u2_word_done_r_reg/P0001  , \u1_u2_word_done_reg/NET0131  , \u1_u2_wr_done_reg/P0001  , \u1_u2_wr_last_reg/P0001  , \u1_u3_abort_reg/P0001  , \u1_u3_adr_r_reg[0]/P0001  , \u1_u3_adr_r_reg[10]/P0001  , \u1_u3_adr_r_reg[11]/P0001  , \u1_u3_adr_r_reg[12]/P0001  , \u1_u3_adr_r_reg[13]/P0001  , \u1_u3_adr_r_reg[14]/P0001  , \u1_u3_adr_r_reg[15]/P0001  , \u1_u3_adr_r_reg[16]/P0001  , \u1_u3_adr_r_reg[1]/P0001  , \u1_u3_adr_r_reg[2]/P0001  , \u1_u3_adr_r_reg[3]/P0001  , \u1_u3_adr_r_reg[4]/P0001  , \u1_u3_adr_r_reg[5]/P0001  , \u1_u3_adr_r_reg[6]/P0001  , \u1_u3_adr_r_reg[7]/P0001  , \u1_u3_adr_r_reg[8]/P0001  , \u1_u3_adr_r_reg[9]/P0001  , \u1_u3_adr_reg[0]/P0001  , \u1_u3_adr_reg[10]/P0001  , \u1_u3_adr_reg[11]/P0001  , \u1_u3_adr_reg[12]/P0001  , \u1_u3_adr_reg[13]/P0001  , \u1_u3_adr_reg[14]/P0001  , \u1_u3_adr_reg[15]/P0001  , \u1_u3_adr_reg[16]/P0001  , \u1_u3_adr_reg[1]/P0001  , \u1_u3_adr_reg[2]/P0001  , \u1_u3_adr_reg[3]/P0001  , \u1_u3_adr_reg[4]/P0001  , \u1_u3_adr_reg[5]/P0001  , \u1_u3_adr_reg[6]/P0001  , \u1_u3_adr_reg[7]/P0001  , \u1_u3_adr_reg[8]/P0001  , \u1_u3_adr_reg[9]/P0001  , \u1_u3_buf0_na_reg/NET0131  , \u1_u3_buf0_not_aloc_reg/P0001  , \u1_u3_buf0_rl_reg/P0001  , \u1_u3_buf0_set_reg/P0001  , \u1_u3_buf0_st_max_reg/P0001  , \u1_u3_buf1_na_reg/NET0131  , \u1_u3_buf1_not_aloc_reg/P0001  , \u1_u3_buf1_set_reg/P0001  , \u1_u3_buf1_st_max_reg/P0001  , \u1_u3_buffer_done_reg/P0001  , \u1_u3_buffer_empty_reg/P0001  , \u1_u3_buffer_full_reg/P0001  , \u1_u3_buffer_overflow_reg/P0001  , \u1_u3_idin_reg[0]/P0001  , \u1_u3_idin_reg[10]/P0001  , \u1_u3_idin_reg[11]/P0001  , \u1_u3_idin_reg[12]/P0001  , \u1_u3_idin_reg[13]/P0001  , \u1_u3_idin_reg[14]/P0001  , \u1_u3_idin_reg[15]/P0001  , \u1_u3_idin_reg[16]/P0001  , \u1_u3_idin_reg[17]/P0001  , \u1_u3_idin_reg[18]/P0001  , \u1_u3_idin_reg[19]/P0001  , \u1_u3_idin_reg[1]/P0001  , \u1_u3_idin_reg[20]/P0001  , \u1_u3_idin_reg[21]/P0001  , \u1_u3_idin_reg[22]/P0001  , \u1_u3_idin_reg[23]/P0001  , \u1_u3_idin_reg[24]/P0001  , \u1_u3_idin_reg[25]/P0001  , \u1_u3_idin_reg[26]/P0001  , \u1_u3_idin_reg[27]/P0001  , \u1_u3_idin_reg[28]/P0001  , \u1_u3_idin_reg[29]/P0001  , \u1_u3_idin_reg[2]/P0001  , \u1_u3_idin_reg[30]/P0001  , \u1_u3_idin_reg[31]/P0001  , \u1_u3_idin_reg[3]/P0001  , \u1_u3_idin_reg[4]/P0001  , \u1_u3_idin_reg[5]/P0001  , \u1_u3_idin_reg[6]/P0001  , \u1_u3_idin_reg[7]/P0001  , \u1_u3_idin_reg[8]/P0001  , \u1_u3_idin_reg[9]/P0001  , \u1_u3_in_token_reg/NET0131  , \u1_u3_int_seqerr_set_reg/P0001  , \u1_u3_int_upid_set_reg/P0001  , \u1_u3_match_r_reg/P0001  , \u1_u3_new_size_reg[0]/P0001  , \u1_u3_new_size_reg[10]/P0001  , \u1_u3_new_size_reg[11]/P0001  , \u1_u3_new_size_reg[12]/P0001  , \u1_u3_new_size_reg[13]/P0001  , \u1_u3_new_size_reg[1]/P0001  , \u1_u3_new_size_reg[2]/P0001  , \u1_u3_new_size_reg[3]/P0001  , \u1_u3_new_size_reg[4]/P0001  , \u1_u3_new_size_reg[5]/P0001  , \u1_u3_new_size_reg[6]/P0001  , \u1_u3_new_size_reg[7]/P0001  , \u1_u3_new_size_reg[8]/P0001  , \u1_u3_new_size_reg[9]/P0001  , \u1_u3_new_sizeb_reg[0]/P0001  , \u1_u3_new_sizeb_reg[10]/P0001  , \u1_u3_new_sizeb_reg[1]/P0001  , \u1_u3_new_sizeb_reg[2]/P0001  , \u1_u3_new_sizeb_reg[3]/P0001  , \u1_u3_new_sizeb_reg[4]/P0001  , \u1_u3_new_sizeb_reg[5]/P0001  , \u1_u3_new_sizeb_reg[6]/P0001  , \u1_u3_new_sizeb_reg[7]/P0001  , \u1_u3_new_sizeb_reg[8]/P0001  , \u1_u3_new_sizeb_reg[9]/P0001  , \u1_u3_next_dpid_reg[0]/P0001  , \u1_u3_next_dpid_reg[1]/P0001  , \u1_u3_no_bufs0_reg/P0001  , \u1_u3_no_bufs1_reg/P0001  , \u1_u3_out_to_small_r_reg/P0001  , \u1_u3_out_to_small_reg/P0001  , \u1_u3_out_token_reg/NET0131  , \u1_u3_pid_IN_r_reg/P0001  , \u1_u3_pid_OUT_r_reg/P0001  , \u1_u3_pid_PING_r_reg/P0001  , \u1_u3_pid_SETUP_r_reg/P0001  , \u1_u3_pid_seq_err_reg/P0001  , \u1_u3_rx_ack_to_clr_reg/P0001  , \u1_u3_rx_ack_to_cnt_reg[0]/P0001  , \u1_u3_rx_ack_to_cnt_reg[1]/P0001  , \u1_u3_rx_ack_to_cnt_reg[2]/P0001  , \u1_u3_rx_ack_to_cnt_reg[3]/P0001  , \u1_u3_rx_ack_to_cnt_reg[4]/P0001  , \u1_u3_rx_ack_to_cnt_reg[5]/P0001  , \u1_u3_rx_ack_to_cnt_reg[6]/P0001  , \u1_u3_rx_ack_to_cnt_reg[7]/P0001  , \u1_u3_rx_ack_to_reg/P0001  , \u1_u3_send_token_reg/P0001  , \u1_u3_setup_token_reg/P0001  , \u1_u3_size_next_r_reg[0]/P0001  , \u1_u3_size_next_r_reg[10]/P0001  , \u1_u3_size_next_r_reg[1]/P0001  , \u1_u3_size_next_r_reg[2]/P0001  , \u1_u3_size_next_r_reg[3]/P0001  , \u1_u3_size_next_r_reg[4]/P0001  , \u1_u3_size_next_r_reg[5]/P0001  , \u1_u3_size_next_r_reg[6]/P0001  , \u1_u3_size_next_r_reg[7]/P0001  , \u1_u3_size_next_r_reg[8]/P0001  , \u1_u3_size_next_r_reg[9]/P0001  , \u1_u3_state_reg[0]/P0001  , \u1_u3_state_reg[1]/P0001  , \u1_u3_state_reg[2]/P0001  , \u1_u3_state_reg[3]/P0001  , \u1_u3_state_reg[4]/P0001  , \u1_u3_state_reg[5]/P0001  , \u1_u3_state_reg[6]/P0001  , \u1_u3_state_reg[7]/P0001  , \u1_u3_state_reg[8]/P0001  , \u1_u3_state_reg[9]/P0001  , \u1_u3_this_dpid_reg[0]/P0001  , \u1_u3_this_dpid_reg[1]/P0001  , \u1_u3_to_large_reg/P0001  , \u1_u3_to_small_reg/P0001  , \u1_u3_token_pid_sel_reg[0]/P0001  , \u1_u3_token_pid_sel_reg[1]/P0001  , \u1_u3_tx_data_to_cnt_reg[0]/P0001  , \u1_u3_tx_data_to_cnt_reg[1]/P0001  , \u1_u3_tx_data_to_cnt_reg[2]/P0001  , \u1_u3_tx_data_to_cnt_reg[3]/P0001  , \u1_u3_tx_data_to_cnt_reg[4]/P0001  , \u1_u3_tx_data_to_cnt_reg[5]/P0001  , \u1_u3_tx_data_to_cnt_reg[6]/P0001  , \u1_u3_tx_data_to_cnt_reg[7]/P0001  , \u1_u3_tx_data_to_reg/P0001  , \u1_u3_uc_bsel_set_reg/P0001  , \u2_wack_r_reg/P0001  , \u4_attach_r1_reg/P0001  , \u4_attach_r_reg/P0001  , \u4_buf0_reg[0]/P0001  , \u4_buf0_reg[10]/P0001  , \u4_buf0_reg[11]/P0001  , \u4_buf0_reg[12]/P0001  , \u4_buf0_reg[13]/P0001  , \u4_buf0_reg[14]/P0001  , \u4_buf0_reg[15]/P0001  , \u4_buf0_reg[16]/P0001  , \u4_buf0_reg[17]/NET0131  , \u4_buf0_reg[18]/P0001  , \u4_buf0_reg[19]/NET0131  , \u4_buf0_reg[1]/P0001  , \u4_buf0_reg[20]/NET0131  , \u4_buf0_reg[21]/NET0131  , \u4_buf0_reg[22]/NET0131  , \u4_buf0_reg[23]/NET0131  , \u4_buf0_reg[24]/NET0131  , \u4_buf0_reg[25]/NET0131  , \u4_buf0_reg[26]/NET0131  , \u4_buf0_reg[27]/P0001  , \u4_buf0_reg[28]/P0001  , \u4_buf0_reg[29]/P0001  , \u4_buf0_reg[2]/P0001  , \u4_buf0_reg[30]/P0001  , \u4_buf0_reg[31]/P0001  , \u4_buf0_reg[3]/P0001  , \u4_buf0_reg[4]/P0001  , \u4_buf0_reg[5]/P0001  , \u4_buf0_reg[6]/P0001  , \u4_buf0_reg[7]/P0001  , \u4_buf0_reg[8]/P0001  , \u4_buf0_reg[9]/P0001  , \u4_buf1_reg[0]/P0001  , \u4_buf1_reg[10]/P0001  , \u4_buf1_reg[11]/P0001  , \u4_buf1_reg[12]/P0001  , \u4_buf1_reg[13]/P0001  , \u4_buf1_reg[14]/P0001  , \u4_buf1_reg[15]/P0001  , \u4_buf1_reg[16]/P0001  , \u4_buf1_reg[17]/NET0131  , \u4_buf1_reg[18]/P0001  , \u4_buf1_reg[19]/NET0131  , \u4_buf1_reg[1]/P0001  , \u4_buf1_reg[20]/NET0131  , \u4_buf1_reg[21]/NET0131  , \u4_buf1_reg[22]/NET0131  , \u4_buf1_reg[23]/NET0131  , \u4_buf1_reg[24]/NET0131  , \u4_buf1_reg[25]/NET0131  , \u4_buf1_reg[26]/NET0131  , \u4_buf1_reg[27]/P0001  , \u4_buf1_reg[28]/P0001  , \u4_buf1_reg[29]/P0001  , \u4_buf1_reg[2]/P0001  , \u4_buf1_reg[30]/P0001  , \u4_buf1_reg[31]/P0001  , \u4_buf1_reg[3]/P0001  , \u4_buf1_reg[4]/P0001  , \u4_buf1_reg[5]/P0001  , \u4_buf1_reg[6]/P0001  , \u4_buf1_reg[7]/P0001  , \u4_buf1_reg[8]/P0001  , \u4_buf1_reg[9]/P0001  , \u4_crc5_err_r_reg/P0001  , \u4_csr_reg[0]/P0001  , \u4_csr_reg[10]/P0001  , \u4_csr_reg[11]/P0001  , \u4_csr_reg[12]/P0001  , \u4_csr_reg[15]/NET0131  , \u4_csr_reg[16]/P0001  , \u4_csr_reg[17]/P0001  , \u4_csr_reg[1]/P0001  , \u4_csr_reg[22]/P0001  , \u4_csr_reg[23]/P0001  , \u4_csr_reg[24]/P0001  , \u4_csr_reg[25]/P0001  , \u4_csr_reg[26]/NET0131  , \u4_csr_reg[27]/NET0131  , \u4_csr_reg[28]/P0001  , \u4_csr_reg[29]/P0001  , \u4_csr_reg[2]/NET0131  , \u4_csr_reg[30]/NET0131  , \u4_csr_reg[31]/P0001  , \u4_csr_reg[3]/P0001  , \u4_csr_reg[4]/NET0131  , \u4_csr_reg[5]/NET0131  , \u4_csr_reg[6]/NET0131  , \u4_csr_reg[7]/P0001  , \u4_csr_reg[8]/P0001  , \u4_csr_reg[9]/NET0131  , \u4_dma_in_buf_sz1_reg/P0001  , \u4_dma_out_buf_avail_reg/P0001  , \u4_dout_reg[0]/P0001  , \u4_dout_reg[10]/P0001  , \u4_dout_reg[11]/P0001  , \u4_dout_reg[12]/P0001  , \u4_dout_reg[13]/P0001  , \u4_dout_reg[14]/P0001  , \u4_dout_reg[15]/P0001  , \u4_dout_reg[16]/P0001  , \u4_dout_reg[17]/P0001  , \u4_dout_reg[18]/P0001  , \u4_dout_reg[19]/P0001  , \u4_dout_reg[1]/P0001  , \u4_dout_reg[20]/P0001  , \u4_dout_reg[21]/P0001  , \u4_dout_reg[22]/P0001  , \u4_dout_reg[23]/P0001  , \u4_dout_reg[24]/P0001  , \u4_dout_reg[25]/P0001  , \u4_dout_reg[26]/P0001  , \u4_dout_reg[27]/P0001  , \u4_dout_reg[28]/P0001  , \u4_dout_reg[29]/P0001  , \u4_dout_reg[2]/P0001  , \u4_dout_reg[30]/P0001  , \u4_dout_reg[31]/P0001  , \u4_dout_reg[3]/P0001  , \u4_dout_reg[4]/P0001  , \u4_dout_reg[5]/P0001  , \u4_dout_reg[6]/P0001  , \u4_dout_reg[7]/P0001  , \u4_dout_reg[8]/P0001  , \u4_dout_reg[9]/P0001  , \u4_funct_adr_reg[0]/P0001  , \u4_funct_adr_reg[1]/P0001  , \u4_funct_adr_reg[2]/P0001  , \u4_funct_adr_reg[3]/P0001  , \u4_funct_adr_reg[4]/P0001  , \u4_funct_adr_reg[5]/P0001  , \u4_funct_adr_reg[6]/P0001  , \u4_int_src_re_reg/P0001  , \u4_int_srca_reg[0]/P0001  , \u4_int_srca_reg[1]/P0001  , \u4_int_srca_reg[2]/P0001  , \u4_int_srca_reg[3]/P0001  , \u4_int_srcb_reg[0]/P0001  , \u4_int_srcb_reg[1]/P0001  , \u4_int_srcb_reg[2]/P0001  , \u4_int_srcb_reg[3]/P0001  , \u4_int_srcb_reg[4]/P0001  , \u4_int_srcb_reg[5]/P0001  , \u4_int_srcb_reg[6]/P0001  , \u4_int_srcb_reg[7]/P0001  , \u4_int_srcb_reg[8]/P0001  , \u4_inta_msk_reg[0]/P0001  , \u4_inta_msk_reg[1]/P0001  , \u4_inta_msk_reg[2]/P0001  , \u4_inta_msk_reg[3]/P0001  , \u4_inta_msk_reg[4]/P0001  , \u4_inta_msk_reg[5]/P0001  , \u4_inta_msk_reg[6]/P0001  , \u4_inta_msk_reg[7]/P0001  , \u4_inta_msk_reg[8]/P0001  , \u4_intb_msk_reg[0]/P0001  , \u4_intb_msk_reg[1]/P0001  , \u4_intb_msk_reg[2]/P0001  , \u4_intb_msk_reg[3]/P0001  , \u4_intb_msk_reg[4]/P0001  , \u4_intb_msk_reg[5]/P0001  , \u4_intb_msk_reg[6]/P0001  , \u4_intb_msk_reg[7]/P0001  , \u4_intb_msk_reg[8]/P0001  , \u4_match_r1_reg/P0001  , \u4_nse_err_r_reg/P0001  , \u4_pid_cs_err_r_reg/P0001  , \u4_rx_err_r_reg/P0001  , \u4_suspend_r1_reg/P0001  , \u4_u0_buf0_orig_m3_reg[0]/P0001  , \u4_u0_buf0_orig_m3_reg[10]/P0001  , \u4_u0_buf0_orig_m3_reg[11]/P0001  , \u4_u0_buf0_orig_m3_reg[1]/P0001  , \u4_u0_buf0_orig_m3_reg[2]/P0001  , \u4_u0_buf0_orig_m3_reg[3]/P0001  , \u4_u0_buf0_orig_m3_reg[4]/P0001  , \u4_u0_buf0_orig_m3_reg[5]/P0001  , \u4_u0_buf0_orig_m3_reg[6]/P0001  , \u4_u0_buf0_orig_m3_reg[7]/P0001  , \u4_u0_buf0_orig_m3_reg[8]/P0001  , \u4_u0_buf0_orig_m3_reg[9]/P0001  , \u4_u0_buf0_orig_reg[0]/P0001  , \u4_u0_buf0_orig_reg[10]/P0001  , \u4_u0_buf0_orig_reg[11]/P0001  , \u4_u0_buf0_orig_reg[12]/P0001  , \u4_u0_buf0_orig_reg[13]/P0001  , \u4_u0_buf0_orig_reg[14]/P0001  , \u4_u0_buf0_orig_reg[15]/P0001  , \u4_u0_buf0_orig_reg[16]/P0001  , \u4_u0_buf0_orig_reg[17]/P0001  , \u4_u0_buf0_orig_reg[18]/P0001  , \u4_u0_buf0_orig_reg[19]/P0001  , \u4_u0_buf0_orig_reg[1]/P0001  , \u4_u0_buf0_orig_reg[20]/P0001  , \u4_u0_buf0_orig_reg[21]/P0001  , \u4_u0_buf0_orig_reg[22]/P0001  , \u4_u0_buf0_orig_reg[23]/P0001  , \u4_u0_buf0_orig_reg[24]/P0001  , \u4_u0_buf0_orig_reg[25]/P0001  , \u4_u0_buf0_orig_reg[26]/P0001  , \u4_u0_buf0_orig_reg[27]/P0001  , \u4_u0_buf0_orig_reg[28]/P0001  , \u4_u0_buf0_orig_reg[29]/NET0131  , \u4_u0_buf0_orig_reg[2]/P0001  , \u4_u0_buf0_orig_reg[30]/NET0131  , \u4_u0_buf0_orig_reg[31]/P0001  , \u4_u0_buf0_orig_reg[3]/P0001  , \u4_u0_buf0_orig_reg[4]/P0001  , \u4_u0_buf0_orig_reg[5]/P0001  , \u4_u0_buf0_orig_reg[6]/P0001  , \u4_u0_buf0_orig_reg[7]/P0001  , \u4_u0_buf0_orig_reg[8]/P0001  , \u4_u0_buf0_orig_reg[9]/P0001  , \u4_u0_buf0_reg[0]/P0001  , \u4_u0_buf0_reg[10]/P0001  , \u4_u0_buf0_reg[11]/P0001  , \u4_u0_buf0_reg[12]/P0001  , \u4_u0_buf0_reg[13]/P0001  , \u4_u0_buf0_reg[14]/P0001  , \u4_u0_buf0_reg[15]/P0001  , \u4_u0_buf0_reg[16]/P0001  , \u4_u0_buf0_reg[17]/P0001  , \u4_u0_buf0_reg[18]/P0001  , \u4_u0_buf0_reg[19]/P0001  , \u4_u0_buf0_reg[1]/P0001  , \u4_u0_buf0_reg[20]/P0001  , \u4_u0_buf0_reg[21]/P0001  , \u4_u0_buf0_reg[22]/P0001  , \u4_u0_buf0_reg[23]/P0001  , \u4_u0_buf0_reg[24]/P0001  , \u4_u0_buf0_reg[25]/P0001  , \u4_u0_buf0_reg[26]/P0001  , \u4_u0_buf0_reg[27]/P0001  , \u4_u0_buf0_reg[28]/P0001  , \u4_u0_buf0_reg[29]/P0001  , \u4_u0_buf0_reg[2]/P0001  , \u4_u0_buf0_reg[30]/P0001  , \u4_u0_buf0_reg[31]/P0001  , \u4_u0_buf0_reg[3]/P0001  , \u4_u0_buf0_reg[4]/P0001  , \u4_u0_buf0_reg[5]/P0001  , \u4_u0_buf0_reg[6]/P0001  , \u4_u0_buf0_reg[7]/P0001  , \u4_u0_buf0_reg[8]/P0001  , \u4_u0_buf0_reg[9]/P0001  , \u4_u0_buf1_reg[0]/P0001  , \u4_u0_buf1_reg[10]/P0001  , \u4_u0_buf1_reg[11]/P0001  , \u4_u0_buf1_reg[12]/P0001  , \u4_u0_buf1_reg[13]/P0001  , \u4_u0_buf1_reg[14]/P0001  , \u4_u0_buf1_reg[15]/P0001  , \u4_u0_buf1_reg[16]/P0001  , \u4_u0_buf1_reg[17]/P0001  , \u4_u0_buf1_reg[18]/P0001  , \u4_u0_buf1_reg[19]/P0001  , \u4_u0_buf1_reg[1]/P0001  , \u4_u0_buf1_reg[20]/P0001  , \u4_u0_buf1_reg[21]/P0001  , \u4_u0_buf1_reg[22]/P0001  , \u4_u0_buf1_reg[23]/P0001  , \u4_u0_buf1_reg[24]/P0001  , \u4_u0_buf1_reg[25]/P0001  , \u4_u0_buf1_reg[26]/P0001  , \u4_u0_buf1_reg[27]/P0001  , \u4_u0_buf1_reg[28]/P0001  , \u4_u0_buf1_reg[29]/P0001  , \u4_u0_buf1_reg[2]/P0001  , \u4_u0_buf1_reg[30]/P0001  , \u4_u0_buf1_reg[31]/P0001  , \u4_u0_buf1_reg[3]/P0001  , \u4_u0_buf1_reg[4]/P0001  , \u4_u0_buf1_reg[5]/P0001  , \u4_u0_buf1_reg[6]/P0001  , \u4_u0_buf1_reg[7]/P0001  , \u4_u0_buf1_reg[8]/P0001  , \u4_u0_buf1_reg[9]/P0001  , \u4_u0_csr0_reg[0]/P0001  , \u4_u0_csr0_reg[10]/P0001  , \u4_u0_csr0_reg[11]/P0001  , \u4_u0_csr0_reg[12]/P0001  , \u4_u0_csr0_reg[1]/P0001  , \u4_u0_csr0_reg[2]/P0001  , \u4_u0_csr0_reg[3]/NET0131  , \u4_u0_csr0_reg[4]/P0001  , \u4_u0_csr0_reg[5]/P0001  , \u4_u0_csr0_reg[6]/P0001  , \u4_u0_csr0_reg[7]/P0001  , \u4_u0_csr0_reg[8]/P0001  , \u4_u0_csr0_reg[9]/P0001  , \u4_u0_csr1_reg[0]/P0001  , \u4_u0_csr1_reg[10]/P0001  , \u4_u0_csr1_reg[11]/P0001  , \u4_u0_csr1_reg[12]/P0001  , \u4_u0_csr1_reg[1]/P0001  , \u4_u0_csr1_reg[2]/P0001  , \u4_u0_csr1_reg[3]/P0001  , \u4_u0_csr1_reg[4]/P0001  , \u4_u0_csr1_reg[5]/P0001  , \u4_u0_csr1_reg[6]/P0001  , \u4_u0_csr1_reg[7]/P0001  , \u4_u0_csr1_reg[8]/P0001  , \u4_u0_csr1_reg[9]/P0001  , \u4_u0_dma_ack_clr1_reg/P0001  , \u4_u0_dma_ack_wr1_reg/P0001  , \u4_u0_dma_in_buf_sz1_reg/P0001  , \u4_u0_dma_in_cnt_reg[0]/P0001  , \u4_u0_dma_in_cnt_reg[10]/P0001  , \u4_u0_dma_in_cnt_reg[11]/P0001  , \u4_u0_dma_in_cnt_reg[1]/P0001  , \u4_u0_dma_in_cnt_reg[2]/P0001  , \u4_u0_dma_in_cnt_reg[3]/P0001  , \u4_u0_dma_in_cnt_reg[4]/P0001  , \u4_u0_dma_in_cnt_reg[5]/P0001  , \u4_u0_dma_in_cnt_reg[6]/P0001  , \u4_u0_dma_in_cnt_reg[7]/P0001  , \u4_u0_dma_in_cnt_reg[8]/P0001  , \u4_u0_dma_in_cnt_reg[9]/P0001  , \u4_u0_dma_out_buf_avail_reg/P0001  , \u4_u0_dma_out_cnt_reg[10]/P0001  , \u4_u0_dma_out_cnt_reg[11]/P0001  , \u4_u0_dma_out_cnt_reg[1]/P0001  , \u4_u0_dma_out_cnt_reg[2]/P0001  , \u4_u0_dma_out_cnt_reg[3]/P0001  , \u4_u0_dma_out_cnt_reg[4]/P0001  , \u4_u0_dma_out_cnt_reg[5]/P0001  , \u4_u0_dma_out_cnt_reg[6]/P0001  , \u4_u0_dma_out_cnt_reg[7]/P0001  , \u4_u0_dma_out_cnt_reg[8]/P0001  , \u4_u0_dma_out_cnt_reg[9]/P0001  , \u4_u0_dma_out_left_reg[0]/P0001  , \u4_u0_dma_out_left_reg[10]/P0001  , \u4_u0_dma_out_left_reg[11]/P0001  , \u4_u0_dma_out_left_reg[1]/P0001  , \u4_u0_dma_out_left_reg[2]/P0001  , \u4_u0_dma_out_left_reg[3]/P0001  , \u4_u0_dma_out_left_reg[4]/P0001  , \u4_u0_dma_out_left_reg[5]/P0001  , \u4_u0_dma_out_left_reg[6]/P0001  , \u4_u0_dma_out_left_reg[7]/P0001  , \u4_u0_dma_out_left_reg[8]/P0001  , \u4_u0_dma_out_left_reg[9]/P0001  , \u4_u0_dma_req_in_hold2_reg/P0001  , \u4_u0_dma_req_in_hold_reg/P0001  , \u4_u0_dma_req_out_hold_reg/P0001  , \u4_u0_ep_match_r_reg/P0001  , \u4_u0_iena_reg[0]/P0001  , \u4_u0_iena_reg[1]/P0001  , \u4_u0_iena_reg[2]/P0001  , \u4_u0_iena_reg[3]/P0001  , \u4_u0_iena_reg[4]/P0001  , \u4_u0_iena_reg[5]/P0001  , \u4_u0_ienb_reg[0]/P0001  , \u4_u0_ienb_reg[1]/P0001  , \u4_u0_ienb_reg[2]/P0001  , \u4_u0_ienb_reg[3]/P0001  , \u4_u0_ienb_reg[4]/P0001  , \u4_u0_ienb_reg[5]/P0001  , \u4_u0_int_re_reg/P0001  , \u4_u0_int_stat_reg[0]/P0001  , \u4_u0_int_stat_reg[1]/P0001  , \u4_u0_int_stat_reg[2]/P0001  , \u4_u0_int_stat_reg[3]/P0001  , \u4_u0_int_stat_reg[4]/P0001  , \u4_u0_int_stat_reg[5]/P0001  , \u4_u0_int_stat_reg[6]/P0001  , \u4_u0_inta_reg/P0001  , \u4_u0_intb_reg/P0001  , \u4_u0_ots_stop_reg/P0001  , \u4_u0_r1_reg/P0001  , \u4_u0_r2_reg/P0001  , \u4_u0_r4_reg/P0001  , \u4_u0_r5_reg/NET0131  , \u4_u0_set_r_reg/P0001  , \u4_u0_uc_bsel_reg[0]/P0001  , \u4_u0_uc_bsel_reg[1]/P0001  , \u4_u0_uc_dpd_reg[0]/P0001  , \u4_u0_uc_dpd_reg[1]/P0001  , \u4_u1_buf0_orig_m3_reg[0]/P0001  , \u4_u1_buf0_orig_m3_reg[10]/P0001  , \u4_u1_buf0_orig_m3_reg[11]/P0001  , \u4_u1_buf0_orig_m3_reg[1]/P0001  , \u4_u1_buf0_orig_m3_reg[2]/P0001  , \u4_u1_buf0_orig_m3_reg[3]/P0001  , \u4_u1_buf0_orig_m3_reg[4]/P0001  , \u4_u1_buf0_orig_m3_reg[5]/P0001  , \u4_u1_buf0_orig_m3_reg[6]/P0001  , \u4_u1_buf0_orig_m3_reg[7]/P0001  , \u4_u1_buf0_orig_m3_reg[8]/P0001  , \u4_u1_buf0_orig_m3_reg[9]/P0001  , \u4_u1_buf0_orig_reg[0]/P0001  , \u4_u1_buf0_orig_reg[10]/P0001  , \u4_u1_buf0_orig_reg[11]/P0001  , \u4_u1_buf0_orig_reg[12]/P0001  , \u4_u1_buf0_orig_reg[13]/P0001  , \u4_u1_buf0_orig_reg[14]/P0001  , \u4_u1_buf0_orig_reg[15]/P0001  , \u4_u1_buf0_orig_reg[16]/P0001  , \u4_u1_buf0_orig_reg[17]/P0001  , \u4_u1_buf0_orig_reg[18]/P0001  , \u4_u1_buf0_orig_reg[19]/P0001  , \u4_u1_buf0_orig_reg[1]/P0001  , \u4_u1_buf0_orig_reg[20]/P0001  , \u4_u1_buf0_orig_reg[21]/P0001  , \u4_u1_buf0_orig_reg[22]/P0001  , \u4_u1_buf0_orig_reg[23]/P0001  , \u4_u1_buf0_orig_reg[24]/P0001  , \u4_u1_buf0_orig_reg[25]/P0001  , \u4_u1_buf0_orig_reg[26]/P0001  , \u4_u1_buf0_orig_reg[27]/P0001  , \u4_u1_buf0_orig_reg[28]/P0001  , \u4_u1_buf0_orig_reg[29]/NET0131  , \u4_u1_buf0_orig_reg[2]/P0001  , \u4_u1_buf0_orig_reg[30]/NET0131  , \u4_u1_buf0_orig_reg[31]/P0001  , \u4_u1_buf0_orig_reg[3]/P0001  , \u4_u1_buf0_orig_reg[4]/P0001  , \u4_u1_buf0_orig_reg[5]/P0001  , \u4_u1_buf0_orig_reg[6]/P0001  , \u4_u1_buf0_orig_reg[7]/P0001  , \u4_u1_buf0_orig_reg[8]/P0001  , \u4_u1_buf0_orig_reg[9]/P0001  , \u4_u1_buf0_reg[0]/P0001  , \u4_u1_buf0_reg[10]/P0001  , \u4_u1_buf0_reg[11]/P0001  , \u4_u1_buf0_reg[12]/P0001  , \u4_u1_buf0_reg[13]/P0001  , \u4_u1_buf0_reg[14]/P0001  , \u4_u1_buf0_reg[15]/P0001  , \u4_u1_buf0_reg[16]/P0001  , \u4_u1_buf0_reg[17]/P0001  , \u4_u1_buf0_reg[18]/P0001  , \u4_u1_buf0_reg[19]/P0001  , \u4_u1_buf0_reg[1]/P0001  , \u4_u1_buf0_reg[20]/P0001  , \u4_u1_buf0_reg[21]/P0001  , \u4_u1_buf0_reg[22]/P0001  , \u4_u1_buf0_reg[23]/P0001  , \u4_u1_buf0_reg[24]/P0001  , \u4_u1_buf0_reg[25]/P0001  , \u4_u1_buf0_reg[26]/P0001  , \u4_u1_buf0_reg[27]/P0001  , \u4_u1_buf0_reg[28]/P0001  , \u4_u1_buf0_reg[29]/P0001  , \u4_u1_buf0_reg[2]/P0001  , \u4_u1_buf0_reg[30]/P0001  , \u4_u1_buf0_reg[31]/P0001  , \u4_u1_buf0_reg[3]/P0001  , \u4_u1_buf0_reg[4]/P0001  , \u4_u1_buf0_reg[5]/P0001  , \u4_u1_buf0_reg[6]/P0001  , \u4_u1_buf0_reg[7]/P0001  , \u4_u1_buf0_reg[8]/P0001  , \u4_u1_buf0_reg[9]/P0001  , \u4_u1_buf1_reg[0]/P0001  , \u4_u1_buf1_reg[10]/P0001  , \u4_u1_buf1_reg[11]/P0001  , \u4_u1_buf1_reg[12]/P0001  , \u4_u1_buf1_reg[13]/P0001  , \u4_u1_buf1_reg[14]/P0001  , \u4_u1_buf1_reg[15]/P0001  , \u4_u1_buf1_reg[16]/P0001  , \u4_u1_buf1_reg[17]/P0001  , \u4_u1_buf1_reg[18]/P0001  , \u4_u1_buf1_reg[19]/P0001  , \u4_u1_buf1_reg[1]/P0001  , \u4_u1_buf1_reg[20]/P0001  , \u4_u1_buf1_reg[21]/P0001  , \u4_u1_buf1_reg[22]/P0001  , \u4_u1_buf1_reg[23]/P0001  , \u4_u1_buf1_reg[24]/P0001  , \u4_u1_buf1_reg[25]/P0001  , \u4_u1_buf1_reg[26]/P0001  , \u4_u1_buf1_reg[27]/P0001  , \u4_u1_buf1_reg[28]/P0001  , \u4_u1_buf1_reg[29]/P0001  , \u4_u1_buf1_reg[2]/P0001  , \u4_u1_buf1_reg[30]/P0001  , \u4_u1_buf1_reg[31]/P0001  , \u4_u1_buf1_reg[3]/P0001  , \u4_u1_buf1_reg[4]/P0001  , \u4_u1_buf1_reg[5]/P0001  , \u4_u1_buf1_reg[6]/P0001  , \u4_u1_buf1_reg[7]/P0001  , \u4_u1_buf1_reg[8]/P0001  , \u4_u1_buf1_reg[9]/P0001  , \u4_u1_csr0_reg[0]/P0001  , \u4_u1_csr0_reg[10]/P0001  , \u4_u1_csr0_reg[11]/P0001  , \u4_u1_csr0_reg[12]/P0001  , \u4_u1_csr0_reg[1]/P0001  , \u4_u1_csr0_reg[2]/P0001  , \u4_u1_csr0_reg[3]/NET0131  , \u4_u1_csr0_reg[4]/P0001  , \u4_u1_csr0_reg[5]/P0001  , \u4_u1_csr0_reg[6]/P0001  , \u4_u1_csr0_reg[7]/P0001  , \u4_u1_csr0_reg[8]/P0001  , \u4_u1_csr0_reg[9]/P0001  , \u4_u1_csr1_reg[0]/P0001  , \u4_u1_csr1_reg[10]/P0001  , \u4_u1_csr1_reg[11]/P0001  , \u4_u1_csr1_reg[12]/P0001  , \u4_u1_csr1_reg[1]/P0001  , \u4_u1_csr1_reg[2]/P0001  , \u4_u1_csr1_reg[3]/P0001  , \u4_u1_csr1_reg[4]/P0001  , \u4_u1_csr1_reg[5]/P0001  , \u4_u1_csr1_reg[6]/P0001  , \u4_u1_csr1_reg[7]/P0001  , \u4_u1_csr1_reg[8]/P0001  , \u4_u1_csr1_reg[9]/P0001  , \u4_u1_dma_ack_clr1_reg/P0001  , \u4_u1_dma_ack_wr1_reg/P0001  , \u4_u1_dma_in_buf_sz1_reg/P0001  , \u4_u1_dma_in_cnt_reg[0]/P0001  , \u4_u1_dma_in_cnt_reg[10]/P0001  , \u4_u1_dma_in_cnt_reg[11]/P0001  , \u4_u1_dma_in_cnt_reg[1]/P0001  , \u4_u1_dma_in_cnt_reg[2]/P0001  , \u4_u1_dma_in_cnt_reg[3]/P0001  , \u4_u1_dma_in_cnt_reg[4]/P0001  , \u4_u1_dma_in_cnt_reg[5]/P0001  , \u4_u1_dma_in_cnt_reg[6]/P0001  , \u4_u1_dma_in_cnt_reg[7]/P0001  , \u4_u1_dma_in_cnt_reg[8]/P0001  , \u4_u1_dma_in_cnt_reg[9]/P0001  , \u4_u1_dma_out_buf_avail_reg/P0001  , \u4_u1_dma_out_cnt_reg[10]/P0001  , \u4_u1_dma_out_cnt_reg[11]/P0001  , \u4_u1_dma_out_cnt_reg[1]/P0001  , \u4_u1_dma_out_cnt_reg[2]/P0001  , \u4_u1_dma_out_cnt_reg[3]/P0001  , \u4_u1_dma_out_cnt_reg[4]/P0001  , \u4_u1_dma_out_cnt_reg[5]/P0001  , \u4_u1_dma_out_cnt_reg[6]/P0001  , \u4_u1_dma_out_cnt_reg[7]/P0001  , \u4_u1_dma_out_cnt_reg[8]/P0001  , \u4_u1_dma_out_cnt_reg[9]/P0001  , \u4_u1_dma_out_left_reg[0]/P0001  , \u4_u1_dma_out_left_reg[10]/P0001  , \u4_u1_dma_out_left_reg[11]/P0001  , \u4_u1_dma_out_left_reg[1]/P0001  , \u4_u1_dma_out_left_reg[2]/P0001  , \u4_u1_dma_out_left_reg[3]/P0001  , \u4_u1_dma_out_left_reg[4]/P0001  , \u4_u1_dma_out_left_reg[5]/P0001  , \u4_u1_dma_out_left_reg[6]/P0001  , \u4_u1_dma_out_left_reg[7]/P0001  , \u4_u1_dma_out_left_reg[8]/P0001  , \u4_u1_dma_out_left_reg[9]/P0001  , \u4_u1_dma_req_in_hold2_reg/P0001  , \u4_u1_dma_req_in_hold_reg/P0001  , \u4_u1_dma_req_out_hold_reg/P0001  , \u4_u1_ep_match_r_reg/P0001  , \u4_u1_iena_reg[0]/P0001  , \u4_u1_iena_reg[1]/P0001  , \u4_u1_iena_reg[2]/P0001  , \u4_u1_iena_reg[3]/P0001  , \u4_u1_iena_reg[4]/P0001  , \u4_u1_iena_reg[5]/P0001  , \u4_u1_ienb_reg[0]/P0001  , \u4_u1_ienb_reg[1]/P0001  , \u4_u1_ienb_reg[2]/P0001  , \u4_u1_ienb_reg[3]/P0001  , \u4_u1_ienb_reg[4]/P0001  , \u4_u1_ienb_reg[5]/P0001  , \u4_u1_int_re_reg/P0001  , \u4_u1_int_stat_reg[0]/P0001  , \u4_u1_int_stat_reg[1]/P0001  , \u4_u1_int_stat_reg[2]/P0001  , \u4_u1_int_stat_reg[3]/P0001  , \u4_u1_int_stat_reg[4]/P0001  , \u4_u1_int_stat_reg[5]/P0001  , \u4_u1_int_stat_reg[6]/P0001  , \u4_u1_inta_reg/P0001  , \u4_u1_intb_reg/P0001  , \u4_u1_ots_stop_reg/P0001  , \u4_u1_r1_reg/P0001  , \u4_u1_r2_reg/P0001  , \u4_u1_r4_reg/P0001  , \u4_u1_r5_reg/NET0131  , \u4_u1_set_r_reg/P0001  , \u4_u1_uc_bsel_reg[0]/P0001  , \u4_u1_uc_bsel_reg[1]/P0001  , \u4_u1_uc_dpd_reg[0]/P0001  , \u4_u1_uc_dpd_reg[1]/P0001  , \u4_u2_buf0_orig_m3_reg[0]/P0001  , \u4_u2_buf0_orig_m3_reg[10]/P0001  , \u4_u2_buf0_orig_m3_reg[11]/P0001  , \u4_u2_buf0_orig_m3_reg[1]/P0001  , \u4_u2_buf0_orig_m3_reg[2]/P0001  , \u4_u2_buf0_orig_m3_reg[3]/P0001  , \u4_u2_buf0_orig_m3_reg[4]/P0001  , \u4_u2_buf0_orig_m3_reg[5]/P0001  , \u4_u2_buf0_orig_m3_reg[6]/P0001  , \u4_u2_buf0_orig_m3_reg[7]/P0001  , \u4_u2_buf0_orig_m3_reg[8]/P0001  , \u4_u2_buf0_orig_m3_reg[9]/P0001  , \u4_u2_buf0_orig_reg[0]/P0001  , \u4_u2_buf0_orig_reg[10]/P0001  , \u4_u2_buf0_orig_reg[11]/P0001  , \u4_u2_buf0_orig_reg[12]/P0001  , \u4_u2_buf0_orig_reg[13]/P0001  , \u4_u2_buf0_orig_reg[14]/P0001  , \u4_u2_buf0_orig_reg[15]/P0001  , \u4_u2_buf0_orig_reg[16]/P0001  , \u4_u2_buf0_orig_reg[17]/P0001  , \u4_u2_buf0_orig_reg[18]/P0001  , \u4_u2_buf0_orig_reg[19]/P0001  , \u4_u2_buf0_orig_reg[1]/P0001  , \u4_u2_buf0_orig_reg[20]/P0001  , \u4_u2_buf0_orig_reg[21]/P0001  , \u4_u2_buf0_orig_reg[22]/P0001  , \u4_u2_buf0_orig_reg[23]/P0001  , \u4_u2_buf0_orig_reg[24]/P0001  , \u4_u2_buf0_orig_reg[25]/P0001  , \u4_u2_buf0_orig_reg[26]/P0001  , \u4_u2_buf0_orig_reg[27]/P0001  , \u4_u2_buf0_orig_reg[28]/P0001  , \u4_u2_buf0_orig_reg[29]/NET0131  , \u4_u2_buf0_orig_reg[2]/P0001  , \u4_u2_buf0_orig_reg[30]/NET0131  , \u4_u2_buf0_orig_reg[31]/P0001  , \u4_u2_buf0_orig_reg[3]/P0001  , \u4_u2_buf0_orig_reg[4]/P0001  , \u4_u2_buf0_orig_reg[5]/P0001  , \u4_u2_buf0_orig_reg[6]/P0001  , \u4_u2_buf0_orig_reg[7]/P0001  , \u4_u2_buf0_orig_reg[8]/P0001  , \u4_u2_buf0_orig_reg[9]/P0001  , \u4_u2_buf0_reg[0]/P0001  , \u4_u2_buf0_reg[10]/P0001  , \u4_u2_buf0_reg[11]/P0001  , \u4_u2_buf0_reg[12]/P0001  , \u4_u2_buf0_reg[13]/P0001  , \u4_u2_buf0_reg[14]/P0001  , \u4_u2_buf0_reg[15]/P0001  , \u4_u2_buf0_reg[16]/P0001  , \u4_u2_buf0_reg[17]/P0001  , \u4_u2_buf0_reg[18]/P0001  , \u4_u2_buf0_reg[19]/P0001  , \u4_u2_buf0_reg[1]/P0001  , \u4_u2_buf0_reg[20]/P0001  , \u4_u2_buf0_reg[21]/P0001  , \u4_u2_buf0_reg[22]/P0001  , \u4_u2_buf0_reg[23]/P0001  , \u4_u2_buf0_reg[24]/P0001  , \u4_u2_buf0_reg[25]/P0001  , \u4_u2_buf0_reg[26]/P0001  , \u4_u2_buf0_reg[27]/P0001  , \u4_u2_buf0_reg[28]/P0001  , \u4_u2_buf0_reg[29]/P0001  , \u4_u2_buf0_reg[2]/P0001  , \u4_u2_buf0_reg[30]/P0001  , \u4_u2_buf0_reg[31]/P0001  , \u4_u2_buf0_reg[3]/P0001  , \u4_u2_buf0_reg[4]/P0001  , \u4_u2_buf0_reg[5]/P0001  , \u4_u2_buf0_reg[6]/P0001  , \u4_u2_buf0_reg[7]/P0001  , \u4_u2_buf0_reg[8]/P0001  , \u4_u2_buf0_reg[9]/P0001  , \u4_u2_buf1_reg[0]/P0001  , \u4_u2_buf1_reg[10]/P0001  , \u4_u2_buf1_reg[11]/P0001  , \u4_u2_buf1_reg[12]/P0001  , \u4_u2_buf1_reg[13]/P0001  , \u4_u2_buf1_reg[14]/P0001  , \u4_u2_buf1_reg[15]/P0001  , \u4_u2_buf1_reg[16]/P0001  , \u4_u2_buf1_reg[17]/P0001  , \u4_u2_buf1_reg[18]/P0001  , \u4_u2_buf1_reg[19]/P0001  , \u4_u2_buf1_reg[1]/P0001  , \u4_u2_buf1_reg[20]/P0001  , \u4_u2_buf1_reg[21]/P0001  , \u4_u2_buf1_reg[22]/P0001  , \u4_u2_buf1_reg[23]/P0001  , \u4_u2_buf1_reg[24]/P0001  , \u4_u2_buf1_reg[25]/P0001  , \u4_u2_buf1_reg[26]/P0001  , \u4_u2_buf1_reg[27]/P0001  , \u4_u2_buf1_reg[28]/P0001  , \u4_u2_buf1_reg[29]/P0001  , \u4_u2_buf1_reg[2]/P0001  , \u4_u2_buf1_reg[30]/P0001  , \u4_u2_buf1_reg[31]/P0001  , \u4_u2_buf1_reg[3]/P0001  , \u4_u2_buf1_reg[4]/P0001  , \u4_u2_buf1_reg[5]/P0001  , \u4_u2_buf1_reg[6]/P0001  , \u4_u2_buf1_reg[7]/P0001  , \u4_u2_buf1_reg[8]/P0001  , \u4_u2_buf1_reg[9]/P0001  , \u4_u2_csr0_reg[0]/P0001  , \u4_u2_csr0_reg[10]/P0001  , \u4_u2_csr0_reg[11]/P0001  , \u4_u2_csr0_reg[12]/P0001  , \u4_u2_csr0_reg[1]/P0001  , \u4_u2_csr0_reg[2]/P0001  , \u4_u2_csr0_reg[3]/NET0131  , \u4_u2_csr0_reg[4]/P0001  , \u4_u2_csr0_reg[5]/P0001  , \u4_u2_csr0_reg[6]/P0001  , \u4_u2_csr0_reg[7]/P0001  , \u4_u2_csr0_reg[8]/P0001  , \u4_u2_csr0_reg[9]/P0001  , \u4_u2_csr1_reg[0]/P0001  , \u4_u2_csr1_reg[10]/P0001  , \u4_u2_csr1_reg[11]/P0001  , \u4_u2_csr1_reg[12]/P0001  , \u4_u2_csr1_reg[1]/P0001  , \u4_u2_csr1_reg[2]/P0001  , \u4_u2_csr1_reg[3]/P0001  , \u4_u2_csr1_reg[4]/P0001  , \u4_u2_csr1_reg[5]/P0001  , \u4_u2_csr1_reg[6]/P0001  , \u4_u2_csr1_reg[7]/P0001  , \u4_u2_csr1_reg[8]/P0001  , \u4_u2_csr1_reg[9]/P0001  , \u4_u2_dma_ack_clr1_reg/P0001  , \u4_u2_dma_ack_wr1_reg/P0001  , \u4_u2_dma_in_buf_sz1_reg/P0001  , \u4_u2_dma_in_cnt_reg[0]/P0001  , \u4_u2_dma_in_cnt_reg[10]/P0001  , \u4_u2_dma_in_cnt_reg[11]/P0001  , \u4_u2_dma_in_cnt_reg[1]/P0001  , \u4_u2_dma_in_cnt_reg[2]/P0001  , \u4_u2_dma_in_cnt_reg[3]/P0001  , \u4_u2_dma_in_cnt_reg[4]/P0001  , \u4_u2_dma_in_cnt_reg[5]/P0001  , \u4_u2_dma_in_cnt_reg[6]/P0001  , \u4_u2_dma_in_cnt_reg[7]/P0001  , \u4_u2_dma_in_cnt_reg[8]/P0001  , \u4_u2_dma_in_cnt_reg[9]/P0001  , \u4_u2_dma_out_buf_avail_reg/P0001  , \u4_u2_dma_out_cnt_reg[10]/P0001  , \u4_u2_dma_out_cnt_reg[11]/P0001  , \u4_u2_dma_out_cnt_reg[1]/P0001  , \u4_u2_dma_out_cnt_reg[2]/P0001  , \u4_u2_dma_out_cnt_reg[3]/P0001  , \u4_u2_dma_out_cnt_reg[4]/P0001  , \u4_u2_dma_out_cnt_reg[5]/P0001  , \u4_u2_dma_out_cnt_reg[6]/P0001  , \u4_u2_dma_out_cnt_reg[7]/P0001  , \u4_u2_dma_out_cnt_reg[8]/P0001  , \u4_u2_dma_out_cnt_reg[9]/P0001  , \u4_u2_dma_out_left_reg[0]/P0001  , \u4_u2_dma_out_left_reg[10]/P0001  , \u4_u2_dma_out_left_reg[11]/P0001  , \u4_u2_dma_out_left_reg[1]/P0001  , \u4_u2_dma_out_left_reg[2]/P0001  , \u4_u2_dma_out_left_reg[3]/P0001  , \u4_u2_dma_out_left_reg[4]/P0001  , \u4_u2_dma_out_left_reg[5]/P0001  , \u4_u2_dma_out_left_reg[6]/P0001  , \u4_u2_dma_out_left_reg[7]/P0001  , \u4_u2_dma_out_left_reg[8]/P0001  , \u4_u2_dma_out_left_reg[9]/P0001  , \u4_u2_dma_req_in_hold2_reg/P0001  , \u4_u2_dma_req_in_hold_reg/P0001  , \u4_u2_dma_req_out_hold_reg/P0001  , \u4_u2_ep_match_r_reg/P0001  , \u4_u2_iena_reg[0]/P0001  , \u4_u2_iena_reg[1]/P0001  , \u4_u2_iena_reg[2]/P0001  , \u4_u2_iena_reg[3]/P0001  , \u4_u2_iena_reg[4]/P0001  , \u4_u2_iena_reg[5]/P0001  , \u4_u2_ienb_reg[0]/P0001  , \u4_u2_ienb_reg[1]/P0001  , \u4_u2_ienb_reg[2]/P0001  , \u4_u2_ienb_reg[3]/P0001  , \u4_u2_ienb_reg[4]/P0001  , \u4_u2_ienb_reg[5]/P0001  , \u4_u2_int_re_reg/P0001  , \u4_u2_int_stat_reg[0]/P0001  , \u4_u2_int_stat_reg[1]/P0001  , \u4_u2_int_stat_reg[2]/P0001  , \u4_u2_int_stat_reg[3]/P0001  , \u4_u2_int_stat_reg[4]/P0001  , \u4_u2_int_stat_reg[5]/P0001  , \u4_u2_int_stat_reg[6]/P0001  , \u4_u2_inta_reg/P0001  , \u4_u2_intb_reg/P0001  , \u4_u2_ots_stop_reg/P0001  , \u4_u2_r1_reg/P0001  , \u4_u2_r2_reg/P0001  , \u4_u2_r4_reg/P0001  , \u4_u2_r5_reg/NET0131  , \u4_u2_set_r_reg/P0001  , \u4_u2_uc_bsel_reg[0]/P0001  , \u4_u2_uc_bsel_reg[1]/P0001  , \u4_u2_uc_dpd_reg[0]/P0001  , \u4_u2_uc_dpd_reg[1]/P0001  , \u4_u3_buf0_orig_m3_reg[0]/P0001  , \u4_u3_buf0_orig_m3_reg[10]/P0001  , \u4_u3_buf0_orig_m3_reg[11]/P0001  , \u4_u3_buf0_orig_m3_reg[1]/P0001  , \u4_u3_buf0_orig_m3_reg[2]/P0001  , \u4_u3_buf0_orig_m3_reg[3]/P0001  , \u4_u3_buf0_orig_m3_reg[4]/P0001  , \u4_u3_buf0_orig_m3_reg[5]/P0001  , \u4_u3_buf0_orig_m3_reg[6]/P0001  , \u4_u3_buf0_orig_m3_reg[7]/P0001  , \u4_u3_buf0_orig_m3_reg[8]/P0001  , \u4_u3_buf0_orig_m3_reg[9]/P0001  , \u4_u3_buf0_orig_reg[0]/P0001  , \u4_u3_buf0_orig_reg[10]/P0001  , \u4_u3_buf0_orig_reg[11]/P0001  , \u4_u3_buf0_orig_reg[12]/P0001  , \u4_u3_buf0_orig_reg[13]/P0001  , \u4_u3_buf0_orig_reg[14]/P0001  , \u4_u3_buf0_orig_reg[15]/P0001  , \u4_u3_buf0_orig_reg[16]/P0001  , \u4_u3_buf0_orig_reg[17]/P0001  , \u4_u3_buf0_orig_reg[18]/P0001  , \u4_u3_buf0_orig_reg[19]/P0001  , \u4_u3_buf0_orig_reg[1]/P0001  , \u4_u3_buf0_orig_reg[20]/P0001  , \u4_u3_buf0_orig_reg[21]/P0001  , \u4_u3_buf0_orig_reg[22]/P0001  , \u4_u3_buf0_orig_reg[23]/P0001  , \u4_u3_buf0_orig_reg[24]/P0001  , \u4_u3_buf0_orig_reg[25]/P0001  , \u4_u3_buf0_orig_reg[26]/P0001  , \u4_u3_buf0_orig_reg[27]/P0001  , \u4_u3_buf0_orig_reg[28]/P0001  , \u4_u3_buf0_orig_reg[29]/NET0131  , \u4_u3_buf0_orig_reg[2]/P0001  , \u4_u3_buf0_orig_reg[30]/NET0131  , \u4_u3_buf0_orig_reg[31]/P0001  , \u4_u3_buf0_orig_reg[3]/P0001  , \u4_u3_buf0_orig_reg[4]/P0001  , \u4_u3_buf0_orig_reg[5]/P0001  , \u4_u3_buf0_orig_reg[6]/P0001  , \u4_u3_buf0_orig_reg[7]/P0001  , \u4_u3_buf0_orig_reg[8]/P0001  , \u4_u3_buf0_orig_reg[9]/P0001  , \u4_u3_buf0_reg[0]/P0001  , \u4_u3_buf0_reg[10]/P0001  , \u4_u3_buf0_reg[11]/P0001  , \u4_u3_buf0_reg[12]/P0001  , \u4_u3_buf0_reg[13]/P0001  , \u4_u3_buf0_reg[14]/P0001  , \u4_u3_buf0_reg[15]/P0001  , \u4_u3_buf0_reg[16]/P0001  , \u4_u3_buf0_reg[17]/P0001  , \u4_u3_buf0_reg[18]/P0001  , \u4_u3_buf0_reg[19]/P0001  , \u4_u3_buf0_reg[1]/P0001  , \u4_u3_buf0_reg[20]/P0001  , \u4_u3_buf0_reg[21]/P0001  , \u4_u3_buf0_reg[22]/P0001  , \u4_u3_buf0_reg[23]/P0001  , \u4_u3_buf0_reg[24]/P0001  , \u4_u3_buf0_reg[25]/P0001  , \u4_u3_buf0_reg[26]/P0001  , \u4_u3_buf0_reg[27]/P0001  , \u4_u3_buf0_reg[28]/P0001  , \u4_u3_buf0_reg[29]/P0001  , \u4_u3_buf0_reg[2]/P0001  , \u4_u3_buf0_reg[30]/P0001  , \u4_u3_buf0_reg[31]/P0001  , \u4_u3_buf0_reg[3]/P0001  , \u4_u3_buf0_reg[4]/P0001  , \u4_u3_buf0_reg[5]/P0001  , \u4_u3_buf0_reg[6]/P0001  , \u4_u3_buf0_reg[7]/P0001  , \u4_u3_buf0_reg[8]/P0001  , \u4_u3_buf0_reg[9]/P0001  , \u4_u3_buf1_reg[0]/P0001  , \u4_u3_buf1_reg[10]/P0001  , \u4_u3_buf1_reg[11]/P0001  , \u4_u3_buf1_reg[12]/P0001  , \u4_u3_buf1_reg[13]/P0001  , \u4_u3_buf1_reg[14]/P0001  , \u4_u3_buf1_reg[15]/P0001  , \u4_u3_buf1_reg[16]/P0001  , \u4_u3_buf1_reg[17]/P0001  , \u4_u3_buf1_reg[18]/P0001  , \u4_u3_buf1_reg[19]/P0001  , \u4_u3_buf1_reg[1]/P0001  , \u4_u3_buf1_reg[20]/P0001  , \u4_u3_buf1_reg[21]/P0001  , \u4_u3_buf1_reg[22]/P0001  , \u4_u3_buf1_reg[23]/P0001  , \u4_u3_buf1_reg[24]/P0001  , \u4_u3_buf1_reg[25]/P0001  , \u4_u3_buf1_reg[26]/P0001  , \u4_u3_buf1_reg[27]/P0001  , \u4_u3_buf1_reg[28]/P0001  , \u4_u3_buf1_reg[29]/P0001  , \u4_u3_buf1_reg[2]/P0001  , \u4_u3_buf1_reg[30]/P0001  , \u4_u3_buf1_reg[31]/P0001  , \u4_u3_buf1_reg[3]/P0001  , \u4_u3_buf1_reg[4]/P0001  , \u4_u3_buf1_reg[5]/P0001  , \u4_u3_buf1_reg[6]/P0001  , \u4_u3_buf1_reg[7]/P0001  , \u4_u3_buf1_reg[8]/P0001  , \u4_u3_buf1_reg[9]/P0001  , \u4_u3_csr0_reg[0]/P0001  , \u4_u3_csr0_reg[10]/P0001  , \u4_u3_csr0_reg[11]/P0001  , \u4_u3_csr0_reg[12]/P0001  , \u4_u3_csr0_reg[1]/P0001  , \u4_u3_csr0_reg[2]/P0001  , \u4_u3_csr0_reg[3]/NET0131  , \u4_u3_csr0_reg[4]/P0001  , \u4_u3_csr0_reg[5]/P0001  , \u4_u3_csr0_reg[6]/P0001  , \u4_u3_csr0_reg[7]/P0001  , \u4_u3_csr0_reg[8]/P0001  , \u4_u3_csr0_reg[9]/P0001  , \u4_u3_csr1_reg[0]/P0001  , \u4_u3_csr1_reg[10]/P0001  , \u4_u3_csr1_reg[11]/P0001  , \u4_u3_csr1_reg[12]/P0001  , \u4_u3_csr1_reg[1]/P0001  , \u4_u3_csr1_reg[2]/P0001  , \u4_u3_csr1_reg[3]/P0001  , \u4_u3_csr1_reg[4]/P0001  , \u4_u3_csr1_reg[5]/P0001  , \u4_u3_csr1_reg[6]/P0001  , \u4_u3_csr1_reg[7]/P0001  , \u4_u3_csr1_reg[8]/P0001  , \u4_u3_csr1_reg[9]/P0001  , \u4_u3_dma_ack_clr1_reg/P0001  , \u4_u3_dma_ack_wr1_reg/P0001  , \u4_u3_dma_in_buf_sz1_reg/P0001  , \u4_u3_dma_in_cnt_reg[0]/P0001  , \u4_u3_dma_in_cnt_reg[10]/P0001  , \u4_u3_dma_in_cnt_reg[11]/P0001  , \u4_u3_dma_in_cnt_reg[1]/P0001  , \u4_u3_dma_in_cnt_reg[2]/P0001  , \u4_u3_dma_in_cnt_reg[3]/P0001  , \u4_u3_dma_in_cnt_reg[4]/P0001  , \u4_u3_dma_in_cnt_reg[5]/P0001  , \u4_u3_dma_in_cnt_reg[6]/P0001  , \u4_u3_dma_in_cnt_reg[7]/P0001  , \u4_u3_dma_in_cnt_reg[8]/P0001  , \u4_u3_dma_in_cnt_reg[9]/P0001  , \u4_u3_dma_out_buf_avail_reg/P0001  , \u4_u3_dma_out_cnt_reg[10]/P0001  , \u4_u3_dma_out_cnt_reg[11]/P0001  , \u4_u3_dma_out_cnt_reg[1]/P0001  , \u4_u3_dma_out_cnt_reg[2]/P0001  , \u4_u3_dma_out_cnt_reg[3]/P0001  , \u4_u3_dma_out_cnt_reg[4]/P0001  , \u4_u3_dma_out_cnt_reg[5]/P0001  , \u4_u3_dma_out_cnt_reg[6]/P0001  , \u4_u3_dma_out_cnt_reg[7]/P0001  , \u4_u3_dma_out_cnt_reg[8]/P0001  , \u4_u3_dma_out_cnt_reg[9]/P0001  , \u4_u3_dma_out_left_reg[0]/P0001  , \u4_u3_dma_out_left_reg[10]/P0001  , \u4_u3_dma_out_left_reg[11]/P0001  , \u4_u3_dma_out_left_reg[1]/P0001  , \u4_u3_dma_out_left_reg[2]/P0001  , \u4_u3_dma_out_left_reg[3]/P0001  , \u4_u3_dma_out_left_reg[4]/P0001  , \u4_u3_dma_out_left_reg[5]/P0001  , \u4_u3_dma_out_left_reg[6]/P0001  , \u4_u3_dma_out_left_reg[7]/P0001  , \u4_u3_dma_out_left_reg[8]/P0001  , \u4_u3_dma_out_left_reg[9]/P0001  , \u4_u3_dma_req_in_hold2_reg/P0001  , \u4_u3_dma_req_in_hold_reg/P0001  , \u4_u3_dma_req_out_hold_reg/P0001  , \u4_u3_ep_match_r_reg/P0001  , \u4_u3_iena_reg[0]/P0001  , \u4_u3_iena_reg[1]/P0001  , \u4_u3_iena_reg[2]/P0001  , \u4_u3_iena_reg[3]/P0001  , \u4_u3_iena_reg[4]/P0001  , \u4_u3_iena_reg[5]/P0001  , \u4_u3_ienb_reg[0]/P0001  , \u4_u3_ienb_reg[1]/P0001  , \u4_u3_ienb_reg[2]/P0001  , \u4_u3_ienb_reg[3]/P0001  , \u4_u3_ienb_reg[4]/P0001  , \u4_u3_ienb_reg[5]/P0001  , \u4_u3_int_re_reg/P0001  , \u4_u3_int_stat_reg[0]/P0001  , \u4_u3_int_stat_reg[1]/P0001  , \u4_u3_int_stat_reg[2]/P0001  , \u4_u3_int_stat_reg[3]/P0001  , \u4_u3_int_stat_reg[4]/P0001  , \u4_u3_int_stat_reg[5]/P0001  , \u4_u3_int_stat_reg[6]/P0001  , \u4_u3_inta_reg/P0001  , \u4_u3_intb_reg/P0001  , \u4_u3_ots_stop_reg/P0001  , \u4_u3_r1_reg/P0001  , \u4_u3_r2_reg/P0001  , \u4_u3_r4_reg/P0001  , \u4_u3_r5_reg/NET0131  , \u4_u3_set_r_reg/P0001  , \u4_u3_uc_bsel_reg[0]/P0001  , \u4_u3_uc_bsel_reg[1]/P0001  , \u4_u3_uc_dpd_reg[0]/P0001  , \u4_u3_uc_dpd_reg[1]/P0001  , \u4_usb_reset_r_reg/P0001  , \u4_utmi_vend_ctrl_r_reg[0]/P0001  , \u4_utmi_vend_ctrl_r_reg[1]/P0001  , \u4_utmi_vend_ctrl_r_reg[2]/P0001  , \u4_utmi_vend_ctrl_r_reg[3]/P0001  , \u4_utmi_vend_stat_r_reg[0]/P0001  , \u4_utmi_vend_stat_r_reg[1]/P0001  , \u4_utmi_vend_stat_r_reg[2]/P0001  , \u4_utmi_vend_stat_r_reg[3]/P0001  , \u4_utmi_vend_stat_r_reg[4]/P0001  , \u4_utmi_vend_stat_r_reg[5]/P0001  , \u4_utmi_vend_stat_r_reg[6]/P0001  , \u4_utmi_vend_stat_r_reg[7]/P0001  , \u4_utmi_vend_wr_r_reg/P0001  , \u5_state_reg[0]/P0001  , \u5_state_reg[1]/P0001  , \u5_state_reg[2]/P0001  , \u5_state_reg[3]/P0001  , \u5_state_reg[4]/P0001  , \u5_state_reg[5]/NET0131  , \u5_wb_ack_s1_reg/P0001  , \u5_wb_ack_s2_reg/P0001  , \u5_wb_req_s1_reg/P0001  , usb_vbus_pad_i_pad , wb_ack_o_pad , \wb_addr_i[10]_pad  , \wb_addr_i[11]_pad  , \wb_addr_i[12]_pad  , \wb_addr_i[13]_pad  , \wb_addr_i[14]_pad  , \wb_addr_i[15]_pad  , \wb_addr_i[16]_pad  , \wb_addr_i[17]_pad  , \wb_addr_i[2]_pad  , \wb_addr_i[3]_pad  , \wb_addr_i[4]_pad  , \wb_addr_i[5]_pad  , \wb_addr_i[6]_pad  , \wb_addr_i[7]_pad  , \wb_addr_i[8]_pad  , \wb_addr_i[9]_pad  , wb_cyc_i_pad , \wb_data_i[0]_pad  , \wb_data_i[10]_pad  , \wb_data_i[11]_pad  , \wb_data_i[12]_pad  , \wb_data_i[13]_pad  , \wb_data_i[14]_pad  , \wb_data_i[15]_pad  , \wb_data_i[16]_pad  , \wb_data_i[17]_pad  , \wb_data_i[18]_pad  , \wb_data_i[19]_pad  , \wb_data_i[1]_pad  , \wb_data_i[20]_pad  , \wb_data_i[21]_pad  , \wb_data_i[22]_pad  , \wb_data_i[23]_pad  , \wb_data_i[24]_pad  , \wb_data_i[25]_pad  , \wb_data_i[26]_pad  , \wb_data_i[27]_pad  , \wb_data_i[28]_pad  , \wb_data_i[29]_pad  , \wb_data_i[2]_pad  , \wb_data_i[30]_pad  , \wb_data_i[31]_pad  , \wb_data_i[3]_pad  , \wb_data_i[4]_pad  , \wb_data_i[5]_pad  , \wb_data_i[6]_pad  , \wb_data_i[7]_pad  , \wb_data_i[8]_pad  , \wb_data_i[9]_pad  , wb_stb_i_pad , wb_we_i_pad , \dma_req_o[6]_pad  , \g37425/_0_  , \g37426/_0_  , \g37432/_0_  , \g37433/_0_  , \g37439/_0_  , \g37440/_0_  , \g37444/_00_  , \g37448/_0_  , \g37450/_0_  , \g37454/_0_  , \g37473/_0_  , \g37474/_0_  , \g37475/_0_  , \g37476/_0_  , \g37477/_0_  , \g37478/_0_  , \g37479/_0_  , \g37488/_0_  , \g37489/_0_  , \g37490/_0_  , \g37491/_0_  , \g37492/_0_  , \g37517/_0_  , \g37518/_0_  , \g37519/_0_  , \g37520/_0_  , \g37521/_0_  , \g37522/_0_  , \g37540/_0_  , \g37542/_0_  , \g37543/_0_  , \g37545/_0_  , \g37546/_0_  , \g37548/_0_  , \g37549/_0_  , \g37550/_0_  , \g37551/_0_  , \g37556/_0_  , \g37589/_0_  , \g37591/_0_  , \g37592/_0_  , \g37593/_0_  , \g37594/_0_  , \g37596/_0_  , \g37597/_0_  , \g37598/_0_  , \g37599/_0_  , \g37601/_0_  , \g37603/_0_  , \g37604/_0_  , \g37605/_0_  , \g37607/_0_  , \g37608/_0_  , \g37609/_0_  , \g37610/_0_  , \g37645/_0_  , \g37648/_0_  , \g37650/_0_  , \g37653/_0_  , \g37664/_3_  , \g37703/_0_  , \g37704/_0_  , \g37706/_0_  , \g37708/_0_  , \g37709/_0_  , \g37711/_0_  , \g37714/_0_  , \g37715/_0_  , \g37717/_0_  , \g37718/_0_  , \g37719/_0_  , \g37720/_0_  , \g37723/_0_  , \g37724/_0_  , \g37726/_0_  , \g37728/_0_  , \g37729/_0_  , \g37730/_0_  , \g37731/_0_  , \g37732/_0_  , \g37733/_0_  , \g37735/_0_  , \g37736/_0_  , \g37737/_0_  , \g37856/_0_  , \g37857/_0_  , \g37859/_0_  , \g37868/_0_  , \g37869/_0_  , \g37870/_0_  , \g37872/_0_  , \g37886/_0_  , \g37887/_0_  , \g37889/_0_  , \g37897/_0_  , \g37899/_0_  , \g37900/_0_  , \g37907/_0_  , \g37925/_0_  , \g37927/_0_  , \g37928/_0_  , \g37929/_0_  , \g37930/_0_  , \g37932/_0_  , \g37933/_0_  , \g37934/_0_  , \g37935/_0_  , \g37936/_0_  , \g37937/_0_  , \g37938/_0_  , \g37939/_0_  , \g37941/_0_  , \g37942/_0_  , \g37943/_0_  , \g37944/_0_  , \g37945/_0_  , \g38030/_3_  , \g38035/_0_  , \g38036/_0_  , \g38054/_0_  , \g38129/_0_  , \g38130/_0_  , \g38148/_3_  , \g38149/_3_  , \g38150/_3_  , \g38166/_0_  , \g38198/_0_  , \g38201/_0_  , \g38257/_0_  , \g38286/_0_  , \g38294/_3_  , \g38295/_3_  , \g38296/_3_  , \g38297/_3_  , \g38332/_0_  , \g38350/_0_  , \g38365/_3_  , \g38366/_3_  , \g38367/_3_  , \g38389/_0_  , \g38397/_0_  , \g38398/_0_  , \g38399/_0_  , \g38400/_0_  , \g38417/_3_  , \g38418/_3_  , \g38422/_0_  , \g38440/_0_  , \g38443/_0_  , \g38448/_3_  , \g38449/_0_  , \g38450/_0_  , \g38460/_0_  , \g38466/_0_  , \g38467/_0_  , \g38468/_0_  , \g38469/_0_  , \g38470/_0_  , \g38471/_0_  , \g38472/_0_  , \g38473/_0_  , \g38474/_0_  , \g38475/_0_  , \g38476/_0_  , \g38477/_0_  , \g38478/_0_  , \g38479/_0_  , \g38528/_0_  , \g38533/_0_  , \g38534/_0_  , \g38536/_0_  , \g38545/_0_  , \g38551/_0_  , \g38554/_0_  , \g38555/_0_  , \g38556/_0_  , \g38575/_0_  , \g38616/_0_  , \g38653/_0_  , \g38656/_0_  , \g38657/_0_  , \g38658/_0_  , \g38660/_0_  , \g38706/_0_  , \g38716/_0_  , \g38717/_0_  , \g38738/_1_  , \g38763/_0_  , \g38790/_0_  , \g38792/_0_  , \g38801/_0_  , \g38803/_0_  , \g38804/_0_  , \g38805/_0_  , \g38806/_0_  , \g38807/_0_  , \g38808/_0_  , \g38809/_0_  , \g38810/_0_  , \g38814/_0_  , \g38833/_0_  , \g38834/_0_  , \g38839/_0_  , \g38840/_0_  , \g38841/_0_  , \g38842/_0_  , \g38846/_0_  , \g38847/_0_  , \g38848/_0_  , \g38849/_0_  , \g38853/_0_  , \g38857/_0_  , \g38872/_0_  , \g38882/_0_  , \g38884/_0_  , \g38885/_0_  , \g38886/_0_  , \g38887/_0_  , \g38931/_0_  , \g38952/_0_  , \g38960/_0_  , \g38971/_0_  , \g38973/_0_  , \g38974/_0_  , \g38975/_0_  , \g38976/_0_  , \g38978/_0_  , \g38981/_0_  , \g38986/_0_  , \g38987/_0_  , \g39001/_3_  , \g39003/_3_  , \g39009/_3_  , \g39011/_3_  , \g39013/_3_  , \g39015/_2_  , \g39017/_2_  , \g39019/_2_  , \g39021/_2_  , \g39060/_0_  , \g39061/_3_  , \g39062/_0_  , \g39063/_0_  , \g39065/_0_  , \g39066/_0_  , \g39093/_0_  , \g39099/_2_  , \g39118/_0_  , \g39123/_0_  , \g39174/_0_  , \g39175/_0_  , \g39176/_0_  , \g39177/_0_  , \g39178/_0_  , \g39185/_0_  , \g39186/_0_  , \g39187/_0_  , \g39188/_0_  , \g39194/_0_  , \g39195/_0_  , \g39196/_0_  , \g39197/_0_  , \g39198/_0_  , \g39199/_0_  , \g39200/_0_  , \g39201/_0_  , \g39202/_0_  , \g39203/_0_  , \g39204/_0_  , \g39216/_3_  , \g39217/_3_  , \g39218/_0_  , \g39219/_0_  , \g39220/_0_  , \g39221/_0_  , \g39299/_0_  , \g39300/_0_  , \g39301/_0_  , \g39302/_0_  , \g39303/_0_  , \g39304/_0_  , \g39305/_0_  , \g39306/_0_  , \g39307/_0_  , \g39308/_0_  , \g39309/_0_  , \g39310/_0_  , \g39311/_0_  , \g39315/_0_  , \g39318/_0_  , \g39321/_0_  , \g39322/_0_  , \g39323/_0_  , \g39333/_0_  , \g39334/_0_  , \g39336/_0_  , \g39338/_0_  , \g39339/_0_  , \g39340/_0_  , \g39341/_0_  , \g39342/_0_  , \g39343/_0_  , \g39344/_0_  , \g39345/_0_  , \g39346/_0_  , \g39349/_0_  , \g39352/_3_  , \g39354/_3_  , \g39371/_3_  , \g39372/_3_  , \g39373/_3_  , \g39374/_3_  , \g39376/_0_  , \g39377/_0_  , \g39471/_0_  , \g39472/_0_  , \g39473/_0_  , \g39474/_0_  , \g39475/_0_  , \g39476/_0_  , \g39477/_0_  , \g39478/_0_  , \g39479/_0_  , \g39480/_0_  , \g39481/_0_  , \g39482/_0_  , \g39483/_0_  , \g39484/_0_  , \g39485/_0_  , \g39486/_0_  , \g39487/_0_  , \g39488/_0_  , \g39492/_0_  , \g39497/_0_  , \g39501/_0_  , \g39502/_0_  , \g39503/_0_  , \g39504/_0_  , \g39505/_0_  , \g39506/_0_  , \g39539/_0_  , \g39541/_0_  , \g39542/_0_  , \g39543/_0_  , \g39544/_0_  , \g39545/_0_  , \g39546/_0_  , \g39547/_0_  , \g39550/_0_  , \g39551/_0_  , \g39563/_0_  , \g39568/_00_  , \g39617/_0_  , \g39618/_0_  , \g39621/_0_  , \g39622/_0_  , \g39623/_0_  , \g39624/_00_  , \g39685/_0_  , \g39690/_0_  , \g39693/_0_  , \g39695/_0_  , \g39697/_0_  , \g39706/_0_  , \g39749/_0_  , \g39750/_0_  , \g39751/_0_  , \g39752/_0_  , \g39753/_0_  , \g39754/_0_  , \g39755/_0_  , \g39756/_0_  , \g39757/_0_  , \g39758/_0_  , \g39759/_0_  , \g39760/_0_  , \g39761/_0_  , \g39762/_0_  , \g39763/_0_  , \g39764/_0_  , \g39765/_0_  , \g39766/_0_  , \g39767/_0_  , \g39768/_0_  , \g39769/_0_  , \g39770/_0_  , \g39772/_0_  , \g39773/_0_  , \g39775/_3_  , \g39776/_3_  , \g39777/_3_  , \g39778/_3_  , \g39779/_3_  , \g39780/_3_  , \g39781/_3_  , \g39782/_3_  , \g39788/_3_  , \g39799/_0_  , \g39800/_0_  , \g39801/_0_  , \g39802/_0_  , \g39927/_0_  , \g39928/_0_  , \g39929/_0_  , \g39930/_0_  , \g39931/_0_  , \g39932/_0_  , \g39933/_0_  , \g39934/_0_  , \g39935/_0_  , \g39936/_0_  , \g39937/_0_  , \g39938/_0_  , \g39939/_0_  , \g39940/_0_  , \g39942/_0_  , \g39943/_0_  , \g39944/_0_  , \g39945/_0_  , \g39956/_0_  , \g39957/_0_  , \g39958/_0_  , \g39959/_0_  , \g39960/_0_  , \g39961/_0_  , \g39962/_0_  , \g39963/_0_  , \g39964/_0_  , \g39969/_0_  , \g39974/_0_  , \g39975/_0_  , \g39993/_0_  , \g39994/_0_  , \g40003/_0_  , \g40004/_0_  , \g40005/_0_  , \g40006/_0_  , \g40016/_0_  , \g40023/_3_  , \g40033/_0_  , \g40034/_0_  , \g40035/_0_  , \g40036/_0_  , \g40037/_0_  , \g40038/_0_  , \g40199/_0_  , \g40200/_0_  , \g40201/_0_  , \g40202/_0_  , \g40203/_0_  , \g40204/_0_  , \g40205/_0_  , \g40206/_0_  , \g40207/_0_  , \g40208/_0_  , \g40209/_0_  , \g40210/_0_  , \g40224/_0_  , \g40225/_0_  , \g40226/_0_  , \g40227/_0_  , \g40234/_0_  , \g40235/_0_  , \g40236/_0_  , \g40237/_0_  , \g40238/_0_  , \g40239/_0_  , \g40240/_0_  , \g40241/_0_  , \g40242/_0_  , \g40243/_0_  , \g40244/_0_  , \g40246/_0_  , \g40247/_0_  , \g40248/_0_  , \g40249/_0_  , \g40250/_0_  , \g40251/_0_  , \g40252/_0_  , \g40253/_0_  , \g40254/_0_  , \g40255/_0_  , \g40257/_0_  , \g40258/_0_  , \g40262/_0_  , \g40264/_0_  , \g40265/_0_  , \g40266/_0_  , \g40267/_0_  , \g40268/_0_  , \g40269/_0_  , \g40270/_0_  , \g40271/_0_  , \g40272/_0_  , \g40273/_0_  , \g40274/_0_  , \g40275/_0_  , \g40276/_0_  , \g40277/_0_  , \g40278/_0_  , \g40280/_2_  , \g40281/_0_  , \g40282/_0_  , \g40283/_0_  , \g40284/_0_  , \g40285/_0_  , \g40286/_0_  , \g40287/_0_  , \g40288/_0_  , \g40289/_0_  , \g40290/_0_  , \g40291/_0_  , \g40297/_0_  , \g40298/_0_  , \g40299/_0_  , \g40300/_0_  , \g40301/_0_  , \g40302/_0_  , \g40303/_0_  , \g40304/_0_  , \g40306/_0_  , \g40307/_0_  , \g40308/_0_  , \g40309/_0_  , \g40310/_0_  , \g40311/_0_  , \g40312/_0_  , \g40313/_0_  , \g40314/_0_  , \g40315/_0_  , \g40316/_0_  , \g40317/_0_  , \g40318/_0_  , \g40319/_0_  , \g40320/_0_  , \g40324/_0_  , \g40325/_0_  , \g40326/_0_  , \g40327/_0_  , \g40328/_0_  , \g40329/_0_  , \g40330/_0_  , \g40331/_0_  , \g40332/_0_  , \g40333/_0_  , \g40334/_0_  , \g40335/_0_  , \g40336/_0_  , \g40337/_0_  , \g40338/_0_  , \g40339/_0_  , \g40340/_0_  , \g40341/_0_  , \g40342/_0_  , \g40343/_0_  , \g40344/_0_  , \g40345/_0_  , \g40346/_0_  , \g40347/_0_  , \g40350/_0_  , \g40353/_0_  , \g40354/_0_  , \g40355/_0_  , \g40374/_0_  , \g40457/_0_  , \g40458/_0_  , \g40549/_0_  , \g40550/_0_  , \g40551/_0_  , \g40552/_0_  , \g40553/_0_  , \g40554/_0_  , \g40556/_0_  , \g40557/_0_  , \g40558/_0_  , \g40559/_0_  , \g40561/_0_  , \g40562/_0_  , \g40563/_0_  , \g40565/_0_  , \g40566/_0_  , \g40567/_0_  , \g40569/_0_  , \g40570/_0_  , \g40571/_0_  , \g40572/_0_  , \g40573/_0_  , \g40574/_0_  , \g40575/_0_  , \g40576/_0_  , \g40577/_0_  , \g40578/_0_  , \g40579/_0_  , \g40580/_0_  , \g40581/_0_  , \g40582/_0_  , \g40583/_0_  , \g40584/_0_  , \g40586/_0_  , \g40587/_0_  , \g40588/_0_  , \g40589/_0_  , \g40591/_0_  , \g40592/_0_  , \g40593/_0_  , \g40594/_0_  , \g40595/_0_  , \g40596/_0_  , \g40597/_0_  , \g40598/_0_  , \g40599/_0_  , \g40600/_0_  , \g40601/_0_  , \g40602/_0_  , \g40603/_0_  , \g40604/_0_  , \g40605/_0_  , \g40606/_0_  , \g40607/_0_  , \g40608/_0_  , \g40609/_0_  , \g40610/_0_  , \g40611/_0_  , \g40612/_0_  , \g40613/_0_  , \g40614/_0_  , \g40617/_0_  , \g40629/_0_  , \g40632/_0_  , \g40633/_0_  , \g40634/_0_  , \g40635/_0_  , \g40636/_0_  , \g40637/_0_  , \g40638/_0_  , \g40639/_0_  , \g40640/_0_  , \g40641/_0_  , \g40642/_0_  , \g40643/_0_  , \g40644/_0_  , \g40645/_0_  , \g40646/_0_  , \g40647/_0_  , \g40648/_0_  , \g40649/_0_  , \g40650/_0_  , \g40651/_0_  , \g40652/_0_  , \g40653/_0_  , \g40654/_0_  , \g40655/_0_  , \g40661/_0_  , \g40663/_0_  , \g40664/_0_  , \g40665/_0_  , \g40666/_0_  , \g40667/_0_  , \g40668/_0_  , \g40669/_0_  , \g40670/_0_  , \g40671/_0_  , \g40672/_0_  , \g40673/_0_  , \g40674/_0_  , \g40675/_0_  , \g40676/_0_  , \g40677/_0_  , \g40678/_0_  , \g40679/_0_  , \g40680/_0_  , \g40681/_0_  , \g40682/_0_  , \g40683/_0_  , \g40684/_0_  , \g40685/_0_  , \g40689/_0_  , \g40690/_0_  , \g40691/_0_  , \g40692/_0_  , \g40693/_0_  , \g40694/_0_  , \g40695/_0_  , \g40696/_0_  , \g40697/_0_  , \g40698/_0_  , \g40699/_0_  , \g40700/_0_  , \g40701/_0_  , \g40702/_0_  , \g40703/_0_  , \g40704/_0_  , \g40705/_0_  , \g40706/_0_  , \g40707/_0_  , \g40708/_0_  , \g40709/_0_  , \g40710/_0_  , \g40711/_0_  , \g40712/_0_  , \g40758/_00_  , \g40759/_0_  , \g40812/_0_  , \g40816/_0_  , \g40817/_0_  , \g40818/_0_  , \g40819/_0_  , \g40820/_0_  , \g40822/_3_  , \g40823/_3_  , \g40824/_3_  , \g40825/_3_  , \g40849/_3_  , \g40915/_0_  , \g40916/_0_  , \g40917/_0_  , \g40920/_0_  , \g40923/_0_  , \g40926/_0_  , \g40927/_0_  , \g40930/_0_  , \g40931/_0_  , \g41138/_0_  , \g41152/_0_  , \g41180/_0_  , \g41185/_0_  , \g41186/_0_  , \g41187/_0_  , \g41189/_0_  , \g41190/_0_  , \g41191/_0_  , \g41192/_0_  , \g41193/_0_  , \g41195/_0_  , \g41199/_0_  , \g41207/_0_  , \g41221/_0_  , \g41226/_0_  , \g41227/_0_  , \g41230/_0_  , \g41231/_0_  , \g41234/_0_  , \g41238/_0_  , \g41239/_0_  , \g41275/_0_  , \g41277/_0_  , \g41278/_0_  , \g41279/_0_  , \g41280/_0_  , \g41281/_0_  , \g41282/_0_  , \g41283/_0_  , \g41284/_0_  , \g41285/_0_  , \g41286/_0_  , \g41287/_0_  , \g41288/_0_  , \g41289/_0_  , \g41291/_3_  , \g41330/_0_  , \g41332/_0_  , \g41334/_0_  , \g41340/_0_  , \g41343/_0_  , \g41345/_0_  , \g41348/_0_  , \g41349/_0_  , \g41350/_0_  , \g41351/_0_  , \g41356/_0_  , \g41394/_0_  , \g41423/_0_  , \g41426/_3_  , \g41427/_3_  , \g41428/_3_  , \g41429/_3_  , \g41430/_3_  , \g41431/_3_  , \g41432/_3_  , \g41433/_3_  , \g41434/_3_  , \g41435/_3_  , \g41436/_3_  , \g41437/_3_  , \g41438/_3_  , \g41439/_3_  , \g41440/_3_  , \g41441/_3_  , \g41442/_0_  , \g41445/_3_  , \g41446/_0_  , \g41449/_0_  , \g41464/_0_  , \g41466/_0_  , \g41468/_0_  , \g41469/_0_  , \g41471/_0_  , \g41795/_0_  , \g41799/_0_  , \g41800/_0_  , \g41801/_0_  , \g41802/_0_  , \g41803/_0_  , \g41804/_0_  , \g41805/_0_  , \g41806/_0_  , \g41807/_0_  , \g41808/_0_  , \g41809/_0_  , \g41810/_0_  , \g41811/_0_  , \g41812/_0_  , \g41814/_0_  , \g41815/_0_  , \g41816/_0_  , \g41817/_0_  , \g41818/_0_  , \g41819/_0_  , \g41820/_0_  , \g41821/_0_  , \g41822/_0_  , \g41823/_0_  , \g41825/_0_  , \g41826/_0_  , \g41827/_0_  , \g41828/_0_  , \g41829/_0_  , \g41830/_0_  , \g41831/_0_  , \g41832/_0_  , \g41833/_0_  , \g41834/_0_  , \g41835/_0_  , \g41836/_0_  , \g41837/_0_  , \g41838/_0_  , \g41839/_0_  , \g41840/_0_  , \g41841/_0_  , \g41842/_0_  , \g41843/_0_  , \g41844/_0_  , \g41845/_0_  , \g41846/_0_  , \g41847/_0_  , \g41848/_0_  , \g41849/_0_  , \g41850/_0_  , \g41851/_0_  , \g41852/_0_  , \g41853/_0_  , \g41854/_0_  , \g41855/_0_  , \g41856/_0_  , \g41857/_0_  , \g41858/_0_  , \g41859/_0_  , \g41860/_0_  , \g41861/_0_  , \g41862/_0_  , \g41863/_0_  , \g41864/_0_  , \g41865/_0_  , \g41866/_0_  , \g41867/_0_  , \g41868/_0_  , \g41869/_0_  , \g41870/_0_  , \g41871/_0_  , \g41872/_0_  , \g41873/_0_  , \g41874/_0_  , \g41875/_0_  , \g41876/_0_  , \g41877/_0_  , \g41878/_0_  , \g41879/_0_  , \g41880/_0_  , \g41881/_0_  , \g41882/_0_  , \g41883/_0_  , \g41884/_0_  , \g41885/_0_  , \g41886/_0_  , \g41887/_0_  , \g41888/_0_  , \g41889/_0_  , \g41890/_0_  , \g41891/_0_  , \g41902/_0_  , \g41904/_0_  , \g41906/_0_  , \g41907/_0_  , \g41954/_0_  , \g41955/_0_  , \g41956/_0_  , \g41957/_0_  , \g41958/_0_  , \g41959/_0_  , \g41960/_0_  , \g41962/_0_  , \g41963/_0_  , \g41964/_0_  , \g41965/_0_  , \g41966/_0_  , \g41967/_0_  , \g41968/_0_  , \g41969/_0_  , \g41970/_0_  , \g41971/_0_  , \g41972/_0_  , \g41973/_0_  , \g41974/_0_  , \g41975/_0_  , \g41976/_0_  , \g41977/_0_  , \g41978/_0_  , \g41979/_0_  , \g42062/_0_  , \g42079/_0_  , \g42142/_0_  , \g42143/_0_  , \g42144/_0_  , \g42154/_0_  , \g42157/_0_  , \g42160/_0_  , \g42181/_0_  , \g42203/_0_  , \g42204/_3_  , \g42205/_3_  , \g42206/_3_  , \g42208/_0_  , \g42220/_0_  , \g42225/_0_  , \g42251/_0_  , \g42273/_0_  , \g42335/_0_  , \g42357/_0_  , \g42380/_0_  , \g42381/_0_  , \g42383/_0_  , \g42386/_0_  , \g42388/_0_  , \g42475/_0_  , \g42476/_0_  , \g42477/_0_  , \g42478/_0_  , \g42479/_0_  , \g42480/_0_  , \g42481/_0_  , \g42482/_0_  , \g42483/_0_  , \g42484/_0_  , \g42485/_0_  , \g42486/_0_  , \g42487/_0_  , \g42488/_0_  , \g42490/_0_  , \g42491/_0_  , \g42493/_0_  , \g42494/_0_  , \g42495/_0_  , \g42496/_0_  , \g42497/_0_  , \g42498/_0_  , \g42499/_0_  , \g42500/_0_  , \g42501/_0_  , \g42502/_0_  , \g42503/_0_  , \g42504/_0_  , \g42505/_0_  , \g42506/_0_  , \g42507/_0_  , \g42508/_0_  , \g42509/_0_  , \g42510/_0_  , \g42511/_0_  , \g42512/_0_  , \g42513/_0_  , \g42514/_0_  , \g42515/_0_  , \g42516/_0_  , \g42517/_0_  , \g42518/_0_  , \g42519/_0_  , \g42521/_0_  , \g42522/_0_  , \g42523/_0_  , \g42524/_0_  , \g42525/_0_  , \g42526/_0_  , \g42527/_0_  , \g42528/_0_  , \g42529/_0_  , \g42530/_0_  , \g42531/_0_  , \g42532/_0_  , \g42533/_0_  , \g42534/_0_  , \g42535/_0_  , \g42536/_0_  , \g42537/_0_  , \g42538/_0_  , \g42539/_0_  , \g42540/_0_  , \g42541/_0_  , \g42542/_0_  , \g42543/_0_  , \g42544/_0_  , \g42545/_0_  , \g42548/_0_  , \g42557/_0_  , \g42564/_0_  , \g42565/_0_  , \g42566/_0_  , \g42567/_0_  , \g42568/_0_  , \g42569/_0_  , \g42570/_0_  , \g42571/_0_  , \g42572/_0_  , \g42573/_0_  , \g42574/_0_  , \g42575/_0_  , \g42576/_0_  , \g42577/_0_  , \g42578/_0_  , \g42581/_0_  , \g42589/_0_  , \g42590/_0_  , \g42591/_0_  , \g42592/_0_  , \g42593/_0_  , \g42594/_0_  , \g42595/_0_  , \g42596/_0_  , \g42597/_0_  , \g42598/_0_  , \g42599/_0_  , \g42600/_0_  , \g42601/_0_  , \g42602/_0_  , \g42603/_0_  , \g42604/_0_  , \g42605/_0_  , \g42606/_0_  , \g42607/_0_  , \g42608/_0_  , \g42609/_0_  , \g42610/_0_  , \g42611/_0_  , \g42612/_0_  , \g42613/_0_  , \g42614/_0_  , \g42615/_0_  , \g42616/_0_  , \g42617/_0_  , \g42618/_0_  , \g42619/_0_  , \g42620/_0_  , \g42622/_0_  , \g42623/_0_  , \g42627/_0_  , \g42628/_0_  , \g42629/_0_  , \g42630/_0_  , \g42631/_0_  , \g42632/_0_  , \g42633/_0_  , \g42634/_0_  , \g42635/_0_  , \g42636/_0_  , \g42637/_0_  , \g42638/_0_  , \g42639/_0_  , \g42640/_0_  , \g42641/_0_  , \g42642/_0_  , \g42643/_0_  , \g42644/_0_  , \g42645/_0_  , \g42646/_0_  , \g42647/_0_  , \g42648/_0_  , \g42649/_0_  , \g42650/_0_  , \g42666/_0_  , \g42667/_0_  , \g42668/_0_  , \g42669/_0_  , \g42670/_0_  , \g42671/_0_  , \g42672/_0_  , \g42673/_0_  , \g42674/_0_  , \g42675/_0_  , \g42676/_0_  , \g42677/_0_  , \g42678/_0_  , \g42680/_0_  , \g42681/_0_  , \g42685/_0_  , \g42686/_0_  , \g42688/_0_  , \g42689/_0_  , \g42690/_0_  , \g42691/_0_  , \g42692/_0_  , \g42693/_0_  , \g42694/_0_  , \g42695/_0_  , \g42696/_0_  , \g42697/_0_  , \g42698/_0_  , \g42699/_0_  , \g42700/_0_  , \g42701/_0_  , \g42702/_0_  , \g42703/_0_  , \g42704/_0_  , \g42705/_0_  , \g42706/_0_  , \g42707/_0_  , \g42708/_0_  , \g42709/_0_  , \g42710/_0_  , \g42711/_0_  , \g42712/_0_  , \g42713/_0_  , \g42715/_0_  , \g42716/_0_  , \g42717/_0_  , \g42718/_0_  , \g42723/_1_  , \g42727/_0_  , \g42728/_0_  , \g42729/_0_  , \g42730/_0_  , \g42731/_0_  , \g42732/_0_  , \g42733/_0_  , \g42734/_0_  , \g42735/_0_  , \g42736/_0_  , \g42737/_0_  , \g42738/_0_  , \g42739/_0_  , \g42740/_0_  , \g42741/_0_  , \g42742/_0_  , \g42743/_0_  , \g42744/_0_  , \g42745/_0_  , \g42746/_0_  , \g42747/_0_  , \g42748/_0_  , \g42749/_0_  , \g42750/_0_  , \g42751/_0_  , \g42754/_0_  , \g42767/_0_  , \g42768/_0_  , \g42772/_0_  , \g42773/_0_  , \g42774/_0_  , \g42775/_0_  , \g42776/_0_  , \g42777/_0_  , \g42778/_0_  , \g42779/_0_  , \g42780/_0_  , \g42781/_0_  , \g42782/_0_  , \g42783/_0_  , \g42784/_0_  , \g42785/_0_  , \g42790/_0_  , \g42791/_0_  , \g42792/_0_  , \g42793/_0_  , \g42794/_0_  , \g42795/_0_  , \g42796/_0_  , \g42797/_0_  , \g42798/_0_  , \g42799/_0_  , \g42800/_0_  , \g42801/_0_  , \g42802/_0_  , \g42803/_0_  , \g42804/_0_  , \g42805/_0_  , \g42806/_0_  , \g42807/_0_  , \g42808/_0_  , \g42809/_0_  , \g42810/_0_  , \g42811/_0_  , \g42812/_0_  , \g42813/_0_  , \g42814/_0_  , \g42815/_0_  , \g42816/_0_  , \g42817/_0_  , \g42818/_0_  , \g42819/_0_  , \g42820/_0_  , \g42821/_0_  , \g42824/_0_  , \g42825/_0_  , \g42826/_0_  , \g42827/_0_  , \g42828/_0_  , \g42829/_0_  , \g42830/_0_  , \g42831/_0_  , \g42832/_0_  , \g42833/_0_  , \g42834/_0_  , \g42835/_0_  , \g42836/_0_  , \g42837/_0_  , \g42838/_0_  , \g42839/_0_  , \g42840/_0_  , \g42841/_0_  , \g42842/_0_  , \g42843/_0_  , \g42844/_0_  , \g42845/_0_  , \g42846/_0_  , \g42907/_0_  , \g42914/_0_  , \g42924/_0_  , \g42925/_0_  , \g42926/_0_  , \g42927/_0_  , \g42928/_0_  , \g42929/_0_  , \g42930/_0_  , \g42931/_0_  , \g42933/_0_  , \g42941/_0_  , \g42947/_0_  , \g42950/_0_  , \g42955/_0_  , \g42956/_0_  , \g42972/_3_  , \g42973/_3_  , \g42974/_3_  , \g43178/_0_  , \g43179/_0_  , \g43184/_0_  , \g43186/_0_  , \g43187/_0_  , \g43190/_0_  , \g43191/_0_  , \g43192/_0_  , \g43202/_0_  , \g43205/_0_  , \g43206/_0_  , \g43207/_0_  , \g43209/_2_  , \g43228/_0_  , \g43233/_0_  , \g43235/_0_  , \g43236/_0_  , \g43237/_0_  , \g43238/_0_  , \g43280/_0_  , \g43287/_0_  , \g43289/_0_  , \g43290/_0_  , \g43291/_0_  , \g43292/_0_  , \g43303/_0_  , \g43311/_0_  , \g43312/_0_  , \g43363/_0_  , \g43364/_0_  , \g43366/_0_  , \g43367/_0_  , \g43370/_0_  , \g43371/_0_  , \g43374/_0_  , \g43413/_0_  , \g43414/_0_  , \g43415/_0_  , \g43416/_0_  , \g43422/_0_  , \g43427/_0_  , \g43428/_0_  , \g43528/_1__syn_2  , \g43630/_0_  , \g43633/_3_  , \g43647/_0_  , \g43648/_0_  , \g43656/_0_  , \g43657/_0_  , \g43667/_0_  , \g43668/_0_  , \g43675/_0_  , \g43678/_0_  , \g43787/_0_  , \g44055/_0_  , \g44092/_0_  , \g44093/_0_  , \g44176/_0_  , \g44181/_0_  , \g44433/_0_  , \g44510/_0_  , \g44515/_2_  , \g44522/_0_  , \g44529/_2_  , \g44537/_2_  , \g44544/_2_  , \g44594/_0_  , \g44695/_0_  , \g44697/_0_  , \g44699/_0_  , \g44700/_0_  , \g44843/_0_  , \g44844/_0_  , \g44879/_0_  , \g44880/_0_  , \g44881/_0_  , \g44882/_0_  , \g44906/_2_  , \g44910/_0_  , \g44912/_0_  , \g44954/_0_  , \g45000/_0_  , \g45001/_0_  , \g45002/_0_  , \g45003/_0_  , \g45021/_1_  , \g45025/_0_  , \g45051/_0_  , \g45104/_0_  , \g45111/_0_  , \g45112/_0_  , \g45116/_0_  , \g45155/_0_  , \g45238/_0_  , \g45239/_0_  , \g45240/_0_  , \g45241/_0_  , \g45249/_0_  , \g45257/_0_  , \g45332/_0_  , \g45334/_0_  , \g45336/_0_  , \g45337/_0_  , \g45342/_0_  , \g45459/_0_  , \g45460/_0_  , \g45466/_0_  , \g45469/_0_  , \g45470/_0_  , \g45474/_0_  , \g45475/_0_  , \g45477/_0_  , \g45481/_0_  , \g45482/_0_  , \g45487/_0_  , \g45488/_0_  , \g45518/_3_  , \g45519/_3_  , \g45520/_3_  , \g45521/_3_  , \g45522/_3_  , \g45523/_3_  , \g45524/_3_  , \g45525/_3_  , \g45526/_3_  , \g45530/_3_  , \g45531/_3_  , \g45532/_3_  , \g45533/_3_  , \g45534/_3_  , \g45535/_3_  , \g45536/_3_  , \g45559/_3_  , \g45596/_0_  , \g45605/_0_  , \g45622/_0_  , \g45623/_0_  , \g45630/_0_  , \g45747/_0_  , \g45753/_0_  , \g45796/_0_  , \g45837/_0_  , \g45882/_0_  , \g45903/_0_  , \g45912/_0_  , \g45946/_0_  , \g45999/_0_  , \g46000/_0_  , \g46001/_0_  , \g46002/_0_  , \g46012/_0_  , \g46014/_0_  , \g46017/_0_  , \g46018/_0_  , \g46021/_0_  , \g46024/_0_  , \g46026/_0_  , \g46029/_0_  , \g46053/_0_  , \g46083/_0_  , \g46093/_0_  , \g46142/_0_  , \g46154/_1__syn_2  , \g46265/_0_  , \g46266/_0_  , \g46268/_0_  , \g46270/_0_  , \g46273/_0_  , \g46274/_0_  , \g46275/_0_  , \g46276/_0_  , \g46278/_0_  , \g46385/_0_  , \g46411/_0_  , \g46414/_0_  , \g46479/_0_  , \g46520/_0_  , \g46521/_0_  , \g46530/_0_  , \g46531/_0_  , \g46597/_0_  , \g46610/_0_  , \g46617/_0_  , \g46632/_0_  , \g46637/_0_  , \g46722/_0_  , \g46723/_0_  , \g46724/_0_  , \g46725/_0_  , \g46813/_0_  , \g46842/_0_  , \g46888/_0_  , \g46891/_0_  , \g46894/_0_  , \g46905/_0_  , \g46940/_0_  , \g46992/_0_  , \g46995/_0_  , \g47037/_3_  , \g47053/_0_  , \g47140/_0_  , \g47155/_3_  , \g47209/_0_  , \g47211/_0_  , \g47213/_0_  , \g47215/_0_  , \g47337/_0_  , \g47433/_0_  , \g47972/_0_  , \g47976/_0_  , \g48081/_0_  , \g48171/_0_  , \g48227/_0_  , \g48234/_1_  , \g48257/_1_  , \g48266/_0_  , \g48281/_0_  , \g48291/_1_  , \g48322/_0_  , \g48345/_0_  , \g48429/_0_  , \g48495/_1_  , \g48549/_0_  , \g48589/_0_  , \g48642/_0_  , \g48722/_0_  , \g48748/_0_  , \g48749/_0_  , \g48763/_0_  , \g48867/_0_  , \g48876/_0_  , \g48880/_0_  , \g49023/_0_  , \g49205/_0_  , \g49314/_0_  , \g49432/_0__syn_2  , \g49512/_0_  , \g49707/_0_  , \g49737/_0_  , \g49831/_0_  , \g49922/_1_  , \g50132/_0_  , \g51376/_0_  , \g51412/_0_  , \g51822/_0_  , \g52114/_0_  , \g52156/_0_  , \g54427/_0_  , \g54557/_0_  , \g54561/_3_  , \g55079/_0_  , \sram_adr_o[0]_pad  , \sram_adr_o[10]_pad  , \sram_adr_o[11]_pad  , \sram_adr_o[12]_pad  , \sram_adr_o[13]_pad  , \sram_adr_o[14]_pad  , \sram_adr_o[1]_pad  , \sram_adr_o[2]_pad  , \sram_adr_o[3]_pad  , \sram_adr_o[4]_pad  , \sram_adr_o[5]_pad  , \sram_adr_o[6]_pad  , \sram_adr_o[7]_pad  , \sram_adr_o[8]_pad  , \sram_adr_o[9]_pad  , \sram_data_o[0]_pad  , \sram_data_o[10]_pad  , \sram_data_o[11]_pad  , \sram_data_o[12]_pad  , \sram_data_o[13]_pad  , \sram_data_o[14]_pad  , \sram_data_o[15]_pad  , \sram_data_o[16]_pad  , \sram_data_o[17]_pad  , \sram_data_o[18]_pad  , \sram_data_o[19]_pad  , \sram_data_o[1]_pad  , \sram_data_o[20]_pad  , \sram_data_o[21]_pad  , \sram_data_o[22]_pad  , \sram_data_o[23]_pad  , \sram_data_o[24]_pad  , \sram_data_o[25]_pad  , \sram_data_o[26]_pad  , \sram_data_o[27]_pad  , \sram_data_o[28]_pad  , \sram_data_o[29]_pad  , \sram_data_o[2]_pad  , \sram_data_o[30]_pad  , \sram_data_o[31]_pad  , \sram_data_o[3]_pad  , \sram_data_o[4]_pad  , \sram_data_o[5]_pad  , \sram_data_o[6]_pad  , \sram_data_o[7]_pad  , \sram_data_o[8]_pad  , \sram_data_o[9]_pad  , sram_re_o_pad , sram_we_o_pad , \u4_utmi_vend_ctrl_r_reg[0]/P0001_reg_syn_3  , \u4_utmi_vend_ctrl_r_reg[1]/P0001_reg_syn_3  , \u4_utmi_vend_ctrl_r_reg[2]/P0001_reg_syn_3  , \u4_utmi_vend_ctrl_r_reg[3]/P0001_reg_syn_3  );
  input \DataOut_pad_o[0]_pad  ;
  input \DataOut_pad_o[1]_pad  ;
  input \DataOut_pad_o[2]_pad  ;
  input \DataOut_pad_o[3]_pad  ;
  input \DataOut_pad_o[4]_pad  ;
  input \DataOut_pad_o[5]_pad  ;
  input \DataOut_pad_o[6]_pad  ;
  input \DataOut_pad_o[7]_pad  ;
  input \LineState_pad_i[0]_pad  ;
  input \LineState_pad_i[1]_pad  ;
  input \LineState_r_reg[0]/P0001  ;
  input \LineState_r_reg[1]/P0001  ;
  input \OpMode_pad_o[1]_pad  ;
  input RxActive_pad_i_pad ;
  input RxError_pad_i_pad ;
  input RxValid_pad_i_pad ;
  input TermSel_pad_o_pad ;
  input TxReady_pad_i_pad ;
  input TxValid_pad_o_pad ;
  input VControl_Load_pad_o_pad ;
  input XcvSelect_pad_o_pad ;
  input \dma_ack_i[0]_pad  ;
  input \dma_ack_i[1]_pad  ;
  input \dma_ack_i[2]_pad  ;
  input \dma_ack_i[3]_pad  ;
  input \dma_req_o[0]_pad  ;
  input \dma_req_o[1]_pad  ;
  input \dma_req_o[2]_pad  ;
  input \dma_req_o[3]_pad  ;
  input resume_req_i_pad ;
  input \resume_req_r_reg/P0001  ;
  input rst_i_pad ;
  input \sram_data_i[0]_pad  ;
  input \sram_data_i[10]_pad  ;
  input \sram_data_i[11]_pad  ;
  input \sram_data_i[12]_pad  ;
  input \sram_data_i[13]_pad  ;
  input \sram_data_i[14]_pad  ;
  input \sram_data_i[15]_pad  ;
  input \sram_data_i[16]_pad  ;
  input \sram_data_i[17]_pad  ;
  input \sram_data_i[18]_pad  ;
  input \sram_data_i[19]_pad  ;
  input \sram_data_i[1]_pad  ;
  input \sram_data_i[20]_pad  ;
  input \sram_data_i[21]_pad  ;
  input \sram_data_i[22]_pad  ;
  input \sram_data_i[23]_pad  ;
  input \sram_data_i[24]_pad  ;
  input \sram_data_i[25]_pad  ;
  input \sram_data_i[26]_pad  ;
  input \sram_data_i[27]_pad  ;
  input \sram_data_i[28]_pad  ;
  input \sram_data_i[29]_pad  ;
  input \sram_data_i[2]_pad  ;
  input \sram_data_i[30]_pad  ;
  input \sram_data_i[31]_pad  ;
  input \sram_data_i[3]_pad  ;
  input \sram_data_i[4]_pad  ;
  input \sram_data_i[5]_pad  ;
  input \sram_data_i[6]_pad  ;
  input \sram_data_i[7]_pad  ;
  input \sram_data_i[8]_pad  ;
  input \sram_data_i[9]_pad  ;
  input susp_o_pad ;
  input \suspend_clr_wr_reg/P0001  ;
  input \u0_drive_k_r_reg/P0001  ;
  input \u0_rx_active_reg/P0001  ;
  input \u0_rx_data_reg[0]/P0001  ;
  input \u0_rx_data_reg[1]/P0001  ;
  input \u0_rx_data_reg[2]/P0001  ;
  input \u0_rx_data_reg[3]/P0001  ;
  input \u0_rx_data_reg[4]/P0001  ;
  input \u0_rx_data_reg[5]/P0001  ;
  input \u0_rx_data_reg[6]/P0001  ;
  input \u0_rx_data_reg[7]/P0001  ;
  input \u0_rx_err_reg/P0001  ;
  input \u0_rx_valid_reg/P0001  ;
  input \u0_tx_ready_reg/NET0131  ;
  input \u0_u0_T1_gt_2_5_uS_reg/P0001  ;
  input \u0_u0_T1_gt_3_0_mS_reg/P0001  ;
  input \u0_u0_T1_gt_5_0_mS_reg/P0001  ;
  input \u0_u0_T1_st_3_0_mS_reg/P0001  ;
  input \u0_u0_T2_gt_100_uS_reg/P0001  ;
  input \u0_u0_T2_gt_1_0_mS_reg/P0001  ;
  input \u0_u0_T2_wakeup_reg/P0001  ;
  input \u0_u0_chirp_cnt_is_6_reg/P0001  ;
  input \u0_u0_chirp_cnt_reg[0]/P0001  ;
  input \u0_u0_chirp_cnt_reg[1]/P0001  ;
  input \u0_u0_chirp_cnt_reg[2]/P0001  ;
  input \u0_u0_drive_k_reg/P0001  ;
  input \u0_u0_idle_cnt1_clr_reg/P0001  ;
  input \u0_u0_idle_cnt1_next_reg[0]/P0001  ;
  input \u0_u0_idle_cnt1_next_reg[1]/P0001  ;
  input \u0_u0_idle_cnt1_next_reg[2]/P0001  ;
  input \u0_u0_idle_cnt1_next_reg[3]/P0001  ;
  input \u0_u0_idle_cnt1_next_reg[4]/P0001  ;
  input \u0_u0_idle_cnt1_next_reg[5]/P0001  ;
  input \u0_u0_idle_cnt1_next_reg[6]/P0001  ;
  input \u0_u0_idle_cnt1_next_reg[7]/P0001  ;
  input \u0_u0_idle_cnt1_reg[0]/P0001  ;
  input \u0_u0_idle_cnt1_reg[1]/P0001  ;
  input \u0_u0_idle_cnt1_reg[2]/P0001  ;
  input \u0_u0_idle_cnt1_reg[3]/P0001  ;
  input \u0_u0_idle_cnt1_reg[4]/P0001  ;
  input \u0_u0_idle_cnt1_reg[5]/P0001  ;
  input \u0_u0_idle_cnt1_reg[6]/P0001  ;
  input \u0_u0_idle_cnt1_reg[7]/P0001  ;
  input \u0_u0_idle_long_reg/P0001  ;
  input \u0_u0_ls_idle_r_reg/P0001  ;
  input \u0_u0_ls_j_r_reg/P0001  ;
  input \u0_u0_ls_k_r_reg/P0001  ;
  input \u0_u0_ls_se0_r_reg/P0001  ;
  input \u0_u0_me_cnt_100_ms_reg/P0001  ;
  input \u0_u0_me_cnt_reg[0]/P0001  ;
  input \u0_u0_me_cnt_reg[1]/P0001  ;
  input \u0_u0_me_cnt_reg[2]/P0001  ;
  input \u0_u0_me_cnt_reg[3]/P0001  ;
  input \u0_u0_me_cnt_reg[4]/P0001  ;
  input \u0_u0_me_cnt_reg[5]/P0001  ;
  input \u0_u0_me_cnt_reg[6]/P0001  ;
  input \u0_u0_me_cnt_reg[7]/P0001  ;
  input \u0_u0_me_ps2_0_5_ms_reg/P0001  ;
  input \u0_u0_me_ps2_reg[0]/P0001  ;
  input \u0_u0_me_ps2_reg[1]/P0001  ;
  input \u0_u0_me_ps2_reg[2]/P0001  ;
  input \u0_u0_me_ps2_reg[3]/P0001  ;
  input \u0_u0_me_ps2_reg[4]/P0001  ;
  input \u0_u0_me_ps2_reg[5]/P0001  ;
  input \u0_u0_me_ps2_reg[6]/P0001  ;
  input \u0_u0_me_ps2_reg[7]/P0001  ;
  input \u0_u0_me_ps_2_5_us_reg/P0001  ;
  input \u0_u0_me_ps_reg[0]/P0001  ;
  input \u0_u0_me_ps_reg[1]/P0001  ;
  input \u0_u0_me_ps_reg[2]/P0001  ;
  input \u0_u0_me_ps_reg[3]/P0001  ;
  input \u0_u0_me_ps_reg[4]/P0001  ;
  input \u0_u0_me_ps_reg[5]/P0001  ;
  input \u0_u0_me_ps_reg[6]/P0001  ;
  input \u0_u0_me_ps_reg[7]/P0001  ;
  input \u0_u0_mode_hs_reg/P0001  ;
  input \u0_u0_ps_cnt_clr_reg/P0001  ;
  input \u0_u0_ps_cnt_reg[0]/P0001  ;
  input \u0_u0_ps_cnt_reg[1]/P0001  ;
  input \u0_u0_ps_cnt_reg[2]/P0001  ;
  input \u0_u0_ps_cnt_reg[3]/P0001  ;
  input \u0_u0_resume_req_s_reg/P0001  ;
  input \u0_u0_state_reg[0]/NET0131  ;
  input \u0_u0_state_reg[10]/P0001  ;
  input \u0_u0_state_reg[11]/NET0131  ;
  input \u0_u0_state_reg[12]/NET0131  ;
  input \u0_u0_state_reg[13]/NET0131  ;
  input \u0_u0_state_reg[14]/P0001  ;
  input \u0_u0_state_reg[1]/P0001  ;
  input \u0_u0_state_reg[2]/NET0131  ;
  input \u0_u0_state_reg[3]/P0001  ;
  input \u0_u0_state_reg[4]/NET0131  ;
  input \u0_u0_state_reg[5]/P0001  ;
  input \u0_u0_state_reg[6]/NET0131  ;
  input \u0_u0_state_reg[7]/NET0131  ;
  input \u0_u0_state_reg[8]/NET0131  ;
  input \u0_u0_state_reg[9]/P0001  ;
  input \u0_u0_usb_attached_reg/P0001  ;
  input \u0_u0_usb_suspend_reg/P0001  ;
  input \u1_clr_sof_time_reg/P0001  ;
  input \u1_frame_no_r_reg[0]/P0001  ;
  input \u1_frame_no_r_reg[10]/P0001  ;
  input \u1_frame_no_r_reg[1]/P0001  ;
  input \u1_frame_no_r_reg[2]/P0001  ;
  input \u1_frame_no_r_reg[3]/P0001  ;
  input \u1_frame_no_r_reg[4]/P0001  ;
  input \u1_frame_no_r_reg[5]/P0001  ;
  input \u1_frame_no_r_reg[6]/P0001  ;
  input \u1_frame_no_r_reg[7]/P0001  ;
  input \u1_frame_no_r_reg[8]/P0001  ;
  input \u1_frame_no_r_reg[9]/P0001  ;
  input \u1_frame_no_same_reg/P0001  ;
  input \u1_hms_clk_reg/P0001  ;
  input \u1_hms_cnt_reg[0]/P0001  ;
  input \u1_hms_cnt_reg[1]/P0001  ;
  input \u1_hms_cnt_reg[2]/P0001  ;
  input \u1_hms_cnt_reg[3]/P0001  ;
  input \u1_hms_cnt_reg[4]/P0001  ;
  input \u1_mfm_cnt_reg[0]/P0001  ;
  input \u1_mfm_cnt_reg[1]/P0001  ;
  input \u1_mfm_cnt_reg[2]/P0001  ;
  input \u1_mfm_cnt_reg[3]/P0001  ;
  input \u1_sof_time_reg[0]/P0001  ;
  input \u1_sof_time_reg[10]/P0001  ;
  input \u1_sof_time_reg[11]/P0001  ;
  input \u1_sof_time_reg[1]/P0001  ;
  input \u1_sof_time_reg[2]/P0001  ;
  input \u1_sof_time_reg[3]/P0001  ;
  input \u1_sof_time_reg[4]/P0001  ;
  input \u1_sof_time_reg[5]/P0001  ;
  input \u1_sof_time_reg[6]/P0001  ;
  input \u1_sof_time_reg[7]/P0001  ;
  input \u1_sof_time_reg[8]/P0001  ;
  input \u1_sof_time_reg[9]/P0001  ;
  input \u1_u0_crc16_sum_reg[0]/P0001  ;
  input \u1_u0_crc16_sum_reg[10]/P0001  ;
  input \u1_u0_crc16_sum_reg[11]/P0001  ;
  input \u1_u0_crc16_sum_reg[12]/P0001  ;
  input \u1_u0_crc16_sum_reg[13]/P0001  ;
  input \u1_u0_crc16_sum_reg[14]/P0001  ;
  input \u1_u0_crc16_sum_reg[15]/P0001  ;
  input \u1_u0_crc16_sum_reg[1]/P0001  ;
  input \u1_u0_crc16_sum_reg[2]/P0001  ;
  input \u1_u0_crc16_sum_reg[3]/P0001  ;
  input \u1_u0_crc16_sum_reg[4]/P0001  ;
  input \u1_u0_crc16_sum_reg[5]/P0001  ;
  input \u1_u0_crc16_sum_reg[6]/P0001  ;
  input \u1_u0_crc16_sum_reg[7]/P0001  ;
  input \u1_u0_crc16_sum_reg[8]/P0001  ;
  input \u1_u0_crc16_sum_reg[9]/P0001  ;
  input \u1_u0_data_valid0_reg/P0001  ;
  input \u1_u0_pid_reg[0]/NET0131  ;
  input \u1_u0_pid_reg[1]/NET0131  ;
  input \u1_u0_pid_reg[2]/NET0131  ;
  input \u1_u0_pid_reg[3]/NET0131  ;
  input \u1_u0_pid_reg[4]/P0001  ;
  input \u1_u0_pid_reg[5]/P0001  ;
  input \u1_u0_pid_reg[6]/P0001  ;
  input \u1_u0_pid_reg[7]/P0001  ;
  input \u1_u0_rx_active_r_reg/P0001  ;
  input \u1_u0_rxv1_reg/P0001  ;
  input \u1_u0_rxv2_reg/P0001  ;
  input \u1_u0_state_reg[0]/P0001  ;
  input \u1_u0_state_reg[1]/P0001  ;
  input \u1_u0_state_reg[2]/P0001  ;
  input \u1_u0_state_reg[3]/P0001  ;
  input \u1_u0_token0_reg[0]/NET0131  ;
  input \u1_u0_token0_reg[1]/P0001  ;
  input \u1_u0_token0_reg[2]/NET0131  ;
  input \u1_u0_token0_reg[3]/NET0131  ;
  input \u1_u0_token0_reg[4]/P0001  ;
  input \u1_u0_token0_reg[5]/NET0131  ;
  input \u1_u0_token0_reg[6]/P0001  ;
  input \u1_u0_token0_reg[7]/P0001  ;
  input \u1_u0_token1_reg[0]/P0001  ;
  input \u1_u0_token1_reg[1]/P0001  ;
  input \u1_u0_token1_reg[2]/P0001  ;
  input \u1_u0_token1_reg[3]/P0001  ;
  input \u1_u0_token1_reg[4]/P0001  ;
  input \u1_u0_token1_reg[5]/P0001  ;
  input \u1_u0_token1_reg[6]/P0001  ;
  input \u1_u0_token1_reg[7]/P0001  ;
  input \u1_u0_token_valid_r1_reg/P0001  ;
  input \u1_u0_token_valid_str1_reg/P0001  ;
  input \u1_u1_crc16_reg[0]/P0001  ;
  input \u1_u1_crc16_reg[10]/P0001  ;
  input \u1_u1_crc16_reg[11]/P0001  ;
  input \u1_u1_crc16_reg[12]/P0001  ;
  input \u1_u1_crc16_reg[13]/P0001  ;
  input \u1_u1_crc16_reg[14]/P0001  ;
  input \u1_u1_crc16_reg[15]/P0001  ;
  input \u1_u1_crc16_reg[1]/P0001  ;
  input \u1_u1_crc16_reg[2]/P0001  ;
  input \u1_u1_crc16_reg[3]/P0001  ;
  input \u1_u1_crc16_reg[4]/P0001  ;
  input \u1_u1_crc16_reg[5]/P0001  ;
  input \u1_u1_crc16_reg[6]/P0001  ;
  input \u1_u1_crc16_reg[7]/P0001  ;
  input \u1_u1_crc16_reg[8]/P0001  ;
  input \u1_u1_crc16_reg[9]/P0001  ;
  input \u1_u1_send_data_r2_reg/P0001  ;
  input \u1_u1_send_data_r_reg/P0001  ;
  input \u1_u1_send_token_r_reg/P0001  ;
  input \u1_u1_send_zero_length_r_reg/P0001  ;
  input \u1_u1_state_reg[0]/NET0131  ;
  input \u1_u1_state_reg[1]/NET0131  ;
  input \u1_u1_state_reg[2]/NET0131  ;
  input \u1_u1_state_reg[3]/NET0131  ;
  input \u1_u1_state_reg[4]/NET0131  ;
  input \u1_u1_tx_first_r_reg/P0001  ;
  input \u1_u1_tx_valid_r_reg/NET0131  ;
  input \u1_u1_zero_length_r_reg/P0001  ;
  input \u1_u2_adr_cb_reg[0]/NET0131  ;
  input \u1_u2_adr_cb_reg[1]/NET0131  ;
  input \u1_u2_adr_cb_reg[2]/NET0131  ;
  input \u1_u2_adr_cw_reg[0]/NET0131  ;
  input \u1_u2_adr_cw_reg[10]/P0001  ;
  input \u1_u2_adr_cw_reg[11]/P0001  ;
  input \u1_u2_adr_cw_reg[12]/P0001  ;
  input \u1_u2_adr_cw_reg[13]/P0001  ;
  input \u1_u2_adr_cw_reg[14]/P0001  ;
  input \u1_u2_adr_cw_reg[1]/P0001  ;
  input \u1_u2_adr_cw_reg[2]/P0001  ;
  input \u1_u2_adr_cw_reg[3]/NET0131  ;
  input \u1_u2_adr_cw_reg[4]/P0001  ;
  input \u1_u2_adr_cw_reg[5]/NET0131  ;
  input \u1_u2_adr_cw_reg[6]/NET0131  ;
  input \u1_u2_adr_cw_reg[7]/NET0131  ;
  input \u1_u2_adr_cw_reg[8]/P0001  ;
  input \u1_u2_adr_cw_reg[9]/NET0131  ;
  input \u1_u2_dout_r_reg[0]/P0001  ;
  input \u1_u2_dout_r_reg[10]/P0001  ;
  input \u1_u2_dout_r_reg[11]/P0001  ;
  input \u1_u2_dout_r_reg[12]/P0001  ;
  input \u1_u2_dout_r_reg[13]/P0001  ;
  input \u1_u2_dout_r_reg[14]/P0001  ;
  input \u1_u2_dout_r_reg[15]/P0001  ;
  input \u1_u2_dout_r_reg[16]/P0001  ;
  input \u1_u2_dout_r_reg[17]/P0001  ;
  input \u1_u2_dout_r_reg[18]/P0001  ;
  input \u1_u2_dout_r_reg[19]/P0001  ;
  input \u1_u2_dout_r_reg[1]/P0001  ;
  input \u1_u2_dout_r_reg[20]/P0001  ;
  input \u1_u2_dout_r_reg[21]/P0001  ;
  input \u1_u2_dout_r_reg[22]/P0001  ;
  input \u1_u2_dout_r_reg[23]/P0001  ;
  input \u1_u2_dout_r_reg[24]/P0001  ;
  input \u1_u2_dout_r_reg[25]/P0001  ;
  input \u1_u2_dout_r_reg[26]/P0001  ;
  input \u1_u2_dout_r_reg[27]/P0001  ;
  input \u1_u2_dout_r_reg[28]/P0001  ;
  input \u1_u2_dout_r_reg[29]/P0001  ;
  input \u1_u2_dout_r_reg[2]/P0001  ;
  input \u1_u2_dout_r_reg[30]/P0001  ;
  input \u1_u2_dout_r_reg[31]/P0001  ;
  input \u1_u2_dout_r_reg[3]/P0001  ;
  input \u1_u2_dout_r_reg[4]/P0001  ;
  input \u1_u2_dout_r_reg[5]/P0001  ;
  input \u1_u2_dout_r_reg[6]/P0001  ;
  input \u1_u2_dout_r_reg[7]/P0001  ;
  input \u1_u2_dout_r_reg[8]/P0001  ;
  input \u1_u2_dout_r_reg[9]/P0001  ;
  input \u1_u2_dtmp_r_reg[0]/P0001  ;
  input \u1_u2_dtmp_r_reg[10]/P0001  ;
  input \u1_u2_dtmp_r_reg[11]/P0001  ;
  input \u1_u2_dtmp_r_reg[12]/P0001  ;
  input \u1_u2_dtmp_r_reg[13]/P0001  ;
  input \u1_u2_dtmp_r_reg[14]/P0001  ;
  input \u1_u2_dtmp_r_reg[15]/P0001  ;
  input \u1_u2_dtmp_r_reg[16]/P0001  ;
  input \u1_u2_dtmp_r_reg[17]/P0001  ;
  input \u1_u2_dtmp_r_reg[18]/P0001  ;
  input \u1_u2_dtmp_r_reg[19]/P0001  ;
  input \u1_u2_dtmp_r_reg[1]/P0001  ;
  input \u1_u2_dtmp_r_reg[20]/P0001  ;
  input \u1_u2_dtmp_r_reg[21]/P0001  ;
  input \u1_u2_dtmp_r_reg[22]/P0001  ;
  input \u1_u2_dtmp_r_reg[23]/P0001  ;
  input \u1_u2_dtmp_r_reg[24]/P0001  ;
  input \u1_u2_dtmp_r_reg[25]/P0001  ;
  input \u1_u2_dtmp_r_reg[26]/P0001  ;
  input \u1_u2_dtmp_r_reg[27]/P0001  ;
  input \u1_u2_dtmp_r_reg[28]/P0001  ;
  input \u1_u2_dtmp_r_reg[29]/P0001  ;
  input \u1_u2_dtmp_r_reg[2]/P0001  ;
  input \u1_u2_dtmp_r_reg[30]/P0001  ;
  input \u1_u2_dtmp_r_reg[31]/P0001  ;
  input \u1_u2_dtmp_r_reg[3]/P0001  ;
  input \u1_u2_dtmp_r_reg[4]/P0001  ;
  input \u1_u2_dtmp_r_reg[5]/P0001  ;
  input \u1_u2_dtmp_r_reg[6]/P0001  ;
  input \u1_u2_dtmp_r_reg[7]/P0001  ;
  input \u1_u2_dtmp_r_reg[8]/P0001  ;
  input \u1_u2_dtmp_r_reg[9]/P0001  ;
  input \u1_u2_dtmp_sel_r_reg/P0001  ;
  input \u1_u2_idma_done_reg/P0001  ;
  input \u1_u2_last_buf_adr_reg[0]/P0001  ;
  input \u1_u2_last_buf_adr_reg[10]/P0001  ;
  input \u1_u2_last_buf_adr_reg[11]/P0001  ;
  input \u1_u2_last_buf_adr_reg[12]/P0001  ;
  input \u1_u2_last_buf_adr_reg[13]/P0001  ;
  input \u1_u2_last_buf_adr_reg[14]/P0001  ;
  input \u1_u2_last_buf_adr_reg[1]/P0001  ;
  input \u1_u2_last_buf_adr_reg[2]/P0001  ;
  input \u1_u2_last_buf_adr_reg[3]/P0001  ;
  input \u1_u2_last_buf_adr_reg[4]/P0001  ;
  input \u1_u2_last_buf_adr_reg[5]/P0001  ;
  input \u1_u2_last_buf_adr_reg[6]/P0001  ;
  input \u1_u2_last_buf_adr_reg[7]/P0001  ;
  input \u1_u2_last_buf_adr_reg[8]/P0001  ;
  input \u1_u2_last_buf_adr_reg[9]/P0001  ;
  input \u1_u2_mack_r_reg/P0001  ;
  input \u1_u2_mwe_reg/P0001  ;
  input \u1_u2_rd_buf0_reg[0]/NET0131  ;
  input \u1_u2_rd_buf0_reg[10]/NET0131  ;
  input \u1_u2_rd_buf0_reg[11]/NET0131  ;
  input \u1_u2_rd_buf0_reg[12]/P0001  ;
  input \u1_u2_rd_buf0_reg[13]/P0001  ;
  input \u1_u2_rd_buf0_reg[14]/P0001  ;
  input \u1_u2_rd_buf0_reg[15]/P0001  ;
  input \u1_u2_rd_buf0_reg[16]/NET0131  ;
  input \u1_u2_rd_buf0_reg[17]/NET0131  ;
  input \u1_u2_rd_buf0_reg[18]/NET0131  ;
  input \u1_u2_rd_buf0_reg[19]/NET0131  ;
  input \u1_u2_rd_buf0_reg[1]/NET0131  ;
  input \u1_u2_rd_buf0_reg[20]/P0001  ;
  input \u1_u2_rd_buf0_reg[21]/P0001  ;
  input \u1_u2_rd_buf0_reg[22]/P0001  ;
  input \u1_u2_rd_buf0_reg[23]/P0001  ;
  input \u1_u2_rd_buf0_reg[24]/NET0131  ;
  input \u1_u2_rd_buf0_reg[25]/NET0131  ;
  input \u1_u2_rd_buf0_reg[26]/NET0131  ;
  input \u1_u2_rd_buf0_reg[27]/NET0131  ;
  input \u1_u2_rd_buf0_reg[28]/P0001  ;
  input \u1_u2_rd_buf0_reg[29]/P0001  ;
  input \u1_u2_rd_buf0_reg[2]/NET0131  ;
  input \u1_u2_rd_buf0_reg[30]/P0001  ;
  input \u1_u2_rd_buf0_reg[31]/P0001  ;
  input \u1_u2_rd_buf0_reg[3]/NET0131  ;
  input \u1_u2_rd_buf0_reg[4]/P0001  ;
  input \u1_u2_rd_buf0_reg[5]/P0001  ;
  input \u1_u2_rd_buf0_reg[6]/P0001  ;
  input \u1_u2_rd_buf0_reg[7]/P0001  ;
  input \u1_u2_rd_buf0_reg[8]/NET0131  ;
  input \u1_u2_rd_buf0_reg[9]/NET0131  ;
  input \u1_u2_rd_buf1_reg[0]/NET0131  ;
  input \u1_u2_rd_buf1_reg[10]/NET0131  ;
  input \u1_u2_rd_buf1_reg[11]/NET0131  ;
  input \u1_u2_rd_buf1_reg[12]/P0001  ;
  input \u1_u2_rd_buf1_reg[13]/P0001  ;
  input \u1_u2_rd_buf1_reg[14]/P0001  ;
  input \u1_u2_rd_buf1_reg[15]/P0001  ;
  input \u1_u2_rd_buf1_reg[16]/NET0131  ;
  input \u1_u2_rd_buf1_reg[17]/NET0131  ;
  input \u1_u2_rd_buf1_reg[18]/NET0131  ;
  input \u1_u2_rd_buf1_reg[19]/NET0131  ;
  input \u1_u2_rd_buf1_reg[1]/NET0131  ;
  input \u1_u2_rd_buf1_reg[20]/P0001  ;
  input \u1_u2_rd_buf1_reg[21]/P0001  ;
  input \u1_u2_rd_buf1_reg[22]/P0001  ;
  input \u1_u2_rd_buf1_reg[23]/P0001  ;
  input \u1_u2_rd_buf1_reg[24]/NET0131  ;
  input \u1_u2_rd_buf1_reg[25]/NET0131  ;
  input \u1_u2_rd_buf1_reg[26]/NET0131  ;
  input \u1_u2_rd_buf1_reg[27]/NET0131  ;
  input \u1_u2_rd_buf1_reg[28]/P0001  ;
  input \u1_u2_rd_buf1_reg[29]/P0001  ;
  input \u1_u2_rd_buf1_reg[2]/NET0131  ;
  input \u1_u2_rd_buf1_reg[30]/P0001  ;
  input \u1_u2_rd_buf1_reg[31]/P0001  ;
  input \u1_u2_rd_buf1_reg[3]/NET0131  ;
  input \u1_u2_rd_buf1_reg[4]/P0001  ;
  input \u1_u2_rd_buf1_reg[5]/P0001  ;
  input \u1_u2_rd_buf1_reg[6]/P0001  ;
  input \u1_u2_rd_buf1_reg[7]/P0001  ;
  input \u1_u2_rd_buf1_reg[8]/NET0131  ;
  input \u1_u2_rd_buf1_reg[9]/NET0131  ;
  input \u1_u2_rx_data_done_r2_reg/P0001  ;
  input \u1_u2_rx_data_done_r_reg/P0001  ;
  input \u1_u2_rx_data_st_r_reg[0]/P0001  ;
  input \u1_u2_rx_data_st_r_reg[1]/P0001  ;
  input \u1_u2_rx_data_st_r_reg[2]/P0001  ;
  input \u1_u2_rx_data_st_r_reg[3]/P0001  ;
  input \u1_u2_rx_data_st_r_reg[4]/P0001  ;
  input \u1_u2_rx_data_st_r_reg[5]/P0001  ;
  input \u1_u2_rx_data_st_r_reg[6]/P0001  ;
  input \u1_u2_rx_data_st_r_reg[7]/P0001  ;
  input \u1_u2_rx_data_valid_r_reg/NET0131  ;
  input \u1_u2_rx_dma_en_r_reg/P0001  ;
  input \u1_u2_send_data_r_reg/NET0131  ;
  input \u1_u2_sizd_c_reg[0]/P0001  ;
  input \u1_u2_sizd_c_reg[10]/P0001  ;
  input \u1_u2_sizd_c_reg[11]/P0001  ;
  input \u1_u2_sizd_c_reg[12]/P0001  ;
  input \u1_u2_sizd_c_reg[13]/P0001  ;
  input \u1_u2_sizd_c_reg[1]/P0001  ;
  input \u1_u2_sizd_c_reg[2]/P0001  ;
  input \u1_u2_sizd_c_reg[3]/P0001  ;
  input \u1_u2_sizd_c_reg[4]/P0001  ;
  input \u1_u2_sizd_c_reg[5]/P0001  ;
  input \u1_u2_sizd_c_reg[6]/P0001  ;
  input \u1_u2_sizd_c_reg[7]/P0001  ;
  input \u1_u2_sizd_c_reg[8]/P0001  ;
  input \u1_u2_sizd_c_reg[9]/P0001  ;
  input \u1_u2_sizd_is_zero_reg/P0001  ;
  input \u1_u2_sizu_c_reg[0]/P0001  ;
  input \u1_u2_sizu_c_reg[10]/P0001  ;
  input \u1_u2_sizu_c_reg[1]/P0001  ;
  input \u1_u2_sizu_c_reg[2]/P0001  ;
  input \u1_u2_sizu_c_reg[3]/P0001  ;
  input \u1_u2_sizu_c_reg[4]/P0001  ;
  input \u1_u2_sizu_c_reg[5]/P0001  ;
  input \u1_u2_sizu_c_reg[6]/P0001  ;
  input \u1_u2_sizu_c_reg[7]/P0001  ;
  input \u1_u2_sizu_c_reg[8]/NET0131  ;
  input \u1_u2_sizu_c_reg[9]/P0001  ;
  input \u1_u2_state_reg[0]/P0001  ;
  input \u1_u2_state_reg[1]/NET0131  ;
  input \u1_u2_state_reg[2]/NET0131  ;
  input \u1_u2_state_reg[3]/NET0131  ;
  input \u1_u2_state_reg[4]/NET0131  ;
  input \u1_u2_state_reg[5]/NET0131  ;
  input \u1_u2_state_reg[6]/NET0131  ;
  input \u1_u2_state_reg[7]/NET0131  ;
  input \u1_u2_tx_dma_en_r_reg/P0001  ;
  input \u1_u2_word_done_r_reg/P0001  ;
  input \u1_u2_word_done_reg/NET0131  ;
  input \u1_u2_wr_done_reg/P0001  ;
  input \u1_u2_wr_last_reg/P0001  ;
  input \u1_u3_abort_reg/P0001  ;
  input \u1_u3_adr_r_reg[0]/P0001  ;
  input \u1_u3_adr_r_reg[10]/P0001  ;
  input \u1_u3_adr_r_reg[11]/P0001  ;
  input \u1_u3_adr_r_reg[12]/P0001  ;
  input \u1_u3_adr_r_reg[13]/P0001  ;
  input \u1_u3_adr_r_reg[14]/P0001  ;
  input \u1_u3_adr_r_reg[15]/P0001  ;
  input \u1_u3_adr_r_reg[16]/P0001  ;
  input \u1_u3_adr_r_reg[1]/P0001  ;
  input \u1_u3_adr_r_reg[2]/P0001  ;
  input \u1_u3_adr_r_reg[3]/P0001  ;
  input \u1_u3_adr_r_reg[4]/P0001  ;
  input \u1_u3_adr_r_reg[5]/P0001  ;
  input \u1_u3_adr_r_reg[6]/P0001  ;
  input \u1_u3_adr_r_reg[7]/P0001  ;
  input \u1_u3_adr_r_reg[8]/P0001  ;
  input \u1_u3_adr_r_reg[9]/P0001  ;
  input \u1_u3_adr_reg[0]/P0001  ;
  input \u1_u3_adr_reg[10]/P0001  ;
  input \u1_u3_adr_reg[11]/P0001  ;
  input \u1_u3_adr_reg[12]/P0001  ;
  input \u1_u3_adr_reg[13]/P0001  ;
  input \u1_u3_adr_reg[14]/P0001  ;
  input \u1_u3_adr_reg[15]/P0001  ;
  input \u1_u3_adr_reg[16]/P0001  ;
  input \u1_u3_adr_reg[1]/P0001  ;
  input \u1_u3_adr_reg[2]/P0001  ;
  input \u1_u3_adr_reg[3]/P0001  ;
  input \u1_u3_adr_reg[4]/P0001  ;
  input \u1_u3_adr_reg[5]/P0001  ;
  input \u1_u3_adr_reg[6]/P0001  ;
  input \u1_u3_adr_reg[7]/P0001  ;
  input \u1_u3_adr_reg[8]/P0001  ;
  input \u1_u3_adr_reg[9]/P0001  ;
  input \u1_u3_buf0_na_reg/NET0131  ;
  input \u1_u3_buf0_not_aloc_reg/P0001  ;
  input \u1_u3_buf0_rl_reg/P0001  ;
  input \u1_u3_buf0_set_reg/P0001  ;
  input \u1_u3_buf0_st_max_reg/P0001  ;
  input \u1_u3_buf1_na_reg/NET0131  ;
  input \u1_u3_buf1_not_aloc_reg/P0001  ;
  input \u1_u3_buf1_set_reg/P0001  ;
  input \u1_u3_buf1_st_max_reg/P0001  ;
  input \u1_u3_buffer_done_reg/P0001  ;
  input \u1_u3_buffer_empty_reg/P0001  ;
  input \u1_u3_buffer_full_reg/P0001  ;
  input \u1_u3_buffer_overflow_reg/P0001  ;
  input \u1_u3_idin_reg[0]/P0001  ;
  input \u1_u3_idin_reg[10]/P0001  ;
  input \u1_u3_idin_reg[11]/P0001  ;
  input \u1_u3_idin_reg[12]/P0001  ;
  input \u1_u3_idin_reg[13]/P0001  ;
  input \u1_u3_idin_reg[14]/P0001  ;
  input \u1_u3_idin_reg[15]/P0001  ;
  input \u1_u3_idin_reg[16]/P0001  ;
  input \u1_u3_idin_reg[17]/P0001  ;
  input \u1_u3_idin_reg[18]/P0001  ;
  input \u1_u3_idin_reg[19]/P0001  ;
  input \u1_u3_idin_reg[1]/P0001  ;
  input \u1_u3_idin_reg[20]/P0001  ;
  input \u1_u3_idin_reg[21]/P0001  ;
  input \u1_u3_idin_reg[22]/P0001  ;
  input \u1_u3_idin_reg[23]/P0001  ;
  input \u1_u3_idin_reg[24]/P0001  ;
  input \u1_u3_idin_reg[25]/P0001  ;
  input \u1_u3_idin_reg[26]/P0001  ;
  input \u1_u3_idin_reg[27]/P0001  ;
  input \u1_u3_idin_reg[28]/P0001  ;
  input \u1_u3_idin_reg[29]/P0001  ;
  input \u1_u3_idin_reg[2]/P0001  ;
  input \u1_u3_idin_reg[30]/P0001  ;
  input \u1_u3_idin_reg[31]/P0001  ;
  input \u1_u3_idin_reg[3]/P0001  ;
  input \u1_u3_idin_reg[4]/P0001  ;
  input \u1_u3_idin_reg[5]/P0001  ;
  input \u1_u3_idin_reg[6]/P0001  ;
  input \u1_u3_idin_reg[7]/P0001  ;
  input \u1_u3_idin_reg[8]/P0001  ;
  input \u1_u3_idin_reg[9]/P0001  ;
  input \u1_u3_in_token_reg/NET0131  ;
  input \u1_u3_int_seqerr_set_reg/P0001  ;
  input \u1_u3_int_upid_set_reg/P0001  ;
  input \u1_u3_match_r_reg/P0001  ;
  input \u1_u3_new_size_reg[0]/P0001  ;
  input \u1_u3_new_size_reg[10]/P0001  ;
  input \u1_u3_new_size_reg[11]/P0001  ;
  input \u1_u3_new_size_reg[12]/P0001  ;
  input \u1_u3_new_size_reg[13]/P0001  ;
  input \u1_u3_new_size_reg[1]/P0001  ;
  input \u1_u3_new_size_reg[2]/P0001  ;
  input \u1_u3_new_size_reg[3]/P0001  ;
  input \u1_u3_new_size_reg[4]/P0001  ;
  input \u1_u3_new_size_reg[5]/P0001  ;
  input \u1_u3_new_size_reg[6]/P0001  ;
  input \u1_u3_new_size_reg[7]/P0001  ;
  input \u1_u3_new_size_reg[8]/P0001  ;
  input \u1_u3_new_size_reg[9]/P0001  ;
  input \u1_u3_new_sizeb_reg[0]/P0001  ;
  input \u1_u3_new_sizeb_reg[10]/P0001  ;
  input \u1_u3_new_sizeb_reg[1]/P0001  ;
  input \u1_u3_new_sizeb_reg[2]/P0001  ;
  input \u1_u3_new_sizeb_reg[3]/P0001  ;
  input \u1_u3_new_sizeb_reg[4]/P0001  ;
  input \u1_u3_new_sizeb_reg[5]/P0001  ;
  input \u1_u3_new_sizeb_reg[6]/P0001  ;
  input \u1_u3_new_sizeb_reg[7]/P0001  ;
  input \u1_u3_new_sizeb_reg[8]/P0001  ;
  input \u1_u3_new_sizeb_reg[9]/P0001  ;
  input \u1_u3_next_dpid_reg[0]/P0001  ;
  input \u1_u3_next_dpid_reg[1]/P0001  ;
  input \u1_u3_no_bufs0_reg/P0001  ;
  input \u1_u3_no_bufs1_reg/P0001  ;
  input \u1_u3_out_to_small_r_reg/P0001  ;
  input \u1_u3_out_to_small_reg/P0001  ;
  input \u1_u3_out_token_reg/NET0131  ;
  input \u1_u3_pid_IN_r_reg/P0001  ;
  input \u1_u3_pid_OUT_r_reg/P0001  ;
  input \u1_u3_pid_PING_r_reg/P0001  ;
  input \u1_u3_pid_SETUP_r_reg/P0001  ;
  input \u1_u3_pid_seq_err_reg/P0001  ;
  input \u1_u3_rx_ack_to_clr_reg/P0001  ;
  input \u1_u3_rx_ack_to_cnt_reg[0]/P0001  ;
  input \u1_u3_rx_ack_to_cnt_reg[1]/P0001  ;
  input \u1_u3_rx_ack_to_cnt_reg[2]/P0001  ;
  input \u1_u3_rx_ack_to_cnt_reg[3]/P0001  ;
  input \u1_u3_rx_ack_to_cnt_reg[4]/P0001  ;
  input \u1_u3_rx_ack_to_cnt_reg[5]/P0001  ;
  input \u1_u3_rx_ack_to_cnt_reg[6]/P0001  ;
  input \u1_u3_rx_ack_to_cnt_reg[7]/P0001  ;
  input \u1_u3_rx_ack_to_reg/P0001  ;
  input \u1_u3_send_token_reg/P0001  ;
  input \u1_u3_setup_token_reg/P0001  ;
  input \u1_u3_size_next_r_reg[0]/P0001  ;
  input \u1_u3_size_next_r_reg[10]/P0001  ;
  input \u1_u3_size_next_r_reg[1]/P0001  ;
  input \u1_u3_size_next_r_reg[2]/P0001  ;
  input \u1_u3_size_next_r_reg[3]/P0001  ;
  input \u1_u3_size_next_r_reg[4]/P0001  ;
  input \u1_u3_size_next_r_reg[5]/P0001  ;
  input \u1_u3_size_next_r_reg[6]/P0001  ;
  input \u1_u3_size_next_r_reg[7]/P0001  ;
  input \u1_u3_size_next_r_reg[8]/P0001  ;
  input \u1_u3_size_next_r_reg[9]/P0001  ;
  input \u1_u3_state_reg[0]/P0001  ;
  input \u1_u3_state_reg[1]/P0001  ;
  input \u1_u3_state_reg[2]/P0001  ;
  input \u1_u3_state_reg[3]/P0001  ;
  input \u1_u3_state_reg[4]/P0001  ;
  input \u1_u3_state_reg[5]/P0001  ;
  input \u1_u3_state_reg[6]/P0001  ;
  input \u1_u3_state_reg[7]/P0001  ;
  input \u1_u3_state_reg[8]/P0001  ;
  input \u1_u3_state_reg[9]/P0001  ;
  input \u1_u3_this_dpid_reg[0]/P0001  ;
  input \u1_u3_this_dpid_reg[1]/P0001  ;
  input \u1_u3_to_large_reg/P0001  ;
  input \u1_u3_to_small_reg/P0001  ;
  input \u1_u3_token_pid_sel_reg[0]/P0001  ;
  input \u1_u3_token_pid_sel_reg[1]/P0001  ;
  input \u1_u3_tx_data_to_cnt_reg[0]/P0001  ;
  input \u1_u3_tx_data_to_cnt_reg[1]/P0001  ;
  input \u1_u3_tx_data_to_cnt_reg[2]/P0001  ;
  input \u1_u3_tx_data_to_cnt_reg[3]/P0001  ;
  input \u1_u3_tx_data_to_cnt_reg[4]/P0001  ;
  input \u1_u3_tx_data_to_cnt_reg[5]/P0001  ;
  input \u1_u3_tx_data_to_cnt_reg[6]/P0001  ;
  input \u1_u3_tx_data_to_cnt_reg[7]/P0001  ;
  input \u1_u3_tx_data_to_reg/P0001  ;
  input \u1_u3_uc_bsel_set_reg/P0001  ;
  input \u2_wack_r_reg/P0001  ;
  input \u4_attach_r1_reg/P0001  ;
  input \u4_attach_r_reg/P0001  ;
  input \u4_buf0_reg[0]/P0001  ;
  input \u4_buf0_reg[10]/P0001  ;
  input \u4_buf0_reg[11]/P0001  ;
  input \u4_buf0_reg[12]/P0001  ;
  input \u4_buf0_reg[13]/P0001  ;
  input \u4_buf0_reg[14]/P0001  ;
  input \u4_buf0_reg[15]/P0001  ;
  input \u4_buf0_reg[16]/P0001  ;
  input \u4_buf0_reg[17]/NET0131  ;
  input \u4_buf0_reg[18]/P0001  ;
  input \u4_buf0_reg[19]/NET0131  ;
  input \u4_buf0_reg[1]/P0001  ;
  input \u4_buf0_reg[20]/NET0131  ;
  input \u4_buf0_reg[21]/NET0131  ;
  input \u4_buf0_reg[22]/NET0131  ;
  input \u4_buf0_reg[23]/NET0131  ;
  input \u4_buf0_reg[24]/NET0131  ;
  input \u4_buf0_reg[25]/NET0131  ;
  input \u4_buf0_reg[26]/NET0131  ;
  input \u4_buf0_reg[27]/P0001  ;
  input \u4_buf0_reg[28]/P0001  ;
  input \u4_buf0_reg[29]/P0001  ;
  input \u4_buf0_reg[2]/P0001  ;
  input \u4_buf0_reg[30]/P0001  ;
  input \u4_buf0_reg[31]/P0001  ;
  input \u4_buf0_reg[3]/P0001  ;
  input \u4_buf0_reg[4]/P0001  ;
  input \u4_buf0_reg[5]/P0001  ;
  input \u4_buf0_reg[6]/P0001  ;
  input \u4_buf0_reg[7]/P0001  ;
  input \u4_buf0_reg[8]/P0001  ;
  input \u4_buf0_reg[9]/P0001  ;
  input \u4_buf1_reg[0]/P0001  ;
  input \u4_buf1_reg[10]/P0001  ;
  input \u4_buf1_reg[11]/P0001  ;
  input \u4_buf1_reg[12]/P0001  ;
  input \u4_buf1_reg[13]/P0001  ;
  input \u4_buf1_reg[14]/P0001  ;
  input \u4_buf1_reg[15]/P0001  ;
  input \u4_buf1_reg[16]/P0001  ;
  input \u4_buf1_reg[17]/NET0131  ;
  input \u4_buf1_reg[18]/P0001  ;
  input \u4_buf1_reg[19]/NET0131  ;
  input \u4_buf1_reg[1]/P0001  ;
  input \u4_buf1_reg[20]/NET0131  ;
  input \u4_buf1_reg[21]/NET0131  ;
  input \u4_buf1_reg[22]/NET0131  ;
  input \u4_buf1_reg[23]/NET0131  ;
  input \u4_buf1_reg[24]/NET0131  ;
  input \u4_buf1_reg[25]/NET0131  ;
  input \u4_buf1_reg[26]/NET0131  ;
  input \u4_buf1_reg[27]/P0001  ;
  input \u4_buf1_reg[28]/P0001  ;
  input \u4_buf1_reg[29]/P0001  ;
  input \u4_buf1_reg[2]/P0001  ;
  input \u4_buf1_reg[30]/P0001  ;
  input \u4_buf1_reg[31]/P0001  ;
  input \u4_buf1_reg[3]/P0001  ;
  input \u4_buf1_reg[4]/P0001  ;
  input \u4_buf1_reg[5]/P0001  ;
  input \u4_buf1_reg[6]/P0001  ;
  input \u4_buf1_reg[7]/P0001  ;
  input \u4_buf1_reg[8]/P0001  ;
  input \u4_buf1_reg[9]/P0001  ;
  input \u4_crc5_err_r_reg/P0001  ;
  input \u4_csr_reg[0]/P0001  ;
  input \u4_csr_reg[10]/P0001  ;
  input \u4_csr_reg[11]/P0001  ;
  input \u4_csr_reg[12]/P0001  ;
  input \u4_csr_reg[15]/NET0131  ;
  input \u4_csr_reg[16]/P0001  ;
  input \u4_csr_reg[17]/P0001  ;
  input \u4_csr_reg[1]/P0001  ;
  input \u4_csr_reg[22]/P0001  ;
  input \u4_csr_reg[23]/P0001  ;
  input \u4_csr_reg[24]/P0001  ;
  input \u4_csr_reg[25]/P0001  ;
  input \u4_csr_reg[26]/NET0131  ;
  input \u4_csr_reg[27]/NET0131  ;
  input \u4_csr_reg[28]/P0001  ;
  input \u4_csr_reg[29]/P0001  ;
  input \u4_csr_reg[2]/NET0131  ;
  input \u4_csr_reg[30]/NET0131  ;
  input \u4_csr_reg[31]/P0001  ;
  input \u4_csr_reg[3]/P0001  ;
  input \u4_csr_reg[4]/NET0131  ;
  input \u4_csr_reg[5]/NET0131  ;
  input \u4_csr_reg[6]/NET0131  ;
  input \u4_csr_reg[7]/P0001  ;
  input \u4_csr_reg[8]/P0001  ;
  input \u4_csr_reg[9]/NET0131  ;
  input \u4_dma_in_buf_sz1_reg/P0001  ;
  input \u4_dma_out_buf_avail_reg/P0001  ;
  input \u4_dout_reg[0]/P0001  ;
  input \u4_dout_reg[10]/P0001  ;
  input \u4_dout_reg[11]/P0001  ;
  input \u4_dout_reg[12]/P0001  ;
  input \u4_dout_reg[13]/P0001  ;
  input \u4_dout_reg[14]/P0001  ;
  input \u4_dout_reg[15]/P0001  ;
  input \u4_dout_reg[16]/P0001  ;
  input \u4_dout_reg[17]/P0001  ;
  input \u4_dout_reg[18]/P0001  ;
  input \u4_dout_reg[19]/P0001  ;
  input \u4_dout_reg[1]/P0001  ;
  input \u4_dout_reg[20]/P0001  ;
  input \u4_dout_reg[21]/P0001  ;
  input \u4_dout_reg[22]/P0001  ;
  input \u4_dout_reg[23]/P0001  ;
  input \u4_dout_reg[24]/P0001  ;
  input \u4_dout_reg[25]/P0001  ;
  input \u4_dout_reg[26]/P0001  ;
  input \u4_dout_reg[27]/P0001  ;
  input \u4_dout_reg[28]/P0001  ;
  input \u4_dout_reg[29]/P0001  ;
  input \u4_dout_reg[2]/P0001  ;
  input \u4_dout_reg[30]/P0001  ;
  input \u4_dout_reg[31]/P0001  ;
  input \u4_dout_reg[3]/P0001  ;
  input \u4_dout_reg[4]/P0001  ;
  input \u4_dout_reg[5]/P0001  ;
  input \u4_dout_reg[6]/P0001  ;
  input \u4_dout_reg[7]/P0001  ;
  input \u4_dout_reg[8]/P0001  ;
  input \u4_dout_reg[9]/P0001  ;
  input \u4_funct_adr_reg[0]/P0001  ;
  input \u4_funct_adr_reg[1]/P0001  ;
  input \u4_funct_adr_reg[2]/P0001  ;
  input \u4_funct_adr_reg[3]/P0001  ;
  input \u4_funct_adr_reg[4]/P0001  ;
  input \u4_funct_adr_reg[5]/P0001  ;
  input \u4_funct_adr_reg[6]/P0001  ;
  input \u4_int_src_re_reg/P0001  ;
  input \u4_int_srca_reg[0]/P0001  ;
  input \u4_int_srca_reg[1]/P0001  ;
  input \u4_int_srca_reg[2]/P0001  ;
  input \u4_int_srca_reg[3]/P0001  ;
  input \u4_int_srcb_reg[0]/P0001  ;
  input \u4_int_srcb_reg[1]/P0001  ;
  input \u4_int_srcb_reg[2]/P0001  ;
  input \u4_int_srcb_reg[3]/P0001  ;
  input \u4_int_srcb_reg[4]/P0001  ;
  input \u4_int_srcb_reg[5]/P0001  ;
  input \u4_int_srcb_reg[6]/P0001  ;
  input \u4_int_srcb_reg[7]/P0001  ;
  input \u4_int_srcb_reg[8]/P0001  ;
  input \u4_inta_msk_reg[0]/P0001  ;
  input \u4_inta_msk_reg[1]/P0001  ;
  input \u4_inta_msk_reg[2]/P0001  ;
  input \u4_inta_msk_reg[3]/P0001  ;
  input \u4_inta_msk_reg[4]/P0001  ;
  input \u4_inta_msk_reg[5]/P0001  ;
  input \u4_inta_msk_reg[6]/P0001  ;
  input \u4_inta_msk_reg[7]/P0001  ;
  input \u4_inta_msk_reg[8]/P0001  ;
  input \u4_intb_msk_reg[0]/P0001  ;
  input \u4_intb_msk_reg[1]/P0001  ;
  input \u4_intb_msk_reg[2]/P0001  ;
  input \u4_intb_msk_reg[3]/P0001  ;
  input \u4_intb_msk_reg[4]/P0001  ;
  input \u4_intb_msk_reg[5]/P0001  ;
  input \u4_intb_msk_reg[6]/P0001  ;
  input \u4_intb_msk_reg[7]/P0001  ;
  input \u4_intb_msk_reg[8]/P0001  ;
  input \u4_match_r1_reg/P0001  ;
  input \u4_nse_err_r_reg/P0001  ;
  input \u4_pid_cs_err_r_reg/P0001  ;
  input \u4_rx_err_r_reg/P0001  ;
  input \u4_suspend_r1_reg/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[0]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[10]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[11]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[1]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[2]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[3]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[4]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[5]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[6]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[7]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[8]/P0001  ;
  input \u4_u0_buf0_orig_m3_reg[9]/P0001  ;
  input \u4_u0_buf0_orig_reg[0]/P0001  ;
  input \u4_u0_buf0_orig_reg[10]/P0001  ;
  input \u4_u0_buf0_orig_reg[11]/P0001  ;
  input \u4_u0_buf0_orig_reg[12]/P0001  ;
  input \u4_u0_buf0_orig_reg[13]/P0001  ;
  input \u4_u0_buf0_orig_reg[14]/P0001  ;
  input \u4_u0_buf0_orig_reg[15]/P0001  ;
  input \u4_u0_buf0_orig_reg[16]/P0001  ;
  input \u4_u0_buf0_orig_reg[17]/P0001  ;
  input \u4_u0_buf0_orig_reg[18]/P0001  ;
  input \u4_u0_buf0_orig_reg[19]/P0001  ;
  input \u4_u0_buf0_orig_reg[1]/P0001  ;
  input \u4_u0_buf0_orig_reg[20]/P0001  ;
  input \u4_u0_buf0_orig_reg[21]/P0001  ;
  input \u4_u0_buf0_orig_reg[22]/P0001  ;
  input \u4_u0_buf0_orig_reg[23]/P0001  ;
  input \u4_u0_buf0_orig_reg[24]/P0001  ;
  input \u4_u0_buf0_orig_reg[25]/P0001  ;
  input \u4_u0_buf0_orig_reg[26]/P0001  ;
  input \u4_u0_buf0_orig_reg[27]/P0001  ;
  input \u4_u0_buf0_orig_reg[28]/P0001  ;
  input \u4_u0_buf0_orig_reg[29]/NET0131  ;
  input \u4_u0_buf0_orig_reg[2]/P0001  ;
  input \u4_u0_buf0_orig_reg[30]/NET0131  ;
  input \u4_u0_buf0_orig_reg[31]/P0001  ;
  input \u4_u0_buf0_orig_reg[3]/P0001  ;
  input \u4_u0_buf0_orig_reg[4]/P0001  ;
  input \u4_u0_buf0_orig_reg[5]/P0001  ;
  input \u4_u0_buf0_orig_reg[6]/P0001  ;
  input \u4_u0_buf0_orig_reg[7]/P0001  ;
  input \u4_u0_buf0_orig_reg[8]/P0001  ;
  input \u4_u0_buf0_orig_reg[9]/P0001  ;
  input \u4_u0_buf0_reg[0]/P0001  ;
  input \u4_u0_buf0_reg[10]/P0001  ;
  input \u4_u0_buf0_reg[11]/P0001  ;
  input \u4_u0_buf0_reg[12]/P0001  ;
  input \u4_u0_buf0_reg[13]/P0001  ;
  input \u4_u0_buf0_reg[14]/P0001  ;
  input \u4_u0_buf0_reg[15]/P0001  ;
  input \u4_u0_buf0_reg[16]/P0001  ;
  input \u4_u0_buf0_reg[17]/P0001  ;
  input \u4_u0_buf0_reg[18]/P0001  ;
  input \u4_u0_buf0_reg[19]/P0001  ;
  input \u4_u0_buf0_reg[1]/P0001  ;
  input \u4_u0_buf0_reg[20]/P0001  ;
  input \u4_u0_buf0_reg[21]/P0001  ;
  input \u4_u0_buf0_reg[22]/P0001  ;
  input \u4_u0_buf0_reg[23]/P0001  ;
  input \u4_u0_buf0_reg[24]/P0001  ;
  input \u4_u0_buf0_reg[25]/P0001  ;
  input \u4_u0_buf0_reg[26]/P0001  ;
  input \u4_u0_buf0_reg[27]/P0001  ;
  input \u4_u0_buf0_reg[28]/P0001  ;
  input \u4_u0_buf0_reg[29]/P0001  ;
  input \u4_u0_buf0_reg[2]/P0001  ;
  input \u4_u0_buf0_reg[30]/P0001  ;
  input \u4_u0_buf0_reg[31]/P0001  ;
  input \u4_u0_buf0_reg[3]/P0001  ;
  input \u4_u0_buf0_reg[4]/P0001  ;
  input \u4_u0_buf0_reg[5]/P0001  ;
  input \u4_u0_buf0_reg[6]/P0001  ;
  input \u4_u0_buf0_reg[7]/P0001  ;
  input \u4_u0_buf0_reg[8]/P0001  ;
  input \u4_u0_buf0_reg[9]/P0001  ;
  input \u4_u0_buf1_reg[0]/P0001  ;
  input \u4_u0_buf1_reg[10]/P0001  ;
  input \u4_u0_buf1_reg[11]/P0001  ;
  input \u4_u0_buf1_reg[12]/P0001  ;
  input \u4_u0_buf1_reg[13]/P0001  ;
  input \u4_u0_buf1_reg[14]/P0001  ;
  input \u4_u0_buf1_reg[15]/P0001  ;
  input \u4_u0_buf1_reg[16]/P0001  ;
  input \u4_u0_buf1_reg[17]/P0001  ;
  input \u4_u0_buf1_reg[18]/P0001  ;
  input \u4_u0_buf1_reg[19]/P0001  ;
  input \u4_u0_buf1_reg[1]/P0001  ;
  input \u4_u0_buf1_reg[20]/P0001  ;
  input \u4_u0_buf1_reg[21]/P0001  ;
  input \u4_u0_buf1_reg[22]/P0001  ;
  input \u4_u0_buf1_reg[23]/P0001  ;
  input \u4_u0_buf1_reg[24]/P0001  ;
  input \u4_u0_buf1_reg[25]/P0001  ;
  input \u4_u0_buf1_reg[26]/P0001  ;
  input \u4_u0_buf1_reg[27]/P0001  ;
  input \u4_u0_buf1_reg[28]/P0001  ;
  input \u4_u0_buf1_reg[29]/P0001  ;
  input \u4_u0_buf1_reg[2]/P0001  ;
  input \u4_u0_buf1_reg[30]/P0001  ;
  input \u4_u0_buf1_reg[31]/P0001  ;
  input \u4_u0_buf1_reg[3]/P0001  ;
  input \u4_u0_buf1_reg[4]/P0001  ;
  input \u4_u0_buf1_reg[5]/P0001  ;
  input \u4_u0_buf1_reg[6]/P0001  ;
  input \u4_u0_buf1_reg[7]/P0001  ;
  input \u4_u0_buf1_reg[8]/P0001  ;
  input \u4_u0_buf1_reg[9]/P0001  ;
  input \u4_u0_csr0_reg[0]/P0001  ;
  input \u4_u0_csr0_reg[10]/P0001  ;
  input \u4_u0_csr0_reg[11]/P0001  ;
  input \u4_u0_csr0_reg[12]/P0001  ;
  input \u4_u0_csr0_reg[1]/P0001  ;
  input \u4_u0_csr0_reg[2]/P0001  ;
  input \u4_u0_csr0_reg[3]/NET0131  ;
  input \u4_u0_csr0_reg[4]/P0001  ;
  input \u4_u0_csr0_reg[5]/P0001  ;
  input \u4_u0_csr0_reg[6]/P0001  ;
  input \u4_u0_csr0_reg[7]/P0001  ;
  input \u4_u0_csr0_reg[8]/P0001  ;
  input \u4_u0_csr0_reg[9]/P0001  ;
  input \u4_u0_csr1_reg[0]/P0001  ;
  input \u4_u0_csr1_reg[10]/P0001  ;
  input \u4_u0_csr1_reg[11]/P0001  ;
  input \u4_u0_csr1_reg[12]/P0001  ;
  input \u4_u0_csr1_reg[1]/P0001  ;
  input \u4_u0_csr1_reg[2]/P0001  ;
  input \u4_u0_csr1_reg[3]/P0001  ;
  input \u4_u0_csr1_reg[4]/P0001  ;
  input \u4_u0_csr1_reg[5]/P0001  ;
  input \u4_u0_csr1_reg[6]/P0001  ;
  input \u4_u0_csr1_reg[7]/P0001  ;
  input \u4_u0_csr1_reg[8]/P0001  ;
  input \u4_u0_csr1_reg[9]/P0001  ;
  input \u4_u0_dma_ack_clr1_reg/P0001  ;
  input \u4_u0_dma_ack_wr1_reg/P0001  ;
  input \u4_u0_dma_in_buf_sz1_reg/P0001  ;
  input \u4_u0_dma_in_cnt_reg[0]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[10]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[11]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[1]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[2]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[3]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[4]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[5]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[6]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[7]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[8]/P0001  ;
  input \u4_u0_dma_in_cnt_reg[9]/P0001  ;
  input \u4_u0_dma_out_buf_avail_reg/P0001  ;
  input \u4_u0_dma_out_cnt_reg[10]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[11]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[1]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[2]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[3]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[4]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[5]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[6]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[7]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[8]/P0001  ;
  input \u4_u0_dma_out_cnt_reg[9]/P0001  ;
  input \u4_u0_dma_out_left_reg[0]/P0001  ;
  input \u4_u0_dma_out_left_reg[10]/P0001  ;
  input \u4_u0_dma_out_left_reg[11]/P0001  ;
  input \u4_u0_dma_out_left_reg[1]/P0001  ;
  input \u4_u0_dma_out_left_reg[2]/P0001  ;
  input \u4_u0_dma_out_left_reg[3]/P0001  ;
  input \u4_u0_dma_out_left_reg[4]/P0001  ;
  input \u4_u0_dma_out_left_reg[5]/P0001  ;
  input \u4_u0_dma_out_left_reg[6]/P0001  ;
  input \u4_u0_dma_out_left_reg[7]/P0001  ;
  input \u4_u0_dma_out_left_reg[8]/P0001  ;
  input \u4_u0_dma_out_left_reg[9]/P0001  ;
  input \u4_u0_dma_req_in_hold2_reg/P0001  ;
  input \u4_u0_dma_req_in_hold_reg/P0001  ;
  input \u4_u0_dma_req_out_hold_reg/P0001  ;
  input \u4_u0_ep_match_r_reg/P0001  ;
  input \u4_u0_iena_reg[0]/P0001  ;
  input \u4_u0_iena_reg[1]/P0001  ;
  input \u4_u0_iena_reg[2]/P0001  ;
  input \u4_u0_iena_reg[3]/P0001  ;
  input \u4_u0_iena_reg[4]/P0001  ;
  input \u4_u0_iena_reg[5]/P0001  ;
  input \u4_u0_ienb_reg[0]/P0001  ;
  input \u4_u0_ienb_reg[1]/P0001  ;
  input \u4_u0_ienb_reg[2]/P0001  ;
  input \u4_u0_ienb_reg[3]/P0001  ;
  input \u4_u0_ienb_reg[4]/P0001  ;
  input \u4_u0_ienb_reg[5]/P0001  ;
  input \u4_u0_int_re_reg/P0001  ;
  input \u4_u0_int_stat_reg[0]/P0001  ;
  input \u4_u0_int_stat_reg[1]/P0001  ;
  input \u4_u0_int_stat_reg[2]/P0001  ;
  input \u4_u0_int_stat_reg[3]/P0001  ;
  input \u4_u0_int_stat_reg[4]/P0001  ;
  input \u4_u0_int_stat_reg[5]/P0001  ;
  input \u4_u0_int_stat_reg[6]/P0001  ;
  input \u4_u0_inta_reg/P0001  ;
  input \u4_u0_intb_reg/P0001  ;
  input \u4_u0_ots_stop_reg/P0001  ;
  input \u4_u0_r1_reg/P0001  ;
  input \u4_u0_r2_reg/P0001  ;
  input \u4_u0_r4_reg/P0001  ;
  input \u4_u0_r5_reg/NET0131  ;
  input \u4_u0_set_r_reg/P0001  ;
  input \u4_u0_uc_bsel_reg[0]/P0001  ;
  input \u4_u0_uc_bsel_reg[1]/P0001  ;
  input \u4_u0_uc_dpd_reg[0]/P0001  ;
  input \u4_u0_uc_dpd_reg[1]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[0]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[10]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[11]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[1]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[2]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[3]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[4]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[5]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[6]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[7]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[8]/P0001  ;
  input \u4_u1_buf0_orig_m3_reg[9]/P0001  ;
  input \u4_u1_buf0_orig_reg[0]/P0001  ;
  input \u4_u1_buf0_orig_reg[10]/P0001  ;
  input \u4_u1_buf0_orig_reg[11]/P0001  ;
  input \u4_u1_buf0_orig_reg[12]/P0001  ;
  input \u4_u1_buf0_orig_reg[13]/P0001  ;
  input \u4_u1_buf0_orig_reg[14]/P0001  ;
  input \u4_u1_buf0_orig_reg[15]/P0001  ;
  input \u4_u1_buf0_orig_reg[16]/P0001  ;
  input \u4_u1_buf0_orig_reg[17]/P0001  ;
  input \u4_u1_buf0_orig_reg[18]/P0001  ;
  input \u4_u1_buf0_orig_reg[19]/P0001  ;
  input \u4_u1_buf0_orig_reg[1]/P0001  ;
  input \u4_u1_buf0_orig_reg[20]/P0001  ;
  input \u4_u1_buf0_orig_reg[21]/P0001  ;
  input \u4_u1_buf0_orig_reg[22]/P0001  ;
  input \u4_u1_buf0_orig_reg[23]/P0001  ;
  input \u4_u1_buf0_orig_reg[24]/P0001  ;
  input \u4_u1_buf0_orig_reg[25]/P0001  ;
  input \u4_u1_buf0_orig_reg[26]/P0001  ;
  input \u4_u1_buf0_orig_reg[27]/P0001  ;
  input \u4_u1_buf0_orig_reg[28]/P0001  ;
  input \u4_u1_buf0_orig_reg[29]/NET0131  ;
  input \u4_u1_buf0_orig_reg[2]/P0001  ;
  input \u4_u1_buf0_orig_reg[30]/NET0131  ;
  input \u4_u1_buf0_orig_reg[31]/P0001  ;
  input \u4_u1_buf0_orig_reg[3]/P0001  ;
  input \u4_u1_buf0_orig_reg[4]/P0001  ;
  input \u4_u1_buf0_orig_reg[5]/P0001  ;
  input \u4_u1_buf0_orig_reg[6]/P0001  ;
  input \u4_u1_buf0_orig_reg[7]/P0001  ;
  input \u4_u1_buf0_orig_reg[8]/P0001  ;
  input \u4_u1_buf0_orig_reg[9]/P0001  ;
  input \u4_u1_buf0_reg[0]/P0001  ;
  input \u4_u1_buf0_reg[10]/P0001  ;
  input \u4_u1_buf0_reg[11]/P0001  ;
  input \u4_u1_buf0_reg[12]/P0001  ;
  input \u4_u1_buf0_reg[13]/P0001  ;
  input \u4_u1_buf0_reg[14]/P0001  ;
  input \u4_u1_buf0_reg[15]/P0001  ;
  input \u4_u1_buf0_reg[16]/P0001  ;
  input \u4_u1_buf0_reg[17]/P0001  ;
  input \u4_u1_buf0_reg[18]/P0001  ;
  input \u4_u1_buf0_reg[19]/P0001  ;
  input \u4_u1_buf0_reg[1]/P0001  ;
  input \u4_u1_buf0_reg[20]/P0001  ;
  input \u4_u1_buf0_reg[21]/P0001  ;
  input \u4_u1_buf0_reg[22]/P0001  ;
  input \u4_u1_buf0_reg[23]/P0001  ;
  input \u4_u1_buf0_reg[24]/P0001  ;
  input \u4_u1_buf0_reg[25]/P0001  ;
  input \u4_u1_buf0_reg[26]/P0001  ;
  input \u4_u1_buf0_reg[27]/P0001  ;
  input \u4_u1_buf0_reg[28]/P0001  ;
  input \u4_u1_buf0_reg[29]/P0001  ;
  input \u4_u1_buf0_reg[2]/P0001  ;
  input \u4_u1_buf0_reg[30]/P0001  ;
  input \u4_u1_buf0_reg[31]/P0001  ;
  input \u4_u1_buf0_reg[3]/P0001  ;
  input \u4_u1_buf0_reg[4]/P0001  ;
  input \u4_u1_buf0_reg[5]/P0001  ;
  input \u4_u1_buf0_reg[6]/P0001  ;
  input \u4_u1_buf0_reg[7]/P0001  ;
  input \u4_u1_buf0_reg[8]/P0001  ;
  input \u4_u1_buf0_reg[9]/P0001  ;
  input \u4_u1_buf1_reg[0]/P0001  ;
  input \u4_u1_buf1_reg[10]/P0001  ;
  input \u4_u1_buf1_reg[11]/P0001  ;
  input \u4_u1_buf1_reg[12]/P0001  ;
  input \u4_u1_buf1_reg[13]/P0001  ;
  input \u4_u1_buf1_reg[14]/P0001  ;
  input \u4_u1_buf1_reg[15]/P0001  ;
  input \u4_u1_buf1_reg[16]/P0001  ;
  input \u4_u1_buf1_reg[17]/P0001  ;
  input \u4_u1_buf1_reg[18]/P0001  ;
  input \u4_u1_buf1_reg[19]/P0001  ;
  input \u4_u1_buf1_reg[1]/P0001  ;
  input \u4_u1_buf1_reg[20]/P0001  ;
  input \u4_u1_buf1_reg[21]/P0001  ;
  input \u4_u1_buf1_reg[22]/P0001  ;
  input \u4_u1_buf1_reg[23]/P0001  ;
  input \u4_u1_buf1_reg[24]/P0001  ;
  input \u4_u1_buf1_reg[25]/P0001  ;
  input \u4_u1_buf1_reg[26]/P0001  ;
  input \u4_u1_buf1_reg[27]/P0001  ;
  input \u4_u1_buf1_reg[28]/P0001  ;
  input \u4_u1_buf1_reg[29]/P0001  ;
  input \u4_u1_buf1_reg[2]/P0001  ;
  input \u4_u1_buf1_reg[30]/P0001  ;
  input \u4_u1_buf1_reg[31]/P0001  ;
  input \u4_u1_buf1_reg[3]/P0001  ;
  input \u4_u1_buf1_reg[4]/P0001  ;
  input \u4_u1_buf1_reg[5]/P0001  ;
  input \u4_u1_buf1_reg[6]/P0001  ;
  input \u4_u1_buf1_reg[7]/P0001  ;
  input \u4_u1_buf1_reg[8]/P0001  ;
  input \u4_u1_buf1_reg[9]/P0001  ;
  input \u4_u1_csr0_reg[0]/P0001  ;
  input \u4_u1_csr0_reg[10]/P0001  ;
  input \u4_u1_csr0_reg[11]/P0001  ;
  input \u4_u1_csr0_reg[12]/P0001  ;
  input \u4_u1_csr0_reg[1]/P0001  ;
  input \u4_u1_csr0_reg[2]/P0001  ;
  input \u4_u1_csr0_reg[3]/NET0131  ;
  input \u4_u1_csr0_reg[4]/P0001  ;
  input \u4_u1_csr0_reg[5]/P0001  ;
  input \u4_u1_csr0_reg[6]/P0001  ;
  input \u4_u1_csr0_reg[7]/P0001  ;
  input \u4_u1_csr0_reg[8]/P0001  ;
  input \u4_u1_csr0_reg[9]/P0001  ;
  input \u4_u1_csr1_reg[0]/P0001  ;
  input \u4_u1_csr1_reg[10]/P0001  ;
  input \u4_u1_csr1_reg[11]/P0001  ;
  input \u4_u1_csr1_reg[12]/P0001  ;
  input \u4_u1_csr1_reg[1]/P0001  ;
  input \u4_u1_csr1_reg[2]/P0001  ;
  input \u4_u1_csr1_reg[3]/P0001  ;
  input \u4_u1_csr1_reg[4]/P0001  ;
  input \u4_u1_csr1_reg[5]/P0001  ;
  input \u4_u1_csr1_reg[6]/P0001  ;
  input \u4_u1_csr1_reg[7]/P0001  ;
  input \u4_u1_csr1_reg[8]/P0001  ;
  input \u4_u1_csr1_reg[9]/P0001  ;
  input \u4_u1_dma_ack_clr1_reg/P0001  ;
  input \u4_u1_dma_ack_wr1_reg/P0001  ;
  input \u4_u1_dma_in_buf_sz1_reg/P0001  ;
  input \u4_u1_dma_in_cnt_reg[0]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[10]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[11]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[1]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[2]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[3]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[4]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[5]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[6]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[7]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[8]/P0001  ;
  input \u4_u1_dma_in_cnt_reg[9]/P0001  ;
  input \u4_u1_dma_out_buf_avail_reg/P0001  ;
  input \u4_u1_dma_out_cnt_reg[10]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[11]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[1]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[2]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[3]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[4]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[5]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[6]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[7]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[8]/P0001  ;
  input \u4_u1_dma_out_cnt_reg[9]/P0001  ;
  input \u4_u1_dma_out_left_reg[0]/P0001  ;
  input \u4_u1_dma_out_left_reg[10]/P0001  ;
  input \u4_u1_dma_out_left_reg[11]/P0001  ;
  input \u4_u1_dma_out_left_reg[1]/P0001  ;
  input \u4_u1_dma_out_left_reg[2]/P0001  ;
  input \u4_u1_dma_out_left_reg[3]/P0001  ;
  input \u4_u1_dma_out_left_reg[4]/P0001  ;
  input \u4_u1_dma_out_left_reg[5]/P0001  ;
  input \u4_u1_dma_out_left_reg[6]/P0001  ;
  input \u4_u1_dma_out_left_reg[7]/P0001  ;
  input \u4_u1_dma_out_left_reg[8]/P0001  ;
  input \u4_u1_dma_out_left_reg[9]/P0001  ;
  input \u4_u1_dma_req_in_hold2_reg/P0001  ;
  input \u4_u1_dma_req_in_hold_reg/P0001  ;
  input \u4_u1_dma_req_out_hold_reg/P0001  ;
  input \u4_u1_ep_match_r_reg/P0001  ;
  input \u4_u1_iena_reg[0]/P0001  ;
  input \u4_u1_iena_reg[1]/P0001  ;
  input \u4_u1_iena_reg[2]/P0001  ;
  input \u4_u1_iena_reg[3]/P0001  ;
  input \u4_u1_iena_reg[4]/P0001  ;
  input \u4_u1_iena_reg[5]/P0001  ;
  input \u4_u1_ienb_reg[0]/P0001  ;
  input \u4_u1_ienb_reg[1]/P0001  ;
  input \u4_u1_ienb_reg[2]/P0001  ;
  input \u4_u1_ienb_reg[3]/P0001  ;
  input \u4_u1_ienb_reg[4]/P0001  ;
  input \u4_u1_ienb_reg[5]/P0001  ;
  input \u4_u1_int_re_reg/P0001  ;
  input \u4_u1_int_stat_reg[0]/P0001  ;
  input \u4_u1_int_stat_reg[1]/P0001  ;
  input \u4_u1_int_stat_reg[2]/P0001  ;
  input \u4_u1_int_stat_reg[3]/P0001  ;
  input \u4_u1_int_stat_reg[4]/P0001  ;
  input \u4_u1_int_stat_reg[5]/P0001  ;
  input \u4_u1_int_stat_reg[6]/P0001  ;
  input \u4_u1_inta_reg/P0001  ;
  input \u4_u1_intb_reg/P0001  ;
  input \u4_u1_ots_stop_reg/P0001  ;
  input \u4_u1_r1_reg/P0001  ;
  input \u4_u1_r2_reg/P0001  ;
  input \u4_u1_r4_reg/P0001  ;
  input \u4_u1_r5_reg/NET0131  ;
  input \u4_u1_set_r_reg/P0001  ;
  input \u4_u1_uc_bsel_reg[0]/P0001  ;
  input \u4_u1_uc_bsel_reg[1]/P0001  ;
  input \u4_u1_uc_dpd_reg[0]/P0001  ;
  input \u4_u1_uc_dpd_reg[1]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[0]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[10]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[11]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[1]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[2]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[3]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[4]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[5]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[6]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[7]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[8]/P0001  ;
  input \u4_u2_buf0_orig_m3_reg[9]/P0001  ;
  input \u4_u2_buf0_orig_reg[0]/P0001  ;
  input \u4_u2_buf0_orig_reg[10]/P0001  ;
  input \u4_u2_buf0_orig_reg[11]/P0001  ;
  input \u4_u2_buf0_orig_reg[12]/P0001  ;
  input \u4_u2_buf0_orig_reg[13]/P0001  ;
  input \u4_u2_buf0_orig_reg[14]/P0001  ;
  input \u4_u2_buf0_orig_reg[15]/P0001  ;
  input \u4_u2_buf0_orig_reg[16]/P0001  ;
  input \u4_u2_buf0_orig_reg[17]/P0001  ;
  input \u4_u2_buf0_orig_reg[18]/P0001  ;
  input \u4_u2_buf0_orig_reg[19]/P0001  ;
  input \u4_u2_buf0_orig_reg[1]/P0001  ;
  input \u4_u2_buf0_orig_reg[20]/P0001  ;
  input \u4_u2_buf0_orig_reg[21]/P0001  ;
  input \u4_u2_buf0_orig_reg[22]/P0001  ;
  input \u4_u2_buf0_orig_reg[23]/P0001  ;
  input \u4_u2_buf0_orig_reg[24]/P0001  ;
  input \u4_u2_buf0_orig_reg[25]/P0001  ;
  input \u4_u2_buf0_orig_reg[26]/P0001  ;
  input \u4_u2_buf0_orig_reg[27]/P0001  ;
  input \u4_u2_buf0_orig_reg[28]/P0001  ;
  input \u4_u2_buf0_orig_reg[29]/NET0131  ;
  input \u4_u2_buf0_orig_reg[2]/P0001  ;
  input \u4_u2_buf0_orig_reg[30]/NET0131  ;
  input \u4_u2_buf0_orig_reg[31]/P0001  ;
  input \u4_u2_buf0_orig_reg[3]/P0001  ;
  input \u4_u2_buf0_orig_reg[4]/P0001  ;
  input \u4_u2_buf0_orig_reg[5]/P0001  ;
  input \u4_u2_buf0_orig_reg[6]/P0001  ;
  input \u4_u2_buf0_orig_reg[7]/P0001  ;
  input \u4_u2_buf0_orig_reg[8]/P0001  ;
  input \u4_u2_buf0_orig_reg[9]/P0001  ;
  input \u4_u2_buf0_reg[0]/P0001  ;
  input \u4_u2_buf0_reg[10]/P0001  ;
  input \u4_u2_buf0_reg[11]/P0001  ;
  input \u4_u2_buf0_reg[12]/P0001  ;
  input \u4_u2_buf0_reg[13]/P0001  ;
  input \u4_u2_buf0_reg[14]/P0001  ;
  input \u4_u2_buf0_reg[15]/P0001  ;
  input \u4_u2_buf0_reg[16]/P0001  ;
  input \u4_u2_buf0_reg[17]/P0001  ;
  input \u4_u2_buf0_reg[18]/P0001  ;
  input \u4_u2_buf0_reg[19]/P0001  ;
  input \u4_u2_buf0_reg[1]/P0001  ;
  input \u4_u2_buf0_reg[20]/P0001  ;
  input \u4_u2_buf0_reg[21]/P0001  ;
  input \u4_u2_buf0_reg[22]/P0001  ;
  input \u4_u2_buf0_reg[23]/P0001  ;
  input \u4_u2_buf0_reg[24]/P0001  ;
  input \u4_u2_buf0_reg[25]/P0001  ;
  input \u4_u2_buf0_reg[26]/P0001  ;
  input \u4_u2_buf0_reg[27]/P0001  ;
  input \u4_u2_buf0_reg[28]/P0001  ;
  input \u4_u2_buf0_reg[29]/P0001  ;
  input \u4_u2_buf0_reg[2]/P0001  ;
  input \u4_u2_buf0_reg[30]/P0001  ;
  input \u4_u2_buf0_reg[31]/P0001  ;
  input \u4_u2_buf0_reg[3]/P0001  ;
  input \u4_u2_buf0_reg[4]/P0001  ;
  input \u4_u2_buf0_reg[5]/P0001  ;
  input \u4_u2_buf0_reg[6]/P0001  ;
  input \u4_u2_buf0_reg[7]/P0001  ;
  input \u4_u2_buf0_reg[8]/P0001  ;
  input \u4_u2_buf0_reg[9]/P0001  ;
  input \u4_u2_buf1_reg[0]/P0001  ;
  input \u4_u2_buf1_reg[10]/P0001  ;
  input \u4_u2_buf1_reg[11]/P0001  ;
  input \u4_u2_buf1_reg[12]/P0001  ;
  input \u4_u2_buf1_reg[13]/P0001  ;
  input \u4_u2_buf1_reg[14]/P0001  ;
  input \u4_u2_buf1_reg[15]/P0001  ;
  input \u4_u2_buf1_reg[16]/P0001  ;
  input \u4_u2_buf1_reg[17]/P0001  ;
  input \u4_u2_buf1_reg[18]/P0001  ;
  input \u4_u2_buf1_reg[19]/P0001  ;
  input \u4_u2_buf1_reg[1]/P0001  ;
  input \u4_u2_buf1_reg[20]/P0001  ;
  input \u4_u2_buf1_reg[21]/P0001  ;
  input \u4_u2_buf1_reg[22]/P0001  ;
  input \u4_u2_buf1_reg[23]/P0001  ;
  input \u4_u2_buf1_reg[24]/P0001  ;
  input \u4_u2_buf1_reg[25]/P0001  ;
  input \u4_u2_buf1_reg[26]/P0001  ;
  input \u4_u2_buf1_reg[27]/P0001  ;
  input \u4_u2_buf1_reg[28]/P0001  ;
  input \u4_u2_buf1_reg[29]/P0001  ;
  input \u4_u2_buf1_reg[2]/P0001  ;
  input \u4_u2_buf1_reg[30]/P0001  ;
  input \u4_u2_buf1_reg[31]/P0001  ;
  input \u4_u2_buf1_reg[3]/P0001  ;
  input \u4_u2_buf1_reg[4]/P0001  ;
  input \u4_u2_buf1_reg[5]/P0001  ;
  input \u4_u2_buf1_reg[6]/P0001  ;
  input \u4_u2_buf1_reg[7]/P0001  ;
  input \u4_u2_buf1_reg[8]/P0001  ;
  input \u4_u2_buf1_reg[9]/P0001  ;
  input \u4_u2_csr0_reg[0]/P0001  ;
  input \u4_u2_csr0_reg[10]/P0001  ;
  input \u4_u2_csr0_reg[11]/P0001  ;
  input \u4_u2_csr0_reg[12]/P0001  ;
  input \u4_u2_csr0_reg[1]/P0001  ;
  input \u4_u2_csr0_reg[2]/P0001  ;
  input \u4_u2_csr0_reg[3]/NET0131  ;
  input \u4_u2_csr0_reg[4]/P0001  ;
  input \u4_u2_csr0_reg[5]/P0001  ;
  input \u4_u2_csr0_reg[6]/P0001  ;
  input \u4_u2_csr0_reg[7]/P0001  ;
  input \u4_u2_csr0_reg[8]/P0001  ;
  input \u4_u2_csr0_reg[9]/P0001  ;
  input \u4_u2_csr1_reg[0]/P0001  ;
  input \u4_u2_csr1_reg[10]/P0001  ;
  input \u4_u2_csr1_reg[11]/P0001  ;
  input \u4_u2_csr1_reg[12]/P0001  ;
  input \u4_u2_csr1_reg[1]/P0001  ;
  input \u4_u2_csr1_reg[2]/P0001  ;
  input \u4_u2_csr1_reg[3]/P0001  ;
  input \u4_u2_csr1_reg[4]/P0001  ;
  input \u4_u2_csr1_reg[5]/P0001  ;
  input \u4_u2_csr1_reg[6]/P0001  ;
  input \u4_u2_csr1_reg[7]/P0001  ;
  input \u4_u2_csr1_reg[8]/P0001  ;
  input \u4_u2_csr1_reg[9]/P0001  ;
  input \u4_u2_dma_ack_clr1_reg/P0001  ;
  input \u4_u2_dma_ack_wr1_reg/P0001  ;
  input \u4_u2_dma_in_buf_sz1_reg/P0001  ;
  input \u4_u2_dma_in_cnt_reg[0]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[10]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[11]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[1]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[2]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[3]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[4]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[5]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[6]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[7]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[8]/P0001  ;
  input \u4_u2_dma_in_cnt_reg[9]/P0001  ;
  input \u4_u2_dma_out_buf_avail_reg/P0001  ;
  input \u4_u2_dma_out_cnt_reg[10]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[11]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[1]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[2]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[3]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[4]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[5]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[6]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[7]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[8]/P0001  ;
  input \u4_u2_dma_out_cnt_reg[9]/P0001  ;
  input \u4_u2_dma_out_left_reg[0]/P0001  ;
  input \u4_u2_dma_out_left_reg[10]/P0001  ;
  input \u4_u2_dma_out_left_reg[11]/P0001  ;
  input \u4_u2_dma_out_left_reg[1]/P0001  ;
  input \u4_u2_dma_out_left_reg[2]/P0001  ;
  input \u4_u2_dma_out_left_reg[3]/P0001  ;
  input \u4_u2_dma_out_left_reg[4]/P0001  ;
  input \u4_u2_dma_out_left_reg[5]/P0001  ;
  input \u4_u2_dma_out_left_reg[6]/P0001  ;
  input \u4_u2_dma_out_left_reg[7]/P0001  ;
  input \u4_u2_dma_out_left_reg[8]/P0001  ;
  input \u4_u2_dma_out_left_reg[9]/P0001  ;
  input \u4_u2_dma_req_in_hold2_reg/P0001  ;
  input \u4_u2_dma_req_in_hold_reg/P0001  ;
  input \u4_u2_dma_req_out_hold_reg/P0001  ;
  input \u4_u2_ep_match_r_reg/P0001  ;
  input \u4_u2_iena_reg[0]/P0001  ;
  input \u4_u2_iena_reg[1]/P0001  ;
  input \u4_u2_iena_reg[2]/P0001  ;
  input \u4_u2_iena_reg[3]/P0001  ;
  input \u4_u2_iena_reg[4]/P0001  ;
  input \u4_u2_iena_reg[5]/P0001  ;
  input \u4_u2_ienb_reg[0]/P0001  ;
  input \u4_u2_ienb_reg[1]/P0001  ;
  input \u4_u2_ienb_reg[2]/P0001  ;
  input \u4_u2_ienb_reg[3]/P0001  ;
  input \u4_u2_ienb_reg[4]/P0001  ;
  input \u4_u2_ienb_reg[5]/P0001  ;
  input \u4_u2_int_re_reg/P0001  ;
  input \u4_u2_int_stat_reg[0]/P0001  ;
  input \u4_u2_int_stat_reg[1]/P0001  ;
  input \u4_u2_int_stat_reg[2]/P0001  ;
  input \u4_u2_int_stat_reg[3]/P0001  ;
  input \u4_u2_int_stat_reg[4]/P0001  ;
  input \u4_u2_int_stat_reg[5]/P0001  ;
  input \u4_u2_int_stat_reg[6]/P0001  ;
  input \u4_u2_inta_reg/P0001  ;
  input \u4_u2_intb_reg/P0001  ;
  input \u4_u2_ots_stop_reg/P0001  ;
  input \u4_u2_r1_reg/P0001  ;
  input \u4_u2_r2_reg/P0001  ;
  input \u4_u2_r4_reg/P0001  ;
  input \u4_u2_r5_reg/NET0131  ;
  input \u4_u2_set_r_reg/P0001  ;
  input \u4_u2_uc_bsel_reg[0]/P0001  ;
  input \u4_u2_uc_bsel_reg[1]/P0001  ;
  input \u4_u2_uc_dpd_reg[0]/P0001  ;
  input \u4_u2_uc_dpd_reg[1]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[0]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[10]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[11]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[1]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[2]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[3]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[4]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[5]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[6]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[7]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[8]/P0001  ;
  input \u4_u3_buf0_orig_m3_reg[9]/P0001  ;
  input \u4_u3_buf0_orig_reg[0]/P0001  ;
  input \u4_u3_buf0_orig_reg[10]/P0001  ;
  input \u4_u3_buf0_orig_reg[11]/P0001  ;
  input \u4_u3_buf0_orig_reg[12]/P0001  ;
  input \u4_u3_buf0_orig_reg[13]/P0001  ;
  input \u4_u3_buf0_orig_reg[14]/P0001  ;
  input \u4_u3_buf0_orig_reg[15]/P0001  ;
  input \u4_u3_buf0_orig_reg[16]/P0001  ;
  input \u4_u3_buf0_orig_reg[17]/P0001  ;
  input \u4_u3_buf0_orig_reg[18]/P0001  ;
  input \u4_u3_buf0_orig_reg[19]/P0001  ;
  input \u4_u3_buf0_orig_reg[1]/P0001  ;
  input \u4_u3_buf0_orig_reg[20]/P0001  ;
  input \u4_u3_buf0_orig_reg[21]/P0001  ;
  input \u4_u3_buf0_orig_reg[22]/P0001  ;
  input \u4_u3_buf0_orig_reg[23]/P0001  ;
  input \u4_u3_buf0_orig_reg[24]/P0001  ;
  input \u4_u3_buf0_orig_reg[25]/P0001  ;
  input \u4_u3_buf0_orig_reg[26]/P0001  ;
  input \u4_u3_buf0_orig_reg[27]/P0001  ;
  input \u4_u3_buf0_orig_reg[28]/P0001  ;
  input \u4_u3_buf0_orig_reg[29]/NET0131  ;
  input \u4_u3_buf0_orig_reg[2]/P0001  ;
  input \u4_u3_buf0_orig_reg[30]/NET0131  ;
  input \u4_u3_buf0_orig_reg[31]/P0001  ;
  input \u4_u3_buf0_orig_reg[3]/P0001  ;
  input \u4_u3_buf0_orig_reg[4]/P0001  ;
  input \u4_u3_buf0_orig_reg[5]/P0001  ;
  input \u4_u3_buf0_orig_reg[6]/P0001  ;
  input \u4_u3_buf0_orig_reg[7]/P0001  ;
  input \u4_u3_buf0_orig_reg[8]/P0001  ;
  input \u4_u3_buf0_orig_reg[9]/P0001  ;
  input \u4_u3_buf0_reg[0]/P0001  ;
  input \u4_u3_buf0_reg[10]/P0001  ;
  input \u4_u3_buf0_reg[11]/P0001  ;
  input \u4_u3_buf0_reg[12]/P0001  ;
  input \u4_u3_buf0_reg[13]/P0001  ;
  input \u4_u3_buf0_reg[14]/P0001  ;
  input \u4_u3_buf0_reg[15]/P0001  ;
  input \u4_u3_buf0_reg[16]/P0001  ;
  input \u4_u3_buf0_reg[17]/P0001  ;
  input \u4_u3_buf0_reg[18]/P0001  ;
  input \u4_u3_buf0_reg[19]/P0001  ;
  input \u4_u3_buf0_reg[1]/P0001  ;
  input \u4_u3_buf0_reg[20]/P0001  ;
  input \u4_u3_buf0_reg[21]/P0001  ;
  input \u4_u3_buf0_reg[22]/P0001  ;
  input \u4_u3_buf0_reg[23]/P0001  ;
  input \u4_u3_buf0_reg[24]/P0001  ;
  input \u4_u3_buf0_reg[25]/P0001  ;
  input \u4_u3_buf0_reg[26]/P0001  ;
  input \u4_u3_buf0_reg[27]/P0001  ;
  input \u4_u3_buf0_reg[28]/P0001  ;
  input \u4_u3_buf0_reg[29]/P0001  ;
  input \u4_u3_buf0_reg[2]/P0001  ;
  input \u4_u3_buf0_reg[30]/P0001  ;
  input \u4_u3_buf0_reg[31]/P0001  ;
  input \u4_u3_buf0_reg[3]/P0001  ;
  input \u4_u3_buf0_reg[4]/P0001  ;
  input \u4_u3_buf0_reg[5]/P0001  ;
  input \u4_u3_buf0_reg[6]/P0001  ;
  input \u4_u3_buf0_reg[7]/P0001  ;
  input \u4_u3_buf0_reg[8]/P0001  ;
  input \u4_u3_buf0_reg[9]/P0001  ;
  input \u4_u3_buf1_reg[0]/P0001  ;
  input \u4_u3_buf1_reg[10]/P0001  ;
  input \u4_u3_buf1_reg[11]/P0001  ;
  input \u4_u3_buf1_reg[12]/P0001  ;
  input \u4_u3_buf1_reg[13]/P0001  ;
  input \u4_u3_buf1_reg[14]/P0001  ;
  input \u4_u3_buf1_reg[15]/P0001  ;
  input \u4_u3_buf1_reg[16]/P0001  ;
  input \u4_u3_buf1_reg[17]/P0001  ;
  input \u4_u3_buf1_reg[18]/P0001  ;
  input \u4_u3_buf1_reg[19]/P0001  ;
  input \u4_u3_buf1_reg[1]/P0001  ;
  input \u4_u3_buf1_reg[20]/P0001  ;
  input \u4_u3_buf1_reg[21]/P0001  ;
  input \u4_u3_buf1_reg[22]/P0001  ;
  input \u4_u3_buf1_reg[23]/P0001  ;
  input \u4_u3_buf1_reg[24]/P0001  ;
  input \u4_u3_buf1_reg[25]/P0001  ;
  input \u4_u3_buf1_reg[26]/P0001  ;
  input \u4_u3_buf1_reg[27]/P0001  ;
  input \u4_u3_buf1_reg[28]/P0001  ;
  input \u4_u3_buf1_reg[29]/P0001  ;
  input \u4_u3_buf1_reg[2]/P0001  ;
  input \u4_u3_buf1_reg[30]/P0001  ;
  input \u4_u3_buf1_reg[31]/P0001  ;
  input \u4_u3_buf1_reg[3]/P0001  ;
  input \u4_u3_buf1_reg[4]/P0001  ;
  input \u4_u3_buf1_reg[5]/P0001  ;
  input \u4_u3_buf1_reg[6]/P0001  ;
  input \u4_u3_buf1_reg[7]/P0001  ;
  input \u4_u3_buf1_reg[8]/P0001  ;
  input \u4_u3_buf1_reg[9]/P0001  ;
  input \u4_u3_csr0_reg[0]/P0001  ;
  input \u4_u3_csr0_reg[10]/P0001  ;
  input \u4_u3_csr0_reg[11]/P0001  ;
  input \u4_u3_csr0_reg[12]/P0001  ;
  input \u4_u3_csr0_reg[1]/P0001  ;
  input \u4_u3_csr0_reg[2]/P0001  ;
  input \u4_u3_csr0_reg[3]/NET0131  ;
  input \u4_u3_csr0_reg[4]/P0001  ;
  input \u4_u3_csr0_reg[5]/P0001  ;
  input \u4_u3_csr0_reg[6]/P0001  ;
  input \u4_u3_csr0_reg[7]/P0001  ;
  input \u4_u3_csr0_reg[8]/P0001  ;
  input \u4_u3_csr0_reg[9]/P0001  ;
  input \u4_u3_csr1_reg[0]/P0001  ;
  input \u4_u3_csr1_reg[10]/P0001  ;
  input \u4_u3_csr1_reg[11]/P0001  ;
  input \u4_u3_csr1_reg[12]/P0001  ;
  input \u4_u3_csr1_reg[1]/P0001  ;
  input \u4_u3_csr1_reg[2]/P0001  ;
  input \u4_u3_csr1_reg[3]/P0001  ;
  input \u4_u3_csr1_reg[4]/P0001  ;
  input \u4_u3_csr1_reg[5]/P0001  ;
  input \u4_u3_csr1_reg[6]/P0001  ;
  input \u4_u3_csr1_reg[7]/P0001  ;
  input \u4_u3_csr1_reg[8]/P0001  ;
  input \u4_u3_csr1_reg[9]/P0001  ;
  input \u4_u3_dma_ack_clr1_reg/P0001  ;
  input \u4_u3_dma_ack_wr1_reg/P0001  ;
  input \u4_u3_dma_in_buf_sz1_reg/P0001  ;
  input \u4_u3_dma_in_cnt_reg[0]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[10]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[11]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[1]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[2]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[3]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[4]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[5]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[6]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[7]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[8]/P0001  ;
  input \u4_u3_dma_in_cnt_reg[9]/P0001  ;
  input \u4_u3_dma_out_buf_avail_reg/P0001  ;
  input \u4_u3_dma_out_cnt_reg[10]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[11]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[1]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[2]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[3]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[4]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[5]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[6]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[7]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[8]/P0001  ;
  input \u4_u3_dma_out_cnt_reg[9]/P0001  ;
  input \u4_u3_dma_out_left_reg[0]/P0001  ;
  input \u4_u3_dma_out_left_reg[10]/P0001  ;
  input \u4_u3_dma_out_left_reg[11]/P0001  ;
  input \u4_u3_dma_out_left_reg[1]/P0001  ;
  input \u4_u3_dma_out_left_reg[2]/P0001  ;
  input \u4_u3_dma_out_left_reg[3]/P0001  ;
  input \u4_u3_dma_out_left_reg[4]/P0001  ;
  input \u4_u3_dma_out_left_reg[5]/P0001  ;
  input \u4_u3_dma_out_left_reg[6]/P0001  ;
  input \u4_u3_dma_out_left_reg[7]/P0001  ;
  input \u4_u3_dma_out_left_reg[8]/P0001  ;
  input \u4_u3_dma_out_left_reg[9]/P0001  ;
  input \u4_u3_dma_req_in_hold2_reg/P0001  ;
  input \u4_u3_dma_req_in_hold_reg/P0001  ;
  input \u4_u3_dma_req_out_hold_reg/P0001  ;
  input \u4_u3_ep_match_r_reg/P0001  ;
  input \u4_u3_iena_reg[0]/P0001  ;
  input \u4_u3_iena_reg[1]/P0001  ;
  input \u4_u3_iena_reg[2]/P0001  ;
  input \u4_u3_iena_reg[3]/P0001  ;
  input \u4_u3_iena_reg[4]/P0001  ;
  input \u4_u3_iena_reg[5]/P0001  ;
  input \u4_u3_ienb_reg[0]/P0001  ;
  input \u4_u3_ienb_reg[1]/P0001  ;
  input \u4_u3_ienb_reg[2]/P0001  ;
  input \u4_u3_ienb_reg[3]/P0001  ;
  input \u4_u3_ienb_reg[4]/P0001  ;
  input \u4_u3_ienb_reg[5]/P0001  ;
  input \u4_u3_int_re_reg/P0001  ;
  input \u4_u3_int_stat_reg[0]/P0001  ;
  input \u4_u3_int_stat_reg[1]/P0001  ;
  input \u4_u3_int_stat_reg[2]/P0001  ;
  input \u4_u3_int_stat_reg[3]/P0001  ;
  input \u4_u3_int_stat_reg[4]/P0001  ;
  input \u4_u3_int_stat_reg[5]/P0001  ;
  input \u4_u3_int_stat_reg[6]/P0001  ;
  input \u4_u3_inta_reg/P0001  ;
  input \u4_u3_intb_reg/P0001  ;
  input \u4_u3_ots_stop_reg/P0001  ;
  input \u4_u3_r1_reg/P0001  ;
  input \u4_u3_r2_reg/P0001  ;
  input \u4_u3_r4_reg/P0001  ;
  input \u4_u3_r5_reg/NET0131  ;
  input \u4_u3_set_r_reg/P0001  ;
  input \u4_u3_uc_bsel_reg[0]/P0001  ;
  input \u4_u3_uc_bsel_reg[1]/P0001  ;
  input \u4_u3_uc_dpd_reg[0]/P0001  ;
  input \u4_u3_uc_dpd_reg[1]/P0001  ;
  input \u4_usb_reset_r_reg/P0001  ;
  input \u4_utmi_vend_ctrl_r_reg[0]/P0001  ;
  input \u4_utmi_vend_ctrl_r_reg[1]/P0001  ;
  input \u4_utmi_vend_ctrl_r_reg[2]/P0001  ;
  input \u4_utmi_vend_ctrl_r_reg[3]/P0001  ;
  input \u4_utmi_vend_stat_r_reg[0]/P0001  ;
  input \u4_utmi_vend_stat_r_reg[1]/P0001  ;
  input \u4_utmi_vend_stat_r_reg[2]/P0001  ;
  input \u4_utmi_vend_stat_r_reg[3]/P0001  ;
  input \u4_utmi_vend_stat_r_reg[4]/P0001  ;
  input \u4_utmi_vend_stat_r_reg[5]/P0001  ;
  input \u4_utmi_vend_stat_r_reg[6]/P0001  ;
  input \u4_utmi_vend_stat_r_reg[7]/P0001  ;
  input \u4_utmi_vend_wr_r_reg/P0001  ;
  input \u5_state_reg[0]/P0001  ;
  input \u5_state_reg[1]/P0001  ;
  input \u5_state_reg[2]/P0001  ;
  input \u5_state_reg[3]/P0001  ;
  input \u5_state_reg[4]/P0001  ;
  input \u5_state_reg[5]/NET0131  ;
  input \u5_wb_ack_s1_reg/P0001  ;
  input \u5_wb_ack_s2_reg/P0001  ;
  input \u5_wb_req_s1_reg/P0001  ;
  input usb_vbus_pad_i_pad ;
  input wb_ack_o_pad ;
  input \wb_addr_i[10]_pad  ;
  input \wb_addr_i[11]_pad  ;
  input \wb_addr_i[12]_pad  ;
  input \wb_addr_i[13]_pad  ;
  input \wb_addr_i[14]_pad  ;
  input \wb_addr_i[15]_pad  ;
  input \wb_addr_i[16]_pad  ;
  input \wb_addr_i[17]_pad  ;
  input \wb_addr_i[2]_pad  ;
  input \wb_addr_i[3]_pad  ;
  input \wb_addr_i[4]_pad  ;
  input \wb_addr_i[5]_pad  ;
  input \wb_addr_i[6]_pad  ;
  input \wb_addr_i[7]_pad  ;
  input \wb_addr_i[8]_pad  ;
  input \wb_addr_i[9]_pad  ;
  input wb_cyc_i_pad ;
  input \wb_data_i[0]_pad  ;
  input \wb_data_i[10]_pad  ;
  input \wb_data_i[11]_pad  ;
  input \wb_data_i[12]_pad  ;
  input \wb_data_i[13]_pad  ;
  input \wb_data_i[14]_pad  ;
  input \wb_data_i[15]_pad  ;
  input \wb_data_i[16]_pad  ;
  input \wb_data_i[17]_pad  ;
  input \wb_data_i[18]_pad  ;
  input \wb_data_i[19]_pad  ;
  input \wb_data_i[1]_pad  ;
  input \wb_data_i[20]_pad  ;
  input \wb_data_i[21]_pad  ;
  input \wb_data_i[22]_pad  ;
  input \wb_data_i[23]_pad  ;
  input \wb_data_i[24]_pad  ;
  input \wb_data_i[25]_pad  ;
  input \wb_data_i[26]_pad  ;
  input \wb_data_i[27]_pad  ;
  input \wb_data_i[28]_pad  ;
  input \wb_data_i[29]_pad  ;
  input \wb_data_i[2]_pad  ;
  input \wb_data_i[30]_pad  ;
  input \wb_data_i[31]_pad  ;
  input \wb_data_i[3]_pad  ;
  input \wb_data_i[4]_pad  ;
  input \wb_data_i[5]_pad  ;
  input \wb_data_i[6]_pad  ;
  input \wb_data_i[7]_pad  ;
  input \wb_data_i[8]_pad  ;
  input \wb_data_i[9]_pad  ;
  input wb_stb_i_pad ;
  input wb_we_i_pad ;
  output \dma_req_o[6]_pad  ;
  output \g37425/_0_  ;
  output \g37426/_0_  ;
  output \g37432/_0_  ;
  output \g37433/_0_  ;
  output \g37439/_0_  ;
  output \g37440/_0_  ;
  output \g37444/_00_  ;
  output \g37448/_0_  ;
  output \g37450/_0_  ;
  output \g37454/_0_  ;
  output \g37473/_0_  ;
  output \g37474/_0_  ;
  output \g37475/_0_  ;
  output \g37476/_0_  ;
  output \g37477/_0_  ;
  output \g37478/_0_  ;
  output \g37479/_0_  ;
  output \g37488/_0_  ;
  output \g37489/_0_  ;
  output \g37490/_0_  ;
  output \g37491/_0_  ;
  output \g37492/_0_  ;
  output \g37517/_0_  ;
  output \g37518/_0_  ;
  output \g37519/_0_  ;
  output \g37520/_0_  ;
  output \g37521/_0_  ;
  output \g37522/_0_  ;
  output \g37540/_0_  ;
  output \g37542/_0_  ;
  output \g37543/_0_  ;
  output \g37545/_0_  ;
  output \g37546/_0_  ;
  output \g37548/_0_  ;
  output \g37549/_0_  ;
  output \g37550/_0_  ;
  output \g37551/_0_  ;
  output \g37556/_0_  ;
  output \g37589/_0_  ;
  output \g37591/_0_  ;
  output \g37592/_0_  ;
  output \g37593/_0_  ;
  output \g37594/_0_  ;
  output \g37596/_0_  ;
  output \g37597/_0_  ;
  output \g37598/_0_  ;
  output \g37599/_0_  ;
  output \g37601/_0_  ;
  output \g37603/_0_  ;
  output \g37604/_0_  ;
  output \g37605/_0_  ;
  output \g37607/_0_  ;
  output \g37608/_0_  ;
  output \g37609/_0_  ;
  output \g37610/_0_  ;
  output \g37645/_0_  ;
  output \g37648/_0_  ;
  output \g37650/_0_  ;
  output \g37653/_0_  ;
  output \g37664/_3_  ;
  output \g37703/_0_  ;
  output \g37704/_0_  ;
  output \g37706/_0_  ;
  output \g37708/_0_  ;
  output \g37709/_0_  ;
  output \g37711/_0_  ;
  output \g37714/_0_  ;
  output \g37715/_0_  ;
  output \g37717/_0_  ;
  output \g37718/_0_  ;
  output \g37719/_0_  ;
  output \g37720/_0_  ;
  output \g37723/_0_  ;
  output \g37724/_0_  ;
  output \g37726/_0_  ;
  output \g37728/_0_  ;
  output \g37729/_0_  ;
  output \g37730/_0_  ;
  output \g37731/_0_  ;
  output \g37732/_0_  ;
  output \g37733/_0_  ;
  output \g37735/_0_  ;
  output \g37736/_0_  ;
  output \g37737/_0_  ;
  output \g37856/_0_  ;
  output \g37857/_0_  ;
  output \g37859/_0_  ;
  output \g37868/_0_  ;
  output \g37869/_0_  ;
  output \g37870/_0_  ;
  output \g37872/_0_  ;
  output \g37886/_0_  ;
  output \g37887/_0_  ;
  output \g37889/_0_  ;
  output \g37897/_0_  ;
  output \g37899/_0_  ;
  output \g37900/_0_  ;
  output \g37907/_0_  ;
  output \g37925/_0_  ;
  output \g37927/_0_  ;
  output \g37928/_0_  ;
  output \g37929/_0_  ;
  output \g37930/_0_  ;
  output \g37932/_0_  ;
  output \g37933/_0_  ;
  output \g37934/_0_  ;
  output \g37935/_0_  ;
  output \g37936/_0_  ;
  output \g37937/_0_  ;
  output \g37938/_0_  ;
  output \g37939/_0_  ;
  output \g37941/_0_  ;
  output \g37942/_0_  ;
  output \g37943/_0_  ;
  output \g37944/_0_  ;
  output \g37945/_0_  ;
  output \g38030/_3_  ;
  output \g38035/_0_  ;
  output \g38036/_0_  ;
  output \g38054/_0_  ;
  output \g38129/_0_  ;
  output \g38130/_0_  ;
  output \g38148/_3_  ;
  output \g38149/_3_  ;
  output \g38150/_3_  ;
  output \g38166/_0_  ;
  output \g38198/_0_  ;
  output \g38201/_0_  ;
  output \g38257/_0_  ;
  output \g38286/_0_  ;
  output \g38294/_3_  ;
  output \g38295/_3_  ;
  output \g38296/_3_  ;
  output \g38297/_3_  ;
  output \g38332/_0_  ;
  output \g38350/_0_  ;
  output \g38365/_3_  ;
  output \g38366/_3_  ;
  output \g38367/_3_  ;
  output \g38389/_0_  ;
  output \g38397/_0_  ;
  output \g38398/_0_  ;
  output \g38399/_0_  ;
  output \g38400/_0_  ;
  output \g38417/_3_  ;
  output \g38418/_3_  ;
  output \g38422/_0_  ;
  output \g38440/_0_  ;
  output \g38443/_0_  ;
  output \g38448/_3_  ;
  output \g38449/_0_  ;
  output \g38450/_0_  ;
  output \g38460/_0_  ;
  output \g38466/_0_  ;
  output \g38467/_0_  ;
  output \g38468/_0_  ;
  output \g38469/_0_  ;
  output \g38470/_0_  ;
  output \g38471/_0_  ;
  output \g38472/_0_  ;
  output \g38473/_0_  ;
  output \g38474/_0_  ;
  output \g38475/_0_  ;
  output \g38476/_0_  ;
  output \g38477/_0_  ;
  output \g38478/_0_  ;
  output \g38479/_0_  ;
  output \g38528/_0_  ;
  output \g38533/_0_  ;
  output \g38534/_0_  ;
  output \g38536/_0_  ;
  output \g38545/_0_  ;
  output \g38551/_0_  ;
  output \g38554/_0_  ;
  output \g38555/_0_  ;
  output \g38556/_0_  ;
  output \g38575/_0_  ;
  output \g38616/_0_  ;
  output \g38653/_0_  ;
  output \g38656/_0_  ;
  output \g38657/_0_  ;
  output \g38658/_0_  ;
  output \g38660/_0_  ;
  output \g38706/_0_  ;
  output \g38716/_0_  ;
  output \g38717/_0_  ;
  output \g38738/_1_  ;
  output \g38763/_0_  ;
  output \g38790/_0_  ;
  output \g38792/_0_  ;
  output \g38801/_0_  ;
  output \g38803/_0_  ;
  output \g38804/_0_  ;
  output \g38805/_0_  ;
  output \g38806/_0_  ;
  output \g38807/_0_  ;
  output \g38808/_0_  ;
  output \g38809/_0_  ;
  output \g38810/_0_  ;
  output \g38814/_0_  ;
  output \g38833/_0_  ;
  output \g38834/_0_  ;
  output \g38839/_0_  ;
  output \g38840/_0_  ;
  output \g38841/_0_  ;
  output \g38842/_0_  ;
  output \g38846/_0_  ;
  output \g38847/_0_  ;
  output \g38848/_0_  ;
  output \g38849/_0_  ;
  output \g38853/_0_  ;
  output \g38857/_0_  ;
  output \g38872/_0_  ;
  output \g38882/_0_  ;
  output \g38884/_0_  ;
  output \g38885/_0_  ;
  output \g38886/_0_  ;
  output \g38887/_0_  ;
  output \g38931/_0_  ;
  output \g38952/_0_  ;
  output \g38960/_0_  ;
  output \g38971/_0_  ;
  output \g38973/_0_  ;
  output \g38974/_0_  ;
  output \g38975/_0_  ;
  output \g38976/_0_  ;
  output \g38978/_0_  ;
  output \g38981/_0_  ;
  output \g38986/_0_  ;
  output \g38987/_0_  ;
  output \g39001/_3_  ;
  output \g39003/_3_  ;
  output \g39009/_3_  ;
  output \g39011/_3_  ;
  output \g39013/_3_  ;
  output \g39015/_2_  ;
  output \g39017/_2_  ;
  output \g39019/_2_  ;
  output \g39021/_2_  ;
  output \g39060/_0_  ;
  output \g39061/_3_  ;
  output \g39062/_0_  ;
  output \g39063/_0_  ;
  output \g39065/_0_  ;
  output \g39066/_0_  ;
  output \g39093/_0_  ;
  output \g39099/_2_  ;
  output \g39118/_0_  ;
  output \g39123/_0_  ;
  output \g39174/_0_  ;
  output \g39175/_0_  ;
  output \g39176/_0_  ;
  output \g39177/_0_  ;
  output \g39178/_0_  ;
  output \g39185/_0_  ;
  output \g39186/_0_  ;
  output \g39187/_0_  ;
  output \g39188/_0_  ;
  output \g39194/_0_  ;
  output \g39195/_0_  ;
  output \g39196/_0_  ;
  output \g39197/_0_  ;
  output \g39198/_0_  ;
  output \g39199/_0_  ;
  output \g39200/_0_  ;
  output \g39201/_0_  ;
  output \g39202/_0_  ;
  output \g39203/_0_  ;
  output \g39204/_0_  ;
  output \g39216/_3_  ;
  output \g39217/_3_  ;
  output \g39218/_0_  ;
  output \g39219/_0_  ;
  output \g39220/_0_  ;
  output \g39221/_0_  ;
  output \g39299/_0_  ;
  output \g39300/_0_  ;
  output \g39301/_0_  ;
  output \g39302/_0_  ;
  output \g39303/_0_  ;
  output \g39304/_0_  ;
  output \g39305/_0_  ;
  output \g39306/_0_  ;
  output \g39307/_0_  ;
  output \g39308/_0_  ;
  output \g39309/_0_  ;
  output \g39310/_0_  ;
  output \g39311/_0_  ;
  output \g39315/_0_  ;
  output \g39318/_0_  ;
  output \g39321/_0_  ;
  output \g39322/_0_  ;
  output \g39323/_0_  ;
  output \g39333/_0_  ;
  output \g39334/_0_  ;
  output \g39336/_0_  ;
  output \g39338/_0_  ;
  output \g39339/_0_  ;
  output \g39340/_0_  ;
  output \g39341/_0_  ;
  output \g39342/_0_  ;
  output \g39343/_0_  ;
  output \g39344/_0_  ;
  output \g39345/_0_  ;
  output \g39346/_0_  ;
  output \g39349/_0_  ;
  output \g39352/_3_  ;
  output \g39354/_3_  ;
  output \g39371/_3_  ;
  output \g39372/_3_  ;
  output \g39373/_3_  ;
  output \g39374/_3_  ;
  output \g39376/_0_  ;
  output \g39377/_0_  ;
  output \g39471/_0_  ;
  output \g39472/_0_  ;
  output \g39473/_0_  ;
  output \g39474/_0_  ;
  output \g39475/_0_  ;
  output \g39476/_0_  ;
  output \g39477/_0_  ;
  output \g39478/_0_  ;
  output \g39479/_0_  ;
  output \g39480/_0_  ;
  output \g39481/_0_  ;
  output \g39482/_0_  ;
  output \g39483/_0_  ;
  output \g39484/_0_  ;
  output \g39485/_0_  ;
  output \g39486/_0_  ;
  output \g39487/_0_  ;
  output \g39488/_0_  ;
  output \g39492/_0_  ;
  output \g39497/_0_  ;
  output \g39501/_0_  ;
  output \g39502/_0_  ;
  output \g39503/_0_  ;
  output \g39504/_0_  ;
  output \g39505/_0_  ;
  output \g39506/_0_  ;
  output \g39539/_0_  ;
  output \g39541/_0_  ;
  output \g39542/_0_  ;
  output \g39543/_0_  ;
  output \g39544/_0_  ;
  output \g39545/_0_  ;
  output \g39546/_0_  ;
  output \g39547/_0_  ;
  output \g39550/_0_  ;
  output \g39551/_0_  ;
  output \g39563/_0_  ;
  output \g39568/_00_  ;
  output \g39617/_0_  ;
  output \g39618/_0_  ;
  output \g39621/_0_  ;
  output \g39622/_0_  ;
  output \g39623/_0_  ;
  output \g39624/_00_  ;
  output \g39685/_0_  ;
  output \g39690/_0_  ;
  output \g39693/_0_  ;
  output \g39695/_0_  ;
  output \g39697/_0_  ;
  output \g39706/_0_  ;
  output \g39749/_0_  ;
  output \g39750/_0_  ;
  output \g39751/_0_  ;
  output \g39752/_0_  ;
  output \g39753/_0_  ;
  output \g39754/_0_  ;
  output \g39755/_0_  ;
  output \g39756/_0_  ;
  output \g39757/_0_  ;
  output \g39758/_0_  ;
  output \g39759/_0_  ;
  output \g39760/_0_  ;
  output \g39761/_0_  ;
  output \g39762/_0_  ;
  output \g39763/_0_  ;
  output \g39764/_0_  ;
  output \g39765/_0_  ;
  output \g39766/_0_  ;
  output \g39767/_0_  ;
  output \g39768/_0_  ;
  output \g39769/_0_  ;
  output \g39770/_0_  ;
  output \g39772/_0_  ;
  output \g39773/_0_  ;
  output \g39775/_3_  ;
  output \g39776/_3_  ;
  output \g39777/_3_  ;
  output \g39778/_3_  ;
  output \g39779/_3_  ;
  output \g39780/_3_  ;
  output \g39781/_3_  ;
  output \g39782/_3_  ;
  output \g39788/_3_  ;
  output \g39799/_0_  ;
  output \g39800/_0_  ;
  output \g39801/_0_  ;
  output \g39802/_0_  ;
  output \g39927/_0_  ;
  output \g39928/_0_  ;
  output \g39929/_0_  ;
  output \g39930/_0_  ;
  output \g39931/_0_  ;
  output \g39932/_0_  ;
  output \g39933/_0_  ;
  output \g39934/_0_  ;
  output \g39935/_0_  ;
  output \g39936/_0_  ;
  output \g39937/_0_  ;
  output \g39938/_0_  ;
  output \g39939/_0_  ;
  output \g39940/_0_  ;
  output \g39942/_0_  ;
  output \g39943/_0_  ;
  output \g39944/_0_  ;
  output \g39945/_0_  ;
  output \g39956/_0_  ;
  output \g39957/_0_  ;
  output \g39958/_0_  ;
  output \g39959/_0_  ;
  output \g39960/_0_  ;
  output \g39961/_0_  ;
  output \g39962/_0_  ;
  output \g39963/_0_  ;
  output \g39964/_0_  ;
  output \g39969/_0_  ;
  output \g39974/_0_  ;
  output \g39975/_0_  ;
  output \g39993/_0_  ;
  output \g39994/_0_  ;
  output \g40003/_0_  ;
  output \g40004/_0_  ;
  output \g40005/_0_  ;
  output \g40006/_0_  ;
  output \g40016/_0_  ;
  output \g40023/_3_  ;
  output \g40033/_0_  ;
  output \g40034/_0_  ;
  output \g40035/_0_  ;
  output \g40036/_0_  ;
  output \g40037/_0_  ;
  output \g40038/_0_  ;
  output \g40199/_0_  ;
  output \g40200/_0_  ;
  output \g40201/_0_  ;
  output \g40202/_0_  ;
  output \g40203/_0_  ;
  output \g40204/_0_  ;
  output \g40205/_0_  ;
  output \g40206/_0_  ;
  output \g40207/_0_  ;
  output \g40208/_0_  ;
  output \g40209/_0_  ;
  output \g40210/_0_  ;
  output \g40224/_0_  ;
  output \g40225/_0_  ;
  output \g40226/_0_  ;
  output \g40227/_0_  ;
  output \g40234/_0_  ;
  output \g40235/_0_  ;
  output \g40236/_0_  ;
  output \g40237/_0_  ;
  output \g40238/_0_  ;
  output \g40239/_0_  ;
  output \g40240/_0_  ;
  output \g40241/_0_  ;
  output \g40242/_0_  ;
  output \g40243/_0_  ;
  output \g40244/_0_  ;
  output \g40246/_0_  ;
  output \g40247/_0_  ;
  output \g40248/_0_  ;
  output \g40249/_0_  ;
  output \g40250/_0_  ;
  output \g40251/_0_  ;
  output \g40252/_0_  ;
  output \g40253/_0_  ;
  output \g40254/_0_  ;
  output \g40255/_0_  ;
  output \g40257/_0_  ;
  output \g40258/_0_  ;
  output \g40262/_0_  ;
  output \g40264/_0_  ;
  output \g40265/_0_  ;
  output \g40266/_0_  ;
  output \g40267/_0_  ;
  output \g40268/_0_  ;
  output \g40269/_0_  ;
  output \g40270/_0_  ;
  output \g40271/_0_  ;
  output \g40272/_0_  ;
  output \g40273/_0_  ;
  output \g40274/_0_  ;
  output \g40275/_0_  ;
  output \g40276/_0_  ;
  output \g40277/_0_  ;
  output \g40278/_0_  ;
  output \g40280/_2_  ;
  output \g40281/_0_  ;
  output \g40282/_0_  ;
  output \g40283/_0_  ;
  output \g40284/_0_  ;
  output \g40285/_0_  ;
  output \g40286/_0_  ;
  output \g40287/_0_  ;
  output \g40288/_0_  ;
  output \g40289/_0_  ;
  output \g40290/_0_  ;
  output \g40291/_0_  ;
  output \g40297/_0_  ;
  output \g40298/_0_  ;
  output \g40299/_0_  ;
  output \g40300/_0_  ;
  output \g40301/_0_  ;
  output \g40302/_0_  ;
  output \g40303/_0_  ;
  output \g40304/_0_  ;
  output \g40306/_0_  ;
  output \g40307/_0_  ;
  output \g40308/_0_  ;
  output \g40309/_0_  ;
  output \g40310/_0_  ;
  output \g40311/_0_  ;
  output \g40312/_0_  ;
  output \g40313/_0_  ;
  output \g40314/_0_  ;
  output \g40315/_0_  ;
  output \g40316/_0_  ;
  output \g40317/_0_  ;
  output \g40318/_0_  ;
  output \g40319/_0_  ;
  output \g40320/_0_  ;
  output \g40324/_0_  ;
  output \g40325/_0_  ;
  output \g40326/_0_  ;
  output \g40327/_0_  ;
  output \g40328/_0_  ;
  output \g40329/_0_  ;
  output \g40330/_0_  ;
  output \g40331/_0_  ;
  output \g40332/_0_  ;
  output \g40333/_0_  ;
  output \g40334/_0_  ;
  output \g40335/_0_  ;
  output \g40336/_0_  ;
  output \g40337/_0_  ;
  output \g40338/_0_  ;
  output \g40339/_0_  ;
  output \g40340/_0_  ;
  output \g40341/_0_  ;
  output \g40342/_0_  ;
  output \g40343/_0_  ;
  output \g40344/_0_  ;
  output \g40345/_0_  ;
  output \g40346/_0_  ;
  output \g40347/_0_  ;
  output \g40350/_0_  ;
  output \g40353/_0_  ;
  output \g40354/_0_  ;
  output \g40355/_0_  ;
  output \g40374/_0_  ;
  output \g40457/_0_  ;
  output \g40458/_0_  ;
  output \g40549/_0_  ;
  output \g40550/_0_  ;
  output \g40551/_0_  ;
  output \g40552/_0_  ;
  output \g40553/_0_  ;
  output \g40554/_0_  ;
  output \g40556/_0_  ;
  output \g40557/_0_  ;
  output \g40558/_0_  ;
  output \g40559/_0_  ;
  output \g40561/_0_  ;
  output \g40562/_0_  ;
  output \g40563/_0_  ;
  output \g40565/_0_  ;
  output \g40566/_0_  ;
  output \g40567/_0_  ;
  output \g40569/_0_  ;
  output \g40570/_0_  ;
  output \g40571/_0_  ;
  output \g40572/_0_  ;
  output \g40573/_0_  ;
  output \g40574/_0_  ;
  output \g40575/_0_  ;
  output \g40576/_0_  ;
  output \g40577/_0_  ;
  output \g40578/_0_  ;
  output \g40579/_0_  ;
  output \g40580/_0_  ;
  output \g40581/_0_  ;
  output \g40582/_0_  ;
  output \g40583/_0_  ;
  output \g40584/_0_  ;
  output \g40586/_0_  ;
  output \g40587/_0_  ;
  output \g40588/_0_  ;
  output \g40589/_0_  ;
  output \g40591/_0_  ;
  output \g40592/_0_  ;
  output \g40593/_0_  ;
  output \g40594/_0_  ;
  output \g40595/_0_  ;
  output \g40596/_0_  ;
  output \g40597/_0_  ;
  output \g40598/_0_  ;
  output \g40599/_0_  ;
  output \g40600/_0_  ;
  output \g40601/_0_  ;
  output \g40602/_0_  ;
  output \g40603/_0_  ;
  output \g40604/_0_  ;
  output \g40605/_0_  ;
  output \g40606/_0_  ;
  output \g40607/_0_  ;
  output \g40608/_0_  ;
  output \g40609/_0_  ;
  output \g40610/_0_  ;
  output \g40611/_0_  ;
  output \g40612/_0_  ;
  output \g40613/_0_  ;
  output \g40614/_0_  ;
  output \g40617/_0_  ;
  output \g40629/_0_  ;
  output \g40632/_0_  ;
  output \g40633/_0_  ;
  output \g40634/_0_  ;
  output \g40635/_0_  ;
  output \g40636/_0_  ;
  output \g40637/_0_  ;
  output \g40638/_0_  ;
  output \g40639/_0_  ;
  output \g40640/_0_  ;
  output \g40641/_0_  ;
  output \g40642/_0_  ;
  output \g40643/_0_  ;
  output \g40644/_0_  ;
  output \g40645/_0_  ;
  output \g40646/_0_  ;
  output \g40647/_0_  ;
  output \g40648/_0_  ;
  output \g40649/_0_  ;
  output \g40650/_0_  ;
  output \g40651/_0_  ;
  output \g40652/_0_  ;
  output \g40653/_0_  ;
  output \g40654/_0_  ;
  output \g40655/_0_  ;
  output \g40661/_0_  ;
  output \g40663/_0_  ;
  output \g40664/_0_  ;
  output \g40665/_0_  ;
  output \g40666/_0_  ;
  output \g40667/_0_  ;
  output \g40668/_0_  ;
  output \g40669/_0_  ;
  output \g40670/_0_  ;
  output \g40671/_0_  ;
  output \g40672/_0_  ;
  output \g40673/_0_  ;
  output \g40674/_0_  ;
  output \g40675/_0_  ;
  output \g40676/_0_  ;
  output \g40677/_0_  ;
  output \g40678/_0_  ;
  output \g40679/_0_  ;
  output \g40680/_0_  ;
  output \g40681/_0_  ;
  output \g40682/_0_  ;
  output \g40683/_0_  ;
  output \g40684/_0_  ;
  output \g40685/_0_  ;
  output \g40689/_0_  ;
  output \g40690/_0_  ;
  output \g40691/_0_  ;
  output \g40692/_0_  ;
  output \g40693/_0_  ;
  output \g40694/_0_  ;
  output \g40695/_0_  ;
  output \g40696/_0_  ;
  output \g40697/_0_  ;
  output \g40698/_0_  ;
  output \g40699/_0_  ;
  output \g40700/_0_  ;
  output \g40701/_0_  ;
  output \g40702/_0_  ;
  output \g40703/_0_  ;
  output \g40704/_0_  ;
  output \g40705/_0_  ;
  output \g40706/_0_  ;
  output \g40707/_0_  ;
  output \g40708/_0_  ;
  output \g40709/_0_  ;
  output \g40710/_0_  ;
  output \g40711/_0_  ;
  output \g40712/_0_  ;
  output \g40758/_00_  ;
  output \g40759/_0_  ;
  output \g40812/_0_  ;
  output \g40816/_0_  ;
  output \g40817/_0_  ;
  output \g40818/_0_  ;
  output \g40819/_0_  ;
  output \g40820/_0_  ;
  output \g40822/_3_  ;
  output \g40823/_3_  ;
  output \g40824/_3_  ;
  output \g40825/_3_  ;
  output \g40849/_3_  ;
  output \g40915/_0_  ;
  output \g40916/_0_  ;
  output \g40917/_0_  ;
  output \g40920/_0_  ;
  output \g40923/_0_  ;
  output \g40926/_0_  ;
  output \g40927/_0_  ;
  output \g40930/_0_  ;
  output \g40931/_0_  ;
  output \g41138/_0_  ;
  output \g41152/_0_  ;
  output \g41180/_0_  ;
  output \g41185/_0_  ;
  output \g41186/_0_  ;
  output \g41187/_0_  ;
  output \g41189/_0_  ;
  output \g41190/_0_  ;
  output \g41191/_0_  ;
  output \g41192/_0_  ;
  output \g41193/_0_  ;
  output \g41195/_0_  ;
  output \g41199/_0_  ;
  output \g41207/_0_  ;
  output \g41221/_0_  ;
  output \g41226/_0_  ;
  output \g41227/_0_  ;
  output \g41230/_0_  ;
  output \g41231/_0_  ;
  output \g41234/_0_  ;
  output \g41238/_0_  ;
  output \g41239/_0_  ;
  output \g41275/_0_  ;
  output \g41277/_0_  ;
  output \g41278/_0_  ;
  output \g41279/_0_  ;
  output \g41280/_0_  ;
  output \g41281/_0_  ;
  output \g41282/_0_  ;
  output \g41283/_0_  ;
  output \g41284/_0_  ;
  output \g41285/_0_  ;
  output \g41286/_0_  ;
  output \g41287/_0_  ;
  output \g41288/_0_  ;
  output \g41289/_0_  ;
  output \g41291/_3_  ;
  output \g41330/_0_  ;
  output \g41332/_0_  ;
  output \g41334/_0_  ;
  output \g41340/_0_  ;
  output \g41343/_0_  ;
  output \g41345/_0_  ;
  output \g41348/_0_  ;
  output \g41349/_0_  ;
  output \g41350/_0_  ;
  output \g41351/_0_  ;
  output \g41356/_0_  ;
  output \g41394/_0_  ;
  output \g41423/_0_  ;
  output \g41426/_3_  ;
  output \g41427/_3_  ;
  output \g41428/_3_  ;
  output \g41429/_3_  ;
  output \g41430/_3_  ;
  output \g41431/_3_  ;
  output \g41432/_3_  ;
  output \g41433/_3_  ;
  output \g41434/_3_  ;
  output \g41435/_3_  ;
  output \g41436/_3_  ;
  output \g41437/_3_  ;
  output \g41438/_3_  ;
  output \g41439/_3_  ;
  output \g41440/_3_  ;
  output \g41441/_3_  ;
  output \g41442/_0_  ;
  output \g41445/_3_  ;
  output \g41446/_0_  ;
  output \g41449/_0_  ;
  output \g41464/_0_  ;
  output \g41466/_0_  ;
  output \g41468/_0_  ;
  output \g41469/_0_  ;
  output \g41471/_0_  ;
  output \g41795/_0_  ;
  output \g41799/_0_  ;
  output \g41800/_0_  ;
  output \g41801/_0_  ;
  output \g41802/_0_  ;
  output \g41803/_0_  ;
  output \g41804/_0_  ;
  output \g41805/_0_  ;
  output \g41806/_0_  ;
  output \g41807/_0_  ;
  output \g41808/_0_  ;
  output \g41809/_0_  ;
  output \g41810/_0_  ;
  output \g41811/_0_  ;
  output \g41812/_0_  ;
  output \g41814/_0_  ;
  output \g41815/_0_  ;
  output \g41816/_0_  ;
  output \g41817/_0_  ;
  output \g41818/_0_  ;
  output \g41819/_0_  ;
  output \g41820/_0_  ;
  output \g41821/_0_  ;
  output \g41822/_0_  ;
  output \g41823/_0_  ;
  output \g41825/_0_  ;
  output \g41826/_0_  ;
  output \g41827/_0_  ;
  output \g41828/_0_  ;
  output \g41829/_0_  ;
  output \g41830/_0_  ;
  output \g41831/_0_  ;
  output \g41832/_0_  ;
  output \g41833/_0_  ;
  output \g41834/_0_  ;
  output \g41835/_0_  ;
  output \g41836/_0_  ;
  output \g41837/_0_  ;
  output \g41838/_0_  ;
  output \g41839/_0_  ;
  output \g41840/_0_  ;
  output \g41841/_0_  ;
  output \g41842/_0_  ;
  output \g41843/_0_  ;
  output \g41844/_0_  ;
  output \g41845/_0_  ;
  output \g41846/_0_  ;
  output \g41847/_0_  ;
  output \g41848/_0_  ;
  output \g41849/_0_  ;
  output \g41850/_0_  ;
  output \g41851/_0_  ;
  output \g41852/_0_  ;
  output \g41853/_0_  ;
  output \g41854/_0_  ;
  output \g41855/_0_  ;
  output \g41856/_0_  ;
  output \g41857/_0_  ;
  output \g41858/_0_  ;
  output \g41859/_0_  ;
  output \g41860/_0_  ;
  output \g41861/_0_  ;
  output \g41862/_0_  ;
  output \g41863/_0_  ;
  output \g41864/_0_  ;
  output \g41865/_0_  ;
  output \g41866/_0_  ;
  output \g41867/_0_  ;
  output \g41868/_0_  ;
  output \g41869/_0_  ;
  output \g41870/_0_  ;
  output \g41871/_0_  ;
  output \g41872/_0_  ;
  output \g41873/_0_  ;
  output \g41874/_0_  ;
  output \g41875/_0_  ;
  output \g41876/_0_  ;
  output \g41877/_0_  ;
  output \g41878/_0_  ;
  output \g41879/_0_  ;
  output \g41880/_0_  ;
  output \g41881/_0_  ;
  output \g41882/_0_  ;
  output \g41883/_0_  ;
  output \g41884/_0_  ;
  output \g41885/_0_  ;
  output \g41886/_0_  ;
  output \g41887/_0_  ;
  output \g41888/_0_  ;
  output \g41889/_0_  ;
  output \g41890/_0_  ;
  output \g41891/_0_  ;
  output \g41902/_0_  ;
  output \g41904/_0_  ;
  output \g41906/_0_  ;
  output \g41907/_0_  ;
  output \g41954/_0_  ;
  output \g41955/_0_  ;
  output \g41956/_0_  ;
  output \g41957/_0_  ;
  output \g41958/_0_  ;
  output \g41959/_0_  ;
  output \g41960/_0_  ;
  output \g41962/_0_  ;
  output \g41963/_0_  ;
  output \g41964/_0_  ;
  output \g41965/_0_  ;
  output \g41966/_0_  ;
  output \g41967/_0_  ;
  output \g41968/_0_  ;
  output \g41969/_0_  ;
  output \g41970/_0_  ;
  output \g41971/_0_  ;
  output \g41972/_0_  ;
  output \g41973/_0_  ;
  output \g41974/_0_  ;
  output \g41975/_0_  ;
  output \g41976/_0_  ;
  output \g41977/_0_  ;
  output \g41978/_0_  ;
  output \g41979/_0_  ;
  output \g42062/_0_  ;
  output \g42079/_0_  ;
  output \g42142/_0_  ;
  output \g42143/_0_  ;
  output \g42144/_0_  ;
  output \g42154/_0_  ;
  output \g42157/_0_  ;
  output \g42160/_0_  ;
  output \g42181/_0_  ;
  output \g42203/_0_  ;
  output \g42204/_3_  ;
  output \g42205/_3_  ;
  output \g42206/_3_  ;
  output \g42208/_0_  ;
  output \g42220/_0_  ;
  output \g42225/_0_  ;
  output \g42251/_0_  ;
  output \g42273/_0_  ;
  output \g42335/_0_  ;
  output \g42357/_0_  ;
  output \g42380/_0_  ;
  output \g42381/_0_  ;
  output \g42383/_0_  ;
  output \g42386/_0_  ;
  output \g42388/_0_  ;
  output \g42475/_0_  ;
  output \g42476/_0_  ;
  output \g42477/_0_  ;
  output \g42478/_0_  ;
  output \g42479/_0_  ;
  output \g42480/_0_  ;
  output \g42481/_0_  ;
  output \g42482/_0_  ;
  output \g42483/_0_  ;
  output \g42484/_0_  ;
  output \g42485/_0_  ;
  output \g42486/_0_  ;
  output \g42487/_0_  ;
  output \g42488/_0_  ;
  output \g42490/_0_  ;
  output \g42491/_0_  ;
  output \g42493/_0_  ;
  output \g42494/_0_  ;
  output \g42495/_0_  ;
  output \g42496/_0_  ;
  output \g42497/_0_  ;
  output \g42498/_0_  ;
  output \g42499/_0_  ;
  output \g42500/_0_  ;
  output \g42501/_0_  ;
  output \g42502/_0_  ;
  output \g42503/_0_  ;
  output \g42504/_0_  ;
  output \g42505/_0_  ;
  output \g42506/_0_  ;
  output \g42507/_0_  ;
  output \g42508/_0_  ;
  output \g42509/_0_  ;
  output \g42510/_0_  ;
  output \g42511/_0_  ;
  output \g42512/_0_  ;
  output \g42513/_0_  ;
  output \g42514/_0_  ;
  output \g42515/_0_  ;
  output \g42516/_0_  ;
  output \g42517/_0_  ;
  output \g42518/_0_  ;
  output \g42519/_0_  ;
  output \g42521/_0_  ;
  output \g42522/_0_  ;
  output \g42523/_0_  ;
  output \g42524/_0_  ;
  output \g42525/_0_  ;
  output \g42526/_0_  ;
  output \g42527/_0_  ;
  output \g42528/_0_  ;
  output \g42529/_0_  ;
  output \g42530/_0_  ;
  output \g42531/_0_  ;
  output \g42532/_0_  ;
  output \g42533/_0_  ;
  output \g42534/_0_  ;
  output \g42535/_0_  ;
  output \g42536/_0_  ;
  output \g42537/_0_  ;
  output \g42538/_0_  ;
  output \g42539/_0_  ;
  output \g42540/_0_  ;
  output \g42541/_0_  ;
  output \g42542/_0_  ;
  output \g42543/_0_  ;
  output \g42544/_0_  ;
  output \g42545/_0_  ;
  output \g42548/_0_  ;
  output \g42557/_0_  ;
  output \g42564/_0_  ;
  output \g42565/_0_  ;
  output \g42566/_0_  ;
  output \g42567/_0_  ;
  output \g42568/_0_  ;
  output \g42569/_0_  ;
  output \g42570/_0_  ;
  output \g42571/_0_  ;
  output \g42572/_0_  ;
  output \g42573/_0_  ;
  output \g42574/_0_  ;
  output \g42575/_0_  ;
  output \g42576/_0_  ;
  output \g42577/_0_  ;
  output \g42578/_0_  ;
  output \g42581/_0_  ;
  output \g42589/_0_  ;
  output \g42590/_0_  ;
  output \g42591/_0_  ;
  output \g42592/_0_  ;
  output \g42593/_0_  ;
  output \g42594/_0_  ;
  output \g42595/_0_  ;
  output \g42596/_0_  ;
  output \g42597/_0_  ;
  output \g42598/_0_  ;
  output \g42599/_0_  ;
  output \g42600/_0_  ;
  output \g42601/_0_  ;
  output \g42602/_0_  ;
  output \g42603/_0_  ;
  output \g42604/_0_  ;
  output \g42605/_0_  ;
  output \g42606/_0_  ;
  output \g42607/_0_  ;
  output \g42608/_0_  ;
  output \g42609/_0_  ;
  output \g42610/_0_  ;
  output \g42611/_0_  ;
  output \g42612/_0_  ;
  output \g42613/_0_  ;
  output \g42614/_0_  ;
  output \g42615/_0_  ;
  output \g42616/_0_  ;
  output \g42617/_0_  ;
  output \g42618/_0_  ;
  output \g42619/_0_  ;
  output \g42620/_0_  ;
  output \g42622/_0_  ;
  output \g42623/_0_  ;
  output \g42627/_0_  ;
  output \g42628/_0_  ;
  output \g42629/_0_  ;
  output \g42630/_0_  ;
  output \g42631/_0_  ;
  output \g42632/_0_  ;
  output \g42633/_0_  ;
  output \g42634/_0_  ;
  output \g42635/_0_  ;
  output \g42636/_0_  ;
  output \g42637/_0_  ;
  output \g42638/_0_  ;
  output \g42639/_0_  ;
  output \g42640/_0_  ;
  output \g42641/_0_  ;
  output \g42642/_0_  ;
  output \g42643/_0_  ;
  output \g42644/_0_  ;
  output \g42645/_0_  ;
  output \g42646/_0_  ;
  output \g42647/_0_  ;
  output \g42648/_0_  ;
  output \g42649/_0_  ;
  output \g42650/_0_  ;
  output \g42666/_0_  ;
  output \g42667/_0_  ;
  output \g42668/_0_  ;
  output \g42669/_0_  ;
  output \g42670/_0_  ;
  output \g42671/_0_  ;
  output \g42672/_0_  ;
  output \g42673/_0_  ;
  output \g42674/_0_  ;
  output \g42675/_0_  ;
  output \g42676/_0_  ;
  output \g42677/_0_  ;
  output \g42678/_0_  ;
  output \g42680/_0_  ;
  output \g42681/_0_  ;
  output \g42685/_0_  ;
  output \g42686/_0_  ;
  output \g42688/_0_  ;
  output \g42689/_0_  ;
  output \g42690/_0_  ;
  output \g42691/_0_  ;
  output \g42692/_0_  ;
  output \g42693/_0_  ;
  output \g42694/_0_  ;
  output \g42695/_0_  ;
  output \g42696/_0_  ;
  output \g42697/_0_  ;
  output \g42698/_0_  ;
  output \g42699/_0_  ;
  output \g42700/_0_  ;
  output \g42701/_0_  ;
  output \g42702/_0_  ;
  output \g42703/_0_  ;
  output \g42704/_0_  ;
  output \g42705/_0_  ;
  output \g42706/_0_  ;
  output \g42707/_0_  ;
  output \g42708/_0_  ;
  output \g42709/_0_  ;
  output \g42710/_0_  ;
  output \g42711/_0_  ;
  output \g42712/_0_  ;
  output \g42713/_0_  ;
  output \g42715/_0_  ;
  output \g42716/_0_  ;
  output \g42717/_0_  ;
  output \g42718/_0_  ;
  output \g42723/_1_  ;
  output \g42727/_0_  ;
  output \g42728/_0_  ;
  output \g42729/_0_  ;
  output \g42730/_0_  ;
  output \g42731/_0_  ;
  output \g42732/_0_  ;
  output \g42733/_0_  ;
  output \g42734/_0_  ;
  output \g42735/_0_  ;
  output \g42736/_0_  ;
  output \g42737/_0_  ;
  output \g42738/_0_  ;
  output \g42739/_0_  ;
  output \g42740/_0_  ;
  output \g42741/_0_  ;
  output \g42742/_0_  ;
  output \g42743/_0_  ;
  output \g42744/_0_  ;
  output \g42745/_0_  ;
  output \g42746/_0_  ;
  output \g42747/_0_  ;
  output \g42748/_0_  ;
  output \g42749/_0_  ;
  output \g42750/_0_  ;
  output \g42751/_0_  ;
  output \g42754/_0_  ;
  output \g42767/_0_  ;
  output \g42768/_0_  ;
  output \g42772/_0_  ;
  output \g42773/_0_  ;
  output \g42774/_0_  ;
  output \g42775/_0_  ;
  output \g42776/_0_  ;
  output \g42777/_0_  ;
  output \g42778/_0_  ;
  output \g42779/_0_  ;
  output \g42780/_0_  ;
  output \g42781/_0_  ;
  output \g42782/_0_  ;
  output \g42783/_0_  ;
  output \g42784/_0_  ;
  output \g42785/_0_  ;
  output \g42790/_0_  ;
  output \g42791/_0_  ;
  output \g42792/_0_  ;
  output \g42793/_0_  ;
  output \g42794/_0_  ;
  output \g42795/_0_  ;
  output \g42796/_0_  ;
  output \g42797/_0_  ;
  output \g42798/_0_  ;
  output \g42799/_0_  ;
  output \g42800/_0_  ;
  output \g42801/_0_  ;
  output \g42802/_0_  ;
  output \g42803/_0_  ;
  output \g42804/_0_  ;
  output \g42805/_0_  ;
  output \g42806/_0_  ;
  output \g42807/_0_  ;
  output \g42808/_0_  ;
  output \g42809/_0_  ;
  output \g42810/_0_  ;
  output \g42811/_0_  ;
  output \g42812/_0_  ;
  output \g42813/_0_  ;
  output \g42814/_0_  ;
  output \g42815/_0_  ;
  output \g42816/_0_  ;
  output \g42817/_0_  ;
  output \g42818/_0_  ;
  output \g42819/_0_  ;
  output \g42820/_0_  ;
  output \g42821/_0_  ;
  output \g42824/_0_  ;
  output \g42825/_0_  ;
  output \g42826/_0_  ;
  output \g42827/_0_  ;
  output \g42828/_0_  ;
  output \g42829/_0_  ;
  output \g42830/_0_  ;
  output \g42831/_0_  ;
  output \g42832/_0_  ;
  output \g42833/_0_  ;
  output \g42834/_0_  ;
  output \g42835/_0_  ;
  output \g42836/_0_  ;
  output \g42837/_0_  ;
  output \g42838/_0_  ;
  output \g42839/_0_  ;
  output \g42840/_0_  ;
  output \g42841/_0_  ;
  output \g42842/_0_  ;
  output \g42843/_0_  ;
  output \g42844/_0_  ;
  output \g42845/_0_  ;
  output \g42846/_0_  ;
  output \g42907/_0_  ;
  output \g42914/_0_  ;
  output \g42924/_0_  ;
  output \g42925/_0_  ;
  output \g42926/_0_  ;
  output \g42927/_0_  ;
  output \g42928/_0_  ;
  output \g42929/_0_  ;
  output \g42930/_0_  ;
  output \g42931/_0_  ;
  output \g42933/_0_  ;
  output \g42941/_0_  ;
  output \g42947/_0_  ;
  output \g42950/_0_  ;
  output \g42955/_0_  ;
  output \g42956/_0_  ;
  output \g42972/_3_  ;
  output \g42973/_3_  ;
  output \g42974/_3_  ;
  output \g43178/_0_  ;
  output \g43179/_0_  ;
  output \g43184/_0_  ;
  output \g43186/_0_  ;
  output \g43187/_0_  ;
  output \g43190/_0_  ;
  output \g43191/_0_  ;
  output \g43192/_0_  ;
  output \g43202/_0_  ;
  output \g43205/_0_  ;
  output \g43206/_0_  ;
  output \g43207/_0_  ;
  output \g43209/_2_  ;
  output \g43228/_0_  ;
  output \g43233/_0_  ;
  output \g43235/_0_  ;
  output \g43236/_0_  ;
  output \g43237/_0_  ;
  output \g43238/_0_  ;
  output \g43280/_0_  ;
  output \g43287/_0_  ;
  output \g43289/_0_  ;
  output \g43290/_0_  ;
  output \g43291/_0_  ;
  output \g43292/_0_  ;
  output \g43303/_0_  ;
  output \g43311/_0_  ;
  output \g43312/_0_  ;
  output \g43363/_0_  ;
  output \g43364/_0_  ;
  output \g43366/_0_  ;
  output \g43367/_0_  ;
  output \g43370/_0_  ;
  output \g43371/_0_  ;
  output \g43374/_0_  ;
  output \g43413/_0_  ;
  output \g43414/_0_  ;
  output \g43415/_0_  ;
  output \g43416/_0_  ;
  output \g43422/_0_  ;
  output \g43427/_0_  ;
  output \g43428/_0_  ;
  output \g43528/_1__syn_2  ;
  output \g43630/_0_  ;
  output \g43633/_3_  ;
  output \g43647/_0_  ;
  output \g43648/_0_  ;
  output \g43656/_0_  ;
  output \g43657/_0_  ;
  output \g43667/_0_  ;
  output \g43668/_0_  ;
  output \g43675/_0_  ;
  output \g43678/_0_  ;
  output \g43787/_0_  ;
  output \g44055/_0_  ;
  output \g44092/_0_  ;
  output \g44093/_0_  ;
  output \g44176/_0_  ;
  output \g44181/_0_  ;
  output \g44433/_0_  ;
  output \g44510/_0_  ;
  output \g44515/_2_  ;
  output \g44522/_0_  ;
  output \g44529/_2_  ;
  output \g44537/_2_  ;
  output \g44544/_2_  ;
  output \g44594/_0_  ;
  output \g44695/_0_  ;
  output \g44697/_0_  ;
  output \g44699/_0_  ;
  output \g44700/_0_  ;
  output \g44843/_0_  ;
  output \g44844/_0_  ;
  output \g44879/_0_  ;
  output \g44880/_0_  ;
  output \g44881/_0_  ;
  output \g44882/_0_  ;
  output \g44906/_2_  ;
  output \g44910/_0_  ;
  output \g44912/_0_  ;
  output \g44954/_0_  ;
  output \g45000/_0_  ;
  output \g45001/_0_  ;
  output \g45002/_0_  ;
  output \g45003/_0_  ;
  output \g45021/_1_  ;
  output \g45025/_0_  ;
  output \g45051/_0_  ;
  output \g45104/_0_  ;
  output \g45111/_0_  ;
  output \g45112/_0_  ;
  output \g45116/_0_  ;
  output \g45155/_0_  ;
  output \g45238/_0_  ;
  output \g45239/_0_  ;
  output \g45240/_0_  ;
  output \g45241/_0_  ;
  output \g45249/_0_  ;
  output \g45257/_0_  ;
  output \g45332/_0_  ;
  output \g45334/_0_  ;
  output \g45336/_0_  ;
  output \g45337/_0_  ;
  output \g45342/_0_  ;
  output \g45459/_0_  ;
  output \g45460/_0_  ;
  output \g45466/_0_  ;
  output \g45469/_0_  ;
  output \g45470/_0_  ;
  output \g45474/_0_  ;
  output \g45475/_0_  ;
  output \g45477/_0_  ;
  output \g45481/_0_  ;
  output \g45482/_0_  ;
  output \g45487/_0_  ;
  output \g45488/_0_  ;
  output \g45518/_3_  ;
  output \g45519/_3_  ;
  output \g45520/_3_  ;
  output \g45521/_3_  ;
  output \g45522/_3_  ;
  output \g45523/_3_  ;
  output \g45524/_3_  ;
  output \g45525/_3_  ;
  output \g45526/_3_  ;
  output \g45530/_3_  ;
  output \g45531/_3_  ;
  output \g45532/_3_  ;
  output \g45533/_3_  ;
  output \g45534/_3_  ;
  output \g45535/_3_  ;
  output \g45536/_3_  ;
  output \g45559/_3_  ;
  output \g45596/_0_  ;
  output \g45605/_0_  ;
  output \g45622/_0_  ;
  output \g45623/_0_  ;
  output \g45630/_0_  ;
  output \g45747/_0_  ;
  output \g45753/_0_  ;
  output \g45796/_0_  ;
  output \g45837/_0_  ;
  output \g45882/_0_  ;
  output \g45903/_0_  ;
  output \g45912/_0_  ;
  output \g45946/_0_  ;
  output \g45999/_0_  ;
  output \g46000/_0_  ;
  output \g46001/_0_  ;
  output \g46002/_0_  ;
  output \g46012/_0_  ;
  output \g46014/_0_  ;
  output \g46017/_0_  ;
  output \g46018/_0_  ;
  output \g46021/_0_  ;
  output \g46024/_0_  ;
  output \g46026/_0_  ;
  output \g46029/_0_  ;
  output \g46053/_0_  ;
  output \g46083/_0_  ;
  output \g46093/_0_  ;
  output \g46142/_0_  ;
  output \g46154/_1__syn_2  ;
  output \g46265/_0_  ;
  output \g46266/_0_  ;
  output \g46268/_0_  ;
  output \g46270/_0_  ;
  output \g46273/_0_  ;
  output \g46274/_0_  ;
  output \g46275/_0_  ;
  output \g46276/_0_  ;
  output \g46278/_0_  ;
  output \g46385/_0_  ;
  output \g46411/_0_  ;
  output \g46414/_0_  ;
  output \g46479/_0_  ;
  output \g46520/_0_  ;
  output \g46521/_0_  ;
  output \g46530/_0_  ;
  output \g46531/_0_  ;
  output \g46597/_0_  ;
  output \g46610/_0_  ;
  output \g46617/_0_  ;
  output \g46632/_0_  ;
  output \g46637/_0_  ;
  output \g46722/_0_  ;
  output \g46723/_0_  ;
  output \g46724/_0_  ;
  output \g46725/_0_  ;
  output \g46813/_0_  ;
  output \g46842/_0_  ;
  output \g46888/_0_  ;
  output \g46891/_0_  ;
  output \g46894/_0_  ;
  output \g46905/_0_  ;
  output \g46940/_0_  ;
  output \g46992/_0_  ;
  output \g46995/_0_  ;
  output \g47037/_3_  ;
  output \g47053/_0_  ;
  output \g47140/_0_  ;
  output \g47155/_3_  ;
  output \g47209/_0_  ;
  output \g47211/_0_  ;
  output \g47213/_0_  ;
  output \g47215/_0_  ;
  output \g47337/_0_  ;
  output \g47433/_0_  ;
  output \g47972/_0_  ;
  output \g47976/_0_  ;
  output \g48081/_0_  ;
  output \g48171/_0_  ;
  output \g48227/_0_  ;
  output \g48234/_1_  ;
  output \g48257/_1_  ;
  output \g48266/_0_  ;
  output \g48281/_0_  ;
  output \g48291/_1_  ;
  output \g48322/_0_  ;
  output \g48345/_0_  ;
  output \g48429/_0_  ;
  output \g48495/_1_  ;
  output \g48549/_0_  ;
  output \g48589/_0_  ;
  output \g48642/_0_  ;
  output \g48722/_0_  ;
  output \g48748/_0_  ;
  output \g48749/_0_  ;
  output \g48763/_0_  ;
  output \g48867/_0_  ;
  output \g48876/_0_  ;
  output \g48880/_0_  ;
  output \g49023/_0_  ;
  output \g49205/_0_  ;
  output \g49314/_0_  ;
  output \g49432/_0__syn_2  ;
  output \g49512/_0_  ;
  output \g49707/_0_  ;
  output \g49737/_0_  ;
  output \g49831/_0_  ;
  output \g49922/_1_  ;
  output \g50132/_0_  ;
  output \g51376/_0_  ;
  output \g51412/_0_  ;
  output \g51822/_0_  ;
  output \g52114/_0_  ;
  output \g52156/_0_  ;
  output \g54427/_0_  ;
  output \g54557/_0_  ;
  output \g54561/_3_  ;
  output \g55079/_0_  ;
  output \sram_adr_o[0]_pad  ;
  output \sram_adr_o[10]_pad  ;
  output \sram_adr_o[11]_pad  ;
  output \sram_adr_o[12]_pad  ;
  output \sram_adr_o[13]_pad  ;
  output \sram_adr_o[14]_pad  ;
  output \sram_adr_o[1]_pad  ;
  output \sram_adr_o[2]_pad  ;
  output \sram_adr_o[3]_pad  ;
  output \sram_adr_o[4]_pad  ;
  output \sram_adr_o[5]_pad  ;
  output \sram_adr_o[6]_pad  ;
  output \sram_adr_o[7]_pad  ;
  output \sram_adr_o[8]_pad  ;
  output \sram_adr_o[9]_pad  ;
  output \sram_data_o[0]_pad  ;
  output \sram_data_o[10]_pad  ;
  output \sram_data_o[11]_pad  ;
  output \sram_data_o[12]_pad  ;
  output \sram_data_o[13]_pad  ;
  output \sram_data_o[14]_pad  ;
  output \sram_data_o[15]_pad  ;
  output \sram_data_o[16]_pad  ;
  output \sram_data_o[17]_pad  ;
  output \sram_data_o[18]_pad  ;
  output \sram_data_o[19]_pad  ;
  output \sram_data_o[1]_pad  ;
  output \sram_data_o[20]_pad  ;
  output \sram_data_o[21]_pad  ;
  output \sram_data_o[22]_pad  ;
  output \sram_data_o[23]_pad  ;
  output \sram_data_o[24]_pad  ;
  output \sram_data_o[25]_pad  ;
  output \sram_data_o[26]_pad  ;
  output \sram_data_o[27]_pad  ;
  output \sram_data_o[28]_pad  ;
  output \sram_data_o[29]_pad  ;
  output \sram_data_o[2]_pad  ;
  output \sram_data_o[30]_pad  ;
  output \sram_data_o[31]_pad  ;
  output \sram_data_o[3]_pad  ;
  output \sram_data_o[4]_pad  ;
  output \sram_data_o[5]_pad  ;
  output \sram_data_o[6]_pad  ;
  output \sram_data_o[7]_pad  ;
  output \sram_data_o[8]_pad  ;
  output \sram_data_o[9]_pad  ;
  output sram_re_o_pad ;
  output sram_we_o_pad ;
  output \u4_utmi_vend_ctrl_r_reg[0]/P0001_reg_syn_3  ;
  output \u4_utmi_vend_ctrl_r_reg[1]/P0001_reg_syn_3  ;
  output \u4_utmi_vend_ctrl_r_reg[2]/P0001_reg_syn_3  ;
  output \u4_utmi_vend_ctrl_r_reg[3]/P0001_reg_syn_3  ;
  wire n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 ;
  assign n1749 = ~TxReady_pad_i_pad & \u1_u1_tx_first_r_reg/P0001  ;
  assign n1750 = ~\u1_u1_send_zero_length_r_reg/P0001  & ~\u1_u2_send_data_r_reg/NET0131  ;
  assign n1751 = ~TxReady_pad_i_pad & ~\u1_u3_send_token_reg/P0001  ;
  assign n1752 = n1750 & n1751 ;
  assign n1753 = ~n1749 & ~n1752 ;
  assign n1754 = \DataOut_pad_o[3]_pad  & ~\u0_u0_drive_k_reg/P0001  ;
  assign n1755 = ~n1753 & n1754 ;
  assign n1756 = \u0_tx_ready_reg/NET0131  & \u1_u1_tx_valid_r_reg/NET0131  ;
  assign n1757 = \u1_u1_state_reg[1]/NET0131  & n1756 ;
  assign n1758 = \u1_u2_adr_cb_reg[1]/NET0131  & ~\u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n1759 = \u1_u2_adr_cb_reg[0]/NET0131  & \u1_u2_adr_cb_reg[2]/NET0131  ;
  assign n1760 = n1758 & n1759 ;
  assign n1761 = ~n1757 & n1760 ;
  assign n1762 = \u1_u2_rd_buf1_reg[27]/NET0131  & n1761 ;
  assign n1763 = ~\u1_u2_rx_data_valid_r_reg/NET0131  & ~n1757 ;
  assign n1764 = ~\u1_u2_adr_cb_reg[0]/NET0131  & \u1_u2_adr_cb_reg[2]/NET0131  ;
  assign n1765 = \u1_u2_adr_cb_reg[1]/NET0131  & n1764 ;
  assign n1766 = \u1_u2_rd_buf1_reg[27]/NET0131  & n1765 ;
  assign n1767 = ~n1763 & n1766 ;
  assign n1768 = ~n1762 & ~n1767 ;
  assign n1769 = ~\u1_u2_adr_cb_reg[1]/NET0131  & ~\u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n1770 = n1759 & n1769 ;
  assign n1771 = ~n1757 & n1770 ;
  assign n1772 = \u1_u2_rd_buf1_reg[11]/NET0131  & n1771 ;
  assign n1773 = ~\u1_u2_adr_cb_reg[1]/NET0131  & n1764 ;
  assign n1774 = \u1_u2_rd_buf1_reg[11]/NET0131  & n1773 ;
  assign n1775 = ~n1763 & n1774 ;
  assign n1776 = ~n1772 & ~n1775 ;
  assign n1777 = n1768 & n1776 ;
  assign n1778 = n1764 & n1769 ;
  assign n1779 = ~n1757 & n1778 ;
  assign n1780 = \u1_u2_rd_buf1_reg[3]/NET0131  & n1779 ;
  assign n1781 = \u1_u2_adr_cb_reg[0]/NET0131  & ~\u1_u2_adr_cb_reg[2]/NET0131  ;
  assign n1782 = \u1_u2_adr_cb_reg[1]/NET0131  & n1781 ;
  assign n1783 = \u1_u2_rd_buf1_reg[3]/NET0131  & n1782 ;
  assign n1784 = ~n1763 & n1783 ;
  assign n1785 = ~n1780 & ~n1784 ;
  assign n1786 = n1758 & n1764 ;
  assign n1787 = ~n1757 & n1786 ;
  assign n1788 = \u1_u2_rd_buf1_reg[19]/NET0131  & n1787 ;
  assign n1789 = ~\u1_u2_adr_cb_reg[1]/NET0131  & n1759 ;
  assign n1790 = \u1_u2_rd_buf1_reg[19]/NET0131  & n1789 ;
  assign n1791 = ~n1763 & n1790 ;
  assign n1792 = ~n1788 & ~n1791 ;
  assign n1793 = n1785 & n1792 ;
  assign n1794 = n1777 & n1793 ;
  assign n1795 = n1758 & n1781 ;
  assign n1796 = ~n1757 & n1795 ;
  assign n1797 = \u1_u2_rd_buf0_reg[27]/NET0131  & n1796 ;
  assign n1798 = ~\u1_u2_adr_cb_reg[0]/NET0131  & ~\u1_u2_adr_cb_reg[2]/NET0131  ;
  assign n1799 = \u1_u2_adr_cb_reg[1]/NET0131  & n1798 ;
  assign n1800 = \u1_u2_rd_buf0_reg[27]/NET0131  & n1799 ;
  assign n1801 = ~n1763 & n1800 ;
  assign n1802 = ~n1797 & ~n1801 ;
  assign n1803 = n1769 & n1781 ;
  assign n1804 = ~n1757 & n1803 ;
  assign n1805 = \u1_u2_rd_buf0_reg[11]/NET0131  & n1804 ;
  assign n1806 = ~\u1_u2_adr_cb_reg[1]/NET0131  & n1798 ;
  assign n1807 = \u1_u2_rd_buf0_reg[11]/NET0131  & n1806 ;
  assign n1808 = ~n1763 & n1807 ;
  assign n1809 = ~n1805 & ~n1808 ;
  assign n1810 = n1802 & n1809 ;
  assign n1811 = n1758 & n1798 ;
  assign n1812 = ~n1757 & n1811 ;
  assign n1813 = \u1_u2_rd_buf0_reg[19]/NET0131  & n1812 ;
  assign n1814 = ~\u1_u2_adr_cb_reg[1]/NET0131  & n1781 ;
  assign n1815 = \u1_u2_rd_buf0_reg[19]/NET0131  & n1814 ;
  assign n1816 = ~n1763 & n1815 ;
  assign n1817 = ~n1813 & ~n1816 ;
  assign n1818 = n1769 & n1798 ;
  assign n1819 = ~n1757 & n1818 ;
  assign n1820 = \u1_u2_rd_buf0_reg[3]/NET0131  & n1819 ;
  assign n1821 = \u1_u2_adr_cb_reg[1]/NET0131  & n1759 ;
  assign n1822 = \u1_u2_rd_buf0_reg[3]/NET0131  & n1821 ;
  assign n1823 = ~n1763 & n1822 ;
  assign n1824 = ~n1820 & ~n1823 ;
  assign n1825 = n1817 & n1824 ;
  assign n1826 = n1810 & n1825 ;
  assign n1827 = n1794 & n1826 ;
  assign n1828 = n1750 & n1756 ;
  assign n1829 = ~\u1_u1_state_reg[2]/NET0131  & ~\u1_u1_state_reg[4]/NET0131  ;
  assign n1830 = ~\u1_u1_state_reg[3]/NET0131  & n1829 ;
  assign n1831 = ~\u1_u1_state_reg[0]/NET0131  & \u1_u1_state_reg[1]/NET0131  ;
  assign n1832 = n1830 & n1831 ;
  assign n1833 = n1828 & n1832 ;
  assign n1834 = ~\u1_u1_state_reg[0]/NET0131  & ~\u1_u1_state_reg[1]/NET0131  ;
  assign n1835 = ~\u1_u1_state_reg[3]/NET0131  & n1834 ;
  assign n1836 = ~\u1_u1_state_reg[2]/NET0131  & \u1_u1_state_reg[4]/NET0131  ;
  assign n1837 = n1835 & n1836 ;
  assign n1838 = \u1_u1_state_reg[3]/NET0131  & n1829 ;
  assign n1839 = n1834 & n1838 ;
  assign n1840 = ~n1837 & ~n1839 ;
  assign n1841 = ~n1833 & n1840 ;
  assign n1842 = ~\u1_u1_send_token_r_reg/P0001  & ~\u1_u3_send_token_reg/P0001  ;
  assign n1843 = \u1_u3_token_pid_sel_reg[0]/P0001  & ~\u1_u3_token_pid_sel_reg[1]/P0001  ;
  assign n1844 = ~\u1_u3_token_pid_sel_reg[0]/P0001  & \u1_u3_token_pid_sel_reg[1]/P0001  ;
  assign n1845 = ~n1843 & ~n1844 ;
  assign n1846 = ~n1842 & ~n1845 ;
  assign n1847 = \u1_u1_state_reg[0]/NET0131  & ~\u1_u1_state_reg[1]/NET0131  ;
  assign n1848 = ~n1750 & n1847 ;
  assign n1849 = n1830 & n1848 ;
  assign n1850 = \u1_u1_state_reg[2]/NET0131  & ~\u1_u1_state_reg[4]/NET0131  ;
  assign n1851 = n1835 & n1850 ;
  assign n1852 = ~n1849 & ~n1851 ;
  assign n1853 = ~n1846 & n1852 ;
  assign n1854 = n1841 & n1853 ;
  assign n1855 = n1827 & n1854 ;
  assign n1856 = ~n1842 & ~n1846 ;
  assign n1857 = ~\u0_tx_ready_reg/NET0131  & n1850 ;
  assign n1858 = n1835 & n1857 ;
  assign n1859 = ~n1837 & ~n1858 ;
  assign n1860 = ~n1833 & n1859 ;
  assign n1861 = ~\u1_u1_crc16_reg[12]/P0001  & ~n1860 ;
  assign n1862 = \u0_tx_ready_reg/NET0131  & \u1_u1_state_reg[2]/NET0131  ;
  assign n1863 = ~\u1_u3_this_dpid_reg[0]/P0001  & ~n1862 ;
  assign n1864 = ~n1839 & n1863 ;
  assign n1865 = \u1_u1_crc16_reg[4]/P0001  & n1862 ;
  assign n1866 = \u1_u1_crc16_reg[4]/P0001  & n1834 ;
  assign n1867 = n1838 & n1866 ;
  assign n1868 = ~n1865 & ~n1867 ;
  assign n1869 = ~n1864 & n1868 ;
  assign n1870 = n1860 & n1869 ;
  assign n1871 = ~n1861 & ~n1870 ;
  assign n1872 = n1841 & n1852 ;
  assign n1873 = ~n1846 & ~n1872 ;
  assign n1874 = n1871 & n1873 ;
  assign n1875 = ~n1856 & ~n1874 ;
  assign n1876 = n1753 & n1875 ;
  assign n1877 = ~n1855 & n1876 ;
  assign n1878 = ~n1755 & ~n1877 ;
  assign n1879 = \u1_u1_crc16_reg[8]/P0001  & ~n1860 ;
  assign n1880 = ~\u1_u1_crc16_reg[0]/P0001  & n1862 ;
  assign n1881 = ~\u1_u1_crc16_reg[0]/P0001  & n1834 ;
  assign n1882 = n1838 & n1881 ;
  assign n1883 = ~n1880 & ~n1882 ;
  assign n1884 = ~n1864 & n1883 ;
  assign n1885 = n1860 & n1884 ;
  assign n1886 = ~n1879 & ~n1885 ;
  assign n1887 = n1873 & n1886 ;
  assign n1888 = ~n1856 & ~n1887 ;
  assign n1889 = n1753 & ~n1888 ;
  assign n1890 = \DataOut_pad_o[7]_pad  & ~\u0_u0_drive_k_reg/P0001  ;
  assign n1891 = ~n1753 & n1890 ;
  assign n1892 = \u1_u2_rd_buf0_reg[15]/P0001  & n1804 ;
  assign n1893 = \u1_u2_rd_buf0_reg[15]/P0001  & n1806 ;
  assign n1894 = ~n1763 & n1893 ;
  assign n1895 = ~n1892 & ~n1894 ;
  assign n1896 = \u1_u2_rd_buf0_reg[23]/P0001  & n1812 ;
  assign n1897 = \u1_u2_rd_buf0_reg[23]/P0001  & n1814 ;
  assign n1898 = ~n1763 & n1897 ;
  assign n1899 = ~n1896 & ~n1898 ;
  assign n1900 = n1895 & n1899 ;
  assign n1901 = \u1_u2_rd_buf1_reg[7]/P0001  & n1779 ;
  assign n1902 = \u1_u2_rd_buf1_reg[7]/P0001  & n1782 ;
  assign n1903 = ~n1763 & n1902 ;
  assign n1904 = ~n1901 & ~n1903 ;
  assign n1905 = \u1_u2_rd_buf1_reg[15]/P0001  & n1771 ;
  assign n1906 = \u1_u2_rd_buf1_reg[15]/P0001  & n1773 ;
  assign n1907 = ~n1763 & n1906 ;
  assign n1908 = ~n1905 & ~n1907 ;
  assign n1909 = n1904 & n1908 ;
  assign n1910 = n1900 & n1909 ;
  assign n1911 = \u1_u2_rd_buf1_reg[23]/P0001  & n1787 ;
  assign n1912 = \u1_u2_rd_buf1_reg[23]/P0001  & n1789 ;
  assign n1913 = ~n1763 & n1912 ;
  assign n1914 = ~n1911 & ~n1913 ;
  assign n1915 = \u1_u2_rd_buf1_reg[31]/P0001  & n1761 ;
  assign n1916 = \u1_u2_rd_buf1_reg[31]/P0001  & n1765 ;
  assign n1917 = ~n1763 & n1916 ;
  assign n1918 = ~n1915 & ~n1917 ;
  assign n1919 = n1914 & n1918 ;
  assign n1920 = \u1_u2_rd_buf0_reg[7]/P0001  & n1819 ;
  assign n1921 = \u1_u2_rd_buf0_reg[7]/P0001  & n1821 ;
  assign n1922 = ~n1763 & n1921 ;
  assign n1923 = ~n1920 & ~n1922 ;
  assign n1924 = \u1_u2_rd_buf0_reg[31]/P0001  & n1796 ;
  assign n1925 = \u1_u2_rd_buf0_reg[31]/P0001  & n1799 ;
  assign n1926 = ~n1763 & n1925 ;
  assign n1927 = ~n1924 & ~n1926 ;
  assign n1928 = n1923 & n1927 ;
  assign n1929 = n1919 & n1928 ;
  assign n1930 = n1910 & n1929 ;
  assign n1931 = n1753 & ~n1846 ;
  assign n1932 = n1852 & n1931 ;
  assign n1933 = n1841 & n1932 ;
  assign n1934 = ~n1930 & n1933 ;
  assign n1935 = ~n1891 & ~n1934 ;
  assign n1936 = ~n1889 & n1935 ;
  assign n1937 = \DataOut_pad_o[2]_pad  & ~\u0_u0_drive_k_reg/P0001  ;
  assign n1938 = ~n1753 & n1937 ;
  assign n1939 = \u1_u2_rd_buf0_reg[2]/NET0131  & n1819 ;
  assign n1940 = \u1_u2_rd_buf0_reg[2]/NET0131  & n1821 ;
  assign n1941 = ~n1763 & n1940 ;
  assign n1942 = ~n1939 & ~n1941 ;
  assign n1943 = \u1_u2_rd_buf1_reg[18]/NET0131  & n1787 ;
  assign n1944 = \u1_u2_rd_buf1_reg[18]/NET0131  & n1789 ;
  assign n1945 = ~n1763 & n1944 ;
  assign n1946 = ~n1943 & ~n1945 ;
  assign n1947 = n1942 & n1946 ;
  assign n1948 = \u1_u2_rd_buf0_reg[18]/NET0131  & n1812 ;
  assign n1949 = \u1_u2_rd_buf0_reg[18]/NET0131  & n1814 ;
  assign n1950 = ~n1763 & n1949 ;
  assign n1951 = ~n1948 & ~n1950 ;
  assign n1952 = \u1_u2_rd_buf1_reg[2]/NET0131  & n1779 ;
  assign n1953 = \u1_u2_rd_buf1_reg[2]/NET0131  & n1782 ;
  assign n1954 = ~n1763 & n1953 ;
  assign n1955 = ~n1952 & ~n1954 ;
  assign n1956 = n1951 & n1955 ;
  assign n1957 = n1947 & n1956 ;
  assign n1958 = \u1_u2_rd_buf0_reg[10]/NET0131  & n1804 ;
  assign n1959 = \u1_u2_rd_buf0_reg[10]/NET0131  & n1806 ;
  assign n1960 = ~n1763 & n1959 ;
  assign n1961 = ~n1958 & ~n1960 ;
  assign n1962 = \u1_u2_rd_buf0_reg[26]/NET0131  & n1796 ;
  assign n1963 = \u1_u2_rd_buf0_reg[26]/NET0131  & n1799 ;
  assign n1964 = ~n1763 & n1963 ;
  assign n1965 = ~n1962 & ~n1964 ;
  assign n1966 = n1961 & n1965 ;
  assign n1967 = \u1_u2_rd_buf1_reg[26]/NET0131  & n1761 ;
  assign n1968 = \u1_u2_rd_buf1_reg[26]/NET0131  & n1765 ;
  assign n1969 = ~n1763 & n1968 ;
  assign n1970 = ~n1967 & ~n1969 ;
  assign n1971 = \u1_u2_rd_buf1_reg[10]/NET0131  & n1771 ;
  assign n1972 = \u1_u2_rd_buf1_reg[10]/NET0131  & n1773 ;
  assign n1973 = ~n1763 & n1972 ;
  assign n1974 = ~n1971 & ~n1973 ;
  assign n1975 = n1970 & n1974 ;
  assign n1976 = n1966 & n1975 ;
  assign n1977 = n1957 & n1976 ;
  assign n1978 = \u1_u3_token_pid_sel_reg[1]/P0001  & ~n1842 ;
  assign n1979 = n1852 & ~n1978 ;
  assign n1980 = n1841 & n1979 ;
  assign n1981 = n1977 & n1980 ;
  assign n1982 = ~n1842 & ~n1978 ;
  assign n1983 = ~\u1_u1_crc16_reg[13]/P0001  & ~n1860 ;
  assign n1984 = \u1_u1_crc16_reg[5]/P0001  & n1862 ;
  assign n1985 = \u1_u1_crc16_reg[5]/P0001  & n1834 ;
  assign n1986 = n1838 & n1985 ;
  assign n1987 = ~n1984 & ~n1986 ;
  assign n1988 = ~\u1_u3_this_dpid_reg[1]/P0001  & ~n1862 ;
  assign n1989 = ~n1839 & n1988 ;
  assign n1990 = n1987 & ~n1989 ;
  assign n1991 = n1860 & n1990 ;
  assign n1992 = ~n1983 & ~n1991 ;
  assign n1993 = ~n1872 & ~n1978 ;
  assign n1994 = n1992 & n1993 ;
  assign n1995 = ~n1982 & ~n1994 ;
  assign n1996 = n1753 & n1995 ;
  assign n1997 = ~n1981 & n1996 ;
  assign n1998 = ~n1938 & ~n1997 ;
  assign n1999 = \u1_u1_crc16_reg[9]/P0001  & ~n1860 ;
  assign n2000 = ~\u1_u1_crc16_reg[1]/P0001  & n1862 ;
  assign n2001 = ~\u1_u1_crc16_reg[1]/P0001  & n1834 ;
  assign n2002 = n1838 & n2001 ;
  assign n2003 = ~n2000 & ~n2002 ;
  assign n2004 = ~n1989 & n2003 ;
  assign n2005 = n1860 & n2004 ;
  assign n2006 = ~n1999 & ~n2005 ;
  assign n2007 = n1993 & n2006 ;
  assign n2008 = ~n1982 & ~n2007 ;
  assign n2009 = n1753 & ~n2008 ;
  assign n2010 = \DataOut_pad_o[6]_pad  & ~\u0_u0_drive_k_reg/P0001  ;
  assign n2011 = ~n1753 & n2010 ;
  assign n2012 = \u1_u2_rd_buf1_reg[6]/P0001  & n1779 ;
  assign n2013 = \u1_u2_rd_buf1_reg[6]/P0001  & n1782 ;
  assign n2014 = ~n1763 & n2013 ;
  assign n2015 = ~n2012 & ~n2014 ;
  assign n2016 = \u1_u2_rd_buf1_reg[14]/P0001  & n1771 ;
  assign n2017 = \u1_u2_rd_buf1_reg[14]/P0001  & n1773 ;
  assign n2018 = ~n1763 & n2017 ;
  assign n2019 = ~n2016 & ~n2018 ;
  assign n2020 = n2015 & n2019 ;
  assign n2021 = \u1_u2_rd_buf0_reg[14]/P0001  & n1804 ;
  assign n2022 = \u1_u2_rd_buf0_reg[14]/P0001  & n1806 ;
  assign n2023 = ~n1763 & n2022 ;
  assign n2024 = ~n2021 & ~n2023 ;
  assign n2025 = \u1_u2_rd_buf1_reg[22]/P0001  & n1787 ;
  assign n2026 = \u1_u2_rd_buf1_reg[22]/P0001  & n1789 ;
  assign n2027 = ~n1763 & n2026 ;
  assign n2028 = ~n2025 & ~n2027 ;
  assign n2029 = n2024 & n2028 ;
  assign n2030 = n2020 & n2029 ;
  assign n2031 = \u1_u2_rd_buf1_reg[30]/P0001  & n1761 ;
  assign n2032 = \u1_u2_rd_buf1_reg[30]/P0001  & n1765 ;
  assign n2033 = ~n1763 & n2032 ;
  assign n2034 = ~n2031 & ~n2033 ;
  assign n2035 = \u1_u2_rd_buf0_reg[30]/P0001  & n1796 ;
  assign n2036 = \u1_u2_rd_buf0_reg[30]/P0001  & n1799 ;
  assign n2037 = ~n1763 & n2036 ;
  assign n2038 = ~n2035 & ~n2037 ;
  assign n2039 = n2034 & n2038 ;
  assign n2040 = \u1_u2_rd_buf0_reg[6]/P0001  & n1819 ;
  assign n2041 = \u1_u2_rd_buf0_reg[6]/P0001  & n1821 ;
  assign n2042 = ~n1763 & n2041 ;
  assign n2043 = ~n2040 & ~n2042 ;
  assign n2044 = \u1_u2_rd_buf0_reg[22]/P0001  & n1812 ;
  assign n2045 = \u1_u2_rd_buf0_reg[22]/P0001  & n1814 ;
  assign n2046 = ~n1763 & n2045 ;
  assign n2047 = ~n2044 & ~n2046 ;
  assign n2048 = n2043 & n2047 ;
  assign n2049 = n2039 & n2048 ;
  assign n2050 = n2030 & n2049 ;
  assign n2051 = n1753 & ~n1978 ;
  assign n2052 = n1852 & n2051 ;
  assign n2053 = n1841 & n2052 ;
  assign n2054 = ~n2050 & n2053 ;
  assign n2055 = ~n2011 & ~n2054 ;
  assign n2056 = ~n2009 & n2055 ;
  assign n2057 = \u1_u2_rd_buf0_reg[4]/P0001  & n1819 ;
  assign n2058 = \u1_u2_rd_buf0_reg[4]/P0001  & n1821 ;
  assign n2059 = ~n1763 & n2058 ;
  assign n2060 = ~n2057 & ~n2059 ;
  assign n2061 = \u1_u2_rd_buf0_reg[12]/P0001  & n1804 ;
  assign n2062 = \u1_u2_rd_buf0_reg[12]/P0001  & n1806 ;
  assign n2063 = ~n1763 & n2062 ;
  assign n2064 = ~n2061 & ~n2063 ;
  assign n2065 = n2060 & n2064 ;
  assign n2066 = \u1_u2_rd_buf1_reg[20]/P0001  & n1787 ;
  assign n2067 = \u1_u2_rd_buf1_reg[20]/P0001  & n1789 ;
  assign n2068 = ~n1763 & n2067 ;
  assign n2069 = ~n2066 & ~n2068 ;
  assign n2070 = \u1_u2_rd_buf1_reg[28]/P0001  & n1761 ;
  assign n2071 = \u1_u2_rd_buf1_reg[28]/P0001  & n1765 ;
  assign n2072 = ~n1763 & n2071 ;
  assign n2073 = ~n2070 & ~n2072 ;
  assign n2074 = n2069 & n2073 ;
  assign n2075 = n2065 & n2074 ;
  assign n2076 = \u1_u2_rd_buf0_reg[20]/P0001  & n1812 ;
  assign n2077 = \u1_u2_rd_buf0_reg[20]/P0001  & n1814 ;
  assign n2078 = ~n1763 & n2077 ;
  assign n2079 = ~n2076 & ~n2078 ;
  assign n2080 = \u1_u2_rd_buf0_reg[28]/P0001  & n1796 ;
  assign n2081 = \u1_u2_rd_buf0_reg[28]/P0001  & n1799 ;
  assign n2082 = ~n1763 & n2081 ;
  assign n2083 = ~n2080 & ~n2082 ;
  assign n2084 = n2079 & n2083 ;
  assign n2085 = \u1_u2_rd_buf1_reg[4]/P0001  & n1779 ;
  assign n2086 = \u1_u2_rd_buf1_reg[4]/P0001  & n1782 ;
  assign n2087 = ~n1763 & n2086 ;
  assign n2088 = ~n2085 & ~n2087 ;
  assign n2089 = \u1_u2_rd_buf1_reg[12]/P0001  & n1771 ;
  assign n2090 = \u1_u2_rd_buf1_reg[12]/P0001  & n1773 ;
  assign n2091 = ~n1763 & n2090 ;
  assign n2092 = ~n2089 & ~n2091 ;
  assign n2093 = n2088 & n2092 ;
  assign n2094 = n2084 & n2093 ;
  assign n2095 = n2075 & n2094 ;
  assign n2096 = \u1_u2_rd_buf1_reg[5]/P0001  & n1779 ;
  assign n2097 = \u1_u2_rd_buf1_reg[5]/P0001  & n1782 ;
  assign n2098 = ~n1763 & n2097 ;
  assign n2099 = ~n2096 & ~n2098 ;
  assign n2100 = \u1_u2_rd_buf1_reg[13]/P0001  & n1771 ;
  assign n2101 = \u1_u2_rd_buf1_reg[13]/P0001  & n1773 ;
  assign n2102 = ~n1763 & n2101 ;
  assign n2103 = ~n2100 & ~n2102 ;
  assign n2104 = n2099 & n2103 ;
  assign n2105 = \u1_u2_rd_buf1_reg[21]/P0001  & n1787 ;
  assign n2106 = \u1_u2_rd_buf1_reg[21]/P0001  & n1789 ;
  assign n2107 = ~n1763 & n2106 ;
  assign n2108 = ~n2105 & ~n2107 ;
  assign n2109 = \u1_u2_rd_buf1_reg[29]/P0001  & n1761 ;
  assign n2110 = \u1_u2_rd_buf1_reg[29]/P0001  & n1765 ;
  assign n2111 = ~n1763 & n2110 ;
  assign n2112 = ~n2109 & ~n2111 ;
  assign n2113 = n2108 & n2112 ;
  assign n2114 = n2104 & n2113 ;
  assign n2115 = \u1_u2_rd_buf0_reg[29]/P0001  & n1796 ;
  assign n2116 = \u1_u2_rd_buf0_reg[29]/P0001  & n1799 ;
  assign n2117 = ~n1763 & n2116 ;
  assign n2118 = ~n2115 & ~n2117 ;
  assign n2119 = \u1_u2_rd_buf0_reg[21]/P0001  & n1812 ;
  assign n2120 = \u1_u2_rd_buf0_reg[21]/P0001  & n1814 ;
  assign n2121 = ~n1763 & n2120 ;
  assign n2122 = ~n2119 & ~n2121 ;
  assign n2123 = n2118 & n2122 ;
  assign n2124 = \u1_u2_rd_buf0_reg[13]/P0001  & n1804 ;
  assign n2125 = \u1_u2_rd_buf0_reg[13]/P0001  & n1806 ;
  assign n2126 = ~n1763 & n2125 ;
  assign n2127 = ~n2124 & ~n2126 ;
  assign n2128 = \u1_u2_rd_buf0_reg[5]/P0001  & n1819 ;
  assign n2129 = \u1_u2_rd_buf0_reg[5]/P0001  & n1821 ;
  assign n2130 = ~n1763 & n2129 ;
  assign n2131 = ~n2128 & ~n2130 ;
  assign n2132 = n2127 & n2131 ;
  assign n2133 = n2123 & n2132 ;
  assign n2134 = n2114 & n2133 ;
  assign n2135 = ~n2095 & ~n2134 ;
  assign n2136 = n2095 & n2134 ;
  assign n2137 = ~n2135 & ~n2136 ;
  assign n2138 = ~n1930 & ~n2050 ;
  assign n2139 = n1930 & n2050 ;
  assign n2140 = ~n2138 & ~n2139 ;
  assign n2141 = ~n2137 & ~n2140 ;
  assign n2142 = n2137 & n2140 ;
  assign n2143 = ~n2141 & ~n2142 ;
  assign n2144 = \u1_u1_crc16_reg[7]/P0001  & ~\u1_u1_crc16_reg[8]/P0001  ;
  assign n2145 = ~\u1_u1_crc16_reg[7]/P0001  & \u1_u1_crc16_reg[8]/P0001  ;
  assign n2146 = ~n2144 & ~n2145 ;
  assign n2147 = n1827 & ~n1977 ;
  assign n2148 = ~n1827 & n1977 ;
  assign n2149 = ~n2147 & ~n2148 ;
  assign n2150 = n2146 & ~n2149 ;
  assign n2151 = ~n2143 & n2150 ;
  assign n2152 = n2146 & n2149 ;
  assign n2153 = n2143 & n2152 ;
  assign n2154 = ~n2151 & ~n2153 ;
  assign n2155 = ~n2146 & ~n2149 ;
  assign n2156 = n2143 & n2155 ;
  assign n2157 = ~n2146 & n2149 ;
  assign n2158 = ~n2143 & n2157 ;
  assign n2159 = ~n2156 & ~n2158 ;
  assign n2160 = n2154 & n2159 ;
  assign n2161 = ~\u1_u1_crc16_reg[13]/P0001  & ~\u1_u1_crc16_reg[14]/P0001  ;
  assign n2162 = \u1_u1_crc16_reg[13]/P0001  & \u1_u1_crc16_reg[14]/P0001  ;
  assign n2163 = ~n2161 & ~n2162 ;
  assign n2164 = \u1_u2_rd_buf0_reg[16]/NET0131  & n1812 ;
  assign n2165 = \u1_u2_rd_buf0_reg[16]/NET0131  & n1814 ;
  assign n2166 = ~n1763 & n2165 ;
  assign n2167 = ~n2164 & ~n2166 ;
  assign n2168 = \u1_u2_rd_buf1_reg[8]/NET0131  & n1771 ;
  assign n2169 = \u1_u2_rd_buf1_reg[8]/NET0131  & n1773 ;
  assign n2170 = ~n1763 & n2169 ;
  assign n2171 = ~n2168 & ~n2170 ;
  assign n2172 = n2167 & n2171 ;
  assign n2173 = \u1_u2_rd_buf1_reg[0]/NET0131  & n1779 ;
  assign n2174 = \u1_u2_rd_buf1_reg[0]/NET0131  & n1782 ;
  assign n2175 = ~n1763 & n2174 ;
  assign n2176 = ~n2173 & ~n2175 ;
  assign n2177 = \u1_u2_rd_buf0_reg[24]/NET0131  & n1796 ;
  assign n2178 = \u1_u2_rd_buf0_reg[24]/NET0131  & n1799 ;
  assign n2179 = ~n1763 & n2178 ;
  assign n2180 = ~n2177 & ~n2179 ;
  assign n2181 = n2176 & n2180 ;
  assign n2182 = n2172 & n2181 ;
  assign n2183 = \u1_u2_rd_buf0_reg[8]/NET0131  & n1804 ;
  assign n2184 = \u1_u2_rd_buf0_reg[8]/NET0131  & n1806 ;
  assign n2185 = ~n1763 & n2184 ;
  assign n2186 = ~n2183 & ~n2185 ;
  assign n2187 = \u1_u2_rd_buf1_reg[24]/NET0131  & n1761 ;
  assign n2188 = \u1_u2_rd_buf1_reg[24]/NET0131  & n1765 ;
  assign n2189 = ~n1763 & n2188 ;
  assign n2190 = ~n2187 & ~n2189 ;
  assign n2191 = n2186 & n2190 ;
  assign n2192 = \u1_u2_rd_buf0_reg[0]/NET0131  & n1819 ;
  assign n2193 = \u1_u2_rd_buf0_reg[0]/NET0131  & n1821 ;
  assign n2194 = ~n1763 & n2193 ;
  assign n2195 = ~n2192 & ~n2194 ;
  assign n2196 = \u1_u2_rd_buf1_reg[16]/NET0131  & n1787 ;
  assign n2197 = \u1_u2_rd_buf1_reg[16]/NET0131  & n1789 ;
  assign n2198 = ~n1763 & n2197 ;
  assign n2199 = ~n2196 & ~n2198 ;
  assign n2200 = n2195 & n2199 ;
  assign n2201 = n2191 & n2200 ;
  assign n2202 = n2182 & n2201 ;
  assign n2203 = \u1_u1_crc16_reg[15]/P0001  & ~n2202 ;
  assign n2204 = ~\u1_u1_crc16_reg[15]/P0001  & n2202 ;
  assign n2205 = ~n2203 & ~n2204 ;
  assign n2206 = \u1_u2_rd_buf1_reg[25]/NET0131  & n1765 ;
  assign n2207 = ~n1763 & n2206 ;
  assign n2208 = \u1_u2_rd_buf1_reg[25]/NET0131  & n1761 ;
  assign n2209 = ~n2207 & ~n2208 ;
  assign n2210 = \u1_u2_rd_buf1_reg[9]/NET0131  & n1771 ;
  assign n2211 = \u1_u2_rd_buf1_reg[9]/NET0131  & n1773 ;
  assign n2212 = ~n1763 & n2211 ;
  assign n2213 = ~n2210 & ~n2212 ;
  assign n2214 = n2209 & n2213 ;
  assign n2215 = \u1_u2_rd_buf1_reg[17]/NET0131  & n1787 ;
  assign n2216 = \u1_u2_rd_buf1_reg[17]/NET0131  & n1789 ;
  assign n2217 = ~n1763 & n2216 ;
  assign n2218 = ~n2215 & ~n2217 ;
  assign n2219 = \u1_u2_rd_buf1_reg[1]/NET0131  & n1779 ;
  assign n2220 = \u1_u2_rd_buf1_reg[1]/NET0131  & n1782 ;
  assign n2221 = ~n1763 & n2220 ;
  assign n2222 = ~n2219 & ~n2221 ;
  assign n2223 = n2218 & n2222 ;
  assign n2224 = n2214 & n2223 ;
  assign n2225 = \u1_u2_rd_buf0_reg[9]/NET0131  & n1804 ;
  assign n2226 = \u1_u2_rd_buf0_reg[9]/NET0131  & n1806 ;
  assign n2227 = ~n1763 & n2226 ;
  assign n2228 = ~n2225 & ~n2227 ;
  assign n2229 = \u1_u2_rd_buf0_reg[25]/NET0131  & n1796 ;
  assign n2230 = \u1_u2_rd_buf0_reg[25]/NET0131  & n1799 ;
  assign n2231 = ~n1763 & n2230 ;
  assign n2232 = ~n2229 & ~n2231 ;
  assign n2233 = n2228 & n2232 ;
  assign n2234 = \u1_u2_rd_buf0_reg[17]/NET0131  & n1812 ;
  assign n2235 = \u1_u2_rd_buf0_reg[17]/NET0131  & n1814 ;
  assign n2236 = ~n1763 & n2235 ;
  assign n2237 = ~n2234 & ~n2236 ;
  assign n2238 = \u1_u2_rd_buf0_reg[1]/NET0131  & n1819 ;
  assign n2239 = \u1_u2_rd_buf0_reg[1]/NET0131  & n1821 ;
  assign n2240 = ~n1763 & n2239 ;
  assign n2241 = ~n2238 & ~n2240 ;
  assign n2242 = n2237 & n2241 ;
  assign n2243 = n2233 & n2242 ;
  assign n2244 = n2224 & n2243 ;
  assign n2245 = \u1_u1_crc16_reg[10]/P0001  & ~\u1_u1_crc16_reg[9]/P0001  ;
  assign n2246 = ~\u1_u1_crc16_reg[10]/P0001  & \u1_u1_crc16_reg[9]/P0001  ;
  assign n2247 = ~n2245 & ~n2246 ;
  assign n2248 = \u1_u1_crc16_reg[11]/P0001  & ~\u1_u1_crc16_reg[12]/P0001  ;
  assign n2249 = ~\u1_u1_crc16_reg[11]/P0001  & \u1_u1_crc16_reg[12]/P0001  ;
  assign n2250 = ~n2248 & ~n2249 ;
  assign n2251 = ~n2247 & n2250 ;
  assign n2252 = ~n2244 & n2251 ;
  assign n2253 = ~n2205 & n2252 ;
  assign n2254 = n2244 & n2251 ;
  assign n2255 = n2205 & n2254 ;
  assign n2256 = ~n2253 & ~n2255 ;
  assign n2257 = n2247 & n2250 ;
  assign n2258 = ~n2244 & n2257 ;
  assign n2259 = n2205 & n2258 ;
  assign n2260 = n2244 & n2257 ;
  assign n2261 = ~n2205 & n2260 ;
  assign n2262 = ~n2259 & ~n2261 ;
  assign n2263 = n2256 & n2262 ;
  assign n2264 = ~n2247 & ~n2250 ;
  assign n2265 = ~n2244 & n2264 ;
  assign n2266 = n2205 & n2265 ;
  assign n2267 = n2244 & n2264 ;
  assign n2268 = ~n2205 & n2267 ;
  assign n2269 = ~n2266 & ~n2268 ;
  assign n2270 = n2247 & ~n2250 ;
  assign n2271 = ~n2244 & n2270 ;
  assign n2272 = ~n2205 & n2271 ;
  assign n2273 = n2244 & n2270 ;
  assign n2274 = n2205 & n2273 ;
  assign n2275 = ~n2272 & ~n2274 ;
  assign n2276 = n2269 & n2275 ;
  assign n2277 = n2263 & n2276 ;
  assign n2278 = ~n2163 & ~n2277 ;
  assign n2279 = n2163 & n2277 ;
  assign n2280 = ~n2278 & ~n2279 ;
  assign n2281 = ~n2160 & n2280 ;
  assign n2282 = n1757 & n1860 ;
  assign n2283 = ~\u1_u1_send_data_r2_reg/P0001  & \u1_u1_send_data_r_reg/P0001  ;
  assign n2284 = ~\u1_u1_zero_length_r_reg/P0001  & n2283 ;
  assign n2285 = ~n2282 & ~n2284 ;
  assign n2286 = ~n2160 & ~n2285 ;
  assign n2287 = n2163 & ~n2285 ;
  assign n2288 = ~n2277 & n2287 ;
  assign n2289 = ~n2163 & ~n2285 ;
  assign n2290 = n2277 & n2289 ;
  assign n2291 = ~n2288 & ~n2290 ;
  assign n2292 = ~n2286 & n2291 ;
  assign n2293 = ~n2281 & ~n2292 ;
  assign n2294 = ~\u1_u1_send_data_r_reg/P0001  & ~n1750 ;
  assign n2295 = \u1_u1_crc16_reg[15]/P0001  & ~n2284 ;
  assign n2296 = ~n2282 & n2295 ;
  assign n2297 = ~n2294 & ~n2296 ;
  assign n2298 = ~n2293 & n2297 ;
  assign n2299 = n2202 & ~n2244 ;
  assign n2300 = ~n2149 & n2299 ;
  assign n2301 = n2202 & n2244 ;
  assign n2302 = n2149 & n2301 ;
  assign n2303 = ~n2300 & ~n2302 ;
  assign n2304 = ~n2202 & n2244 ;
  assign n2305 = ~n2149 & n2304 ;
  assign n2306 = ~n2202 & ~n2244 ;
  assign n2307 = n2149 & n2306 ;
  assign n2308 = ~n2305 & ~n2307 ;
  assign n2309 = n2303 & n2308 ;
  assign n2310 = \u1_u1_crc16_reg[10]/P0001  & ~\u1_u1_crc16_reg[11]/P0001  ;
  assign n2311 = ~\u1_u1_crc16_reg[10]/P0001  & \u1_u1_crc16_reg[11]/P0001  ;
  assign n2312 = ~n2310 & ~n2311 ;
  assign n2313 = \u1_u1_crc16_reg[9]/P0001  & ~n2312 ;
  assign n2314 = ~\u1_u1_crc16_reg[9]/P0001  & n2312 ;
  assign n2315 = ~n2313 & ~n2314 ;
  assign n2316 = n2095 & n2315 ;
  assign n2317 = ~n2095 & ~n2315 ;
  assign n2318 = ~n2316 & ~n2317 ;
  assign n2319 = n2050 & ~n2134 ;
  assign n2320 = ~n2050 & n2134 ;
  assign n2321 = ~n2319 & ~n2320 ;
  assign n2322 = \u1_u1_crc16_reg[12]/P0001  & ~\u1_u1_crc16_reg[13]/P0001  ;
  assign n2323 = ~\u1_u1_crc16_reg[12]/P0001  & \u1_u1_crc16_reg[13]/P0001  ;
  assign n2324 = ~n2322 & ~n2323 ;
  assign n2325 = \u1_u1_crc16_reg[14]/P0001  & ~\u1_u1_crc16_reg[15]/P0001  ;
  assign n2326 = ~\u1_u1_crc16_reg[14]/P0001  & \u1_u1_crc16_reg[15]/P0001  ;
  assign n2327 = ~n2325 & ~n2326 ;
  assign n2328 = n2324 & n2327 ;
  assign n2329 = ~n2324 & ~n2327 ;
  assign n2330 = ~n2328 & ~n2329 ;
  assign n2331 = n2321 & ~n2330 ;
  assign n2332 = ~n2321 & n2330 ;
  assign n2333 = ~n2331 & ~n2332 ;
  assign n2334 = ~n2318 & ~n2333 ;
  assign n2335 = n2309 & n2334 ;
  assign n2336 = ~n2318 & n2333 ;
  assign n2337 = ~n2309 & n2336 ;
  assign n2338 = ~n2335 & ~n2337 ;
  assign n2339 = n2318 & ~n2333 ;
  assign n2340 = ~n2309 & n2339 ;
  assign n2341 = n2318 & n2333 ;
  assign n2342 = n2309 & n2341 ;
  assign n2343 = ~n2340 & ~n2342 ;
  assign n2344 = ~n2285 & n2343 ;
  assign n2345 = n2338 & n2344 ;
  assign n2346 = \u1_u1_crc16_reg[1]/P0001  & ~n2284 ;
  assign n2347 = ~n2282 & n2346 ;
  assign n2348 = ~n2294 & ~n2347 ;
  assign n2349 = ~n2345 & n2348 ;
  assign n2350 = \u1_u0_pid_reg[0]/NET0131  & ~\u1_u0_pid_reg[1]/NET0131  ;
  assign n2351 = ~\u1_u0_pid_reg[2]/NET0131  & \u1_u0_pid_reg[3]/NET0131  ;
  assign n2352 = n2350 & n2351 ;
  assign n2353 = \u1_u3_buf1_na_reg/NET0131  & n2352 ;
  assign n2354 = ~\u1_u0_pid_reg[2]/NET0131  & ~\u1_u0_pid_reg[3]/NET0131  ;
  assign n2355 = n2350 & n2354 ;
  assign n2356 = \u1_u3_buf0_na_reg/NET0131  & n2355 ;
  assign n2357 = ~n2353 & ~n2356 ;
  assign n2358 = ~\u4_csr_reg[26]/NET0131  & ~\u4_csr_reg[27]/NET0131  ;
  assign n2359 = ~n2357 & n2358 ;
  assign n2360 = \u1_u3_buf0_na_reg/NET0131  & \u1_u3_buf1_na_reg/NET0131  ;
  assign n2361 = \u4_csr_reg[26]/NET0131  & ~\u4_csr_reg[27]/NET0131  ;
  assign n2362 = ~\u4_dma_in_buf_sz1_reg/P0001  & n2361 ;
  assign n2363 = ~\u4_csr_reg[26]/NET0131  & \u4_csr_reg[27]/NET0131  ;
  assign n2364 = ~\u4_dma_out_buf_avail_reg/P0001  & n2363 ;
  assign n2365 = ~n2362 & ~n2364 ;
  assign n2366 = \u4_csr_reg[15]/NET0131  & ~n2358 ;
  assign n2367 = ~n2365 & n2366 ;
  assign n2368 = ~n2360 & ~n2367 ;
  assign n2369 = ~n2359 & n2368 ;
  assign n2370 = ~\u1_u3_state_reg[7]/P0001  & ~\u1_u3_state_reg[9]/P0001  ;
  assign n2371 = ~\u1_u3_state_reg[6]/P0001  & ~\u1_u3_state_reg[8]/P0001  ;
  assign n2372 = n2370 & n2371 ;
  assign n2373 = ~\u1_u3_state_reg[2]/P0001  & ~\u1_u3_state_reg[3]/P0001  ;
  assign n2374 = ~\u1_u3_state_reg[4]/P0001  & ~\u1_u3_state_reg[5]/P0001  ;
  assign n2375 = n2373 & n2374 ;
  assign n2376 = n2372 & n2375 ;
  assign n2377 = \u1_u3_match_r_reg/P0001  & ~\u1_u3_state_reg[1]/P0001  ;
  assign n2378 = \u1_u0_pid_reg[2]/NET0131  & ~\u1_u0_pid_reg[3]/NET0131  ;
  assign n2379 = n2350 & n2378 ;
  assign n2380 = n2377 & ~n2379 ;
  assign n2381 = n2376 & n2380 ;
  assign n2382 = ~\u4_csr_reg[22]/P0001  & \u4_csr_reg[23]/P0001  ;
  assign n2383 = \u4_csr_reg[22]/P0001  & ~\u4_csr_reg[23]/P0001  ;
  assign n2384 = ~\u1_u3_state_reg[6]/P0001  & ~n2383 ;
  assign n2385 = ~n2382 & n2384 ;
  assign n2386 = n2381 & n2385 ;
  assign n2387 = ~n2369 & n2386 ;
  assign n2388 = ~\u1_u3_to_large_reg/P0001  & ~\u1_u3_to_small_reg/P0001  ;
  assign n2389 = \u1_u3_no_bufs1_reg/P0001  & ~\u1_u3_pid_seq_err_reg/P0001  ;
  assign n2390 = \u0_u0_mode_hs_reg/P0001  & \u1_u3_no_bufs0_reg/P0001  ;
  assign n2391 = n2389 & n2390 ;
  assign n2392 = n2388 & ~n2391 ;
  assign n2393 = ~\u1_u3_abort_reg/P0001  & \u1_u3_state_reg[6]/P0001  ;
  assign n2394 = ~n2392 & n2393 ;
  assign n2395 = ~n2387 & ~n2394 ;
  assign n2396 = \u1_u1_crc16_reg[8]/P0001  & ~\u1_u1_crc16_reg[9]/P0001  ;
  assign n2397 = ~\u1_u1_crc16_reg[8]/P0001  & \u1_u1_crc16_reg[9]/P0001  ;
  assign n2398 = ~n2396 & ~n2397 ;
  assign n2399 = ~n2312 & ~n2398 ;
  assign n2400 = n2312 & n2398 ;
  assign n2401 = ~n2399 & ~n2400 ;
  assign n2402 = n2330 & ~n2401 ;
  assign n2403 = ~n2143 & n2309 ;
  assign n2404 = ~n2402 & ~n2403 ;
  assign n2405 = ~n2330 & n2401 ;
  assign n2406 = n2143 & ~n2309 ;
  assign n2407 = ~n2405 & ~n2406 ;
  assign n2408 = n2404 & n2407 ;
  assign n2409 = ~n2402 & ~n2405 ;
  assign n2410 = n2143 & ~n2409 ;
  assign n2411 = ~n2309 & n2410 ;
  assign n2412 = ~n2143 & ~n2409 ;
  assign n2413 = n2309 & n2412 ;
  assign n2414 = ~n2411 & ~n2413 ;
  assign n2415 = ~n2285 & n2414 ;
  assign n2416 = ~n2408 & n2415 ;
  assign n2417 = \u1_u1_crc16_reg[0]/P0001  & ~n2284 ;
  assign n2418 = ~n2282 & n2417 ;
  assign n2419 = ~n2294 & ~n2418 ;
  assign n2420 = ~n2416 & n2419 ;
  assign n2421 = n2377 & n2382 ;
  assign n2422 = ~n2379 & n2421 ;
  assign n2423 = n2376 & n2422 ;
  assign n2424 = n2388 & n2393 ;
  assign n2425 = n2391 & n2424 ;
  assign n2426 = ~n2423 & ~n2425 ;
  assign n2427 = \u1_u1_crc16_reg[0]/P0001  & ~\u1_u1_crc16_reg[14]/P0001  ;
  assign n2428 = ~n2244 & n2427 ;
  assign n2429 = ~n2205 & n2428 ;
  assign n2430 = ~\u1_u1_crc16_reg[0]/P0001  & ~\u1_u1_crc16_reg[14]/P0001  ;
  assign n2431 = ~n2244 & n2430 ;
  assign n2432 = n2205 & n2431 ;
  assign n2433 = ~n2429 & ~n2432 ;
  assign n2434 = n2244 & n2427 ;
  assign n2435 = n2205 & n2434 ;
  assign n2436 = n2244 & n2430 ;
  assign n2437 = ~n2205 & n2436 ;
  assign n2438 = ~n2435 & ~n2437 ;
  assign n2439 = n2433 & n2438 ;
  assign n2440 = ~\u1_u1_crc16_reg[0]/P0001  & \u1_u1_crc16_reg[14]/P0001  ;
  assign n2441 = ~n2244 & n2440 ;
  assign n2442 = ~n2205 & n2441 ;
  assign n2443 = \u1_u1_crc16_reg[0]/P0001  & \u1_u1_crc16_reg[14]/P0001  ;
  assign n2444 = ~n2244 & n2443 ;
  assign n2445 = n2205 & n2444 ;
  assign n2446 = ~n2442 & ~n2445 ;
  assign n2447 = n2244 & n2440 ;
  assign n2448 = n2205 & n2447 ;
  assign n2449 = n2244 & n2443 ;
  assign n2450 = ~n2205 & n2449 ;
  assign n2451 = ~n2448 & ~n2450 ;
  assign n2452 = n2446 & n2451 ;
  assign n2453 = ~n2285 & n2452 ;
  assign n2454 = n2439 & n2453 ;
  assign n2455 = \u1_u1_crc16_reg[8]/P0001  & ~n2284 ;
  assign n2456 = ~n2282 & n2455 ;
  assign n2457 = ~n2294 & ~n2456 ;
  assign n2458 = ~n2454 & n2457 ;
  assign n2459 = \u1_u1_crc16_reg[8]/P0001  & \u1_u1_crc16_reg[9]/P0001  ;
  assign n2460 = ~n2140 & n2459 ;
  assign n2461 = ~\u1_u1_crc16_reg[8]/P0001  & ~\u1_u1_crc16_reg[9]/P0001  ;
  assign n2462 = ~n2140 & n2461 ;
  assign n2463 = ~n2285 & ~n2462 ;
  assign n2464 = n2140 & n2397 ;
  assign n2465 = n2140 & n2396 ;
  assign n2466 = ~n2464 & ~n2465 ;
  assign n2467 = n2463 & n2466 ;
  assign n2468 = ~n2460 & n2467 ;
  assign n2469 = \u1_u1_crc16_reg[2]/P0001  & ~n2284 ;
  assign n2470 = ~n2282 & n2469 ;
  assign n2471 = ~n2294 & ~n2470 ;
  assign n2472 = ~n2468 & n2471 ;
  assign n2473 = n2247 & n2284 ;
  assign n2474 = n1757 & n2247 ;
  assign n2475 = n1860 & n2474 ;
  assign n2476 = ~n2473 & ~n2475 ;
  assign n2477 = ~n2321 & ~n2476 ;
  assign n2478 = ~n2247 & n2284 ;
  assign n2479 = n1757 & ~n2247 ;
  assign n2480 = n1860 & n2479 ;
  assign n2481 = ~n2478 & ~n2480 ;
  assign n2482 = n2321 & ~n2481 ;
  assign n2483 = \u1_u1_crc16_reg[3]/P0001  & ~n2284 ;
  assign n2484 = ~n2282 & n2483 ;
  assign n2485 = ~n2294 & ~n2484 ;
  assign n2486 = ~n2482 & n2485 ;
  assign n2487 = ~n2477 & n2486 ;
  assign n2488 = ~n2285 & ~n2312 ;
  assign n2489 = ~n2137 & n2488 ;
  assign n2490 = n2284 & n2312 ;
  assign n2491 = n1757 & n2312 ;
  assign n2492 = n1860 & n2491 ;
  assign n2493 = ~n2490 & ~n2492 ;
  assign n2494 = n2137 & ~n2493 ;
  assign n2495 = ~n2489 & ~n2494 ;
  assign n2496 = \u1_u1_crc16_reg[4]/P0001  & ~n2284 ;
  assign n2497 = ~n2282 & n2496 ;
  assign n2498 = ~n2294 & ~n2497 ;
  assign n2499 = n2495 & n2498 ;
  assign n2500 = n1827 & ~n2095 ;
  assign n2501 = ~n1827 & n2095 ;
  assign n2502 = ~n2500 & ~n2501 ;
  assign n2503 = n2250 & n2284 ;
  assign n2504 = n1757 & n2250 ;
  assign n2505 = n1860 & n2504 ;
  assign n2506 = ~n2503 & ~n2505 ;
  assign n2507 = ~n2502 & ~n2506 ;
  assign n2508 = ~n2250 & n2284 ;
  assign n2509 = n1757 & ~n2250 ;
  assign n2510 = n1860 & n2509 ;
  assign n2511 = ~n2508 & ~n2510 ;
  assign n2512 = n2502 & ~n2511 ;
  assign n2513 = \u1_u1_crc16_reg[5]/P0001  & ~n2284 ;
  assign n2514 = ~n2282 & n2513 ;
  assign n2515 = ~n2294 & ~n2514 ;
  assign n2516 = ~n2512 & n2515 ;
  assign n2517 = ~n2507 & n2516 ;
  assign n2518 = ~n2285 & ~n2324 ;
  assign n2519 = n2149 & n2518 ;
  assign n2520 = n2284 & n2324 ;
  assign n2521 = n1757 & n2324 ;
  assign n2522 = n1860 & n2521 ;
  assign n2523 = ~n2520 & ~n2522 ;
  assign n2524 = ~n2149 & ~n2523 ;
  assign n2525 = ~n2519 & ~n2524 ;
  assign n2526 = \u1_u1_crc16_reg[6]/P0001  & ~n2284 ;
  assign n2527 = ~n2282 & n2526 ;
  assign n2528 = ~n2294 & ~n2527 ;
  assign n2529 = n2525 & n2528 ;
  assign n2530 = ~n1977 & ~n2163 ;
  assign n2531 = n1977 & n2163 ;
  assign n2532 = ~n2530 & ~n2531 ;
  assign n2533 = n2244 & n2532 ;
  assign n2534 = n2244 & ~n2285 ;
  assign n2535 = n1977 & n2289 ;
  assign n2536 = ~n1977 & n2287 ;
  assign n2537 = ~n2535 & ~n2536 ;
  assign n2538 = ~n2534 & n2537 ;
  assign n2539 = ~n2533 & ~n2538 ;
  assign n2540 = \u1_u1_crc16_reg[7]/P0001  & ~n2284 ;
  assign n2541 = ~n2282 & n2540 ;
  assign n2542 = ~n2294 & ~n2541 ;
  assign n2543 = ~n2539 & n2542 ;
  assign n2544 = ~\u1_u1_crc16_reg[15]/P0001  & ~\u1_u1_crc16_reg[1]/P0001  ;
  assign n2545 = \u1_u1_crc16_reg[15]/P0001  & \u1_u1_crc16_reg[1]/P0001  ;
  assign n2546 = ~n2544 & ~n2545 ;
  assign n2547 = ~n2285 & ~n2546 ;
  assign n2548 = ~n2202 & n2547 ;
  assign n2549 = ~n2285 & n2546 ;
  assign n2550 = n2202 & n2549 ;
  assign n2551 = ~n2548 & ~n2550 ;
  assign n2552 = \u1_u1_crc16_reg[9]/P0001  & ~n2284 ;
  assign n2553 = ~n2282 & n2552 ;
  assign n2554 = ~n2294 & ~n2553 ;
  assign n2555 = n2551 & n2554 ;
  assign n2556 = ~\u5_state_reg[4]/P0001  & ~\u5_state_reg[5]/NET0131  ;
  assign n2557 = ~\u5_state_reg[3]/P0001  & n2556 ;
  assign n2558 = ~\u5_state_reg[1]/P0001  & ~\u5_state_reg[2]/P0001  ;
  assign n2559 = ~\wb_addr_i[17]_pad  & n2558 ;
  assign n2560 = n2557 & n2559 ;
  assign n2561 = ~\wb_addr_i[7]_pad  & ~\wb_addr_i[8]_pad  ;
  assign n2562 = \wb_addr_i[4]_pad  & n2561 ;
  assign n2563 = \wb_addr_i[5]_pad  & \wb_addr_i[6]_pad  ;
  assign n2564 = \u5_wb_req_s1_reg/P0001  & wb_we_i_pad ;
  assign n2565 = n2563 & n2564 ;
  assign n2566 = n2562 & n2565 ;
  assign n2567 = n2560 & n2566 ;
  assign n2568 = ~\wb_addr_i[2]_pad  & \wb_addr_i[3]_pad  ;
  assign n2569 = \wb_data_i[14]_pad  & n2568 ;
  assign n2570 = n2567 & n2569 ;
  assign n2571 = rst_i_pad & ~n2570 ;
  assign n2572 = n2567 & n2568 ;
  assign n2573 = \u1_u3_buf0_rl_reg/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n2574 = \u1_u3_buf0_set_reg/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n2575 = ~\u4_u3_buf0_reg[14]/P0001  & ~n2574 ;
  assign n2576 = ~\u1_u3_idin_reg[14]/P0001  & n2574 ;
  assign n2577 = ~n2575 & ~n2576 ;
  assign n2578 = ~n2573 & ~n2577 ;
  assign n2579 = ~\u4_u3_buf0_orig_reg[14]/P0001  & n2573 ;
  assign n2580 = ~n2578 & ~n2579 ;
  assign n2581 = ~n2572 & n2580 ;
  assign n2582 = n2571 & ~n2581 ;
  assign n2583 = ~\wb_addr_i[4]_pad  & n2561 ;
  assign n2584 = ~\wb_addr_i[5]_pad  & \wb_addr_i[6]_pad  ;
  assign n2585 = n2564 & n2584 ;
  assign n2586 = n2583 & n2585 ;
  assign n2587 = n2560 & n2586 ;
  assign n2588 = n2569 & n2587 ;
  assign n2589 = rst_i_pad & ~n2588 ;
  assign n2590 = n2568 & n2587 ;
  assign n2591 = \u1_u3_buf0_rl_reg/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n2592 = \u1_u3_buf0_set_reg/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n2593 = ~\u4_u0_buf0_reg[14]/P0001  & ~n2592 ;
  assign n2594 = ~\u1_u3_idin_reg[14]/P0001  & n2592 ;
  assign n2595 = ~n2593 & ~n2594 ;
  assign n2596 = ~n2591 & ~n2595 ;
  assign n2597 = \u1_u3_buf0_rl_reg/P0001  & ~\u4_u0_buf0_orig_reg[14]/P0001  ;
  assign n2598 = \u4_u0_ep_match_r_reg/P0001  & n2597 ;
  assign n2599 = ~n2596 & ~n2598 ;
  assign n2600 = ~n2590 & n2599 ;
  assign n2601 = n2589 & ~n2600 ;
  assign n2602 = n1753 & n1849 ;
  assign n2603 = ~\u1_u1_crc16_reg[14]/P0001  & ~n1860 ;
  assign n2604 = ~\u1_u1_crc16_reg[6]/P0001  & n1860 ;
  assign n2605 = ~n2603 & ~n2604 ;
  assign n2606 = n1753 & ~n1872 ;
  assign n2607 = ~n2605 & n2606 ;
  assign n2608 = ~n2602 & ~n2607 ;
  assign n2609 = n1753 & n1852 ;
  assign n2610 = n1841 & n2609 ;
  assign n2611 = ~n2244 & n2610 ;
  assign n2612 = n2608 & ~n2611 ;
  assign n2613 = ~n1749 & ~n1842 ;
  assign n2614 = ~n1752 & n2613 ;
  assign n2615 = \DataOut_pad_o[1]_pad  & ~\u0_u0_drive_k_reg/P0001  ;
  assign n2616 = ~n1753 & n2615 ;
  assign n2617 = ~n2614 & ~n2616 ;
  assign n2618 = n2612 & n2617 ;
  assign n2619 = n2562 & n2585 ;
  assign n2620 = n2560 & n2619 ;
  assign n2621 = n2569 & n2620 ;
  assign n2622 = rst_i_pad & ~n2621 ;
  assign n2623 = n2568 & n2620 ;
  assign n2624 = \u1_u3_buf0_rl_reg/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n2625 = \u1_u3_buf0_set_reg/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n2626 = ~\u4_u1_buf0_reg[14]/P0001  & ~n2625 ;
  assign n2627 = ~\u1_u3_idin_reg[14]/P0001  & n2625 ;
  assign n2628 = ~n2626 & ~n2627 ;
  assign n2629 = ~n2624 & ~n2628 ;
  assign n2630 = ~\u4_u1_buf0_orig_reg[14]/P0001  & n2624 ;
  assign n2631 = ~n2629 & ~n2630 ;
  assign n2632 = ~n2623 & n2631 ;
  assign n2633 = n2622 & ~n2632 ;
  assign n2634 = n2565 & n2583 ;
  assign n2635 = n2560 & n2634 ;
  assign n2636 = n2569 & n2635 ;
  assign n2637 = rst_i_pad & ~n2636 ;
  assign n2638 = n2568 & n2635 ;
  assign n2639 = \u1_u3_buf0_rl_reg/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n2640 = \u1_u3_buf0_set_reg/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n2641 = ~\u4_u2_buf0_reg[14]/P0001  & ~n2640 ;
  assign n2642 = ~\u1_u3_idin_reg[14]/P0001  & n2640 ;
  assign n2643 = ~n2641 & ~n2642 ;
  assign n2644 = ~n2639 & ~n2643 ;
  assign n2645 = ~\u4_u2_buf0_orig_reg[14]/P0001  & n2639 ;
  assign n2646 = ~n2644 & ~n2645 ;
  assign n2647 = ~n2638 & n2646 ;
  assign n2648 = n2637 & ~n2647 ;
  assign n2649 = \wb_data_i[10]_pad  & n2568 ;
  assign n2650 = n2567 & n2649 ;
  assign n2651 = rst_i_pad & ~n2650 ;
  assign n2652 = ~\u4_u3_buf0_reg[10]/P0001  & ~n2574 ;
  assign n2653 = ~\u1_u3_idin_reg[10]/P0001  & n2574 ;
  assign n2654 = ~n2652 & ~n2653 ;
  assign n2655 = ~n2573 & ~n2654 ;
  assign n2656 = ~\u4_u3_buf0_orig_reg[10]/P0001  & n2573 ;
  assign n2657 = ~n2655 & ~n2656 ;
  assign n2658 = ~n2572 & n2657 ;
  assign n2659 = n2651 & ~n2658 ;
  assign n2660 = n2587 & n2649 ;
  assign n2661 = rst_i_pad & ~n2660 ;
  assign n2662 = ~\u4_u0_buf0_reg[10]/P0001  & ~n2592 ;
  assign n2663 = ~\u1_u3_idin_reg[10]/P0001  & n2592 ;
  assign n2664 = ~n2662 & ~n2663 ;
  assign n2665 = ~n2591 & ~n2664 ;
  assign n2666 = ~\u4_u0_buf0_orig_reg[10]/P0001  & n2591 ;
  assign n2667 = ~n2665 & ~n2666 ;
  assign n2668 = ~n2590 & n2667 ;
  assign n2669 = n2661 & ~n2668 ;
  assign n2670 = n2620 & n2649 ;
  assign n2671 = rst_i_pad & ~n2670 ;
  assign n2672 = ~\u4_u1_buf0_reg[10]/P0001  & ~n2625 ;
  assign n2673 = ~\u1_u3_idin_reg[10]/P0001  & n2625 ;
  assign n2674 = ~n2672 & ~n2673 ;
  assign n2675 = ~n2624 & ~n2674 ;
  assign n2676 = ~\u4_u1_buf0_orig_reg[10]/P0001  & n2624 ;
  assign n2677 = ~n2675 & ~n2676 ;
  assign n2678 = ~n2623 & n2677 ;
  assign n2679 = n2671 & ~n2678 ;
  assign n2680 = n2635 & n2649 ;
  assign n2681 = rst_i_pad & ~n2680 ;
  assign n2682 = ~\u4_u2_buf0_reg[10]/P0001  & ~n2640 ;
  assign n2683 = ~\u1_u3_idin_reg[10]/P0001  & n2640 ;
  assign n2684 = ~n2682 & ~n2683 ;
  assign n2685 = ~n2639 & ~n2684 ;
  assign n2686 = ~\u4_u2_buf0_orig_reg[10]/P0001  & n2639 ;
  assign n2687 = ~n2685 & ~n2686 ;
  assign n2688 = ~n2638 & n2687 ;
  assign n2689 = n2681 & ~n2688 ;
  assign n2690 = \DataOut_pad_o[0]_pad  & ~\u0_u0_drive_k_reg/P0001  ;
  assign n2691 = ~n1753 & n2690 ;
  assign n2692 = ~n1749 & n1842 ;
  assign n2693 = ~n1752 & n2692 ;
  assign n2694 = ~\u1_u1_crc16_reg[15]/P0001  & ~n1860 ;
  assign n2695 = ~\u1_u1_crc16_reg[7]/P0001  & n1860 ;
  assign n2696 = ~n2694 & ~n2695 ;
  assign n2697 = ~n1872 & ~n2696 ;
  assign n2698 = ~n1849 & ~n2697 ;
  assign n2699 = n1872 & ~n2202 ;
  assign n2700 = n2698 & ~n2699 ;
  assign n2701 = n2693 & ~n2700 ;
  assign n2702 = ~n2691 & ~n2701 ;
  assign n2703 = \DataOut_pad_o[4]_pad  & ~\u0_u0_drive_k_reg/P0001  ;
  assign n2704 = ~n1753 & n2703 ;
  assign n2705 = ~n2614 & ~n2704 ;
  assign n2706 = n1872 & n2705 ;
  assign n2707 = n2095 & n2706 ;
  assign n2708 = ~n1753 & n2705 ;
  assign n2709 = ~\u1_u1_crc16_reg[11]/P0001  & ~n1860 ;
  assign n2710 = ~n1872 & ~n2709 ;
  assign n2711 = ~\u1_u1_crc16_reg[3]/P0001  & n1862 ;
  assign n2712 = ~\u1_u1_crc16_reg[3]/P0001  & n1834 ;
  assign n2713 = n1838 & n2712 ;
  assign n2714 = ~n2711 & ~n2713 ;
  assign n2715 = n1860 & ~n2714 ;
  assign n2716 = n2705 & ~n2715 ;
  assign n2717 = n2710 & n2716 ;
  assign n2718 = ~n2708 & ~n2717 ;
  assign n2719 = ~n2707 & n2718 ;
  assign n2720 = \wb_data_i[13]_pad  & n2568 ;
  assign n2721 = n2567 & n2720 ;
  assign n2722 = rst_i_pad & ~n2721 ;
  assign n2723 = ~\u4_u3_buf0_reg[13]/P0001  & ~n2574 ;
  assign n2724 = ~\u1_u3_idin_reg[13]/P0001  & n2574 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = ~n2573 & ~n2725 ;
  assign n2727 = ~\u4_u3_buf0_orig_reg[13]/P0001  & n2573 ;
  assign n2728 = ~n2726 & ~n2727 ;
  assign n2729 = ~n2572 & n2728 ;
  assign n2730 = n2722 & ~n2729 ;
  assign n2731 = \wb_addr_i[2]_pad  & \wb_addr_i[3]_pad  ;
  assign n2732 = n2567 & n2731 ;
  assign n2733 = ~\u1_u3_buf1_set_reg/P0001  & ~\u1_u3_out_to_small_reg/P0001  ;
  assign n2734 = \u4_u3_ep_match_r_reg/P0001  & ~n2733 ;
  assign n2735 = \u4_u3_buf1_reg[14]/P0001  & ~n2734 ;
  assign n2736 = \u1_u3_idin_reg[14]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n2737 = ~n2733 & n2736 ;
  assign n2738 = ~n2735 & ~n2737 ;
  assign n2739 = ~n2732 & ~n2738 ;
  assign n2740 = \wb_data_i[14]_pad  & n2731 ;
  assign n2741 = n2567 & n2740 ;
  assign n2742 = rst_i_pad & ~n2741 ;
  assign n2743 = ~n2739 & n2742 ;
  assign n2744 = n2587 & n2720 ;
  assign n2745 = rst_i_pad & ~n2744 ;
  assign n2746 = ~\u4_u0_buf0_reg[13]/P0001  & ~n2592 ;
  assign n2747 = ~\u1_u3_idin_reg[13]/P0001  & n2592 ;
  assign n2748 = ~n2746 & ~n2747 ;
  assign n2749 = ~n2591 & ~n2748 ;
  assign n2750 = ~\u4_u0_buf0_orig_reg[13]/P0001  & n2591 ;
  assign n2751 = ~n2749 & ~n2750 ;
  assign n2752 = ~n2590 & n2751 ;
  assign n2753 = n2745 & ~n2752 ;
  assign n2754 = n2587 & n2731 ;
  assign n2755 = \u4_u0_ep_match_r_reg/P0001  & ~n2733 ;
  assign n2756 = \u4_u0_buf1_reg[14]/P0001  & ~n2755 ;
  assign n2757 = \u1_u3_idin_reg[14]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n2758 = ~n2733 & n2757 ;
  assign n2759 = ~n2756 & ~n2758 ;
  assign n2760 = ~n2754 & ~n2759 ;
  assign n2761 = n2587 & n2740 ;
  assign n2762 = rst_i_pad & ~n2761 ;
  assign n2763 = ~n2760 & n2762 ;
  assign n2764 = n2620 & n2720 ;
  assign n2765 = rst_i_pad & ~n2764 ;
  assign n2766 = ~\u4_u1_buf0_reg[13]/P0001  & ~n2625 ;
  assign n2767 = ~\u1_u3_idin_reg[13]/P0001  & n2625 ;
  assign n2768 = ~n2766 & ~n2767 ;
  assign n2769 = ~n2624 & ~n2768 ;
  assign n2770 = ~\u4_u1_buf0_orig_reg[13]/P0001  & n2624 ;
  assign n2771 = ~n2769 & ~n2770 ;
  assign n2772 = ~n2623 & n2771 ;
  assign n2773 = n2765 & ~n2772 ;
  assign n2774 = n2620 & n2731 ;
  assign n2775 = \u4_u1_ep_match_r_reg/P0001  & ~n2733 ;
  assign n2776 = \u4_u1_buf1_reg[14]/P0001  & ~n2775 ;
  assign n2777 = \u1_u3_idin_reg[14]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n2778 = ~n2733 & n2777 ;
  assign n2779 = ~n2776 & ~n2778 ;
  assign n2780 = ~n2774 & ~n2779 ;
  assign n2781 = n2620 & n2740 ;
  assign n2782 = rst_i_pad & ~n2781 ;
  assign n2783 = ~n2780 & n2782 ;
  assign n2784 = ~\u1_u3_buf0_na_reg/NET0131  & ~n2367 ;
  assign n2785 = \u1_u3_buf0_st_max_reg/P0001  & \u1_u3_in_token_reg/NET0131  ;
  assign n2786 = n2358 & n2785 ;
  assign n2787 = ~\u1_u3_buf1_na_reg/NET0131  & ~\u4_csr_reg[15]/NET0131  ;
  assign n2788 = ~n2358 & n2787 ;
  assign n2789 = ~\u1_u3_buf0_na_reg/NET0131  & ~\u4_csr_reg[30]/NET0131  ;
  assign n2790 = \u1_u3_buf0_st_max_reg/P0001  & ~n2789 ;
  assign n2791 = n2788 & n2790 ;
  assign n2792 = ~n2786 & ~n2791 ;
  assign n2793 = \u1_u3_in_token_reg/NET0131  & n2358 ;
  assign n2794 = n2788 & ~n2789 ;
  assign n2795 = ~n2793 & ~n2794 ;
  assign n2796 = \u1_u3_buffer_full_reg/P0001  & ~n2366 ;
  assign n2797 = n2795 & n2796 ;
  assign n2798 = n2792 & ~n2797 ;
  assign n2799 = n2784 & n2798 ;
  assign n2800 = n2635 & n2720 ;
  assign n2801 = rst_i_pad & ~n2800 ;
  assign n2802 = ~\u4_u2_buf0_reg[13]/P0001  & ~n2640 ;
  assign n2803 = ~\u1_u3_idin_reg[13]/P0001  & n2640 ;
  assign n2804 = ~n2802 & ~n2803 ;
  assign n2805 = ~n2639 & ~n2804 ;
  assign n2806 = ~\u4_u2_buf0_orig_reg[13]/P0001  & n2639 ;
  assign n2807 = ~n2805 & ~n2806 ;
  assign n2808 = ~n2638 & n2807 ;
  assign n2809 = n2801 & ~n2808 ;
  assign n2810 = n2635 & n2731 ;
  assign n2811 = \u4_u2_ep_match_r_reg/P0001  & ~n2733 ;
  assign n2812 = \u4_u2_buf1_reg[14]/P0001  & ~n2811 ;
  assign n2813 = \u1_u3_idin_reg[14]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n2814 = ~n2733 & n2813 ;
  assign n2815 = ~n2812 & ~n2814 ;
  assign n2816 = ~n2810 & ~n2815 ;
  assign n2817 = n2635 & n2740 ;
  assign n2818 = rst_i_pad & ~n2817 ;
  assign n2819 = ~n2816 & n2818 ;
  assign n2820 = \DataOut_pad_o[5]_pad  & ~\u0_u0_drive_k_reg/P0001  ;
  assign n2821 = ~n1753 & n2820 ;
  assign n2822 = ~n2693 & ~n2821 ;
  assign n2823 = ~\u1_u1_crc16_reg[10]/P0001  & ~n1860 ;
  assign n2824 = ~n1872 & ~n2823 ;
  assign n2825 = ~\u1_u1_crc16_reg[2]/P0001  & n1862 ;
  assign n2826 = ~\u1_u1_crc16_reg[2]/P0001  & n1834 ;
  assign n2827 = n1838 & n2826 ;
  assign n2828 = ~n2825 & ~n2827 ;
  assign n2829 = n1860 & ~n2828 ;
  assign n2830 = ~n2821 & ~n2829 ;
  assign n2831 = n2824 & n2830 ;
  assign n2832 = ~n2822 & ~n2831 ;
  assign n2833 = n1872 & ~n2821 ;
  assign n2834 = n2134 & n2833 ;
  assign n2835 = n2832 & ~n2834 ;
  assign n2836 = \u1_u3_buffer_full_reg/P0001  & n2793 ;
  assign n2837 = \u1_u3_buffer_full_reg/P0001  & ~n2789 ;
  assign n2838 = n2788 & n2837 ;
  assign n2839 = ~n2836 & ~n2838 ;
  assign n2840 = \u1_u3_buf1_st_max_reg/P0001  & ~n2793 ;
  assign n2841 = ~n2794 & n2840 ;
  assign n2842 = ~\u1_u3_buf1_na_reg/NET0131  & ~n2841 ;
  assign n2843 = n2839 & n2842 ;
  assign n2844 = \wb_data_i[11]_pad  & n2568 ;
  assign n2845 = n2567 & n2844 ;
  assign n2846 = rst_i_pad & ~n2845 ;
  assign n2847 = ~\u4_u3_buf0_reg[11]/P0001  & ~n2574 ;
  assign n2848 = ~\u1_u3_idin_reg[11]/P0001  & n2574 ;
  assign n2849 = ~n2847 & ~n2848 ;
  assign n2850 = ~n2573 & ~n2849 ;
  assign n2851 = ~\u4_u3_buf0_orig_reg[11]/P0001  & n2573 ;
  assign n2852 = ~n2850 & ~n2851 ;
  assign n2853 = ~n2572 & n2852 ;
  assign n2854 = n2846 & ~n2853 ;
  assign n2855 = \wb_data_i[15]_pad  & n2568 ;
  assign n2856 = n2567 & n2855 ;
  assign n2857 = rst_i_pad & ~n2856 ;
  assign n2858 = ~\u4_u3_buf0_reg[15]/P0001  & ~n2574 ;
  assign n2859 = ~\u1_u3_idin_reg[15]/P0001  & n2574 ;
  assign n2860 = ~n2858 & ~n2859 ;
  assign n2861 = ~n2573 & ~n2860 ;
  assign n2862 = ~\u4_u3_buf0_orig_reg[15]/P0001  & n2573 ;
  assign n2863 = ~n2861 & ~n2862 ;
  assign n2864 = ~n2572 & n2863 ;
  assign n2865 = n2857 & ~n2864 ;
  assign n2866 = \u4_u3_buf1_reg[10]/P0001  & ~n2734 ;
  assign n2867 = \u1_u3_idin_reg[10]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n2868 = ~n2733 & n2867 ;
  assign n2869 = ~n2866 & ~n2868 ;
  assign n2870 = ~n2732 & ~n2869 ;
  assign n2871 = \wb_data_i[10]_pad  & n2731 ;
  assign n2872 = n2567 & n2871 ;
  assign n2873 = rst_i_pad & ~n2872 ;
  assign n2874 = ~n2870 & n2873 ;
  assign n2875 = \wb_data_i[6]_pad  & n2568 ;
  assign n2876 = n2567 & n2875 ;
  assign n2877 = rst_i_pad & ~n2876 ;
  assign n2878 = ~\u4_u3_buf0_reg[6]/P0001  & ~n2574 ;
  assign n2879 = ~\u1_u3_idin_reg[6]/P0001  & n2574 ;
  assign n2880 = ~n2878 & ~n2879 ;
  assign n2881 = ~n2573 & ~n2880 ;
  assign n2882 = ~\u4_u3_buf0_orig_reg[6]/P0001  & n2573 ;
  assign n2883 = ~n2881 & ~n2882 ;
  assign n2884 = ~n2572 & n2883 ;
  assign n2885 = n2877 & ~n2884 ;
  assign n2886 = n2587 & n2844 ;
  assign n2887 = rst_i_pad & ~n2886 ;
  assign n2888 = ~\u4_u0_buf0_reg[11]/P0001  & ~n2592 ;
  assign n2889 = ~\u1_u3_idin_reg[11]/P0001  & n2592 ;
  assign n2890 = ~n2888 & ~n2889 ;
  assign n2891 = ~n2591 & ~n2890 ;
  assign n2892 = ~\u4_u0_buf0_orig_reg[11]/P0001  & n2591 ;
  assign n2893 = ~n2891 & ~n2892 ;
  assign n2894 = ~n2590 & n2893 ;
  assign n2895 = n2887 & ~n2894 ;
  assign n2896 = n2587 & n2855 ;
  assign n2897 = rst_i_pad & ~n2896 ;
  assign n2898 = ~\u4_u0_buf0_reg[15]/P0001  & ~n2592 ;
  assign n2899 = ~\u1_u3_idin_reg[15]/P0001  & n2592 ;
  assign n2900 = ~n2898 & ~n2899 ;
  assign n2901 = ~n2591 & ~n2900 ;
  assign n2902 = ~\u4_u0_buf0_orig_reg[15]/P0001  & n2591 ;
  assign n2903 = ~n2901 & ~n2902 ;
  assign n2904 = ~n2590 & n2903 ;
  assign n2905 = n2897 & ~n2904 ;
  assign n2906 = n2587 & n2875 ;
  assign n2907 = rst_i_pad & ~n2906 ;
  assign n2908 = ~\u4_u0_buf0_reg[6]/P0001  & ~n2592 ;
  assign n2909 = ~\u1_u3_idin_reg[6]/P0001  & n2592 ;
  assign n2910 = ~n2908 & ~n2909 ;
  assign n2911 = ~n2591 & ~n2910 ;
  assign n2912 = ~\u4_u0_buf0_orig_reg[6]/P0001  & n2591 ;
  assign n2913 = ~n2911 & ~n2912 ;
  assign n2914 = ~n2590 & n2913 ;
  assign n2915 = n2907 & ~n2914 ;
  assign n2916 = \u4_u0_buf1_reg[10]/P0001  & ~n2755 ;
  assign n2917 = \u1_u3_idin_reg[10]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n2918 = ~n2733 & n2917 ;
  assign n2919 = ~n2916 & ~n2918 ;
  assign n2920 = ~n2754 & ~n2919 ;
  assign n2921 = n2587 & n2871 ;
  assign n2922 = rst_i_pad & ~n2921 ;
  assign n2923 = ~n2920 & n2922 ;
  assign n2924 = n2620 & n2844 ;
  assign n2925 = rst_i_pad & ~n2924 ;
  assign n2926 = ~\u4_u1_buf0_reg[11]/P0001  & ~n2625 ;
  assign n2927 = ~\u1_u3_idin_reg[11]/P0001  & n2625 ;
  assign n2928 = ~n2926 & ~n2927 ;
  assign n2929 = ~n2624 & ~n2928 ;
  assign n2930 = ~\u4_u1_buf0_orig_reg[11]/P0001  & n2624 ;
  assign n2931 = ~n2929 & ~n2930 ;
  assign n2932 = ~n2623 & n2931 ;
  assign n2933 = n2925 & ~n2932 ;
  assign n2934 = n2620 & n2855 ;
  assign n2935 = rst_i_pad & ~n2934 ;
  assign n2936 = ~\u4_u1_buf0_reg[15]/P0001  & ~n2625 ;
  assign n2937 = ~\u1_u3_idin_reg[15]/P0001  & n2625 ;
  assign n2938 = ~n2936 & ~n2937 ;
  assign n2939 = ~n2624 & ~n2938 ;
  assign n2940 = ~\u4_u1_buf0_orig_reg[15]/P0001  & n2624 ;
  assign n2941 = ~n2939 & ~n2940 ;
  assign n2942 = ~n2623 & n2941 ;
  assign n2943 = n2935 & ~n2942 ;
  assign n2944 = \u4_u1_buf1_reg[10]/P0001  & ~n2775 ;
  assign n2945 = \u1_u3_idin_reg[10]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n2946 = ~n2733 & n2945 ;
  assign n2947 = ~n2944 & ~n2946 ;
  assign n2948 = ~n2774 & ~n2947 ;
  assign n2949 = n2620 & n2871 ;
  assign n2950 = rst_i_pad & ~n2949 ;
  assign n2951 = ~n2948 & n2950 ;
  assign n2952 = n2620 & n2875 ;
  assign n2953 = rst_i_pad & ~n2952 ;
  assign n2954 = ~\u4_u1_buf0_reg[6]/P0001  & ~n2625 ;
  assign n2955 = ~\u1_u3_idin_reg[6]/P0001  & n2625 ;
  assign n2956 = ~n2954 & ~n2955 ;
  assign n2957 = ~n2624 & ~n2956 ;
  assign n2958 = ~\u4_u1_buf0_orig_reg[6]/P0001  & n2624 ;
  assign n2959 = ~n2957 & ~n2958 ;
  assign n2960 = ~n2623 & n2959 ;
  assign n2961 = n2953 & ~n2960 ;
  assign n2962 = n2635 & n2844 ;
  assign n2963 = rst_i_pad & ~n2962 ;
  assign n2964 = ~\u4_u2_buf0_reg[11]/P0001  & ~n2640 ;
  assign n2965 = ~\u1_u3_idin_reg[11]/P0001  & n2640 ;
  assign n2966 = ~n2964 & ~n2965 ;
  assign n2967 = ~n2639 & ~n2966 ;
  assign n2968 = ~\u4_u2_buf0_orig_reg[11]/P0001  & n2639 ;
  assign n2969 = ~n2967 & ~n2968 ;
  assign n2970 = ~n2638 & n2969 ;
  assign n2971 = n2963 & ~n2970 ;
  assign n2972 = n2635 & n2855 ;
  assign n2973 = rst_i_pad & ~n2972 ;
  assign n2974 = ~\u4_u2_buf0_reg[15]/P0001  & ~n2640 ;
  assign n2975 = ~\u1_u3_idin_reg[15]/P0001  & n2640 ;
  assign n2976 = ~n2974 & ~n2975 ;
  assign n2977 = ~n2639 & ~n2976 ;
  assign n2978 = ~\u4_u2_buf0_orig_reg[15]/P0001  & n2639 ;
  assign n2979 = ~n2977 & ~n2978 ;
  assign n2980 = ~n2638 & n2979 ;
  assign n2981 = n2973 & ~n2980 ;
  assign n2982 = \u4_u2_buf1_reg[10]/P0001  & ~n2811 ;
  assign n2983 = \u1_u3_idin_reg[10]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n2984 = ~n2733 & n2983 ;
  assign n2985 = ~n2982 & ~n2984 ;
  assign n2986 = ~n2810 & ~n2985 ;
  assign n2987 = n2635 & n2871 ;
  assign n2988 = rst_i_pad & ~n2987 ;
  assign n2989 = ~n2986 & n2988 ;
  assign n2990 = n2635 & n2875 ;
  assign n2991 = rst_i_pad & ~n2990 ;
  assign n2992 = ~\u4_u2_buf0_reg[6]/P0001  & ~n2640 ;
  assign n2993 = ~\u1_u3_idin_reg[6]/P0001  & n2640 ;
  assign n2994 = ~n2992 & ~n2993 ;
  assign n2995 = ~n2639 & ~n2994 ;
  assign n2996 = ~\u4_u2_buf0_orig_reg[6]/P0001  & n2639 ;
  assign n2997 = ~n2995 & ~n2996 ;
  assign n2998 = ~n2638 & n2997 ;
  assign n2999 = n2991 & ~n2998 ;
  assign n3000 = \u4_u3_buf1_reg[13]/P0001  & ~n2734 ;
  assign n3001 = \u1_u3_idin_reg[13]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n3002 = ~n2733 & n3001 ;
  assign n3003 = ~n3000 & ~n3002 ;
  assign n3004 = ~n2732 & ~n3003 ;
  assign n3005 = \wb_data_i[13]_pad  & n2731 ;
  assign n3006 = n2567 & n3005 ;
  assign n3007 = rst_i_pad & ~n3006 ;
  assign n3008 = ~n3004 & n3007 ;
  assign n3009 = \u4_u0_buf1_reg[13]/P0001  & ~n2755 ;
  assign n3010 = \u1_u3_idin_reg[13]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n3011 = ~n2733 & n3010 ;
  assign n3012 = ~n3009 & ~n3011 ;
  assign n3013 = ~n2754 & ~n3012 ;
  assign n3014 = n2587 & n3005 ;
  assign n3015 = rst_i_pad & ~n3014 ;
  assign n3016 = ~n3013 & n3015 ;
  assign n3017 = \u4_u1_buf1_reg[13]/P0001  & ~n2775 ;
  assign n3018 = \u1_u3_idin_reg[13]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n3019 = ~n2733 & n3018 ;
  assign n3020 = ~n3017 & ~n3019 ;
  assign n3021 = ~n2774 & ~n3020 ;
  assign n3022 = n2620 & n3005 ;
  assign n3023 = rst_i_pad & ~n3022 ;
  assign n3024 = ~n3021 & n3023 ;
  assign n3025 = \u4_u2_buf1_reg[13]/P0001  & ~n2811 ;
  assign n3026 = \u1_u3_idin_reg[13]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n3027 = ~n2733 & n3026 ;
  assign n3028 = ~n3025 & ~n3027 ;
  assign n3029 = ~n2810 & ~n3028 ;
  assign n3030 = n2635 & n3005 ;
  assign n3031 = rst_i_pad & ~n3030 ;
  assign n3032 = ~n3029 & n3031 ;
  assign n3033 = ~\u1_u3_in_token_reg/NET0131  & ~\u4_csr_reg[26]/NET0131  ;
  assign n3034 = \u1_u3_buffer_empty_reg/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3035 = ~n3033 & n3034 ;
  assign n3036 = ~\u4_csr_reg[27]/NET0131  & ~n3033 ;
  assign n3037 = \u1_u3_buffer_full_reg/P0001  & ~n3036 ;
  assign n3038 = ~n3035 & ~n3037 ;
  assign n3039 = \wb_data_i[4]_pad  & n2568 ;
  assign n3040 = n2567 & n3039 ;
  assign n3041 = rst_i_pad & ~n3040 ;
  assign n3042 = ~\u4_u3_buf0_reg[4]/P0001  & ~n2574 ;
  assign n3043 = ~\u1_u3_idin_reg[4]/P0001  & n2574 ;
  assign n3044 = ~n3042 & ~n3043 ;
  assign n3045 = ~n2573 & ~n3044 ;
  assign n3046 = ~\u4_u3_buf0_orig_reg[4]/P0001  & n2573 ;
  assign n3047 = ~n3045 & ~n3046 ;
  assign n3048 = ~n2572 & n3047 ;
  assign n3049 = n3041 & ~n3048 ;
  assign n3050 = \wb_data_i[5]_pad  & n2568 ;
  assign n3051 = n2567 & n3050 ;
  assign n3052 = rst_i_pad & ~n3051 ;
  assign n3053 = ~\u4_u3_buf0_reg[5]/P0001  & ~n2574 ;
  assign n3054 = ~\u1_u3_idin_reg[5]/P0001  & n2574 ;
  assign n3055 = ~n3053 & ~n3054 ;
  assign n3056 = ~n2573 & ~n3055 ;
  assign n3057 = ~\u4_u3_buf0_orig_reg[5]/P0001  & n2573 ;
  assign n3058 = ~n3056 & ~n3057 ;
  assign n3059 = ~n2572 & n3058 ;
  assign n3060 = n3052 & ~n3059 ;
  assign n3061 = \wb_data_i[7]_pad  & n2568 ;
  assign n3062 = n2567 & n3061 ;
  assign n3063 = rst_i_pad & ~n3062 ;
  assign n3064 = ~\u4_u3_buf0_reg[7]/P0001  & ~n2574 ;
  assign n3065 = ~\u1_u3_idin_reg[7]/P0001  & n2574 ;
  assign n3066 = ~n3064 & ~n3065 ;
  assign n3067 = ~n2573 & ~n3066 ;
  assign n3068 = ~\u4_u3_buf0_orig_reg[7]/P0001  & n2573 ;
  assign n3069 = ~n3067 & ~n3068 ;
  assign n3070 = ~n2572 & n3069 ;
  assign n3071 = n3063 & ~n3070 ;
  assign n3072 = \u4_u3_buf1_reg[11]/P0001  & ~n2734 ;
  assign n3073 = \u1_u3_idin_reg[11]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n3074 = ~n2733 & n3073 ;
  assign n3075 = ~n3072 & ~n3074 ;
  assign n3076 = ~n2732 & ~n3075 ;
  assign n3077 = \wb_data_i[11]_pad  & n2731 ;
  assign n3078 = n2567 & n3077 ;
  assign n3079 = rst_i_pad & ~n3078 ;
  assign n3080 = ~n3076 & n3079 ;
  assign n3081 = \u4_u3_buf1_reg[15]/P0001  & ~n2734 ;
  assign n3082 = \u1_u3_idin_reg[15]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n3083 = ~n2733 & n3082 ;
  assign n3084 = ~n3081 & ~n3083 ;
  assign n3085 = ~n2732 & ~n3084 ;
  assign n3086 = \wb_data_i[15]_pad  & n2731 ;
  assign n3087 = n2567 & n3086 ;
  assign n3088 = rst_i_pad & ~n3087 ;
  assign n3089 = ~n3085 & n3088 ;
  assign n3090 = \u4_u3_buf1_reg[6]/P0001  & ~n2734 ;
  assign n3091 = \u1_u3_idin_reg[6]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n3092 = ~n2733 & n3091 ;
  assign n3093 = ~n3090 & ~n3092 ;
  assign n3094 = ~n2732 & ~n3093 ;
  assign n3095 = \wb_data_i[6]_pad  & n2731 ;
  assign n3096 = n2567 & n3095 ;
  assign n3097 = rst_i_pad & ~n3096 ;
  assign n3098 = ~n3094 & n3097 ;
  assign n3099 = n2587 & n3039 ;
  assign n3100 = rst_i_pad & ~n3099 ;
  assign n3101 = ~\u4_u0_buf0_reg[4]/P0001  & ~n2592 ;
  assign n3102 = ~\u1_u3_idin_reg[4]/P0001  & n2592 ;
  assign n3103 = ~n3101 & ~n3102 ;
  assign n3104 = ~n2591 & ~n3103 ;
  assign n3105 = ~\u4_u0_buf0_orig_reg[4]/P0001  & n2591 ;
  assign n3106 = ~n3104 & ~n3105 ;
  assign n3107 = ~n2590 & n3106 ;
  assign n3108 = n3100 & ~n3107 ;
  assign n3109 = n2587 & n3050 ;
  assign n3110 = rst_i_pad & ~n3109 ;
  assign n3111 = ~\u4_u0_buf0_reg[5]/P0001  & ~n2592 ;
  assign n3112 = ~\u1_u3_idin_reg[5]/P0001  & n2592 ;
  assign n3113 = ~n3111 & ~n3112 ;
  assign n3114 = ~n2591 & ~n3113 ;
  assign n3115 = ~\u4_u0_buf0_orig_reg[5]/P0001  & n2591 ;
  assign n3116 = ~n3114 & ~n3115 ;
  assign n3117 = ~n2590 & n3116 ;
  assign n3118 = n3110 & ~n3117 ;
  assign n3119 = n2587 & n3061 ;
  assign n3120 = rst_i_pad & ~n3119 ;
  assign n3121 = ~\u4_u0_buf0_reg[7]/P0001  & ~n2592 ;
  assign n3122 = ~\u1_u3_idin_reg[7]/P0001  & n2592 ;
  assign n3123 = ~n3121 & ~n3122 ;
  assign n3124 = ~n2591 & ~n3123 ;
  assign n3125 = ~\u4_u0_buf0_orig_reg[7]/P0001  & n2591 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = ~n2590 & n3126 ;
  assign n3128 = n3120 & ~n3127 ;
  assign n3129 = \u4_u0_buf1_reg[11]/P0001  & ~n2755 ;
  assign n3130 = \u1_u3_idin_reg[11]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n3131 = ~n2733 & n3130 ;
  assign n3132 = ~n3129 & ~n3131 ;
  assign n3133 = ~n2754 & ~n3132 ;
  assign n3134 = n2587 & n3077 ;
  assign n3135 = rst_i_pad & ~n3134 ;
  assign n3136 = ~n3133 & n3135 ;
  assign n3137 = \u4_u0_buf1_reg[15]/P0001  & ~n2755 ;
  assign n3138 = \u1_u3_idin_reg[15]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n3139 = ~n2733 & n3138 ;
  assign n3140 = ~n3137 & ~n3139 ;
  assign n3141 = ~n2754 & ~n3140 ;
  assign n3142 = n2587 & n3086 ;
  assign n3143 = rst_i_pad & ~n3142 ;
  assign n3144 = ~n3141 & n3143 ;
  assign n3145 = \u4_u0_buf1_reg[6]/P0001  & ~n2755 ;
  assign n3146 = \u1_u3_idin_reg[6]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n3147 = ~n2733 & n3146 ;
  assign n3148 = ~n3145 & ~n3147 ;
  assign n3149 = ~n2754 & ~n3148 ;
  assign n3150 = n2587 & n3095 ;
  assign n3151 = rst_i_pad & ~n3150 ;
  assign n3152 = ~n3149 & n3151 ;
  assign n3153 = n2620 & n3039 ;
  assign n3154 = rst_i_pad & ~n3153 ;
  assign n3155 = ~\u4_u1_buf0_reg[4]/P0001  & ~n2625 ;
  assign n3156 = ~\u1_u3_idin_reg[4]/P0001  & n2625 ;
  assign n3157 = ~n3155 & ~n3156 ;
  assign n3158 = ~n2624 & ~n3157 ;
  assign n3159 = ~\u4_u1_buf0_orig_reg[4]/P0001  & n2624 ;
  assign n3160 = ~n3158 & ~n3159 ;
  assign n3161 = ~n2623 & n3160 ;
  assign n3162 = n3154 & ~n3161 ;
  assign n3163 = n2620 & n3050 ;
  assign n3164 = rst_i_pad & ~n3163 ;
  assign n3165 = ~\u4_u1_buf0_reg[5]/P0001  & ~n2625 ;
  assign n3166 = ~\u1_u3_idin_reg[5]/P0001  & n2625 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = ~n2624 & ~n3167 ;
  assign n3169 = ~\u4_u1_buf0_orig_reg[5]/P0001  & n2624 ;
  assign n3170 = ~n3168 & ~n3169 ;
  assign n3171 = ~n2623 & n3170 ;
  assign n3172 = n3164 & ~n3171 ;
  assign n3173 = n2620 & n3061 ;
  assign n3174 = rst_i_pad & ~n3173 ;
  assign n3175 = ~\u4_u1_buf0_reg[7]/P0001  & ~n2625 ;
  assign n3176 = ~\u1_u3_idin_reg[7]/P0001  & n2625 ;
  assign n3177 = ~n3175 & ~n3176 ;
  assign n3178 = ~n2624 & ~n3177 ;
  assign n3179 = ~\u4_u1_buf0_orig_reg[7]/P0001  & n2624 ;
  assign n3180 = ~n3178 & ~n3179 ;
  assign n3181 = ~n2623 & n3180 ;
  assign n3182 = n3174 & ~n3181 ;
  assign n3183 = \u4_u1_buf1_reg[11]/P0001  & ~n2775 ;
  assign n3184 = \u1_u3_idin_reg[11]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n3185 = ~n2733 & n3184 ;
  assign n3186 = ~n3183 & ~n3185 ;
  assign n3187 = ~n2774 & ~n3186 ;
  assign n3188 = n2620 & n3077 ;
  assign n3189 = rst_i_pad & ~n3188 ;
  assign n3190 = ~n3187 & n3189 ;
  assign n3191 = \u4_u1_buf1_reg[15]/P0001  & ~n2775 ;
  assign n3192 = \u1_u3_idin_reg[15]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n3193 = ~n2733 & n3192 ;
  assign n3194 = ~n3191 & ~n3193 ;
  assign n3195 = ~n2774 & ~n3194 ;
  assign n3196 = n2620 & n3086 ;
  assign n3197 = rst_i_pad & ~n3196 ;
  assign n3198 = ~n3195 & n3197 ;
  assign n3199 = \u4_u1_buf1_reg[6]/P0001  & ~n2775 ;
  assign n3200 = \u1_u3_idin_reg[6]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n3201 = ~n2733 & n3200 ;
  assign n3202 = ~n3199 & ~n3201 ;
  assign n3203 = ~n2774 & ~n3202 ;
  assign n3204 = n2620 & n3095 ;
  assign n3205 = rst_i_pad & ~n3204 ;
  assign n3206 = ~n3203 & n3205 ;
  assign n3207 = n2635 & n3039 ;
  assign n3208 = rst_i_pad & ~n3207 ;
  assign n3209 = ~\u4_u2_buf0_reg[4]/P0001  & ~n2640 ;
  assign n3210 = ~\u1_u3_idin_reg[4]/P0001  & n2640 ;
  assign n3211 = ~n3209 & ~n3210 ;
  assign n3212 = ~n2639 & ~n3211 ;
  assign n3213 = ~\u4_u2_buf0_orig_reg[4]/P0001  & n2639 ;
  assign n3214 = ~n3212 & ~n3213 ;
  assign n3215 = ~n2638 & n3214 ;
  assign n3216 = n3208 & ~n3215 ;
  assign n3217 = n2635 & n3050 ;
  assign n3218 = rst_i_pad & ~n3217 ;
  assign n3219 = ~\u4_u2_buf0_reg[5]/P0001  & ~n2640 ;
  assign n3220 = ~\u1_u3_idin_reg[5]/P0001  & n2640 ;
  assign n3221 = ~n3219 & ~n3220 ;
  assign n3222 = ~n2639 & ~n3221 ;
  assign n3223 = ~\u4_u2_buf0_orig_reg[5]/P0001  & n2639 ;
  assign n3224 = ~n3222 & ~n3223 ;
  assign n3225 = ~n2638 & n3224 ;
  assign n3226 = n3218 & ~n3225 ;
  assign n3227 = n2635 & n3061 ;
  assign n3228 = rst_i_pad & ~n3227 ;
  assign n3229 = ~\u4_u2_buf0_reg[7]/P0001  & ~n2640 ;
  assign n3230 = ~\u1_u3_idin_reg[7]/P0001  & n2640 ;
  assign n3231 = ~n3229 & ~n3230 ;
  assign n3232 = ~n2639 & ~n3231 ;
  assign n3233 = ~\u4_u2_buf0_orig_reg[7]/P0001  & n2639 ;
  assign n3234 = ~n3232 & ~n3233 ;
  assign n3235 = ~n2638 & n3234 ;
  assign n3236 = n3228 & ~n3235 ;
  assign n3237 = \u4_u2_buf1_reg[11]/P0001  & ~n2811 ;
  assign n3238 = \u1_u3_idin_reg[11]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n3239 = ~n2733 & n3238 ;
  assign n3240 = ~n3237 & ~n3239 ;
  assign n3241 = ~n2810 & ~n3240 ;
  assign n3242 = n2635 & n3077 ;
  assign n3243 = rst_i_pad & ~n3242 ;
  assign n3244 = ~n3241 & n3243 ;
  assign n3245 = \u4_u2_buf1_reg[15]/P0001  & ~n2811 ;
  assign n3246 = \u1_u3_idin_reg[15]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n3247 = ~n2733 & n3246 ;
  assign n3248 = ~n3245 & ~n3247 ;
  assign n3249 = ~n2810 & ~n3248 ;
  assign n3250 = n2635 & n3086 ;
  assign n3251 = rst_i_pad & ~n3250 ;
  assign n3252 = ~n3249 & n3251 ;
  assign n3253 = \u4_u2_buf1_reg[6]/P0001  & ~n2811 ;
  assign n3254 = \u1_u3_idin_reg[6]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n3255 = ~n2733 & n3254 ;
  assign n3256 = ~n3253 & ~n3255 ;
  assign n3257 = ~n2810 & ~n3256 ;
  assign n3258 = n2635 & n3095 ;
  assign n3259 = rst_i_pad & ~n3258 ;
  assign n3260 = ~n3257 & n3259 ;
  assign n3261 = \u4_u3_buf1_reg[4]/P0001  & ~n2734 ;
  assign n3262 = \u1_u3_idin_reg[4]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n3263 = ~n2733 & n3262 ;
  assign n3264 = ~n3261 & ~n3263 ;
  assign n3265 = ~n2732 & ~n3264 ;
  assign n3266 = \wb_data_i[4]_pad  & n2731 ;
  assign n3267 = n2567 & n3266 ;
  assign n3268 = rst_i_pad & ~n3267 ;
  assign n3269 = ~n3265 & n3268 ;
  assign n3270 = \u4_u3_buf1_reg[5]/P0001  & ~n2734 ;
  assign n3271 = \u1_u3_idin_reg[5]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n3272 = ~n2733 & n3271 ;
  assign n3273 = ~n3270 & ~n3272 ;
  assign n3274 = ~n2732 & ~n3273 ;
  assign n3275 = \wb_data_i[5]_pad  & n2731 ;
  assign n3276 = n2567 & n3275 ;
  assign n3277 = rst_i_pad & ~n3276 ;
  assign n3278 = ~n3274 & n3277 ;
  assign n3279 = \u4_u3_buf1_reg[7]/P0001  & ~n2734 ;
  assign n3280 = \u1_u3_idin_reg[7]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n3281 = ~n2733 & n3280 ;
  assign n3282 = ~n3279 & ~n3281 ;
  assign n3283 = ~n2732 & ~n3282 ;
  assign n3284 = \wb_data_i[7]_pad  & n2731 ;
  assign n3285 = n2567 & n3284 ;
  assign n3286 = rst_i_pad & ~n3285 ;
  assign n3287 = ~n3283 & n3286 ;
  assign n3288 = \u4_u0_buf1_reg[4]/P0001  & ~n2755 ;
  assign n3289 = \u1_u3_idin_reg[4]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n3290 = ~n2733 & n3289 ;
  assign n3291 = ~n3288 & ~n3290 ;
  assign n3292 = ~n2754 & ~n3291 ;
  assign n3293 = n2587 & n3266 ;
  assign n3294 = rst_i_pad & ~n3293 ;
  assign n3295 = ~n3292 & n3294 ;
  assign n3296 = \u4_u0_buf1_reg[5]/P0001  & ~n2755 ;
  assign n3297 = \u1_u3_idin_reg[5]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n3298 = ~n2733 & n3297 ;
  assign n3299 = ~n3296 & ~n3298 ;
  assign n3300 = ~n2754 & ~n3299 ;
  assign n3301 = n2587 & n3275 ;
  assign n3302 = rst_i_pad & ~n3301 ;
  assign n3303 = ~n3300 & n3302 ;
  assign n3304 = \u4_u0_buf1_reg[7]/P0001  & ~n2755 ;
  assign n3305 = \u1_u3_idin_reg[7]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n3306 = ~n2733 & n3305 ;
  assign n3307 = ~n3304 & ~n3306 ;
  assign n3308 = ~n2754 & ~n3307 ;
  assign n3309 = n2587 & n3284 ;
  assign n3310 = rst_i_pad & ~n3309 ;
  assign n3311 = ~n3308 & n3310 ;
  assign n3312 = \u1_u3_new_size_reg[4]/P0001  & ~\u4_csr_reg[4]/NET0131  ;
  assign n3313 = \u1_u3_new_size_reg[5]/P0001  & ~\u4_csr_reg[5]/NET0131  ;
  assign n3314 = ~n3312 & ~n3313 ;
  assign n3315 = ~\u1_u3_new_size_reg[4]/P0001  & \u4_csr_reg[4]/NET0131  ;
  assign n3316 = ~\u1_u3_new_size_reg[3]/P0001  & \u4_csr_reg[3]/P0001  ;
  assign n3317 = ~n3315 & ~n3316 ;
  assign n3318 = n3314 & ~n3317 ;
  assign n3319 = \u1_u3_new_size_reg[1]/P0001  & ~\u4_csr_reg[1]/P0001  ;
  assign n3320 = ~\u1_u3_new_size_reg[0]/P0001  & \u4_csr_reg[0]/P0001  ;
  assign n3321 = ~n3319 & n3320 ;
  assign n3322 = ~\u1_u3_new_size_reg[1]/P0001  & \u4_csr_reg[1]/P0001  ;
  assign n3323 = ~\u1_u3_new_size_reg[2]/P0001  & \u4_csr_reg[2]/NET0131  ;
  assign n3324 = ~n3322 & ~n3323 ;
  assign n3325 = ~n3321 & n3324 ;
  assign n3326 = \u1_u3_new_size_reg[3]/P0001  & ~\u4_csr_reg[3]/P0001  ;
  assign n3327 = \u1_u3_new_size_reg[2]/P0001  & ~\u4_csr_reg[2]/NET0131  ;
  assign n3328 = ~n3326 & ~n3327 ;
  assign n3329 = n3314 & n3328 ;
  assign n3330 = ~n3325 & n3329 ;
  assign n3331 = ~n3318 & ~n3330 ;
  assign n3332 = ~\u1_u3_new_size_reg[9]/P0001  & \u4_csr_reg[9]/NET0131  ;
  assign n3333 = ~\u1_u3_new_size_reg[8]/P0001  & \u4_csr_reg[8]/P0001  ;
  assign n3334 = ~n3332 & ~n3333 ;
  assign n3335 = ~\u1_u3_new_size_reg[10]/P0001  & \u4_csr_reg[10]/P0001  ;
  assign n3336 = ~\u1_u3_new_size_reg[7]/P0001  & \u4_csr_reg[7]/P0001  ;
  assign n3337 = ~n3335 & ~n3336 ;
  assign n3338 = ~\u1_u3_new_size_reg[6]/P0001  & \u4_csr_reg[6]/NET0131  ;
  assign n3339 = ~\u1_u3_new_size_reg[5]/P0001  & \u4_csr_reg[5]/NET0131  ;
  assign n3340 = ~n3338 & ~n3339 ;
  assign n3341 = n3337 & n3340 ;
  assign n3342 = n3334 & n3341 ;
  assign n3343 = n3331 & n3342 ;
  assign n3344 = \u1_u3_new_size_reg[9]/P0001  & ~\u4_csr_reg[9]/NET0131  ;
  assign n3345 = ~n3335 & n3344 ;
  assign n3346 = \u1_u3_new_size_reg[6]/P0001  & ~\u4_csr_reg[6]/NET0131  ;
  assign n3347 = ~n3336 & n3346 ;
  assign n3348 = \u1_u3_new_size_reg[7]/P0001  & ~\u4_csr_reg[7]/P0001  ;
  assign n3349 = \u1_u3_new_size_reg[8]/P0001  & ~\u4_csr_reg[8]/P0001  ;
  assign n3350 = ~n3348 & ~n3349 ;
  assign n3351 = ~n3347 & n3350 ;
  assign n3352 = n3334 & ~n3335 ;
  assign n3353 = ~n3351 & n3352 ;
  assign n3354 = ~n3345 & ~n3353 ;
  assign n3355 = \u1_u3_new_size_reg[10]/P0001  & ~\u4_csr_reg[10]/P0001  ;
  assign n3356 = ~\u1_u3_new_size_reg[11]/P0001  & ~\u1_u3_new_size_reg[12]/P0001  ;
  assign n3357 = ~\u1_u3_new_size_reg[13]/P0001  & n3356 ;
  assign n3358 = ~n3355 & n3357 ;
  assign n3359 = n3354 & n3358 ;
  assign n3360 = ~n3343 & n3359 ;
  assign n3361 = \u4_u1_buf1_reg[4]/P0001  & ~n2775 ;
  assign n3362 = \u1_u3_idin_reg[4]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n3363 = ~n2733 & n3362 ;
  assign n3364 = ~n3361 & ~n3363 ;
  assign n3365 = ~n2774 & ~n3364 ;
  assign n3366 = n2620 & n3266 ;
  assign n3367 = rst_i_pad & ~n3366 ;
  assign n3368 = ~n3365 & n3367 ;
  assign n3369 = \u4_u1_buf1_reg[5]/P0001  & ~n2775 ;
  assign n3370 = \u1_u3_idin_reg[5]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n3371 = ~n2733 & n3370 ;
  assign n3372 = ~n3369 & ~n3371 ;
  assign n3373 = ~n2774 & ~n3372 ;
  assign n3374 = n2620 & n3275 ;
  assign n3375 = rst_i_pad & ~n3374 ;
  assign n3376 = ~n3373 & n3375 ;
  assign n3377 = \u4_u1_buf1_reg[7]/P0001  & ~n2775 ;
  assign n3378 = \u1_u3_idin_reg[7]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n3379 = ~n2733 & n3378 ;
  assign n3380 = ~n3377 & ~n3379 ;
  assign n3381 = ~n2774 & ~n3380 ;
  assign n3382 = n2620 & n3284 ;
  assign n3383 = rst_i_pad & ~n3382 ;
  assign n3384 = ~n3381 & n3383 ;
  assign n3385 = \u4_u2_buf1_reg[5]/P0001  & ~n2811 ;
  assign n3386 = \u1_u3_idin_reg[5]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n3387 = ~n2733 & n3386 ;
  assign n3388 = ~n3385 & ~n3387 ;
  assign n3389 = ~n2810 & ~n3388 ;
  assign n3390 = n2635 & n3275 ;
  assign n3391 = rst_i_pad & ~n3390 ;
  assign n3392 = ~n3389 & n3391 ;
  assign n3393 = \u4_u2_buf1_reg[7]/P0001  & ~n2811 ;
  assign n3394 = \u1_u3_idin_reg[7]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n3395 = ~n2733 & n3394 ;
  assign n3396 = ~n3393 & ~n3395 ;
  assign n3397 = ~n2810 & ~n3396 ;
  assign n3398 = n2635 & n3284 ;
  assign n3399 = rst_i_pad & ~n3398 ;
  assign n3400 = ~n3397 & n3399 ;
  assign n3401 = \u4_u2_buf1_reg[4]/P0001  & ~n2811 ;
  assign n3402 = \u1_u3_idin_reg[4]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n3403 = ~n2733 & n3402 ;
  assign n3404 = ~n3401 & ~n3403 ;
  assign n3405 = ~n2810 & ~n3404 ;
  assign n3406 = n2635 & n3266 ;
  assign n3407 = rst_i_pad & ~n3406 ;
  assign n3408 = ~n3405 & n3407 ;
  assign n3409 = ~\u1_u3_new_size_reg[5]/P0001  & ~\u1_u3_new_size_reg[6]/P0001  ;
  assign n3410 = ~\u1_u3_new_size_reg[3]/P0001  & ~\u1_u3_new_size_reg[4]/P0001  ;
  assign n3411 = n3409 & n3410 ;
  assign n3412 = ~\u1_u3_new_size_reg[1]/P0001  & ~\u1_u3_new_size_reg[2]/P0001  ;
  assign n3413 = ~\u1_u3_new_size_reg[0]/P0001  & ~\u1_u3_new_size_reg[10]/P0001  ;
  assign n3414 = n3412 & n3413 ;
  assign n3415 = n3411 & n3414 ;
  assign n3416 = ~\u1_u3_new_size_reg[13]/P0001  & ~\u1_u3_new_size_reg[9]/P0001  ;
  assign n3417 = n3356 & n3416 ;
  assign n3418 = ~\u1_u3_new_size_reg[7]/P0001  & ~\u1_u3_new_size_reg[8]/P0001  ;
  assign n3419 = n3417 & n3418 ;
  assign n3420 = n3415 & n3419 ;
  assign n3421 = ~\u1_u2_sizd_c_reg[12]/P0001  & ~\u1_u2_tx_dma_en_r_reg/P0001  ;
  assign n3422 = \u1_u2_mack_r_reg/P0001  & \u1_u2_state_reg[5]/NET0131  ;
  assign n3423 = ~\u1_u2_sizd_c_reg[0]/P0001  & n3422 ;
  assign n3424 = ~\u1_u2_sizd_c_reg[1]/P0001  & ~\u1_u2_sizd_c_reg[2]/P0001  ;
  assign n3425 = ~\u1_u2_sizd_c_reg[3]/P0001  & ~\u1_u2_sizd_c_reg[4]/P0001  ;
  assign n3426 = n3424 & n3425 ;
  assign n3427 = ~\u1_u2_sizd_c_reg[5]/P0001  & ~\u1_u2_sizd_c_reg[6]/P0001  ;
  assign n3428 = n3426 & n3427 ;
  assign n3429 = n3423 & n3428 ;
  assign n3430 = ~\u1_u2_sizd_c_reg[7]/P0001  & ~\u1_u2_sizd_c_reg[8]/P0001  ;
  assign n3431 = n3427 & n3430 ;
  assign n3432 = n3426 & n3431 ;
  assign n3433 = ~\u1_u2_sizd_c_reg[10]/P0001  & ~\u1_u2_sizd_c_reg[11]/P0001  ;
  assign n3434 = ~\u1_u2_sizd_c_reg[12]/P0001  & ~\u1_u2_sizd_c_reg[13]/P0001  ;
  assign n3435 = ~\u1_u2_sizd_c_reg[9]/P0001  & n3434 ;
  assign n3436 = n3433 & n3435 ;
  assign n3437 = n3432 & n3436 ;
  assign n3438 = \u1_u1_state_reg[1]/NET0131  & ~\u1_u2_sizd_c_reg[0]/P0001  ;
  assign n3439 = n1756 & n3438 ;
  assign n3440 = n3428 & n3439 ;
  assign n3441 = ~n3437 & n3440 ;
  assign n3442 = ~n3429 & ~n3441 ;
  assign n3443 = ~\u1_u2_sizd_c_reg[9]/P0001  & n3430 ;
  assign n3444 = n3433 & n3443 ;
  assign n3445 = ~n3442 & n3444 ;
  assign n3446 = ~\u1_u0_pid_reg[0]/NET0131  & ~\u1_u0_pid_reg[1]/NET0131  ;
  assign n3447 = n2378 & n3446 ;
  assign n3448 = \u0_u0_mode_hs_reg/P0001  & n3447 ;
  assign n3449 = ~n2360 & ~n3448 ;
  assign n3450 = ~n2367 & n3449 ;
  assign n3451 = ~n2359 & n3450 ;
  assign n3452 = ~\u1_u3_state_reg[1]/P0001  & n2376 ;
  assign n3453 = \u1_u3_match_r_reg/P0001  & ~n2383 ;
  assign n3454 = ~n2379 & n3453 ;
  assign n3455 = ~n2382 & n3454 ;
  assign n3456 = ~\u4_csr_reg[26]/NET0131  & ~n2352 ;
  assign n3457 = ~\u4_csr_reg[27]/NET0131  & ~n3456 ;
  assign n3458 = n3455 & n3457 ;
  assign n3459 = n3452 & n3458 ;
  assign n3460 = n3451 & n3459 ;
  assign n3461 = n3445 & ~n3460 ;
  assign n3462 = n3421 & n3461 ;
  assign n3463 = \u1_u2_sizd_c_reg[12]/P0001  & ~\u1_u2_tx_dma_en_r_reg/P0001  ;
  assign n3464 = ~n3460 & n3463 ;
  assign n3465 = ~n3445 & n3464 ;
  assign n3466 = rst_i_pad & ~n3465 ;
  assign n3467 = ~n3462 & n3466 ;
  assign n3468 = ~\u1_u2_tx_dma_en_r_reg/P0001  & ~n3460 ;
  assign n3469 = \u4_buf1_reg[18]/P0001  & n2793 ;
  assign n3470 = \u4_buf1_reg[18]/P0001  & ~n2789 ;
  assign n3471 = n2788 & n3470 ;
  assign n3472 = ~n3469 & ~n3471 ;
  assign n3473 = \u4_buf0_reg[18]/P0001  & ~n2793 ;
  assign n3474 = ~n2794 & n3473 ;
  assign n3475 = n3472 & ~n3474 ;
  assign n3476 = \u4_csr_reg[1]/P0001  & n3475 ;
  assign n3477 = \u4_buf1_reg[17]/NET0131  & n2793 ;
  assign n3478 = \u4_buf1_reg[17]/NET0131  & ~n2789 ;
  assign n3479 = n2788 & n3478 ;
  assign n3480 = ~n3477 & ~n3479 ;
  assign n3481 = \u4_buf0_reg[17]/NET0131  & ~n2793 ;
  assign n3482 = ~n2794 & n3481 ;
  assign n3483 = n3480 & ~n3482 ;
  assign n3484 = \u4_csr_reg[0]/P0001  & n3483 ;
  assign n3485 = ~n3476 & ~n3484 ;
  assign n3486 = ~\u4_csr_reg[1]/P0001  & ~n3475 ;
  assign n3487 = \u4_buf1_reg[19]/NET0131  & n2793 ;
  assign n3488 = \u4_buf1_reg[19]/NET0131  & ~n2789 ;
  assign n3489 = n2788 & n3488 ;
  assign n3490 = ~n3487 & ~n3489 ;
  assign n3491 = \u4_buf0_reg[19]/NET0131  & ~n2793 ;
  assign n3492 = ~n2794 & n3491 ;
  assign n3493 = n3490 & ~n3492 ;
  assign n3494 = ~\u4_csr_reg[2]/NET0131  & ~n3493 ;
  assign n3495 = ~n3486 & ~n3494 ;
  assign n3496 = ~n3485 & n3495 ;
  assign n3497 = \u4_buf1_reg[21]/NET0131  & n2793 ;
  assign n3498 = \u4_buf1_reg[21]/NET0131  & ~n2789 ;
  assign n3499 = n2788 & n3498 ;
  assign n3500 = ~n3497 & ~n3499 ;
  assign n3501 = \u4_buf0_reg[21]/NET0131  & ~n2793 ;
  assign n3502 = ~n2794 & n3501 ;
  assign n3503 = n3500 & ~n3502 ;
  assign n3504 = \u4_csr_reg[4]/NET0131  & n3503 ;
  assign n3505 = \u4_buf1_reg[20]/NET0131  & n2793 ;
  assign n3506 = \u4_buf1_reg[20]/NET0131  & ~n2789 ;
  assign n3507 = n2788 & n3506 ;
  assign n3508 = ~n3505 & ~n3507 ;
  assign n3509 = \u4_buf0_reg[20]/NET0131  & ~n2793 ;
  assign n3510 = ~n2794 & n3509 ;
  assign n3511 = n3508 & ~n3510 ;
  assign n3512 = \u4_csr_reg[3]/P0001  & n3511 ;
  assign n3513 = ~n3504 & ~n3512 ;
  assign n3514 = \u4_csr_reg[2]/NET0131  & n3493 ;
  assign n3515 = n3513 & ~n3514 ;
  assign n3516 = ~n3496 & n3515 ;
  assign n3517 = ~\u4_csr_reg[3]/P0001  & ~n3511 ;
  assign n3518 = ~n3504 & n3517 ;
  assign n3519 = \u4_buf1_reg[22]/NET0131  & n2793 ;
  assign n3520 = \u4_buf1_reg[22]/NET0131  & ~n2789 ;
  assign n3521 = n2788 & n3520 ;
  assign n3522 = ~n3519 & ~n3521 ;
  assign n3523 = \u4_buf0_reg[22]/NET0131  & ~n2793 ;
  assign n3524 = ~n2794 & n3523 ;
  assign n3525 = n3522 & ~n3524 ;
  assign n3526 = ~\u4_csr_reg[5]/NET0131  & ~n3525 ;
  assign n3527 = ~\u4_csr_reg[4]/NET0131  & ~n3503 ;
  assign n3528 = ~n3526 & ~n3527 ;
  assign n3529 = ~n3518 & n3528 ;
  assign n3530 = ~n3516 & n3529 ;
  assign n3531 = \u4_csr_reg[5]/NET0131  & n3525 ;
  assign n3532 = \u4_buf1_reg[24]/NET0131  & n2793 ;
  assign n3533 = \u4_buf1_reg[24]/NET0131  & ~n2789 ;
  assign n3534 = n2788 & n3533 ;
  assign n3535 = ~n3532 & ~n3534 ;
  assign n3536 = \u4_buf0_reg[24]/NET0131  & ~n2793 ;
  assign n3537 = ~n2794 & n3536 ;
  assign n3538 = n3535 & ~n3537 ;
  assign n3539 = \u4_csr_reg[7]/P0001  & n3538 ;
  assign n3540 = \u4_buf1_reg[25]/NET0131  & n2793 ;
  assign n3541 = \u4_buf1_reg[25]/NET0131  & ~n2789 ;
  assign n3542 = n2788 & n3541 ;
  assign n3543 = ~n3540 & ~n3542 ;
  assign n3544 = \u4_buf0_reg[25]/NET0131  & ~n2793 ;
  assign n3545 = ~n2794 & n3544 ;
  assign n3546 = n3543 & ~n3545 ;
  assign n3547 = \u4_csr_reg[8]/P0001  & n3546 ;
  assign n3548 = ~n3539 & ~n3547 ;
  assign n3549 = \u4_buf1_reg[27]/P0001  & n2793 ;
  assign n3550 = \u4_buf1_reg[27]/P0001  & ~n2789 ;
  assign n3551 = n2788 & n3550 ;
  assign n3552 = ~n3549 & ~n3551 ;
  assign n3553 = \u4_buf0_reg[27]/P0001  & ~n2793 ;
  assign n3554 = ~n2794 & n3553 ;
  assign n3555 = n3552 & ~n3554 ;
  assign n3556 = \u4_csr_reg[10]/P0001  & n3555 ;
  assign n3557 = \u4_buf1_reg[26]/NET0131  & n2793 ;
  assign n3558 = \u4_buf1_reg[26]/NET0131  & ~n2789 ;
  assign n3559 = n2788 & n3558 ;
  assign n3560 = ~n3557 & ~n3559 ;
  assign n3561 = \u4_buf0_reg[26]/NET0131  & ~n2793 ;
  assign n3562 = ~n2794 & n3561 ;
  assign n3563 = n3560 & ~n3562 ;
  assign n3564 = \u4_csr_reg[9]/NET0131  & n3563 ;
  assign n3565 = ~n3556 & ~n3564 ;
  assign n3566 = \u4_buf1_reg[23]/NET0131  & n2793 ;
  assign n3567 = \u4_buf1_reg[23]/NET0131  & ~n2789 ;
  assign n3568 = n2788 & n3567 ;
  assign n3569 = ~n3566 & ~n3568 ;
  assign n3570 = \u4_buf0_reg[23]/NET0131  & ~n2793 ;
  assign n3571 = ~n2794 & n3570 ;
  assign n3572 = n3569 & ~n3571 ;
  assign n3573 = \u4_csr_reg[6]/NET0131  & n3572 ;
  assign n3574 = n3565 & ~n3573 ;
  assign n3575 = n3548 & n3574 ;
  assign n3576 = ~n3531 & n3575 ;
  assign n3577 = ~n3530 & n3576 ;
  assign n3578 = ~\u4_csr_reg[7]/P0001  & ~n3538 ;
  assign n3579 = ~\u4_csr_reg[6]/NET0131  & ~n3572 ;
  assign n3580 = ~n3578 & ~n3579 ;
  assign n3581 = n3548 & ~n3580 ;
  assign n3582 = ~\u4_csr_reg[9]/NET0131  & ~n3563 ;
  assign n3583 = ~\u4_csr_reg[8]/P0001  & ~n3546 ;
  assign n3584 = ~n3582 & ~n3583 ;
  assign n3585 = ~n3581 & n3584 ;
  assign n3586 = n3565 & ~n3585 ;
  assign n3587 = ~\u4_csr_reg[10]/P0001  & ~n3555 ;
  assign n3588 = \u4_buf1_reg[29]/P0001  & n2793 ;
  assign n3589 = \u4_buf1_reg[29]/P0001  & ~n2789 ;
  assign n3590 = n2788 & n3589 ;
  assign n3591 = ~n3588 & ~n3590 ;
  assign n3592 = \u4_buf0_reg[29]/P0001  & ~n2793 ;
  assign n3593 = ~n2794 & n3592 ;
  assign n3594 = n3591 & ~n3593 ;
  assign n3595 = \u4_buf1_reg[28]/P0001  & n2793 ;
  assign n3596 = \u4_buf1_reg[28]/P0001  & ~n2789 ;
  assign n3597 = n2788 & n3596 ;
  assign n3598 = ~n3595 & ~n3597 ;
  assign n3599 = \u4_buf0_reg[28]/P0001  & ~n2793 ;
  assign n3600 = ~n2794 & n3599 ;
  assign n3601 = n3598 & ~n3600 ;
  assign n3602 = n3594 & n3601 ;
  assign n3603 = \u4_buf1_reg[30]/P0001  & n2793 ;
  assign n3604 = \u4_buf1_reg[30]/P0001  & ~n2789 ;
  assign n3605 = n2788 & n3604 ;
  assign n3606 = ~n3603 & ~n3605 ;
  assign n3607 = \u4_buf0_reg[30]/P0001  & ~n2793 ;
  assign n3608 = ~n2794 & n3607 ;
  assign n3609 = n3606 & ~n3608 ;
  assign n3610 = n3602 & n3609 ;
  assign n3611 = ~n3587 & n3610 ;
  assign n3612 = ~n3483 & n3611 ;
  assign n3613 = ~n3586 & n3612 ;
  assign n3614 = ~n3577 & n3613 ;
  assign n3615 = ~n3468 & n3614 ;
  assign n3616 = ~n3586 & n3611 ;
  assign n3617 = ~n3577 & n3616 ;
  assign n3618 = \u4_csr_reg[0]/P0001  & ~n3468 ;
  assign n3619 = ~n3617 & n3618 ;
  assign n3620 = ~n3615 & ~n3619 ;
  assign n3621 = ~\u1_u2_sizd_c_reg[0]/P0001  & ~n3422 ;
  assign n3622 = n3437 & n3621 ;
  assign n3623 = ~n1757 & n3621 ;
  assign n3624 = \u1_u1_state_reg[1]/NET0131  & \u1_u2_sizd_c_reg[0]/P0001  ;
  assign n3625 = n1756 & n3624 ;
  assign n3626 = \u1_u2_sizd_c_reg[0]/P0001  & n3422 ;
  assign n3627 = ~n3625 & ~n3626 ;
  assign n3628 = ~n3623 & n3627 ;
  assign n3629 = ~n3622 & n3628 ;
  assign n3630 = ~\u1_u2_tx_dma_en_r_reg/P0001  & n3629 ;
  assign n3631 = ~n3460 & n3630 ;
  assign n3632 = rst_i_pad & ~n3631 ;
  assign n3633 = n3620 & n3632 ;
  assign n3634 = n3555 & n3609 ;
  assign n3635 = n3602 & n3634 ;
  assign n3636 = ~n3577 & n3635 ;
  assign n3637 = \u4_csr_reg[10]/P0001  & ~n3468 ;
  assign n3638 = ~n3636 & n3637 ;
  assign n3639 = rst_i_pad & ~n3468 ;
  assign n3640 = rst_i_pad & \u1_u2_sizd_c_reg[10]/P0001  ;
  assign n3641 = n3443 & n3640 ;
  assign n3642 = ~n3442 & n3641 ;
  assign n3643 = ~n3442 & n3443 ;
  assign n3644 = rst_i_pad & ~\u1_u2_sizd_c_reg[10]/P0001  ;
  assign n3645 = ~n3643 & n3644 ;
  assign n3646 = ~n3642 & ~n3645 ;
  assign n3647 = ~n3639 & n3646 ;
  assign n3648 = ~n3638 & ~n3647 ;
  assign n3649 = ~\u1_u2_sizd_c_reg[10]/P0001  & ~\u1_u2_sizd_c_reg[9]/P0001  ;
  assign n3650 = n3430 & n3649 ;
  assign n3651 = ~n3442 & n3650 ;
  assign n3652 = rst_i_pad & ~\u1_u2_sizd_c_reg[11]/P0001  ;
  assign n3653 = ~n3651 & n3652 ;
  assign n3654 = rst_i_pad & \u1_u2_sizd_c_reg[11]/P0001  ;
  assign n3655 = n3651 & n3654 ;
  assign n3656 = ~n3653 & ~n3655 ;
  assign n3657 = ~n3639 & n3656 ;
  assign n3658 = ~\u1_u2_sizd_c_reg[11]/P0001  & ~\u1_u2_sizd_c_reg[13]/P0001  ;
  assign n3659 = ~\u1_u2_sizd_c_reg[12]/P0001  & n3658 ;
  assign n3660 = n3651 & n3659 ;
  assign n3661 = n3468 & n3660 ;
  assign n3662 = ~\u1_u2_sizd_c_reg[11]/P0001  & ~\u1_u2_sizd_c_reg[12]/P0001  ;
  assign n3663 = n3651 & n3662 ;
  assign n3664 = \u1_u2_sizd_c_reg[13]/P0001  & ~\u1_u2_tx_dma_en_r_reg/P0001  ;
  assign n3665 = ~n3460 & n3664 ;
  assign n3666 = ~n3663 & n3665 ;
  assign n3667 = rst_i_pad & ~n3666 ;
  assign n3668 = ~n3661 & n3667 ;
  assign n3669 = ~n3493 & n3611 ;
  assign n3670 = ~n3586 & n3669 ;
  assign n3671 = ~n3577 & n3670 ;
  assign n3672 = ~n3468 & n3671 ;
  assign n3673 = \u4_csr_reg[2]/NET0131  & ~n3468 ;
  assign n3674 = ~n3617 & n3673 ;
  assign n3675 = ~n3672 & ~n3674 ;
  assign n3676 = ~\u1_u2_sizd_c_reg[1]/P0001  & n3423 ;
  assign n3677 = ~\u1_u2_sizd_c_reg[1]/P0001  & n3439 ;
  assign n3678 = ~n3437 & n3677 ;
  assign n3679 = ~n3676 & ~n3678 ;
  assign n3680 = \u1_u2_sizd_c_reg[2]/P0001  & n3679 ;
  assign n3681 = n3423 & n3424 ;
  assign n3682 = n3424 & n3439 ;
  assign n3683 = ~n3437 & n3682 ;
  assign n3684 = ~n3681 & ~n3683 ;
  assign n3685 = ~n3680 & n3684 ;
  assign n3686 = n3468 & ~n3685 ;
  assign n3687 = rst_i_pad & ~n3686 ;
  assign n3688 = n3675 & n3687 ;
  assign n3689 = ~n3511 & n3611 ;
  assign n3690 = ~n3586 & n3689 ;
  assign n3691 = ~n3577 & n3690 ;
  assign n3692 = ~n3468 & n3691 ;
  assign n3693 = \u4_csr_reg[3]/P0001  & ~n3468 ;
  assign n3694 = ~n3617 & n3693 ;
  assign n3695 = ~n3692 & ~n3694 ;
  assign n3696 = \u1_u2_sizd_c_reg[3]/P0001  & n3684 ;
  assign n3697 = ~\u1_u2_sizd_c_reg[3]/P0001  & ~n3684 ;
  assign n3698 = ~n3696 & ~n3697 ;
  assign n3699 = n3468 & ~n3698 ;
  assign n3700 = rst_i_pad & ~n3699 ;
  assign n3701 = n3695 & n3700 ;
  assign n3702 = ~n3503 & n3611 ;
  assign n3703 = ~n3586 & n3702 ;
  assign n3704 = ~n3577 & n3703 ;
  assign n3705 = ~n3468 & n3704 ;
  assign n3706 = \u4_csr_reg[4]/NET0131  & ~n3468 ;
  assign n3707 = ~n3617 & n3706 ;
  assign n3708 = ~n3705 & ~n3707 ;
  assign n3709 = \u1_u2_sizd_c_reg[4]/P0001  & ~n3697 ;
  assign n3710 = n3423 & n3426 ;
  assign n3711 = n3426 & n3439 ;
  assign n3712 = ~n3437 & n3711 ;
  assign n3713 = ~n3710 & ~n3712 ;
  assign n3714 = rst_i_pad & n3713 ;
  assign n3715 = ~n3709 & n3714 ;
  assign n3716 = ~n3639 & ~n3715 ;
  assign n3717 = n3708 & ~n3716 ;
  assign n3718 = ~n3525 & n3611 ;
  assign n3719 = ~n3586 & n3718 ;
  assign n3720 = ~n3577 & n3719 ;
  assign n3721 = ~n3468 & n3720 ;
  assign n3722 = \u4_csr_reg[5]/NET0131  & ~n3468 ;
  assign n3723 = ~n3617 & n3722 ;
  assign n3724 = ~n3721 & ~n3723 ;
  assign n3725 = ~\u1_u2_sizd_c_reg[5]/P0001  & ~n3713 ;
  assign n3726 = \u1_u2_sizd_c_reg[5]/P0001  & n3713 ;
  assign n3727 = ~n3725 & ~n3726 ;
  assign n3728 = n3468 & ~n3727 ;
  assign n3729 = rst_i_pad & ~n3728 ;
  assign n3730 = n3724 & n3729 ;
  assign n3731 = ~n3572 & n3611 ;
  assign n3732 = ~n3586 & n3731 ;
  assign n3733 = ~n3577 & n3732 ;
  assign n3734 = ~n3468 & n3733 ;
  assign n3735 = \u4_csr_reg[6]/NET0131  & ~n3468 ;
  assign n3736 = ~n3617 & n3735 ;
  assign n3737 = ~n3734 & ~n3736 ;
  assign n3738 = \u1_u2_sizd_c_reg[6]/P0001  & ~n3725 ;
  assign n3739 = rst_i_pad & n3442 ;
  assign n3740 = ~n3738 & n3739 ;
  assign n3741 = ~n3639 & ~n3740 ;
  assign n3742 = n3737 & ~n3741 ;
  assign n3743 = ~n3538 & n3611 ;
  assign n3744 = ~n3586 & n3743 ;
  assign n3745 = ~n3577 & n3744 ;
  assign n3746 = ~n3468 & n3745 ;
  assign n3747 = \u4_csr_reg[7]/P0001  & ~n3468 ;
  assign n3748 = ~n3617 & n3747 ;
  assign n3749 = ~n3746 & ~n3748 ;
  assign n3750 = ~\u1_u2_sizd_c_reg[7]/P0001  & ~n3442 ;
  assign n3751 = \u1_u2_sizd_c_reg[7]/P0001  & n3442 ;
  assign n3752 = ~n3750 & ~n3751 ;
  assign n3753 = n3468 & ~n3752 ;
  assign n3754 = rst_i_pad & ~n3753 ;
  assign n3755 = n3749 & n3754 ;
  assign n3756 = ~n3546 & n3611 ;
  assign n3757 = ~n3586 & n3756 ;
  assign n3758 = ~n3577 & n3757 ;
  assign n3759 = ~n3468 & n3758 ;
  assign n3760 = \u4_csr_reg[8]/P0001  & ~n3468 ;
  assign n3761 = ~n3617 & n3760 ;
  assign n3762 = ~n3759 & ~n3761 ;
  assign n3763 = \u1_u2_sizd_c_reg[8]/P0001  & ~n3750 ;
  assign n3764 = n3430 & ~n3442 ;
  assign n3765 = rst_i_pad & ~n3764 ;
  assign n3766 = ~n3763 & n3765 ;
  assign n3767 = ~n3639 & ~n3766 ;
  assign n3768 = n3762 & ~n3767 ;
  assign n3769 = ~n3563 & n3611 ;
  assign n3770 = ~n3586 & n3769 ;
  assign n3771 = ~n3577 & n3770 ;
  assign n3772 = ~n3468 & n3771 ;
  assign n3773 = \u4_csr_reg[9]/NET0131  & ~n3468 ;
  assign n3774 = ~n3617 & n3773 ;
  assign n3775 = ~n3772 & ~n3774 ;
  assign n3776 = n3423 & n3432 ;
  assign n3777 = ~n3436 & n3439 ;
  assign n3778 = n3432 & n3777 ;
  assign n3779 = ~n3776 & ~n3778 ;
  assign n3780 = ~\u1_u2_sizd_c_reg[9]/P0001  & ~n3779 ;
  assign n3781 = \u1_u2_sizd_c_reg[9]/P0001  & n3779 ;
  assign n3782 = ~n3780 & ~n3781 ;
  assign n3783 = n3468 & ~n3782 ;
  assign n3784 = rst_i_pad & ~n3783 ;
  assign n3785 = n3775 & n3784 ;
  assign n3786 = \u1_u1_crc16_reg[2]/P0001  & ~\u1_u1_zero_length_r_reg/P0001  ;
  assign n3787 = n2283 & n3786 ;
  assign n3788 = \u1_u1_crc16_reg[2]/P0001  & \u1_u1_state_reg[1]/NET0131  ;
  assign n3789 = n1756 & n3788 ;
  assign n3790 = n1860 & n3789 ;
  assign n3791 = ~n3787 & ~n3790 ;
  assign n3792 = \u1_u1_crc16_reg[10]/P0001  & ~n2284 ;
  assign n3793 = ~n2294 & ~n3792 ;
  assign n3794 = n1757 & ~n2294 ;
  assign n3795 = n1860 & n3794 ;
  assign n3796 = ~n3793 & ~n3795 ;
  assign n3797 = n3791 & ~n3796 ;
  assign n3798 = \u1_u1_crc16_reg[3]/P0001  & n2284 ;
  assign n3799 = \u1_u1_crc16_reg[3]/P0001  & n1757 ;
  assign n3800 = n1860 & n3799 ;
  assign n3801 = ~n3798 & ~n3800 ;
  assign n3802 = \u1_u1_crc16_reg[11]/P0001  & ~n2284 ;
  assign n3803 = ~n2282 & n3802 ;
  assign n3804 = ~n2294 & ~n3803 ;
  assign n3805 = n3801 & n3804 ;
  assign n3806 = \u1_u1_crc16_reg[4]/P0001  & n2284 ;
  assign n3807 = \u1_u1_crc16_reg[4]/P0001  & n1757 ;
  assign n3808 = n1860 & n3807 ;
  assign n3809 = ~n3806 & ~n3808 ;
  assign n3810 = \u1_u1_crc16_reg[12]/P0001  & ~n2284 ;
  assign n3811 = ~n2282 & n3810 ;
  assign n3812 = ~n2294 & ~n3811 ;
  assign n3813 = n3809 & n3812 ;
  assign n3814 = \u1_u1_crc16_reg[5]/P0001  & n2284 ;
  assign n3815 = \u1_u1_crc16_reg[5]/P0001  & n1757 ;
  assign n3816 = n1860 & n3815 ;
  assign n3817 = ~n3814 & ~n3816 ;
  assign n3818 = \u1_u1_crc16_reg[13]/P0001  & ~n2284 ;
  assign n3819 = ~n2282 & n3818 ;
  assign n3820 = ~n2294 & ~n3819 ;
  assign n3821 = n3817 & n3820 ;
  assign n3822 = \u1_u1_crc16_reg[6]/P0001  & n2284 ;
  assign n3823 = \u1_u1_crc16_reg[6]/P0001  & n1757 ;
  assign n3824 = n1860 & n3823 ;
  assign n3825 = ~n3822 & ~n3824 ;
  assign n3826 = \u1_u1_crc16_reg[14]/P0001  & ~n2284 ;
  assign n3827 = ~n2282 & n3826 ;
  assign n3828 = ~n2294 & ~n3827 ;
  assign n3829 = n3825 & n3828 ;
  assign n3830 = \u4_csr_reg[15]/NET0131  & \u4_csr_reg[8]/P0001  ;
  assign n3831 = n2363 & n3830 ;
  assign n3832 = ~\u1_u3_adr_r_reg[8]/P0001  & ~n3831 ;
  assign n3833 = \u4_csr_reg[15]/NET0131  & ~\u4_csr_reg[26]/NET0131  ;
  assign n3834 = \u1_u2_sizu_c_reg[8]/NET0131  & \u4_csr_reg[27]/NET0131  ;
  assign n3835 = ~n3833 & n3834 ;
  assign n3836 = \u1_u2_sizu_c_reg[8]/NET0131  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3837 = n3033 & n3836 ;
  assign n3838 = ~n3835 & ~n3837 ;
  assign n3839 = \u1_u3_in_token_reg/NET0131  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3840 = ~n2361 & ~n3839 ;
  assign n3841 = \u1_u3_size_next_r_reg[8]/P0001  & ~n3840 ;
  assign n3842 = n3838 & ~n3841 ;
  assign n3843 = n3832 & n3842 ;
  assign n3844 = \u1_u2_sizu_c_reg[9]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n3845 = ~n3833 & n3844 ;
  assign n3846 = \u1_u2_sizu_c_reg[9]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3847 = n3033 & n3846 ;
  assign n3848 = ~n3845 & ~n3847 ;
  assign n3849 = \u1_u3_size_next_r_reg[9]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3850 = ~n3033 & n3849 ;
  assign n3851 = \u4_csr_reg[15]/NET0131  & \u4_csr_reg[9]/NET0131  ;
  assign n3852 = n2363 & n3851 ;
  assign n3853 = ~\u1_u3_adr_r_reg[9]/P0001  & ~n3852 ;
  assign n3854 = ~n3850 & n3853 ;
  assign n3855 = n3848 & n3854 ;
  assign n3856 = ~n3843 & ~n3855 ;
  assign n3857 = \u1_u2_sizu_c_reg[7]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n3858 = ~n3833 & n3857 ;
  assign n3859 = \u1_u2_sizu_c_reg[7]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3860 = n3033 & n3859 ;
  assign n3861 = ~n3858 & ~n3860 ;
  assign n3862 = \u1_u3_size_next_r_reg[7]/P0001  & ~n3840 ;
  assign n3863 = \u4_csr_reg[15]/NET0131  & \u4_csr_reg[7]/P0001  ;
  assign n3864 = n2363 & n3863 ;
  assign n3865 = ~\u1_u3_adr_r_reg[7]/P0001  & ~n3864 ;
  assign n3866 = ~n3862 & n3865 ;
  assign n3867 = n3861 & n3866 ;
  assign n3868 = \u1_u2_sizu_c_reg[6]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n3869 = ~n3833 & n3868 ;
  assign n3870 = \u1_u2_sizu_c_reg[6]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3871 = n3033 & n3870 ;
  assign n3872 = ~n3869 & ~n3871 ;
  assign n3873 = \u1_u3_size_next_r_reg[6]/P0001  & ~n3840 ;
  assign n3874 = \u4_csr_reg[15]/NET0131  & \u4_csr_reg[6]/NET0131  ;
  assign n3875 = n2363 & n3874 ;
  assign n3876 = ~n3873 & ~n3875 ;
  assign n3877 = n3872 & n3876 ;
  assign n3878 = \u1_u3_adr_r_reg[6]/P0001  & ~n3877 ;
  assign n3879 = ~n3867 & n3878 ;
  assign n3880 = ~n3831 & n3842 ;
  assign n3881 = \u1_u3_adr_r_reg[8]/P0001  & ~n3880 ;
  assign n3882 = ~n3862 & ~n3864 ;
  assign n3883 = n3861 & n3882 ;
  assign n3884 = \u1_u3_adr_r_reg[7]/P0001  & ~n3883 ;
  assign n3885 = ~n3881 & ~n3884 ;
  assign n3886 = ~n3879 & n3885 ;
  assign n3887 = n3856 & ~n3886 ;
  assign n3888 = \u4_csr_reg[10]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n3889 = n3833 & n3888 ;
  assign n3890 = \u1_u3_adr_r_reg[10]/P0001  & n3889 ;
  assign n3891 = \u1_u3_size_next_r_reg[10]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3892 = ~n3033 & n3891 ;
  assign n3893 = \u1_u2_sizu_c_reg[10]/P0001  & ~n3036 ;
  assign n3894 = ~n3892 & ~n3893 ;
  assign n3895 = \u4_csr_reg[27]/NET0131  & n3833 ;
  assign n3896 = \u1_u3_adr_r_reg[10]/P0001  & ~n3895 ;
  assign n3897 = ~n3894 & n3896 ;
  assign n3898 = ~n3890 & ~n3897 ;
  assign n3899 = ~n3850 & ~n3852 ;
  assign n3900 = n3848 & n3899 ;
  assign n3901 = \u1_u3_adr_r_reg[9]/P0001  & ~n3900 ;
  assign n3902 = n3898 & ~n3901 ;
  assign n3903 = ~n3887 & n3902 ;
  assign n3904 = ~n3894 & ~n3895 ;
  assign n3905 = ~\u1_u3_adr_r_reg[10]/P0001  & ~n3889 ;
  assign n3906 = ~n3904 & n3905 ;
  assign n3907 = ~n3903 & ~n3906 ;
  assign n3908 = \u1_u3_size_next_r_reg[5]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3909 = ~n3033 & n3908 ;
  assign n3910 = \u1_u2_sizu_c_reg[5]/P0001  & ~n3036 ;
  assign n3911 = ~n3909 & ~n3910 ;
  assign n3912 = ~n3895 & ~n3911 ;
  assign n3913 = \u4_csr_reg[15]/NET0131  & \u4_csr_reg[5]/NET0131  ;
  assign n3914 = n2363 & n3913 ;
  assign n3915 = ~\u1_u3_adr_r_reg[5]/P0001  & ~n3914 ;
  assign n3916 = ~n3912 & n3915 ;
  assign n3917 = \u1_u2_sizu_c_reg[4]/P0001  & ~n3036 ;
  assign n3918 = \u1_u3_size_next_r_reg[4]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3919 = ~n3033 & n3918 ;
  assign n3920 = ~n3917 & ~n3919 ;
  assign n3921 = ~n3895 & ~n3920 ;
  assign n3922 = \u4_csr_reg[15]/NET0131  & \u4_csr_reg[4]/NET0131  ;
  assign n3923 = n2363 & n3922 ;
  assign n3924 = ~\u1_u3_adr_r_reg[4]/P0001  & ~n3923 ;
  assign n3925 = ~n3921 & n3924 ;
  assign n3926 = ~n3916 & ~n3925 ;
  assign n3927 = \u4_csr_reg[15]/NET0131  & \u4_csr_reg[3]/P0001  ;
  assign n3928 = n2363 & n3927 ;
  assign n3929 = \u1_u3_adr_r_reg[3]/P0001  & n3928 ;
  assign n3930 = \u1_u3_size_next_r_reg[3]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3931 = ~n3033 & n3930 ;
  assign n3932 = \u1_u2_sizu_c_reg[3]/P0001  & ~n3036 ;
  assign n3933 = ~n3931 & ~n3932 ;
  assign n3934 = \u1_u3_adr_r_reg[3]/P0001  & ~n3895 ;
  assign n3935 = ~n3933 & n3934 ;
  assign n3936 = ~n3929 & ~n3935 ;
  assign n3937 = ~n3895 & ~n3933 ;
  assign n3938 = ~\u1_u3_adr_r_reg[3]/P0001  & ~n3928 ;
  assign n3939 = ~n3937 & n3938 ;
  assign n3940 = \u4_csr_reg[15]/NET0131  & \u4_csr_reg[2]/NET0131  ;
  assign n3941 = n2363 & n3940 ;
  assign n3942 = \u1_u3_adr_r_reg[2]/P0001  & n3941 ;
  assign n3943 = \u1_u3_size_next_r_reg[2]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3944 = ~n3033 & n3943 ;
  assign n3945 = \u1_u2_sizu_c_reg[2]/P0001  & ~n3036 ;
  assign n3946 = ~n3944 & ~n3945 ;
  assign n3947 = \u1_u3_adr_r_reg[2]/P0001  & ~n3895 ;
  assign n3948 = ~n3946 & n3947 ;
  assign n3949 = ~n3942 & ~n3948 ;
  assign n3950 = ~n3939 & ~n3949 ;
  assign n3951 = n3936 & ~n3950 ;
  assign n3952 = n3926 & ~n3951 ;
  assign n3953 = \u4_csr_reg[15]/NET0131  & \u4_csr_reg[1]/P0001  ;
  assign n3954 = n2363 & n3953 ;
  assign n3955 = \u1_u3_adr_r_reg[1]/P0001  & n3954 ;
  assign n3956 = \u1_u3_size_next_r_reg[1]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3957 = ~n3033 & n3956 ;
  assign n3958 = \u1_u2_sizu_c_reg[1]/P0001  & ~n3036 ;
  assign n3959 = ~n3957 & ~n3958 ;
  assign n3960 = \u1_u3_adr_r_reg[1]/P0001  & ~n3895 ;
  assign n3961 = ~n3959 & n3960 ;
  assign n3962 = ~n3955 & ~n3961 ;
  assign n3963 = ~n3895 & ~n3959 ;
  assign n3964 = ~\u1_u3_adr_r_reg[1]/P0001  & ~n3954 ;
  assign n3965 = ~n3963 & n3964 ;
  assign n3966 = \u4_csr_reg[0]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n3967 = n3833 & n3966 ;
  assign n3968 = \u1_u3_adr_r_reg[0]/P0001  & n3967 ;
  assign n3969 = \u1_u3_size_next_r_reg[0]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n3970 = ~n3033 & n3969 ;
  assign n3971 = \u1_u2_sizu_c_reg[0]/P0001  & ~n3036 ;
  assign n3972 = ~n3970 & ~n3971 ;
  assign n3973 = \u1_u3_adr_r_reg[0]/P0001  & ~n3895 ;
  assign n3974 = ~n3972 & n3973 ;
  assign n3975 = ~n3968 & ~n3974 ;
  assign n3976 = ~n3965 & ~n3975 ;
  assign n3977 = n3962 & ~n3976 ;
  assign n3978 = ~n3895 & ~n3946 ;
  assign n3979 = ~\u1_u3_adr_r_reg[2]/P0001  & ~n3941 ;
  assign n3980 = ~n3978 & n3979 ;
  assign n3981 = ~n3939 & ~n3980 ;
  assign n3982 = n3926 & n3981 ;
  assign n3983 = ~n3977 & n3982 ;
  assign n3984 = ~n3952 & ~n3983 ;
  assign n3985 = n3895 & ~n3914 ;
  assign n3986 = ~n3909 & ~n3914 ;
  assign n3987 = ~n3910 & n3986 ;
  assign n3988 = ~n3985 & ~n3987 ;
  assign n3989 = \u1_u3_adr_r_reg[5]/P0001  & n3988 ;
  assign n3990 = n3895 & ~n3923 ;
  assign n3991 = ~n3919 & ~n3923 ;
  assign n3992 = ~n3917 & n3991 ;
  assign n3993 = ~n3990 & ~n3992 ;
  assign n3994 = \u1_u3_adr_r_reg[4]/P0001  & n3993 ;
  assign n3995 = ~n3916 & n3994 ;
  assign n3996 = ~n3989 & ~n3995 ;
  assign n3997 = n3984 & n3996 ;
  assign n3998 = ~\u1_u3_adr_r_reg[6]/P0001  & ~n3875 ;
  assign n3999 = ~n3873 & n3998 ;
  assign n4000 = n3872 & n3999 ;
  assign n4001 = ~n3867 & ~n4000 ;
  assign n4002 = n3856 & n4001 ;
  assign n4003 = ~n3906 & n4002 ;
  assign n4004 = ~n3997 & n4003 ;
  assign n4005 = ~n3907 & ~n4004 ;
  assign n4006 = \u1_u3_adr_r_reg[11]/P0001  & \u1_u3_adr_r_reg[12]/P0001  ;
  assign n4007 = \u1_u3_adr_r_reg[13]/P0001  & n4006 ;
  assign n4008 = ~\u1_u3_adr_r_reg[14]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4009 = n4007 & n4008 ;
  assign n4010 = ~n4005 & n4009 ;
  assign n4011 = \u1_u3_adr_r_reg[14]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4012 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[14]/P0001  ;
  assign n4013 = ~n4011 & ~n4012 ;
  assign n4014 = n4007 & ~n4012 ;
  assign n4015 = ~n4005 & n4014 ;
  assign n4016 = ~n4013 & ~n4015 ;
  assign n4017 = ~n4010 & ~n4016 ;
  assign n4018 = \u1_u2_adr_cb_reg[0]/NET0131  & \u1_u2_adr_cb_reg[1]/NET0131  ;
  assign n4019 = ~\u1_u2_adr_cb_reg[2]/NET0131  & ~n4018 ;
  assign n4020 = \u1_u2_adr_cb_reg[2]/NET0131  & n4018 ;
  assign n4021 = ~n4019 & ~n4020 ;
  assign n4022 = ~n1763 & ~n4021 ;
  assign n4023 = ~\u1_u2_rx_dma_en_r_reg/P0001  & ~\u1_u2_tx_dma_en_r_reg/P0001  ;
  assign n4024 = ~\u1_u2_adr_cb_reg[2]/NET0131  & ~\u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n4025 = ~n1757 & n4024 ;
  assign n4026 = n4023 & ~n4025 ;
  assign n4027 = ~n4022 & n4026 ;
  assign n4028 = \u1_u3_adr_reg[2]/P0001  & ~n4023 ;
  assign n4029 = ~n4027 & ~n4028 ;
  assign n4030 = rst_i_pad & ~n4029 ;
  assign n4031 = ~n1757 & n1769 ;
  assign n4032 = n4023 & n4031 ;
  assign n4033 = \u1_u2_adr_cb_reg[0]/NET0131  & ~\u1_u2_adr_cb_reg[1]/NET0131  ;
  assign n4034 = ~\u1_u2_adr_cb_reg[0]/NET0131  & \u1_u2_adr_cb_reg[1]/NET0131  ;
  assign n4035 = ~n4033 & ~n4034 ;
  assign n4036 = n4023 & n4035 ;
  assign n4037 = ~n1763 & n4036 ;
  assign n4038 = ~n4032 & ~n4037 ;
  assign n4039 = ~\u1_u3_adr_reg[1]/P0001  & ~n4023 ;
  assign n4040 = rst_i_pad & ~n4039 ;
  assign n4041 = n4038 & n4040 ;
  assign n4042 = \u1_u2_adr_cb_reg[0]/NET0131  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n4043 = \u1_u1_state_reg[1]/NET0131  & \u1_u2_adr_cb_reg[0]/NET0131  ;
  assign n4044 = n1756 & n4043 ;
  assign n4045 = ~n4042 & ~n4044 ;
  assign n4046 = ~\u1_u2_adr_cb_reg[0]/NET0131  & ~\u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n4047 = ~n1757 & n4046 ;
  assign n4048 = n4045 & ~n4047 ;
  assign n4049 = n4023 & ~n4048 ;
  assign n4050 = ~\u1_u3_adr_reg[0]/P0001  & ~n4023 ;
  assign n4051 = rst_i_pad & ~n4050 ;
  assign n4052 = ~n4049 & n4051 ;
  assign n4053 = \u1_u2_sizd_c_reg[0]/P0001  & ~n1757 ;
  assign n4054 = ~n3422 & ~n4053 ;
  assign n4055 = n3437 & n4054 ;
  assign n4056 = ~\u1_u2_send_data_r_reg/NET0131  & ~n3422 ;
  assign n4057 = rst_i_pad & ~n4056 ;
  assign n4058 = ~n4055 & n4057 ;
  assign n4059 = ~\u1_u2_mack_r_reg/P0001  & ~\u1_u2_state_reg[0]/P0001  ;
  assign n4060 = ~\u1_u2_state_reg[2]/NET0131  & ~\u1_u2_state_reg[3]/NET0131  ;
  assign n4061 = ~\u1_u2_state_reg[0]/P0001  & ~\u1_u2_state_reg[1]/NET0131  ;
  assign n4062 = n4060 & n4061 ;
  assign n4063 = ~\u1_u2_state_reg[5]/NET0131  & ~\u1_u2_state_reg[7]/NET0131  ;
  assign n4064 = \u1_u2_state_reg[4]/NET0131  & ~\u1_u2_state_reg[6]/NET0131  ;
  assign n4065 = n4063 & n4064 ;
  assign n4066 = n4062 & n4065 ;
  assign n4067 = ~n4059 & n4066 ;
  assign n4068 = rst_i_pad & ~n4067 ;
  assign n4069 = ~\u1_u2_state_reg[4]/NET0131  & ~\u1_u2_state_reg[6]/NET0131  ;
  assign n4070 = n4063 & n4069 ;
  assign n4071 = n4061 & n4070 ;
  assign n4072 = ~\u1_u2_rx_data_done_r2_reg/P0001  & \u1_u2_state_reg[0]/P0001  ;
  assign n4073 = ~\u1_u3_abort_reg/P0001  & ~n4072 ;
  assign n4074 = \u1_u2_state_reg[2]/NET0131  & ~\u1_u2_state_reg[3]/NET0131  ;
  assign n4075 = ~n4073 & n4074 ;
  assign n4076 = n4071 & n4075 ;
  assign n4077 = ~\u1_u2_state_reg[0]/P0001  & ~\u1_u2_wr_done_reg/P0001  ;
  assign n4078 = ~\u1_u2_wr_last_reg/P0001  & ~n4077 ;
  assign n4079 = ~\u1_u3_abort_reg/P0001  & ~n4078 ;
  assign n4080 = ~\u1_u2_state_reg[2]/NET0131  & \u1_u2_state_reg[3]/NET0131  ;
  assign n4081 = n4061 & n4080 ;
  assign n4082 = n4070 & n4081 ;
  assign n4083 = ~n4079 & n4082 ;
  assign n4084 = ~n4076 & ~n4083 ;
  assign n4085 = n4068 & n4084 ;
  assign n4086 = \u1_u2_state_reg[0]/P0001  & ~\u1_u2_state_reg[1]/NET0131  ;
  assign n4087 = n4060 & n4086 ;
  assign n4088 = n4070 & n4087 ;
  assign n4089 = ~\u1_u1_send_zero_length_r_reg/P0001  & \u1_u2_tx_dma_en_r_reg/P0001  ;
  assign n4090 = ~\u1_u3_abort_reg/P0001  & n4089 ;
  assign n4091 = \u1_u2_rx_dma_en_r_reg/P0001  & ~\u1_u3_abort_reg/P0001  ;
  assign n4092 = ~n4090 & ~n4091 ;
  assign n4093 = n4088 & n4092 ;
  assign n4094 = n4085 & ~n4093 ;
  assign n4095 = ~\u1_u2_mack_r_reg/P0001  & \u1_u2_state_reg[0]/P0001  ;
  assign n4096 = ~\u1_u3_abort_reg/P0001  & ~n4095 ;
  assign n4097 = \u1_u2_state_reg[5]/NET0131  & ~\u1_u2_state_reg[7]/NET0131  ;
  assign n4098 = n4069 & n4097 ;
  assign n4099 = n4062 & n4098 ;
  assign n4100 = ~\u1_u2_state_reg[4]/NET0131  & \u1_u2_state_reg[6]/NET0131  ;
  assign n4101 = n4063 & n4100 ;
  assign n4102 = n4062 & n4101 ;
  assign n4103 = ~n4099 & ~n4102 ;
  assign n4104 = ~\u1_u2_state_reg[0]/P0001  & \u1_u2_state_reg[1]/NET0131  ;
  assign n4105 = n4060 & n4104 ;
  assign n4106 = n4070 & n4105 ;
  assign n4107 = n4103 & ~n4106 ;
  assign n4108 = ~n4096 & ~n4107 ;
  assign n4109 = ~\u1_u2_sizd_is_zero_reg/P0001  & ~\u1_u3_abort_reg/P0001  ;
  assign n4110 = ~\u1_u2_state_reg[0]/P0001  & n4109 ;
  assign n4111 = n4018 & n4109 ;
  assign n4112 = n1757 & n4111 ;
  assign n4113 = ~n4110 & ~n4112 ;
  assign n4114 = ~\u1_u2_state_reg[5]/NET0131  & \u1_u2_state_reg[7]/NET0131  ;
  assign n4115 = n4062 & n4114 ;
  assign n4116 = n4069 & n4115 ;
  assign n4117 = n4113 & n4116 ;
  assign n4118 = ~n4108 & ~n4117 ;
  assign n4119 = n4094 & n4118 ;
  assign n4120 = ~n3997 & n4002 ;
  assign n4121 = ~n3887 & ~n3901 ;
  assign n4122 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n3890 ;
  assign n4123 = ~n3897 & n4122 ;
  assign n4124 = ~n3906 & n4123 ;
  assign n4125 = n4121 & n4124 ;
  assign n4126 = ~n4120 & n4125 ;
  assign n4127 = n3898 & ~n3906 ;
  assign n4128 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n4127 ;
  assign n4129 = ~n4121 & n4128 ;
  assign n4130 = n4002 & n4128 ;
  assign n4131 = ~n3997 & n4130 ;
  assign n4132 = ~n4129 & ~n4131 ;
  assign n4133 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[10]/P0001  ;
  assign n4134 = n4132 & ~n4133 ;
  assign n4135 = ~n4126 & n4134 ;
  assign n4136 = ~n3881 & ~n3901 ;
  assign n4137 = ~n3855 & ~n3906 ;
  assign n4138 = ~n4136 & n4137 ;
  assign n4139 = n3898 & ~n4138 ;
  assign n4140 = \u1_u3_adr_r_reg[11]/P0001  & ~\u1_u3_adr_r_reg[12]/P0001  ;
  assign n4141 = ~n4139 & n4140 ;
  assign n4142 = ~n3879 & ~n3884 ;
  assign n4143 = n3996 & n4142 ;
  assign n4144 = n3984 & n4143 ;
  assign n4145 = ~n3884 & ~n4001 ;
  assign n4146 = ~n3879 & n4145 ;
  assign n4147 = n3856 & ~n3906 ;
  assign n4148 = n4140 & n4147 ;
  assign n4149 = ~n4146 & n4148 ;
  assign n4150 = ~n4144 & n4149 ;
  assign n4151 = ~n4141 & ~n4150 ;
  assign n4152 = \u1_u3_adr_r_reg[11]/P0001  & n4147 ;
  assign n4153 = ~n4146 & n4152 ;
  assign n4154 = ~n4144 & n4153 ;
  assign n4155 = ~\u1_u3_adr_r_reg[11]/P0001  & \u1_u3_adr_r_reg[12]/P0001  ;
  assign n4156 = \u1_u3_adr_r_reg[12]/P0001  & n3898 ;
  assign n4157 = ~n4138 & n4156 ;
  assign n4158 = ~n4155 & ~n4157 ;
  assign n4159 = ~n4154 & ~n4158 ;
  assign n4160 = n4151 & ~n4159 ;
  assign n4161 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n4160 ;
  assign n4162 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[12]/P0001  ;
  assign n4163 = ~n4161 & ~n4162 ;
  assign n4164 = \u1_u3_adr_r_reg[13]/P0001  & \u1_u3_adr_r_reg[14]/P0001  ;
  assign n4165 = \u1_u3_adr_r_reg[12]/P0001  & \u1_u3_adr_r_reg[15]/P0001  ;
  assign n4166 = n4164 & n4165 ;
  assign n4167 = \u1_u3_adr_r_reg[16]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4168 = ~n4166 & n4167 ;
  assign n4169 = \u1_u3_adr_r_reg[11]/P0001  & ~n4139 ;
  assign n4170 = n4167 & ~n4169 ;
  assign n4171 = ~n4154 & n4170 ;
  assign n4172 = ~n4168 & ~n4171 ;
  assign n4173 = ~n4154 & ~n4169 ;
  assign n4174 = ~\u1_u3_adr_r_reg[16]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4175 = n4166 & n4174 ;
  assign n4176 = ~n4173 & n4175 ;
  assign n4177 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[16]/P0001  ;
  assign n4178 = ~n4176 & ~n4177 ;
  assign n4179 = n4172 & n4178 ;
  assign n4180 = n1757 & n4018 ;
  assign n4181 = ~\u1_u2_state_reg[6]/NET0131  & ~n4180 ;
  assign n4182 = n4069 & n4114 ;
  assign n4183 = n4062 & n4182 ;
  assign n4184 = n4109 & n4183 ;
  assign n4185 = ~n4181 & n4184 ;
  assign n4186 = ~\u1_u2_mack_r_reg/P0001  & ~\u1_u2_state_reg[6]/NET0131  ;
  assign n4187 = ~\u1_u3_abort_reg/P0001  & ~n4186 ;
  assign n4188 = n4099 & n4187 ;
  assign n4189 = ~\u1_u2_mack_r_reg/P0001  & ~\u1_u3_abort_reg/P0001  ;
  assign n4190 = n4102 & n4189 ;
  assign n4191 = ~n4188 & ~n4190 ;
  assign n4192 = ~n4185 & n4191 ;
  assign n4193 = rst_i_pad & ~n4192 ;
  assign n4194 = ~\u1_u2_mack_r_reg/P0001  & ~\u1_u2_state_reg[7]/NET0131  ;
  assign n4195 = rst_i_pad & ~\u1_u3_abort_reg/P0001  ;
  assign n4196 = ~n4194 & n4195 ;
  assign n4197 = n4102 & n4196 ;
  assign n4198 = rst_i_pad & ~n4180 ;
  assign n4199 = n4184 & n4198 ;
  assign n4200 = ~n4197 & ~n4199 ;
  assign n4201 = n3949 & n3962 ;
  assign n4202 = ~n3976 & n4201 ;
  assign n4203 = n3981 & ~n4202 ;
  assign n4204 = n3936 & ~n3994 ;
  assign n4205 = ~n4203 & n4204 ;
  assign n4206 = ~n3843 & ~n3867 ;
  assign n4207 = n3926 & ~n4000 ;
  assign n4208 = n4206 & n4207 ;
  assign n4209 = ~n4205 & n4208 ;
  assign n4210 = n3989 & ~n4000 ;
  assign n4211 = ~n3878 & ~n4210 ;
  assign n4212 = n4206 & ~n4211 ;
  assign n4213 = n3901 & ~n3906 ;
  assign n4214 = n3898 & ~n4213 ;
  assign n4215 = ~n3843 & n3884 ;
  assign n4216 = ~n3881 & ~n4215 ;
  assign n4217 = n4214 & n4216 ;
  assign n4218 = ~n4212 & n4217 ;
  assign n4219 = ~n4209 & n4218 ;
  assign n4220 = n3898 & n3906 ;
  assign n4221 = n3855 & ~n3901 ;
  assign n4222 = n3898 & n4221 ;
  assign n4223 = ~n4220 & ~n4222 ;
  assign n4224 = n4006 & n4223 ;
  assign n4225 = ~\u1_u3_adr_r_reg[13]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4226 = n4224 & n4225 ;
  assign n4227 = ~n4219 & n4226 ;
  assign n4228 = \u1_u3_adr_r_reg[13]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4229 = ~n4224 & n4228 ;
  assign n4230 = n4218 & n4228 ;
  assign n4231 = ~n4209 & n4230 ;
  assign n4232 = ~n4229 & ~n4231 ;
  assign n4233 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[13]/P0001  ;
  assign n4234 = n4232 & ~n4233 ;
  assign n4235 = ~n4227 & n4234 ;
  assign n4236 = ~\u1_u1_send_zero_length_r_reg/P0001  & \u1_u2_send_data_r_reg/NET0131  ;
  assign n4237 = n1847 & n4236 ;
  assign n4238 = rst_i_pad & ~\u1_u1_state_reg[3]/NET0131  ;
  assign n4239 = n1829 & n4238 ;
  assign n4240 = n4237 & n4239 ;
  assign n4241 = rst_i_pad & ~n1828 ;
  assign n4242 = n1832 & n4241 ;
  assign n4243 = ~n4240 & ~n4242 ;
  assign n4244 = ~n4207 & n4211 ;
  assign n4245 = n4204 & n4211 ;
  assign n4246 = ~n4203 & n4245 ;
  assign n4247 = ~n4244 & ~n4246 ;
  assign n4248 = n4006 & n4164 ;
  assign n4249 = n4206 & n4248 ;
  assign n4250 = n4137 & n4249 ;
  assign n4251 = n4247 & n4250 ;
  assign n4252 = ~n4214 & n4248 ;
  assign n4253 = n4137 & n4248 ;
  assign n4254 = ~n4216 & n4253 ;
  assign n4255 = ~n4252 & ~n4254 ;
  assign n4256 = \u1_u3_adr_r_reg[15]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4257 = n4255 & n4256 ;
  assign n4258 = ~n4251 & n4257 ;
  assign n4259 = ~\u1_u3_adr_r_reg[15]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4260 = ~n4255 & n4259 ;
  assign n4261 = n4250 & n4259 ;
  assign n4262 = n4247 & n4261 ;
  assign n4263 = ~n4260 & ~n4262 ;
  assign n4264 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[15]/P0001  ;
  assign n4265 = n4263 & ~n4264 ;
  assign n4266 = ~n4258 & n4265 ;
  assign n4267 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[11]/P0001  ;
  assign n4268 = ~\u1_u3_adr_r_reg[11]/P0001  & ~n4214 ;
  assign n4269 = ~\u1_u3_adr_r_reg[11]/P0001  & n4137 ;
  assign n4270 = ~n4216 & n4269 ;
  assign n4271 = ~n4268 & ~n4270 ;
  assign n4272 = n4137 & n4206 ;
  assign n4273 = ~\u1_u3_adr_r_reg[11]/P0001  & n4272 ;
  assign n4274 = n4247 & n4273 ;
  assign n4275 = n4271 & ~n4274 ;
  assign n4276 = n4247 & n4272 ;
  assign n4277 = n4137 & ~n4216 ;
  assign n4278 = n4214 & ~n4277 ;
  assign n4279 = \u1_u3_adr_r_reg[11]/P0001  & n4278 ;
  assign n4280 = ~n4276 & n4279 ;
  assign n4281 = n4275 & ~n4280 ;
  assign n4282 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n4281 ;
  assign n4283 = ~n4267 & ~n4282 ;
  assign n4284 = ~n3878 & ~n4000 ;
  assign n4285 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n4284 ;
  assign n4286 = ~n3997 & n4285 ;
  assign n4287 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n4000 ;
  assign n4288 = ~n3878 & n4287 ;
  assign n4289 = n3996 & n4288 ;
  assign n4290 = n3984 & n4289 ;
  assign n4291 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[6]/P0001  ;
  assign n4292 = ~n4290 & ~n4291 ;
  assign n4293 = ~n4286 & n4292 ;
  assign n4294 = ~\u1_u3_out_to_small_r_reg/P0001  & n3843 ;
  assign n4295 = \u1_u3_adr_r_reg[8]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4296 = ~n3880 & n4295 ;
  assign n4297 = ~n4294 & ~n4296 ;
  assign n4298 = ~n4146 & ~n4297 ;
  assign n4299 = ~n4144 & n4298 ;
  assign n4300 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n3843 ;
  assign n4301 = ~n3881 & n4300 ;
  assign n4302 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[8]/P0001  ;
  assign n4303 = ~n4301 & ~n4302 ;
  assign n4304 = ~n4146 & ~n4302 ;
  assign n4305 = ~n4144 & n4304 ;
  assign n4306 = ~n4303 & ~n4305 ;
  assign n4307 = ~n4299 & ~n4306 ;
  assign n4308 = ~n4212 & n4216 ;
  assign n4309 = ~n3855 & ~n3901 ;
  assign n4310 = ~\u1_u3_out_to_small_r_reg/P0001  & n4309 ;
  assign n4311 = n4308 & n4310 ;
  assign n4312 = ~n4209 & n4311 ;
  assign n4313 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n4309 ;
  assign n4314 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[9]/P0001  ;
  assign n4315 = ~n4313 & ~n4314 ;
  assign n4316 = n4308 & ~n4314 ;
  assign n4317 = ~n4209 & n4316 ;
  assign n4318 = ~n4315 & ~n4317 ;
  assign n4319 = ~n4312 & ~n4318 ;
  assign n4320 = rst_i_pad & ~n1860 ;
  assign n4321 = \u1_u3_new_size_reg[12]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4322 = ~n3977 & n3981 ;
  assign n4323 = ~n3925 & ~n3994 ;
  assign n4324 = n3951 & n4323 ;
  assign n4325 = ~n4322 & n4324 ;
  assign n4326 = ~n3951 & ~n4323 ;
  assign n4327 = n3981 & ~n4323 ;
  assign n4328 = ~n3977 & n4327 ;
  assign n4329 = ~n4326 & ~n4328 ;
  assign n4330 = ~n4325 & n4329 ;
  assign n4331 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n4330 ;
  assign n4332 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[4]/P0001  ;
  assign n4333 = ~n4331 & ~n4332 ;
  assign n4334 = ~n3925 & ~n4204 ;
  assign n4335 = ~n3925 & n3981 ;
  assign n4336 = ~n4202 & n4335 ;
  assign n4337 = ~n4334 & ~n4336 ;
  assign n4338 = ~n3916 & ~n3989 ;
  assign n4339 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n4338 ;
  assign n4340 = ~n4337 & n4339 ;
  assign n4341 = ~\u1_u3_out_to_small_r_reg/P0001  & n4338 ;
  assign n4342 = n4337 & n4341 ;
  assign n4343 = ~n4340 & ~n4342 ;
  assign n4344 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[5]/P0001  ;
  assign n4345 = n4343 & ~n4344 ;
  assign n4346 = ~n3867 & ~n3884 ;
  assign n4347 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n4346 ;
  assign n4348 = n4247 & n4347 ;
  assign n4349 = ~\u1_u3_out_to_small_r_reg/P0001  & n4346 ;
  assign n4350 = ~n4247 & n4349 ;
  assign n4351 = ~n4348 & ~n4350 ;
  assign n4352 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[7]/P0001  ;
  assign n4353 = n4351 & ~n4352 ;
  assign n4354 = \u1_u3_new_size_reg[13]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4355 = ~\u4_u2_csr1_reg[11]/P0001  & \u4_u2_csr1_reg[12]/P0001  ;
  assign n4356 = \u4_u2_dma_req_out_hold_reg/P0001  & n4355 ;
  assign n4357 = \dma_ack_i[2]_pad  & ~n4356 ;
  assign n4358 = \u4_u2_r1_reg/P0001  & ~\u4_u2_r2_reg/P0001  ;
  assign n4359 = \u4_u2_dma_req_in_hold2_reg/P0001  & \u4_u2_dma_req_in_hold_reg/P0001  ;
  assign n4360 = ~n4355 & n4359 ;
  assign n4361 = ~n4358 & ~n4360 ;
  assign n4362 = n4357 & n4361 ;
  assign n4363 = ~\dma_req_o[2]_pad  & ~n4358 ;
  assign n4364 = rst_i_pad & ~n4363 ;
  assign n4365 = ~n4362 & n4364 ;
  assign n4366 = ~\u4_u3_csr1_reg[11]/P0001  & \u4_u3_csr1_reg[12]/P0001  ;
  assign n4367 = \u4_u3_dma_req_out_hold_reg/P0001  & n4366 ;
  assign n4368 = \dma_ack_i[3]_pad  & ~n4367 ;
  assign n4369 = \u4_u3_r1_reg/P0001  & ~\u4_u3_r2_reg/P0001  ;
  assign n4370 = \u4_u3_dma_req_in_hold2_reg/P0001  & \u4_u3_dma_req_in_hold_reg/P0001  ;
  assign n4371 = ~n4366 & n4370 ;
  assign n4372 = ~n4369 & ~n4371 ;
  assign n4373 = n4368 & n4372 ;
  assign n4374 = ~\dma_req_o[3]_pad  & ~n4369 ;
  assign n4375 = rst_i_pad & ~n4374 ;
  assign n4376 = ~n4373 & n4375 ;
  assign n4377 = ~\u4_u0_csr1_reg[11]/P0001  & \u4_u0_csr1_reg[12]/P0001  ;
  assign n4378 = \u4_u0_dma_req_out_hold_reg/P0001  & n4377 ;
  assign n4379 = \dma_ack_i[0]_pad  & ~n4378 ;
  assign n4380 = \u4_u0_r1_reg/P0001  & ~\u4_u0_r2_reg/P0001  ;
  assign n4381 = \u4_u0_dma_req_in_hold2_reg/P0001  & \u4_u0_dma_req_in_hold_reg/P0001  ;
  assign n4382 = ~n4377 & n4381 ;
  assign n4383 = ~n4380 & ~n4382 ;
  assign n4384 = n4379 & n4383 ;
  assign n4385 = ~\dma_req_o[0]_pad  & ~n4380 ;
  assign n4386 = rst_i_pad & ~n4385 ;
  assign n4387 = ~n4384 & n4386 ;
  assign n4388 = ~\u4_u1_csr1_reg[11]/P0001  & \u4_u1_csr1_reg[12]/P0001  ;
  assign n4389 = \u4_u1_dma_req_out_hold_reg/P0001  & n4388 ;
  assign n4390 = \dma_ack_i[1]_pad  & ~n4389 ;
  assign n4391 = \u4_u1_r1_reg/P0001  & ~\u4_u1_r2_reg/P0001  ;
  assign n4392 = \u4_u1_dma_req_in_hold2_reg/P0001  & \u4_u1_dma_req_in_hold_reg/P0001  ;
  assign n4393 = ~n4388 & n4392 ;
  assign n4394 = ~n4391 & ~n4393 ;
  assign n4395 = n4390 & n4394 ;
  assign n4396 = ~\dma_req_o[1]_pad  & ~n4391 ;
  assign n4397 = rst_i_pad & ~n4396 ;
  assign n4398 = ~n4395 & n4397 ;
  assign n4399 = \u1_u3_buffer_done_reg/P0001  & \u4_csr_reg[15]/NET0131  ;
  assign n4400 = ~n2358 & n4399 ;
  assign n4401 = \u1_u3_state_reg[8]/P0001  & ~n4400 ;
  assign n4402 = ~\u1_u3_next_dpid_reg[0]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4403 = \u1_u3_out_to_small_r_reg/P0001  & ~\u4_buf0_reg[2]/P0001  ;
  assign n4404 = ~n4402 & ~n4403 ;
  assign n4405 = ~n4401 & n4404 ;
  assign n4406 = n3949 & ~n3980 ;
  assign n4407 = n3977 & ~n4406 ;
  assign n4408 = n4401 & ~n4406 ;
  assign n4409 = n3962 & n4401 ;
  assign n4410 = ~n3976 & n4409 ;
  assign n4411 = ~n4408 & ~n4410 ;
  assign n4412 = ~n4407 & ~n4411 ;
  assign n4413 = ~n4405 & ~n4412 ;
  assign n4414 = ~\u1_u3_next_dpid_reg[1]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4415 = \u1_u3_out_to_small_r_reg/P0001  & ~\u4_buf0_reg[3]/P0001  ;
  assign n4416 = ~n4414 & ~n4415 ;
  assign n4417 = ~n4401 & n4416 ;
  assign n4418 = n3936 & n3981 ;
  assign n4419 = ~n4202 & n4418 ;
  assign n4420 = ~n4417 & n4419 ;
  assign n4421 = ~n3979 & n4401 ;
  assign n4422 = ~n3895 & n4401 ;
  assign n4423 = ~n3946 & n4422 ;
  assign n4424 = ~n4421 & ~n4423 ;
  assign n4425 = ~n4202 & ~n4424 ;
  assign n4426 = ~n3938 & n4401 ;
  assign n4427 = ~n3933 & n4422 ;
  assign n4428 = ~n4426 & ~n4427 ;
  assign n4429 = n3936 & ~n4428 ;
  assign n4430 = ~n4417 & ~n4429 ;
  assign n4431 = ~n4425 & n4430 ;
  assign n4432 = ~n4420 & ~n4431 ;
  assign n4433 = \u1_u3_new_sizeb_reg[3]/P0001  & n3511 ;
  assign n4434 = ~\u1_u3_new_sizeb_reg[3]/P0001  & ~n3511 ;
  assign n4435 = ~\u1_u3_new_sizeb_reg[2]/P0001  & ~n3493 ;
  assign n4436 = ~n4434 & ~n4435 ;
  assign n4437 = ~n4433 & ~n4436 ;
  assign n4438 = ~\u1_u3_new_sizeb_reg[1]/P0001  & ~n3475 ;
  assign n4439 = \u1_u3_new_sizeb_reg[1]/P0001  & n3475 ;
  assign n4440 = \u1_u3_new_sizeb_reg[0]/P0001  & n3483 ;
  assign n4441 = ~n4439 & ~n4440 ;
  assign n4442 = ~n4438 & ~n4441 ;
  assign n4443 = \u1_u3_new_sizeb_reg[2]/P0001  & n3493 ;
  assign n4444 = ~n4433 & ~n4443 ;
  assign n4445 = ~n4442 & n4444 ;
  assign n4446 = ~n4437 & ~n4445 ;
  assign n4447 = \u1_u3_new_sizeb_reg[7]/P0001  & n3538 ;
  assign n4448 = \u1_u3_new_sizeb_reg[6]/P0001  & n3572 ;
  assign n4449 = ~n4447 & ~n4448 ;
  assign n4450 = \u1_u3_new_sizeb_reg[5]/P0001  & n3525 ;
  assign n4451 = \u1_u3_new_sizeb_reg[4]/P0001  & n3503 ;
  assign n4452 = ~n4450 & ~n4451 ;
  assign n4453 = n4449 & n4452 ;
  assign n4454 = ~n4446 & n4453 ;
  assign n4455 = ~\u1_u3_new_sizeb_reg[5]/P0001  & ~n3525 ;
  assign n4456 = ~\u1_u3_new_sizeb_reg[4]/P0001  & ~n3503 ;
  assign n4457 = ~n4450 & n4456 ;
  assign n4458 = ~n4455 & ~n4457 ;
  assign n4459 = n4449 & ~n4458 ;
  assign n4460 = ~\u1_u3_new_sizeb_reg[9]/P0001  & ~n3563 ;
  assign n4461 = \u1_u3_new_sizeb_reg[9]/P0001  & n3563 ;
  assign n4462 = ~\u1_u3_new_sizeb_reg[8]/P0001  & ~n3546 ;
  assign n4463 = ~n4461 & n4462 ;
  assign n4464 = ~n4460 & ~n4463 ;
  assign n4465 = ~\u1_u3_new_sizeb_reg[7]/P0001  & ~n3538 ;
  assign n4466 = ~\u1_u3_new_sizeb_reg[6]/P0001  & ~n3572 ;
  assign n4467 = ~n4447 & n4466 ;
  assign n4468 = ~n4465 & ~n4467 ;
  assign n4469 = n4464 & n4468 ;
  assign n4470 = ~n4459 & n4469 ;
  assign n4471 = ~n4454 & n4470 ;
  assign n4472 = \u1_u3_new_sizeb_reg[10]/P0001  & n3555 ;
  assign n4473 = \u1_u3_new_sizeb_reg[8]/P0001  & n3546 ;
  assign n4474 = n3563 & n4473 ;
  assign n4475 = \u1_u3_new_sizeb_reg[8]/P0001  & \u1_u3_new_sizeb_reg[9]/P0001  ;
  assign n4476 = n3546 & n4475 ;
  assign n4477 = ~n4461 & ~n4476 ;
  assign n4478 = ~n4474 & n4477 ;
  assign n4479 = ~n4472 & n4478 ;
  assign n4480 = ~n4471 & n4479 ;
  assign n4481 = ~\u1_u3_new_sizeb_reg[10]/P0001  & ~n3555 ;
  assign n4482 = n3601 & ~n4481 ;
  assign n4483 = ~n4480 & n4482 ;
  assign n4484 = ~n3594 & ~n4483 ;
  assign n4485 = n3602 & ~n4481 ;
  assign n4486 = ~n4480 & n4485 ;
  assign n4487 = ~n4484 & ~n4486 ;
  assign n4488 = ~n1832 & ~n1837 ;
  assign n4489 = n1852 & n4488 ;
  assign n4490 = ~\u0_u0_drive_k_reg/P0001  & ~\u1_u3_send_token_reg/P0001  ;
  assign n4491 = ~TxReady_pad_i_pad & TxValid_pad_o_pad ;
  assign n4492 = ~\u0_drive_k_r_reg/P0001  & n4491 ;
  assign n4493 = ~\u0_tx_ready_reg/NET0131  & ~n4492 ;
  assign n4494 = ~n1839 & n4493 ;
  assign n4495 = \u0_tx_ready_reg/NET0131  & ~n4492 ;
  assign n4496 = ~n1851 & n4495 ;
  assign n4497 = ~n4494 & ~n4496 ;
  assign n4498 = n4490 & ~n4497 ;
  assign n4499 = n4489 & n4498 ;
  assign n4500 = rst_i_pad & ~n4499 ;
  assign n4501 = n3962 & ~n3965 ;
  assign n4502 = ~n3968 & n4401 ;
  assign n4503 = ~n3974 & n4502 ;
  assign n4504 = n4501 & n4503 ;
  assign n4505 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[1]/P0001  ;
  assign n4506 = ~\u1_u3_out_to_small_r_reg/P0001  & ~n2366 ;
  assign n4507 = \u1_u3_buffer_done_reg/P0001  & \u4_csr_reg[30]/NET0131  ;
  assign n4508 = ~\u4_csr_reg[31]/P0001  & ~n4507 ;
  assign n4509 = \u4_csr_reg[31]/P0001  & n4507 ;
  assign n4510 = ~n4508 & ~n4509 ;
  assign n4511 = n4506 & n4510 ;
  assign n4512 = ~n4505 & ~n4511 ;
  assign n4513 = ~n4401 & ~n4512 ;
  assign n4514 = n3968 & n4401 ;
  assign n4515 = n3973 & n4401 ;
  assign n4516 = ~n3972 & n4515 ;
  assign n4517 = ~n4514 & ~n4516 ;
  assign n4518 = ~n4501 & ~n4517 ;
  assign n4519 = ~n4513 & ~n4518 ;
  assign n4520 = ~n4504 & n4519 ;
  assign n4521 = \u1_u2_sizu_c_reg[10]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n4522 = \u1_u3_new_size_reg[10]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n4523 = ~n4521 & ~n4522 ;
  assign n4524 = ~n3601 & n4481 ;
  assign n4525 = ~n3601 & ~n4472 ;
  assign n4526 = n4478 & n4525 ;
  assign n4527 = ~n4471 & n4526 ;
  assign n4528 = ~n4524 & ~n4527 ;
  assign n4529 = ~n4483 & n4528 ;
  assign n4530 = ~n4461 & ~n4472 ;
  assign n4531 = n4485 & ~n4530 ;
  assign n4532 = ~n3609 & n4531 ;
  assign n4533 = ~n4447 & ~n4473 ;
  assign n4534 = ~n4448 & n4533 ;
  assign n4535 = n4466 & n4534 ;
  assign n4536 = ~n4455 & ~n4456 ;
  assign n4537 = ~n4437 & n4536 ;
  assign n4538 = ~n4445 & n4537 ;
  assign n4539 = ~n4452 & ~n4455 ;
  assign n4540 = n4534 & ~n4539 ;
  assign n4541 = ~n4538 & n4540 ;
  assign n4542 = ~n4535 & ~n4541 ;
  assign n4543 = n4460 & ~n4472 ;
  assign n4544 = n4485 & ~n4543 ;
  assign n4545 = n4465 & ~n4473 ;
  assign n4546 = ~n4462 & ~n4545 ;
  assign n4547 = n4544 & n4546 ;
  assign n4548 = ~n3609 & n4547 ;
  assign n4549 = n4542 & n4548 ;
  assign n4550 = ~n4532 & ~n4549 ;
  assign n4551 = n4542 & n4547 ;
  assign n4552 = n3609 & ~n4531 ;
  assign n4553 = ~n4551 & n4552 ;
  assign n4554 = n4550 & ~n4553 ;
  assign n4555 = ~\u1_u2_dtmp_sel_r_reg/P0001  & \u1_u2_mack_r_reg/P0001  ;
  assign n4556 = \u1_u2_adr_cw_reg[0]/NET0131  & \u1_u2_adr_cw_reg[1]/P0001  ;
  assign n4557 = n4555 & n4556 ;
  assign n4558 = \u1_u2_adr_cw_reg[2]/P0001  & \u1_u2_adr_cw_reg[3]/NET0131  ;
  assign n4559 = n4557 & n4558 ;
  assign n4560 = ~\u1_u2_adr_cw_reg[4]/P0001  & ~\u1_u2_last_buf_adr_reg[4]/P0001  ;
  assign n4561 = ~n4559 & n4560 ;
  assign n4562 = \u1_u2_adr_cw_reg[4]/P0001  & ~\u1_u2_last_buf_adr_reg[4]/P0001  ;
  assign n4563 = n4558 & n4562 ;
  assign n4564 = n4557 & n4563 ;
  assign n4565 = ~n4561 & ~n4564 ;
  assign n4566 = ~\u1_u2_adr_cw_reg[4]/P0001  & ~n4559 ;
  assign n4567 = \u1_u2_adr_cw_reg[2]/P0001  & \u1_u2_adr_cw_reg[4]/P0001  ;
  assign n4568 = \u1_u2_adr_cw_reg[3]/NET0131  & n4567 ;
  assign n4569 = n4557 & n4568 ;
  assign n4570 = \u1_u2_last_buf_adr_reg[4]/P0001  & ~n4569 ;
  assign n4571 = ~n4566 & n4570 ;
  assign n4572 = n4565 & ~n4571 ;
  assign n4573 = \u1_u2_adr_cw_reg[2]/P0001  & n4557 ;
  assign n4574 = ~\u1_u2_adr_cw_reg[3]/NET0131  & ~n4573 ;
  assign n4575 = ~\u1_u2_last_buf_adr_reg[3]/P0001  & ~n4559 ;
  assign n4576 = ~n4574 & n4575 ;
  assign n4577 = ~n4572 & ~n4576 ;
  assign n4578 = \u1_u2_adr_cw_reg[0]/NET0131  & n4555 ;
  assign n4579 = ~\u1_u2_adr_cw_reg[1]/P0001  & ~\u1_u2_last_buf_adr_reg[1]/P0001  ;
  assign n4580 = ~n4578 & n4579 ;
  assign n4581 = \u1_u2_adr_cw_reg[1]/P0001  & ~\u1_u2_last_buf_adr_reg[1]/P0001  ;
  assign n4582 = n4578 & n4581 ;
  assign n4583 = ~n4580 & ~n4582 ;
  assign n4584 = ~\u1_u2_adr_cw_reg[1]/P0001  & ~n4578 ;
  assign n4585 = \u1_u2_last_buf_adr_reg[1]/P0001  & ~n4557 ;
  assign n4586 = ~n4584 & n4585 ;
  assign n4587 = n4583 & ~n4586 ;
  assign n4588 = ~\u1_u2_adr_cw_reg[0]/NET0131  & ~\u1_u2_last_buf_adr_reg[0]/P0001  ;
  assign n4589 = ~n4555 & n4588 ;
  assign n4590 = \u1_u2_adr_cw_reg[0]/NET0131  & ~\u1_u2_last_buf_adr_reg[0]/P0001  ;
  assign n4591 = n4555 & n4590 ;
  assign n4592 = ~n4589 & ~n4591 ;
  assign n4593 = \u1_u2_adr_cw_reg[0]/NET0131  & \u1_u2_last_buf_adr_reg[0]/P0001  ;
  assign n4594 = ~n4555 & n4593 ;
  assign n4595 = ~\u1_u2_adr_cw_reg[0]/NET0131  & \u1_u2_last_buf_adr_reg[0]/P0001  ;
  assign n4596 = n4555 & n4595 ;
  assign n4597 = ~n4594 & ~n4596 ;
  assign n4598 = n4592 & n4597 ;
  assign n4599 = n2366 & ~n4598 ;
  assign n4600 = ~n4587 & n4599 ;
  assign n4601 = ~\u1_u2_adr_cw_reg[3]/NET0131  & \u1_u2_last_buf_adr_reg[3]/P0001  ;
  assign n4602 = ~n4573 & n4601 ;
  assign n4603 = \u1_u2_adr_cw_reg[3]/NET0131  & \u1_u2_last_buf_adr_reg[3]/P0001  ;
  assign n4604 = \u1_u2_adr_cw_reg[2]/P0001  & n4603 ;
  assign n4605 = n4557 & n4604 ;
  assign n4606 = ~n4602 & ~n4605 ;
  assign n4607 = ~\u1_u2_adr_cw_reg[2]/P0001  & ~\u1_u2_last_buf_adr_reg[2]/P0001  ;
  assign n4608 = ~n4557 & n4607 ;
  assign n4609 = \u1_u2_adr_cw_reg[2]/P0001  & ~\u1_u2_last_buf_adr_reg[2]/P0001  ;
  assign n4610 = n4557 & n4609 ;
  assign n4611 = ~n4608 & ~n4610 ;
  assign n4612 = ~\u1_u2_adr_cw_reg[2]/P0001  & \u1_u2_last_buf_adr_reg[2]/P0001  ;
  assign n4613 = n4557 & n4612 ;
  assign n4614 = \u1_u2_adr_cw_reg[2]/P0001  & \u1_u2_last_buf_adr_reg[2]/P0001  ;
  assign n4615 = ~n4557 & n4614 ;
  assign n4616 = ~n4613 & ~n4615 ;
  assign n4617 = n4611 & n4616 ;
  assign n4618 = n4606 & ~n4617 ;
  assign n4619 = n4600 & n4618 ;
  assign n4620 = n4577 & n4619 ;
  assign n4621 = ~\u1_u2_adr_cw_reg[5]/NET0131  & \u1_u2_last_buf_adr_reg[5]/P0001  ;
  assign n4622 = ~n4569 & n4621 ;
  assign n4623 = \u1_u2_adr_cw_reg[5]/NET0131  & \u1_u2_last_buf_adr_reg[5]/P0001  ;
  assign n4624 = n4569 & n4623 ;
  assign n4625 = ~n4622 & ~n4624 ;
  assign n4626 = \u1_u2_adr_cw_reg[3]/NET0131  & ~\u1_u2_adr_cw_reg[5]/NET0131  ;
  assign n4627 = n4567 & n4626 ;
  assign n4628 = n4557 & n4627 ;
  assign n4629 = ~\u1_u2_last_buf_adr_reg[5]/P0001  & n4628 ;
  assign n4630 = \u1_u2_adr_cw_reg[5]/NET0131  & ~\u1_u2_last_buf_adr_reg[5]/P0001  ;
  assign n4631 = ~n4569 & n4630 ;
  assign n4632 = ~n4629 & ~n4631 ;
  assign n4633 = n4625 & n4632 ;
  assign n4634 = \u1_u2_adr_cw_reg[5]/NET0131  & \u1_u2_adr_cw_reg[6]/NET0131  ;
  assign n4635 = n4569 & n4634 ;
  assign n4636 = ~\u1_u2_adr_cw_reg[7]/NET0131  & ~n4635 ;
  assign n4637 = \u1_u2_adr_cw_reg[7]/NET0131  & n4634 ;
  assign n4638 = n4569 & n4637 ;
  assign n4639 = ~\u1_u2_last_buf_adr_reg[7]/P0001  & ~n4638 ;
  assign n4640 = ~n4636 & n4639 ;
  assign n4641 = n4633 & ~n4640 ;
  assign n4642 = n4620 & n4641 ;
  assign n4643 = ~\u1_u2_adr_cw_reg[7]/NET0131  & \u1_u2_last_buf_adr_reg[7]/P0001  ;
  assign n4644 = ~n4635 & n4643 ;
  assign n4645 = \u1_u2_adr_cw_reg[7]/NET0131  & \u1_u2_last_buf_adr_reg[7]/P0001  ;
  assign n4646 = n4634 & n4645 ;
  assign n4647 = n4569 & n4646 ;
  assign n4648 = ~n4644 & ~n4647 ;
  assign n4649 = \u1_u2_adr_cw_reg[5]/NET0131  & n4569 ;
  assign n4650 = ~\u1_u2_adr_cw_reg[6]/NET0131  & ~\u1_u2_last_buf_adr_reg[6]/P0001  ;
  assign n4651 = ~n4649 & n4650 ;
  assign n4652 = \u1_u2_adr_cw_reg[5]/NET0131  & ~\u1_u2_last_buf_adr_reg[6]/P0001  ;
  assign n4653 = \u1_u2_adr_cw_reg[6]/NET0131  & n4652 ;
  assign n4654 = n4569 & n4653 ;
  assign n4655 = ~n4651 & ~n4654 ;
  assign n4656 = ~\u1_u2_adr_cw_reg[6]/NET0131  & ~n4649 ;
  assign n4657 = \u1_u2_last_buf_adr_reg[6]/P0001  & ~n4635 ;
  assign n4658 = ~n4656 & n4657 ;
  assign n4659 = n4655 & ~n4658 ;
  assign n4660 = n4648 & ~n4659 ;
  assign n4661 = ~\u1_u2_adr_cw_reg[8]/P0001  & ~\u1_u2_last_buf_adr_reg[8]/P0001  ;
  assign n4662 = ~n4638 & n4661 ;
  assign n4663 = \u1_u2_adr_cw_reg[5]/NET0131  & \u1_u2_adr_cw_reg[7]/NET0131  ;
  assign n4664 = \u1_u2_adr_cw_reg[6]/NET0131  & n4663 ;
  assign n4665 = \u1_u2_adr_cw_reg[8]/P0001  & ~\u1_u2_last_buf_adr_reg[8]/P0001  ;
  assign n4666 = n4664 & n4665 ;
  assign n4667 = n4569 & n4666 ;
  assign n4668 = ~n4662 & ~n4667 ;
  assign n4669 = n4569 & n4664 ;
  assign n4670 = \u1_u2_adr_cw_reg[8]/P0001  & \u1_u2_last_buf_adr_reg[8]/P0001  ;
  assign n4671 = ~n4669 & n4670 ;
  assign n4672 = ~\u1_u2_adr_cw_reg[8]/P0001  & \u1_u2_last_buf_adr_reg[8]/P0001  ;
  assign n4673 = n4637 & n4672 ;
  assign n4674 = n4569 & n4673 ;
  assign n4675 = ~n4671 & ~n4674 ;
  assign n4676 = n4668 & n4675 ;
  assign n4677 = \u1_u2_adr_cw_reg[7]/NET0131  & \u1_u2_adr_cw_reg[8]/P0001  ;
  assign n4678 = n4634 & n4677 ;
  assign n4679 = n4569 & n4678 ;
  assign n4680 = ~\u1_u2_adr_cw_reg[9]/NET0131  & \u1_u2_last_buf_adr_reg[9]/P0001  ;
  assign n4681 = ~n4679 & n4680 ;
  assign n4682 = \u1_u2_adr_cw_reg[9]/NET0131  & \u1_u2_last_buf_adr_reg[9]/P0001  ;
  assign n4683 = n4679 & n4682 ;
  assign n4684 = ~n4681 & ~n4683 ;
  assign n4685 = ~\u1_u2_adr_cw_reg[9]/NET0131  & ~n4679 ;
  assign n4686 = \u1_u2_adr_cw_reg[8]/P0001  & \u1_u2_adr_cw_reg[9]/NET0131  ;
  assign n4687 = n4664 & n4686 ;
  assign n4688 = n4569 & n4687 ;
  assign n4689 = ~\u1_u2_last_buf_adr_reg[9]/P0001  & ~n4688 ;
  assign n4690 = ~n4685 & n4689 ;
  assign n4691 = n4684 & ~n4690 ;
  assign n4692 = ~n4676 & n4691 ;
  assign n4693 = n4660 & n4692 ;
  assign n4694 = n4642 & n4693 ;
  assign n4695 = \u1_u2_adr_cw_reg[10]/P0001  & \u1_u2_adr_cw_reg[9]/NET0131  ;
  assign n4696 = \u1_u2_adr_cw_reg[8]/P0001  & n4695 ;
  assign n4697 = n4664 & n4696 ;
  assign n4698 = n4569 & n4697 ;
  assign n4699 = \u1_u2_adr_cw_reg[11]/P0001  & n4698 ;
  assign n4700 = ~\u1_u2_adr_cw_reg[12]/P0001  & ~\u1_u2_last_buf_adr_reg[12]/P0001  ;
  assign n4701 = ~n4699 & n4700 ;
  assign n4702 = \u1_u2_adr_cw_reg[11]/P0001  & ~\u1_u2_last_buf_adr_reg[12]/P0001  ;
  assign n4703 = \u1_u2_adr_cw_reg[12]/P0001  & n4702 ;
  assign n4704 = n4698 & n4703 ;
  assign n4705 = ~n4701 & ~n4704 ;
  assign n4706 = ~\u1_u2_adr_cw_reg[12]/P0001  & ~n4699 ;
  assign n4707 = \u1_u2_adr_cw_reg[11]/P0001  & \u1_u2_adr_cw_reg[12]/P0001  ;
  assign n4708 = n4698 & n4707 ;
  assign n4709 = \u1_u2_last_buf_adr_reg[12]/P0001  & ~n4708 ;
  assign n4710 = ~n4706 & n4709 ;
  assign n4711 = n4705 & ~n4710 ;
  assign n4712 = \u1_u2_adr_cw_reg[11]/P0001  & ~\u1_u2_last_buf_adr_reg[11]/P0001  ;
  assign n4713 = ~n4698 & n4712 ;
  assign n4714 = n4637 & n4696 ;
  assign n4715 = n4569 & n4714 ;
  assign n4716 = ~\u1_u2_adr_cw_reg[11]/P0001  & ~\u1_u2_last_buf_adr_reg[11]/P0001  ;
  assign n4717 = n4715 & n4716 ;
  assign n4718 = ~n4713 & ~n4717 ;
  assign n4719 = ~\u1_u2_adr_cw_reg[10]/P0001  & ~\u1_u2_last_buf_adr_reg[10]/P0001  ;
  assign n4720 = ~n4688 & n4719 ;
  assign n4721 = \u1_u2_adr_cw_reg[10]/P0001  & ~\u1_u2_last_buf_adr_reg[10]/P0001  ;
  assign n4722 = n4637 & n4686 ;
  assign n4723 = n4569 & n4722 ;
  assign n4724 = n4721 & n4723 ;
  assign n4725 = ~n4720 & ~n4724 ;
  assign n4726 = ~\u1_u2_adr_cw_reg[10]/P0001  & ~n4688 ;
  assign n4727 = \u1_u2_last_buf_adr_reg[10]/P0001  & ~n4698 ;
  assign n4728 = ~n4726 & n4727 ;
  assign n4729 = n4725 & ~n4728 ;
  assign n4730 = n4718 & ~n4729 ;
  assign n4731 = ~\u1_u2_adr_cw_reg[11]/P0001  & \u1_u2_last_buf_adr_reg[11]/P0001  ;
  assign n4732 = ~n4698 & n4731 ;
  assign n4733 = \u1_u2_adr_cw_reg[11]/P0001  & \u1_u2_last_buf_adr_reg[11]/P0001  ;
  assign n4734 = n4715 & n4733 ;
  assign n4735 = ~n4732 & ~n4734 ;
  assign n4736 = n4730 & n4735 ;
  assign n4737 = ~n4711 & n4736 ;
  assign n4738 = n4694 & n4737 ;
  assign n4739 = ~\u1_u2_adr_cw_reg[13]/P0001  & \u1_u2_last_buf_adr_reg[13]/P0001  ;
  assign n4740 = ~n4708 & n4739 ;
  assign n4741 = \u1_u2_adr_cw_reg[13]/P0001  & \u1_u2_last_buf_adr_reg[13]/P0001  ;
  assign n4742 = n4707 & n4741 ;
  assign n4743 = n4698 & n4742 ;
  assign n4744 = ~n4740 & ~n4743 ;
  assign n4745 = ~\u1_u2_adr_cw_reg[13]/P0001  & ~n4708 ;
  assign n4746 = \u1_u2_adr_cw_reg[11]/P0001  & \u1_u2_adr_cw_reg[13]/P0001  ;
  assign n4747 = \u1_u2_adr_cw_reg[12]/P0001  & n4746 ;
  assign n4748 = n4698 & n4747 ;
  assign n4749 = ~\u1_u2_last_buf_adr_reg[13]/P0001  & ~n4748 ;
  assign n4750 = ~n4745 & n4749 ;
  assign n4751 = \u1_u2_adr_cw_reg[14]/P0001  & ~\u1_u2_last_buf_adr_reg[14]/P0001  ;
  assign n4752 = ~n4748 & n4751 ;
  assign n4753 = ~\u1_u2_adr_cw_reg[14]/P0001  & ~\u1_u2_last_buf_adr_reg[14]/P0001  ;
  assign n4754 = n4747 & n4753 ;
  assign n4755 = n4698 & n4754 ;
  assign n4756 = ~n4752 & ~n4755 ;
  assign n4757 = ~\u1_u2_adr_cw_reg[14]/P0001  & \u1_u2_last_buf_adr_reg[14]/P0001  ;
  assign n4758 = ~n4748 & n4757 ;
  assign n4759 = \u1_u2_adr_cw_reg[14]/P0001  & \u1_u2_last_buf_adr_reg[14]/P0001  ;
  assign n4760 = n4748 & n4759 ;
  assign n4761 = ~n4758 & ~n4760 ;
  assign n4762 = n4756 & n4761 ;
  assign n4763 = ~n4750 & n4762 ;
  assign n4764 = n4744 & n4763 ;
  assign n4765 = n4738 & n4764 ;
  assign n4766 = ~\u1_u2_adr_cw_reg[0]/NET0131  & ~n4555 ;
  assign n4767 = ~n4578 & ~n4766 ;
  assign n4768 = n4023 & n4767 ;
  assign n4769 = ~n4765 & n4768 ;
  assign n4770 = ~n4028 & ~n4769 ;
  assign n4771 = \u1_u3_adr_reg[12]/P0001  & ~n4023 ;
  assign n4772 = ~n4698 & ~n4726 ;
  assign n4773 = n4023 & n4772 ;
  assign n4774 = ~n4765 & n4773 ;
  assign n4775 = ~n4771 & ~n4774 ;
  assign n4776 = \u1_u3_adr_reg[13]/P0001  & ~n4023 ;
  assign n4777 = \u1_u2_adr_cw_reg[11]/P0001  & ~n4698 ;
  assign n4778 = ~\u1_u2_adr_cw_reg[11]/P0001  & n4698 ;
  assign n4779 = ~n4777 & ~n4778 ;
  assign n4780 = n4023 & ~n4779 ;
  assign n4781 = ~n4765 & n4780 ;
  assign n4782 = ~n4776 & ~n4781 ;
  assign n4783 = \u1_u3_adr_reg[14]/P0001  & ~n4023 ;
  assign n4784 = ~n4706 & ~n4708 ;
  assign n4785 = n4023 & n4784 ;
  assign n4786 = ~n4765 & n4785 ;
  assign n4787 = ~n4783 & ~n4786 ;
  assign n4788 = \u1_u3_adr_reg[15]/P0001  & ~n4023 ;
  assign n4789 = ~n4745 & ~n4748 ;
  assign n4790 = n4023 & n4789 ;
  assign n4791 = ~n4765 & n4790 ;
  assign n4792 = ~n4788 & ~n4791 ;
  assign n4793 = \u1_u3_adr_reg[16]/P0001  & ~n4023 ;
  assign n4794 = \u1_u2_adr_cw_reg[14]/P0001  & ~n4748 ;
  assign n4795 = ~\u1_u2_adr_cw_reg[14]/P0001  & n4748 ;
  assign n4796 = ~n4794 & ~n4795 ;
  assign n4797 = n4023 & ~n4796 ;
  assign n4798 = ~n4765 & n4797 ;
  assign n4799 = ~n4793 & ~n4798 ;
  assign n4800 = \u1_u3_adr_reg[3]/P0001  & ~n4023 ;
  assign n4801 = ~n4557 & ~n4584 ;
  assign n4802 = n4023 & n4801 ;
  assign n4803 = ~n4765 & n4802 ;
  assign n4804 = ~n4800 & ~n4803 ;
  assign n4805 = \u1_u3_adr_reg[4]/P0001  & ~n4023 ;
  assign n4806 = ~\u1_u2_adr_cw_reg[2]/P0001  & n4557 ;
  assign n4807 = \u1_u2_adr_cw_reg[2]/P0001  & ~n4557 ;
  assign n4808 = ~n4806 & ~n4807 ;
  assign n4809 = n4023 & ~n4808 ;
  assign n4810 = ~n4765 & n4809 ;
  assign n4811 = ~n4805 & ~n4810 ;
  assign n4812 = \u1_u3_adr_reg[5]/P0001  & ~n4023 ;
  assign n4813 = ~n4559 & ~n4574 ;
  assign n4814 = n4023 & n4813 ;
  assign n4815 = ~n4765 & n4814 ;
  assign n4816 = ~n4812 & ~n4815 ;
  assign n4817 = \u1_u3_adr_reg[6]/P0001  & ~n4023 ;
  assign n4818 = ~n4566 & ~n4569 ;
  assign n4819 = n4023 & n4818 ;
  assign n4820 = ~n4765 & n4819 ;
  assign n4821 = ~n4817 & ~n4820 ;
  assign n4822 = \u1_u3_adr_reg[7]/P0001  & ~n4023 ;
  assign n4823 = \u1_u2_adr_cw_reg[5]/NET0131  & ~n4569 ;
  assign n4824 = ~\u1_u2_adr_cw_reg[5]/NET0131  & n4569 ;
  assign n4825 = ~n4823 & ~n4824 ;
  assign n4826 = n4023 & ~n4825 ;
  assign n4827 = ~n4765 & n4826 ;
  assign n4828 = ~n4822 & ~n4827 ;
  assign n4829 = \u1_u3_adr_reg[8]/P0001  & ~n4023 ;
  assign n4830 = ~n4635 & ~n4656 ;
  assign n4831 = n4023 & n4830 ;
  assign n4832 = ~n4765 & n4831 ;
  assign n4833 = ~n4829 & ~n4832 ;
  assign n4834 = \u1_u3_adr_reg[9]/P0001  & ~n4023 ;
  assign n4835 = ~n4636 & ~n4638 ;
  assign n4836 = n4023 & n4835 ;
  assign n4837 = ~n4765 & n4836 ;
  assign n4838 = ~n4834 & ~n4837 ;
  assign n4839 = \u1_u3_adr_reg[10]/P0001  & ~n4023 ;
  assign n4840 = \u1_u2_adr_cw_reg[8]/P0001  & ~n4638 ;
  assign n4841 = \u1_u2_adr_cw_reg[7]/NET0131  & ~\u1_u2_adr_cw_reg[8]/P0001  ;
  assign n4842 = n4634 & n4841 ;
  assign n4843 = n4569 & n4842 ;
  assign n4844 = ~n4840 & ~n4843 ;
  assign n4845 = n4023 & ~n4844 ;
  assign n4846 = ~n4765 & n4845 ;
  assign n4847 = ~n4839 & ~n4846 ;
  assign n4848 = \u1_u3_adr_reg[11]/P0001  & ~n4023 ;
  assign n4849 = ~n4685 & ~n4688 ;
  assign n4850 = n4023 & n4849 ;
  assign n4851 = ~n4765 & n4850 ;
  assign n4852 = ~n4848 & ~n4851 ;
  assign n4853 = ~n4471 & n4478 ;
  assign n4854 = ~n4472 & ~n4481 ;
  assign n4855 = ~n4853 & ~n4854 ;
  assign n4856 = n4478 & n4854 ;
  assign n4857 = ~n4471 & n4856 ;
  assign n4858 = ~n4855 & ~n4857 ;
  assign n4859 = \u0_tx_ready_reg/NET0131  & n1834 ;
  assign n4860 = n1838 & n4859 ;
  assign n4861 = rst_i_pad & ~n4860 ;
  assign n4862 = ~\u1_u1_send_zero_length_r_reg/P0001  & ~\u1_u1_state_reg[3]/NET0131  ;
  assign n4863 = n1829 & n4862 ;
  assign n4864 = n1750 & n1847 ;
  assign n4865 = n4863 & n4864 ;
  assign n4866 = n4861 & ~n4865 ;
  assign n4867 = n1848 & n4239 ;
  assign n4868 = \u1_u1_send_zero_length_r_reg/P0001  & n4867 ;
  assign n4869 = ~\u0_tx_ready_reg/NET0131  & ~n1839 ;
  assign n4870 = \u0_tx_ready_reg/NET0131  & ~n1851 ;
  assign n4871 = ~n4869 & ~n4870 ;
  assign n4872 = ~\u1_u1_send_zero_length_r_reg/P0001  & ~\u1_u1_zero_length_r_reg/P0001  ;
  assign n4873 = \u1_u1_send_data_r_reg/P0001  & ~\u1_u1_zero_length_r_reg/P0001  ;
  assign n4874 = ~n4872 & ~n4873 ;
  assign n4875 = ~\u1_u1_send_data_r_reg/P0001  & ~\u1_u1_send_zero_length_r_reg/P0001  ;
  assign n4876 = \u1_u2_send_data_r_reg/NET0131  & n4875 ;
  assign n4877 = rst_i_pad & ~n4876 ;
  assign n4878 = n4874 & n4877 ;
  assign n4879 = ~n4871 & n4878 ;
  assign n4880 = \u1_u3_out_to_small_r_reg/P0001  & \u4_buf0_reg[0]/P0001  ;
  assign n4881 = ~\u1_u3_buffer_done_reg/P0001  & ~\u4_csr_reg[30]/NET0131  ;
  assign n4882 = ~n4507 & ~n4881 ;
  assign n4883 = n4506 & n4882 ;
  assign n4884 = ~n4880 & ~n4883 ;
  assign n4885 = ~n4401 & ~n4884 ;
  assign n4886 = ~n3895 & ~n3972 ;
  assign n4887 = ~\u1_u3_adr_r_reg[0]/P0001  & ~n3967 ;
  assign n4888 = ~n4886 & n4887 ;
  assign n4889 = n4503 & ~n4888 ;
  assign n4890 = ~n4885 & ~n4889 ;
  assign n4891 = rst_i_pad & n4091 ;
  assign n4892 = ~n4090 & n4891 ;
  assign n4893 = n4088 & n4892 ;
  assign n4894 = rst_i_pad & \u1_u2_state_reg[1]/NET0131  ;
  assign n4895 = n4189 & n4894 ;
  assign n4896 = ~n4107 & n4895 ;
  assign n4897 = ~n4893 & ~n4896 ;
  assign n4898 = \u1_u2_state_reg[5]/NET0131  & ~n4091 ;
  assign n4899 = ~n4090 & ~n4898 ;
  assign n4900 = n4088 & ~n4899 ;
  assign n4901 = rst_i_pad & n4900 ;
  assign n4902 = \u1_u2_state_reg[5]/NET0131  & n4189 ;
  assign n4903 = rst_i_pad & n4902 ;
  assign n4904 = ~n4103 & n4903 ;
  assign n4905 = ~n4901 & ~n4904 ;
  assign n4906 = ~\u1_u3_state_reg[2]/P0001  & n2372 ;
  assign n4907 = ~\u1_u3_abort_reg/P0001  & ~\u1_u3_tx_data_to_reg/P0001  ;
  assign n4908 = ~\u1_u3_state_reg[0]/P0001  & n4907 ;
  assign n4909 = ~\u1_u0_state_reg[0]/P0001  & ~\u1_u0_state_reg[2]/P0001  ;
  assign n4910 = ~\u1_u0_state_reg[1]/P0001  & \u1_u0_state_reg[3]/P0001  ;
  assign n4911 = n4909 & n4910 ;
  assign n4912 = \u0_rx_active_reg/P0001  & ~\u0_rx_err_reg/P0001  ;
  assign n4913 = n4907 & ~n4912 ;
  assign n4914 = n4911 & n4913 ;
  assign n4915 = ~n4908 & ~n4914 ;
  assign n4916 = ~\u1_u3_state_reg[0]/P0001  & ~\u1_u3_state_reg[1]/P0001  ;
  assign n4917 = ~\u1_u3_state_reg[3]/P0001  & ~\u1_u3_state_reg[5]/P0001  ;
  assign n4918 = n4916 & n4917 ;
  assign n4919 = \u1_u3_state_reg[4]/P0001  & n4918 ;
  assign n4920 = n4915 & n4919 ;
  assign n4921 = ~\u1_u0_crc16_sum_reg[14]/P0001  & \u1_u0_crc16_sum_reg[15]/P0001  ;
  assign n4922 = \u1_u0_crc16_sum_reg[0]/P0001  & ~\u1_u0_crc16_sum_reg[1]/P0001  ;
  assign n4923 = n4921 & n4922 ;
  assign n4924 = ~\u1_u0_crc16_sum_reg[10]/P0001  & ~\u1_u0_crc16_sum_reg[11]/P0001  ;
  assign n4925 = ~\u1_u0_crc16_sum_reg[12]/P0001  & ~\u1_u0_crc16_sum_reg[13]/P0001  ;
  assign n4926 = n4924 & n4925 ;
  assign n4927 = n4923 & n4926 ;
  assign n4928 = ~\u1_u0_crc16_sum_reg[6]/P0001  & ~\u1_u0_crc16_sum_reg[7]/P0001  ;
  assign n4929 = ~\u1_u0_crc16_sum_reg[8]/P0001  & ~\u1_u0_crc16_sum_reg[9]/P0001  ;
  assign n4930 = n4928 & n4929 ;
  assign n4931 = ~\u1_u0_crc16_sum_reg[4]/P0001  & ~\u1_u0_crc16_sum_reg[5]/P0001  ;
  assign n4932 = \u1_u0_crc16_sum_reg[2]/P0001  & \u1_u0_crc16_sum_reg[3]/P0001  ;
  assign n4933 = n4931 & n4932 ;
  assign n4934 = n4930 & n4933 ;
  assign n4935 = n4927 & n4934 ;
  assign n4936 = n4911 & ~n4912 ;
  assign n4937 = n4919 & n4936 ;
  assign n4938 = ~n4935 & n4937 ;
  assign n4939 = ~n4920 & ~n4938 ;
  assign n4940 = n4906 & ~n4939 ;
  assign n4941 = ~\u1_u3_state_reg[0]/P0001  & \u1_u3_state_reg[1]/P0001  ;
  assign n4942 = n2376 & n4941 ;
  assign n4943 = n2371 & n4916 ;
  assign n4944 = n2375 & n4943 ;
  assign n4945 = ~\u1_u3_state_reg[7]/P0001  & \u1_u3_state_reg[9]/P0001  ;
  assign n4946 = n4944 & n4945 ;
  assign n4947 = n2370 & n2375 ;
  assign n4948 = ~\u1_u3_abort_reg/P0001  & ~\u1_u3_pid_seq_err_reg/P0001  ;
  assign n4949 = n2388 & n4948 ;
  assign n4950 = \u1_u3_state_reg[6]/P0001  & ~\u1_u3_state_reg[8]/P0001  ;
  assign n4951 = n4916 & n4950 ;
  assign n4952 = ~n4949 & n4951 ;
  assign n4953 = n4947 & n4952 ;
  assign n4954 = ~n4946 & ~n4953 ;
  assign n4955 = ~n4942 & n4954 ;
  assign n4956 = ~\u1_u3_rx_ack_to_reg/P0001  & ~\u1_u3_state_reg[0]/P0001  ;
  assign n4957 = ~\u1_u0_pid_reg[0]/NET0131  & \u1_u0_pid_reg[1]/NET0131  ;
  assign n4958 = n2354 & n4957 ;
  assign n4959 = \u1_u0_token_valid_str1_reg/P0001  & ~\u1_u3_rx_ack_to_reg/P0001  ;
  assign n4960 = n4958 & n4959 ;
  assign n4961 = ~n4956 & ~n4960 ;
  assign n4962 = \u1_u3_state_reg[3]/P0001  & ~\u1_u3_state_reg[5]/P0001  ;
  assign n4963 = ~\u1_u3_state_reg[2]/P0001  & ~\u1_u3_state_reg[4]/P0001  ;
  assign n4964 = n4916 & n4963 ;
  assign n4965 = n2372 & n4964 ;
  assign n4966 = n4962 & n4965 ;
  assign n4967 = n4961 & n4966 ;
  assign n4968 = ~\u1_u3_state_reg[3]/P0001  & \u1_u3_state_reg[5]/P0001  ;
  assign n4969 = \u1_u3_abort_reg/P0001  & n4968 ;
  assign n4970 = n4965 & n4969 ;
  assign n4971 = ~n4967 & ~n4970 ;
  assign n4972 = n4955 & n4971 ;
  assign n4973 = ~n4940 & n4972 ;
  assign n4974 = ~\u1_u0_token0_reg[2]/NET0131  & ~\u4_funct_adr_reg[2]/P0001  ;
  assign n4975 = \u1_u0_token0_reg[2]/NET0131  & \u4_funct_adr_reg[2]/P0001  ;
  assign n4976 = ~n4974 & ~n4975 ;
  assign n4977 = \u1_u0_token0_reg[3]/NET0131  & ~\u4_funct_adr_reg[3]/P0001  ;
  assign n4978 = \u1_u0_token_valid_str1_reg/P0001  & \u4_match_r1_reg/P0001  ;
  assign n4979 = ~n4977 & n4978 ;
  assign n4980 = ~n4976 & n4979 ;
  assign n4981 = n2351 & n3446 ;
  assign n4982 = ~n4958 & ~n4981 ;
  assign n4983 = n4980 & n4982 ;
  assign n4984 = \u1_u0_token0_reg[5]/NET0131  & ~\u4_funct_adr_reg[5]/P0001  ;
  assign n4985 = ~\u1_u0_token0_reg[5]/NET0131  & \u4_funct_adr_reg[5]/P0001  ;
  assign n4986 = ~n4984 & ~n4985 ;
  assign n4987 = ~\u1_u0_token0_reg[0]/NET0131  & \u4_funct_adr_reg[0]/P0001  ;
  assign n4988 = \u1_u0_token0_reg[4]/P0001  & ~\u4_funct_adr_reg[4]/P0001  ;
  assign n4989 = ~n4987 & ~n4988 ;
  assign n4990 = n4986 & n4989 ;
  assign n4991 = \u1_u0_token0_reg[1]/P0001  & ~\u4_funct_adr_reg[1]/P0001  ;
  assign n4992 = ~\u1_u0_token0_reg[6]/P0001  & \u4_funct_adr_reg[6]/P0001  ;
  assign n4993 = ~n4991 & ~n4992 ;
  assign n4994 = ~\u1_u0_token0_reg[1]/P0001  & \u4_funct_adr_reg[1]/P0001  ;
  assign n4995 = \u1_u0_token0_reg[6]/P0001  & ~\u4_funct_adr_reg[6]/P0001  ;
  assign n4996 = ~n4994 & ~n4995 ;
  assign n4997 = n4993 & n4996 ;
  assign n4998 = n4990 & n4997 ;
  assign n4999 = n4983 & n4998 ;
  assign n5000 = ~\u0_u0_mode_hs_reg/P0001  & n3447 ;
  assign n5001 = \u1_u0_token0_reg[0]/NET0131  & ~\u4_funct_adr_reg[0]/P0001  ;
  assign n5002 = ~\u1_u0_token0_reg[4]/P0001  & \u4_funct_adr_reg[4]/P0001  ;
  assign n5003 = ~\u1_u0_token0_reg[3]/NET0131  & \u4_funct_adr_reg[3]/P0001  ;
  assign n5004 = ~n5002 & ~n5003 ;
  assign n5005 = ~n5001 & n5004 ;
  assign n5006 = ~n5000 & n5005 ;
  assign n5007 = \u1_u0_pid_reg[2]/NET0131  & \u1_u0_pid_reg[3]/NET0131  ;
  assign n5008 = ~\u1_u0_pid_reg[1]/NET0131  & ~n5007 ;
  assign n5009 = ~\u1_u0_pid_reg[0]/NET0131  & ~n2354 ;
  assign n5010 = ~n5008 & n5009 ;
  assign n5011 = n5006 & ~n5010 ;
  assign n5012 = n4999 & n5011 ;
  assign n5013 = rst_i_pad & ~n5012 ;
  assign n5014 = \u1_u3_state_reg[0]/P0001  & ~\u1_u3_state_reg[1]/P0001  ;
  assign n5015 = n2376 & n5014 ;
  assign n5016 = n2350 & n5007 ;
  assign n5017 = ~n2355 & ~n5016 ;
  assign n5018 = ~n2352 & n2358 ;
  assign n5019 = n5017 & n5018 ;
  assign n5020 = \u4_csr_reg[26]/NET0131  & \u4_csr_reg[27]/NET0131  ;
  assign n5021 = ~n5019 & ~n5020 ;
  assign n5022 = ~n2382 & ~n5021 ;
  assign n5023 = n3451 & n5022 ;
  assign n5024 = n3454 & ~n5023 ;
  assign n5025 = n5015 & ~n5024 ;
  assign n5026 = n5013 & ~n5025 ;
  assign n5027 = \u1_u0_token0_reg[7]/P0001  & ~\u1_u0_token1_reg[2]/P0001  ;
  assign n5028 = ~\u1_u0_token0_reg[7]/P0001  & \u1_u0_token1_reg[2]/P0001  ;
  assign n5029 = ~n5027 & ~n5028 ;
  assign n5030 = \u1_u0_token1_reg[0]/P0001  & ~\u1_u0_token1_reg[5]/P0001  ;
  assign n5031 = ~\u1_u0_token1_reg[0]/P0001  & \u1_u0_token1_reg[5]/P0001  ;
  assign n5032 = ~n5030 & ~n5031 ;
  assign n5033 = ~\u1_u0_token0_reg[4]/P0001  & n5032 ;
  assign n5034 = \u1_u0_token0_reg[4]/P0001  & ~n5032 ;
  assign n5035 = ~n5033 & ~n5034 ;
  assign n5036 = ~n5029 & ~n5035 ;
  assign n5037 = n5029 & n5035 ;
  assign n5038 = ~n5036 & ~n5037 ;
  assign n5039 = \u1_u0_token0_reg[0]/NET0131  & ~\u1_u0_token0_reg[1]/P0001  ;
  assign n5040 = ~\u1_u0_token0_reg[0]/NET0131  & \u1_u0_token0_reg[1]/P0001  ;
  assign n5041 = ~n5039 & ~n5040 ;
  assign n5042 = \u1_u0_token0_reg[2]/NET0131  & ~\u1_u0_token0_reg[3]/NET0131  ;
  assign n5043 = ~\u1_u0_token0_reg[2]/NET0131  & \u1_u0_token0_reg[3]/NET0131  ;
  assign n5044 = ~n5042 & ~n5043 ;
  assign n5045 = ~n5041 & ~n5044 ;
  assign n5046 = n5041 & n5044 ;
  assign n5047 = ~n5045 & ~n5046 ;
  assign n5048 = ~n5038 & ~n5047 ;
  assign n5049 = ~\u1_u0_token0_reg[2]/NET0131  & n5041 ;
  assign n5050 = \u1_u0_token0_reg[2]/NET0131  & ~n5041 ;
  assign n5051 = ~n5049 & ~n5050 ;
  assign n5052 = ~\u1_u0_token0_reg[6]/P0001  & ~\u1_u0_token1_reg[0]/P0001  ;
  assign n5053 = \u1_u0_token0_reg[6]/P0001  & \u1_u0_token1_reg[0]/P0001  ;
  assign n5054 = ~n5052 & ~n5053 ;
  assign n5055 = \u1_u0_token0_reg[5]/NET0131  & ~\u1_u0_token1_reg[3]/P0001  ;
  assign n5056 = ~\u1_u0_token0_reg[5]/NET0131  & \u1_u0_token1_reg[3]/P0001  ;
  assign n5057 = ~n5055 & ~n5056 ;
  assign n5058 = n5054 & n5057 ;
  assign n5059 = ~n5051 & n5058 ;
  assign n5060 = n5054 & ~n5057 ;
  assign n5061 = n5051 & n5060 ;
  assign n5062 = ~n5059 & ~n5061 ;
  assign n5063 = ~n5048 & n5062 ;
  assign n5064 = ~\u1_u0_token0_reg[7]/P0001  & ~\u1_u0_token1_reg[1]/P0001  ;
  assign n5065 = \u1_u0_token0_reg[7]/P0001  & \u1_u0_token1_reg[1]/P0001  ;
  assign n5066 = ~n5064 & ~n5065 ;
  assign n5067 = \u1_u0_token0_reg[6]/P0001  & ~\u1_u0_token1_reg[4]/P0001  ;
  assign n5068 = ~\u1_u0_token0_reg[6]/P0001  & \u1_u0_token1_reg[4]/P0001  ;
  assign n5069 = ~n5067 & ~n5068 ;
  assign n5070 = n5066 & n5069 ;
  assign n5071 = ~n5066 & ~n5069 ;
  assign n5072 = ~n5070 & ~n5071 ;
  assign n5073 = n5047 & ~n5072 ;
  assign n5074 = ~n5054 & ~n5057 ;
  assign n5075 = ~n5051 & n5074 ;
  assign n5076 = ~n5054 & n5057 ;
  assign n5077 = n5051 & n5076 ;
  assign n5078 = ~n5075 & ~n5077 ;
  assign n5079 = ~n5073 & n5078 ;
  assign n5080 = n5063 & n5079 ;
  assign n5081 = \u1_u0_token0_reg[4]/P0001  & n5029 ;
  assign n5082 = ~\u1_u0_token0_reg[4]/P0001  & ~n5029 ;
  assign n5083 = ~n5081 & ~n5082 ;
  assign n5084 = \u1_u0_token0_reg[5]/NET0131  & ~\u1_u0_token1_reg[7]/P0001  ;
  assign n5085 = ~\u1_u0_token0_reg[5]/NET0131  & \u1_u0_token1_reg[7]/P0001  ;
  assign n5086 = ~n5084 & ~n5085 ;
  assign n5087 = ~n5041 & n5086 ;
  assign n5088 = ~n5083 & n5087 ;
  assign n5089 = n5041 & n5086 ;
  assign n5090 = n5083 & n5089 ;
  assign n5091 = ~n5088 & ~n5090 ;
  assign n5092 = ~n5041 & ~n5086 ;
  assign n5093 = n5083 & n5092 ;
  assign n5094 = n5041 & ~n5086 ;
  assign n5095 = ~n5083 & n5094 ;
  assign n5096 = ~n5093 & ~n5095 ;
  assign n5097 = n5091 & n5096 ;
  assign n5098 = \u1_u0_token1_reg[1]/P0001  & ~\u1_u0_token1_reg[6]/P0001  ;
  assign n5099 = ~\u1_u0_token1_reg[1]/P0001  & \u1_u0_token1_reg[6]/P0001  ;
  assign n5100 = ~n5098 & ~n5099 ;
  assign n5101 = ~\u1_u0_token0_reg[4]/P0001  & ~\u1_u0_token0_reg[6]/P0001  ;
  assign n5102 = \u1_u0_token0_reg[4]/P0001  & \u1_u0_token0_reg[6]/P0001  ;
  assign n5103 = ~n5101 & ~n5102 ;
  assign n5104 = ~\u1_u0_token0_reg[0]/NET0131  & ~\u1_u0_token0_reg[3]/NET0131  ;
  assign n5105 = \u1_u0_token0_reg[0]/NET0131  & \u1_u0_token0_reg[3]/NET0131  ;
  assign n5106 = ~n5104 & ~n5105 ;
  assign n5107 = n5103 & ~n5106 ;
  assign n5108 = ~n5103 & n5106 ;
  assign n5109 = ~n5107 & ~n5108 ;
  assign n5110 = ~n5100 & ~n5109 ;
  assign n5111 = n5100 & n5109 ;
  assign n5112 = ~n5110 & ~n5111 ;
  assign n5113 = n5038 & n5072 ;
  assign n5114 = ~n5112 & ~n5113 ;
  assign n5115 = ~n5097 & n5114 ;
  assign n5116 = n5080 & n5115 ;
  assign n5117 = rst_i_pad & \u1_u0_token_valid_str1_reg/P0001  ;
  assign n5118 = ~n5025 & n5117 ;
  assign n5119 = ~n5116 & n5118 ;
  assign n5120 = ~n5026 & ~n5119 ;
  assign n5121 = n4973 & ~n5120 ;
  assign n5122 = ~\u0_tx_ready_reg/NET0131  & \u1_u1_send_token_r_reg/P0001  ;
  assign n5123 = ~\u1_u3_send_token_reg/P0001  & ~n5122 ;
  assign n5124 = rst_i_pad & ~n5123 ;
  assign n5125 = ~\u1_u3_send_token_reg/P0001  & n1750 ;
  assign n5126 = ~\u1_u0_token1_reg[1]/P0001  & \u4_u0_csr1_reg[5]/P0001  ;
  assign n5127 = ~\u1_u0_token0_reg[7]/P0001  & \u4_u0_csr1_reg[3]/P0001  ;
  assign n5128 = ~n5126 & ~n5127 ;
  assign n5129 = \u1_u0_token1_reg[1]/P0001  & ~\u4_u0_csr1_reg[5]/P0001  ;
  assign n5130 = \u1_u0_token0_reg[7]/P0001  & ~\u4_u0_csr1_reg[3]/P0001  ;
  assign n5131 = ~n5129 & ~n5130 ;
  assign n5132 = n5128 & n5131 ;
  assign n5133 = ~\u1_u0_token1_reg[0]/P0001  & ~\u4_u0_csr1_reg[4]/P0001  ;
  assign n5134 = \u1_u0_token1_reg[0]/P0001  & \u4_u0_csr1_reg[4]/P0001  ;
  assign n5135 = ~n5133 & ~n5134 ;
  assign n5136 = ~\u1_u0_token1_reg[2]/P0001  & ~\u4_u0_csr1_reg[6]/P0001  ;
  assign n5137 = \u1_u0_token1_reg[2]/P0001  & \u4_u0_csr1_reg[6]/P0001  ;
  assign n5138 = ~n5136 & ~n5137 ;
  assign n5139 = ~n5135 & ~n5138 ;
  assign n5140 = n5132 & n5139 ;
  assign n5141 = ~\u1_u0_token1_reg[2]/P0001  & \u4_u1_csr1_reg[6]/P0001  ;
  assign n5142 = ~\u1_u0_token0_reg[7]/P0001  & \u4_u1_csr1_reg[3]/P0001  ;
  assign n5143 = ~n5141 & ~n5142 ;
  assign n5144 = \u1_u0_token1_reg[2]/P0001  & ~\u4_u1_csr1_reg[6]/P0001  ;
  assign n5145 = \u1_u0_token0_reg[7]/P0001  & ~\u4_u1_csr1_reg[3]/P0001  ;
  assign n5146 = ~n5144 & ~n5145 ;
  assign n5147 = n5143 & n5146 ;
  assign n5148 = ~\u1_u0_token1_reg[0]/P0001  & ~\u4_u1_csr1_reg[4]/P0001  ;
  assign n5149 = \u1_u0_token1_reg[0]/P0001  & \u4_u1_csr1_reg[4]/P0001  ;
  assign n5150 = ~n5148 & ~n5149 ;
  assign n5151 = ~\u1_u0_token1_reg[1]/P0001  & ~\u4_u1_csr1_reg[5]/P0001  ;
  assign n5152 = \u1_u0_token1_reg[1]/P0001  & \u4_u1_csr1_reg[5]/P0001  ;
  assign n5153 = ~n5151 & ~n5152 ;
  assign n5154 = ~n5150 & ~n5153 ;
  assign n5155 = n5147 & n5154 ;
  assign n5156 = ~n5140 & ~n5155 ;
  assign n5157 = ~\u1_u0_token1_reg[2]/P0001  & \u4_u2_csr1_reg[6]/P0001  ;
  assign n5158 = ~\u1_u0_token0_reg[7]/P0001  & \u4_u2_csr1_reg[3]/P0001  ;
  assign n5159 = ~n5157 & ~n5158 ;
  assign n5160 = \u1_u0_token1_reg[2]/P0001  & ~\u4_u2_csr1_reg[6]/P0001  ;
  assign n5161 = \u1_u0_token0_reg[7]/P0001  & ~\u4_u2_csr1_reg[3]/P0001  ;
  assign n5162 = ~n5160 & ~n5161 ;
  assign n5163 = n5159 & n5162 ;
  assign n5164 = ~\u1_u0_token1_reg[0]/P0001  & ~\u4_u2_csr1_reg[4]/P0001  ;
  assign n5165 = \u1_u0_token1_reg[0]/P0001  & \u4_u2_csr1_reg[4]/P0001  ;
  assign n5166 = ~n5164 & ~n5165 ;
  assign n5167 = ~\u1_u0_token1_reg[1]/P0001  & ~\u4_u2_csr1_reg[5]/P0001  ;
  assign n5168 = \u1_u0_token1_reg[1]/P0001  & \u4_u2_csr1_reg[5]/P0001  ;
  assign n5169 = ~n5167 & ~n5168 ;
  assign n5170 = ~n5166 & ~n5169 ;
  assign n5171 = n5163 & n5170 ;
  assign n5172 = \u4_u2_dma_out_buf_avail_reg/P0001  & n5171 ;
  assign n5173 = n5156 & n5172 ;
  assign n5174 = \u4_u0_dma_out_buf_avail_reg/P0001  & n5140 ;
  assign n5175 = ~n5140 & n5155 ;
  assign n5176 = \u4_u1_dma_out_buf_avail_reg/P0001  & n5175 ;
  assign n5177 = ~n5174 & ~n5176 ;
  assign n5178 = ~n5173 & n5177 ;
  assign n5179 = ~\u1_u0_token1_reg[2]/P0001  & \u4_u3_csr1_reg[6]/P0001  ;
  assign n5180 = ~\u1_u0_token0_reg[7]/P0001  & \u4_u3_csr1_reg[3]/P0001  ;
  assign n5181 = ~n5179 & ~n5180 ;
  assign n5182 = \u1_u0_token1_reg[2]/P0001  & ~\u4_u3_csr1_reg[6]/P0001  ;
  assign n5183 = \u1_u0_token0_reg[7]/P0001  & ~\u4_u3_csr1_reg[3]/P0001  ;
  assign n5184 = ~n5182 & ~n5183 ;
  assign n5185 = n5181 & n5184 ;
  assign n5186 = ~\u1_u0_token1_reg[1]/P0001  & ~\u4_u3_csr1_reg[5]/P0001  ;
  assign n5187 = \u1_u0_token1_reg[1]/P0001  & \u4_u3_csr1_reg[5]/P0001  ;
  assign n5188 = ~n5186 & ~n5187 ;
  assign n5189 = ~\u1_u0_token1_reg[0]/P0001  & ~\u4_u3_csr1_reg[4]/P0001  ;
  assign n5190 = \u1_u0_token1_reg[0]/P0001  & \u4_u3_csr1_reg[4]/P0001  ;
  assign n5191 = ~n5189 & ~n5190 ;
  assign n5192 = ~n5188 & ~n5191 ;
  assign n5193 = n5185 & n5192 ;
  assign n5194 = ~n5171 & n5193 ;
  assign n5195 = n5156 & n5194 ;
  assign n5196 = \u4_u3_dma_out_buf_avail_reg/P0001  & n5195 ;
  assign n5197 = ~n5171 & ~n5193 ;
  assign n5198 = n5156 & n5197 ;
  assign n5199 = \u4_dma_out_buf_avail_reg/P0001  & n5198 ;
  assign n5200 = ~n5196 & ~n5199 ;
  assign n5201 = n5178 & n5200 ;
  assign n5202 = ~\u4_u2_buf0_orig_m3_reg[11]/P0001  & \u4_u2_dma_in_cnt_reg[11]/P0001  ;
  assign n5203 = \u4_u2_buf0_orig_m3_reg[11]/P0001  & ~\u4_u2_dma_in_cnt_reg[11]/P0001  ;
  assign n5204 = ~\u4_u2_buf0_orig_m3_reg[10]/P0001  & \u4_u2_dma_in_cnt_reg[10]/P0001  ;
  assign n5205 = ~n5203 & n5204 ;
  assign n5206 = ~n5202 & ~n5205 ;
  assign n5207 = \u4_u2_buf0_orig_m3_reg[9]/P0001  & ~\u4_u2_dma_in_cnt_reg[9]/P0001  ;
  assign n5208 = \u4_u2_buf0_orig_m3_reg[10]/P0001  & ~\u4_u2_dma_in_cnt_reg[10]/P0001  ;
  assign n5209 = ~n5207 & ~n5208 ;
  assign n5210 = ~n5203 & n5209 ;
  assign n5211 = n5206 & ~n5210 ;
  assign n5212 = \u4_u2_buf0_orig_m3_reg[8]/P0001  & ~\u4_u2_dma_in_cnt_reg[8]/P0001  ;
  assign n5213 = \u4_u2_buf0_orig_m3_reg[7]/P0001  & ~\u4_u2_dma_in_cnt_reg[7]/P0001  ;
  assign n5214 = ~n5212 & ~n5213 ;
  assign n5215 = ~\u4_u2_buf0_orig_m3_reg[7]/P0001  & \u4_u2_dma_in_cnt_reg[7]/P0001  ;
  assign n5216 = ~\u4_u2_buf0_orig_m3_reg[6]/P0001  & \u4_u2_dma_in_cnt_reg[6]/P0001  ;
  assign n5217 = ~n5215 & ~n5216 ;
  assign n5218 = n5214 & ~n5217 ;
  assign n5219 = ~\u4_u2_buf0_orig_m3_reg[5]/P0001  & \u4_u2_dma_in_cnt_reg[5]/P0001  ;
  assign n5220 = ~\u4_u2_buf0_orig_m3_reg[4]/P0001  & \u4_u2_dma_in_cnt_reg[4]/P0001  ;
  assign n5221 = ~n5219 & ~n5220 ;
  assign n5222 = \u4_u2_buf0_orig_m3_reg[3]/P0001  & ~\u4_u2_dma_in_cnt_reg[3]/P0001  ;
  assign n5223 = \u4_u2_buf0_orig_m3_reg[4]/P0001  & ~\u4_u2_dma_in_cnt_reg[4]/P0001  ;
  assign n5224 = ~n5222 & ~n5223 ;
  assign n5225 = n5221 & ~n5224 ;
  assign n5226 = ~\u4_u2_buf0_orig_m3_reg[1]/P0001  & \u4_u2_dma_in_cnt_reg[1]/P0001  ;
  assign n5227 = \u4_u2_buf0_orig_m3_reg[0]/P0001  & ~\u4_u2_dma_in_cnt_reg[0]/P0001  ;
  assign n5228 = ~n5226 & n5227 ;
  assign n5229 = \u4_u2_buf0_orig_m3_reg[2]/P0001  & ~\u4_u2_dma_in_cnt_reg[2]/P0001  ;
  assign n5230 = \u4_u2_buf0_orig_m3_reg[1]/P0001  & ~\u4_u2_dma_in_cnt_reg[1]/P0001  ;
  assign n5231 = ~n5229 & ~n5230 ;
  assign n5232 = ~n5228 & n5231 ;
  assign n5233 = ~\u4_u2_buf0_orig_m3_reg[3]/P0001  & \u4_u2_dma_in_cnt_reg[3]/P0001  ;
  assign n5234 = ~\u4_u2_buf0_orig_m3_reg[2]/P0001  & \u4_u2_dma_in_cnt_reg[2]/P0001  ;
  assign n5235 = ~n5233 & ~n5234 ;
  assign n5236 = n5221 & n5235 ;
  assign n5237 = ~n5232 & n5236 ;
  assign n5238 = ~n5225 & ~n5237 ;
  assign n5239 = \u4_u2_buf0_orig_m3_reg[5]/P0001  & ~\u4_u2_dma_in_cnt_reg[5]/P0001  ;
  assign n5240 = \u4_u2_buf0_orig_m3_reg[6]/P0001  & ~\u4_u2_dma_in_cnt_reg[6]/P0001  ;
  assign n5241 = ~n5239 & ~n5240 ;
  assign n5242 = n5214 & n5241 ;
  assign n5243 = n5238 & n5242 ;
  assign n5244 = ~n5218 & ~n5243 ;
  assign n5245 = ~\u4_u2_buf0_orig_m3_reg[8]/P0001  & \u4_u2_dma_in_cnt_reg[8]/P0001  ;
  assign n5246 = ~\u4_u2_buf0_orig_m3_reg[9]/P0001  & \u4_u2_dma_in_cnt_reg[9]/P0001  ;
  assign n5247 = ~n5245 & ~n5246 ;
  assign n5248 = n5206 & n5247 ;
  assign n5249 = n5244 & n5248 ;
  assign n5250 = ~n5211 & ~n5249 ;
  assign n5251 = ~\u4_u3_buf0_orig_m3_reg[11]/P0001  & \u4_u3_dma_in_cnt_reg[11]/P0001  ;
  assign n5252 = \u4_u3_buf0_orig_m3_reg[11]/P0001  & ~\u4_u3_dma_in_cnt_reg[11]/P0001  ;
  assign n5253 = ~\u4_u3_buf0_orig_m3_reg[10]/P0001  & \u4_u3_dma_in_cnt_reg[10]/P0001  ;
  assign n5254 = ~n5252 & n5253 ;
  assign n5255 = ~n5251 & ~n5254 ;
  assign n5256 = \u4_u3_buf0_orig_m3_reg[9]/P0001  & ~\u4_u3_dma_in_cnt_reg[9]/P0001  ;
  assign n5257 = \u4_u3_buf0_orig_m3_reg[10]/P0001  & ~\u4_u3_dma_in_cnt_reg[10]/P0001  ;
  assign n5258 = ~n5256 & ~n5257 ;
  assign n5259 = ~n5252 & n5258 ;
  assign n5260 = n5255 & ~n5259 ;
  assign n5261 = \u4_u3_buf0_orig_m3_reg[8]/P0001  & ~\u4_u3_dma_in_cnt_reg[8]/P0001  ;
  assign n5262 = \u4_u3_buf0_orig_m3_reg[7]/P0001  & ~\u4_u3_dma_in_cnt_reg[7]/P0001  ;
  assign n5263 = ~n5261 & ~n5262 ;
  assign n5264 = ~\u4_u3_buf0_orig_m3_reg[7]/P0001  & \u4_u3_dma_in_cnt_reg[7]/P0001  ;
  assign n5265 = ~\u4_u3_buf0_orig_m3_reg[6]/P0001  & \u4_u3_dma_in_cnt_reg[6]/P0001  ;
  assign n5266 = ~n5264 & ~n5265 ;
  assign n5267 = n5263 & ~n5266 ;
  assign n5268 = ~\u4_u3_buf0_orig_m3_reg[5]/P0001  & \u4_u3_dma_in_cnt_reg[5]/P0001  ;
  assign n5269 = ~\u4_u3_buf0_orig_m3_reg[4]/P0001  & \u4_u3_dma_in_cnt_reg[4]/P0001  ;
  assign n5270 = ~n5268 & ~n5269 ;
  assign n5271 = \u4_u3_buf0_orig_m3_reg[3]/P0001  & ~\u4_u3_dma_in_cnt_reg[3]/P0001  ;
  assign n5272 = \u4_u3_buf0_orig_m3_reg[4]/P0001  & ~\u4_u3_dma_in_cnt_reg[4]/P0001  ;
  assign n5273 = ~n5271 & ~n5272 ;
  assign n5274 = n5270 & ~n5273 ;
  assign n5275 = ~\u4_u3_buf0_orig_m3_reg[1]/P0001  & \u4_u3_dma_in_cnt_reg[1]/P0001  ;
  assign n5276 = \u4_u3_buf0_orig_m3_reg[0]/P0001  & ~\u4_u3_dma_in_cnt_reg[0]/P0001  ;
  assign n5277 = ~n5275 & n5276 ;
  assign n5278 = \u4_u3_buf0_orig_m3_reg[2]/P0001  & ~\u4_u3_dma_in_cnt_reg[2]/P0001  ;
  assign n5279 = \u4_u3_buf0_orig_m3_reg[1]/P0001  & ~\u4_u3_dma_in_cnt_reg[1]/P0001  ;
  assign n5280 = ~n5278 & ~n5279 ;
  assign n5281 = ~n5277 & n5280 ;
  assign n5282 = ~\u4_u3_buf0_orig_m3_reg[3]/P0001  & \u4_u3_dma_in_cnt_reg[3]/P0001  ;
  assign n5283 = ~\u4_u3_buf0_orig_m3_reg[2]/P0001  & \u4_u3_dma_in_cnt_reg[2]/P0001  ;
  assign n5284 = ~n5282 & ~n5283 ;
  assign n5285 = n5270 & n5284 ;
  assign n5286 = ~n5281 & n5285 ;
  assign n5287 = ~n5274 & ~n5286 ;
  assign n5288 = \u4_u3_buf0_orig_m3_reg[5]/P0001  & ~\u4_u3_dma_in_cnt_reg[5]/P0001  ;
  assign n5289 = \u4_u3_buf0_orig_m3_reg[6]/P0001  & ~\u4_u3_dma_in_cnt_reg[6]/P0001  ;
  assign n5290 = ~n5288 & ~n5289 ;
  assign n5291 = n5263 & n5290 ;
  assign n5292 = n5287 & n5291 ;
  assign n5293 = ~n5267 & ~n5292 ;
  assign n5294 = ~\u4_u3_buf0_orig_m3_reg[8]/P0001  & \u4_u3_dma_in_cnt_reg[8]/P0001  ;
  assign n5295 = ~\u4_u3_buf0_orig_m3_reg[9]/P0001  & \u4_u3_dma_in_cnt_reg[9]/P0001  ;
  assign n5296 = ~n5294 & ~n5295 ;
  assign n5297 = n5255 & n5296 ;
  assign n5298 = n5293 & n5297 ;
  assign n5299 = ~n5260 & ~n5298 ;
  assign n5300 = ~\u4_u0_buf0_orig_m3_reg[11]/P0001  & \u4_u0_dma_in_cnt_reg[11]/P0001  ;
  assign n5301 = \u4_u0_buf0_orig_m3_reg[11]/P0001  & ~\u4_u0_dma_in_cnt_reg[11]/P0001  ;
  assign n5302 = ~\u4_u0_buf0_orig_m3_reg[10]/P0001  & \u4_u0_dma_in_cnt_reg[10]/P0001  ;
  assign n5303 = ~n5301 & n5302 ;
  assign n5304 = ~n5300 & ~n5303 ;
  assign n5305 = \u4_u0_buf0_orig_m3_reg[9]/P0001  & ~\u4_u0_dma_in_cnt_reg[9]/P0001  ;
  assign n5306 = \u4_u0_buf0_orig_m3_reg[10]/P0001  & ~\u4_u0_dma_in_cnt_reg[10]/P0001  ;
  assign n5307 = ~n5305 & ~n5306 ;
  assign n5308 = ~n5301 & n5307 ;
  assign n5309 = n5304 & ~n5308 ;
  assign n5310 = \u4_u0_buf0_orig_m3_reg[8]/P0001  & ~\u4_u0_dma_in_cnt_reg[8]/P0001  ;
  assign n5311 = \u4_u0_buf0_orig_m3_reg[7]/P0001  & ~\u4_u0_dma_in_cnt_reg[7]/P0001  ;
  assign n5312 = ~n5310 & ~n5311 ;
  assign n5313 = ~\u4_u0_buf0_orig_m3_reg[7]/P0001  & \u4_u0_dma_in_cnt_reg[7]/P0001  ;
  assign n5314 = ~\u4_u0_buf0_orig_m3_reg[6]/P0001  & \u4_u0_dma_in_cnt_reg[6]/P0001  ;
  assign n5315 = ~n5313 & ~n5314 ;
  assign n5316 = n5312 & ~n5315 ;
  assign n5317 = ~\u4_u0_buf0_orig_m3_reg[5]/P0001  & \u4_u0_dma_in_cnt_reg[5]/P0001  ;
  assign n5318 = ~\u4_u0_buf0_orig_m3_reg[4]/P0001  & \u4_u0_dma_in_cnt_reg[4]/P0001  ;
  assign n5319 = ~n5317 & ~n5318 ;
  assign n5320 = \u4_u0_buf0_orig_m3_reg[3]/P0001  & ~\u4_u0_dma_in_cnt_reg[3]/P0001  ;
  assign n5321 = \u4_u0_buf0_orig_m3_reg[4]/P0001  & ~\u4_u0_dma_in_cnt_reg[4]/P0001  ;
  assign n5322 = ~n5320 & ~n5321 ;
  assign n5323 = n5319 & ~n5322 ;
  assign n5324 = ~\u4_u0_buf0_orig_m3_reg[1]/P0001  & \u4_u0_dma_in_cnt_reg[1]/P0001  ;
  assign n5325 = \u4_u0_buf0_orig_m3_reg[0]/P0001  & ~\u4_u0_dma_in_cnt_reg[0]/P0001  ;
  assign n5326 = ~n5324 & n5325 ;
  assign n5327 = \u4_u0_buf0_orig_m3_reg[2]/P0001  & ~\u4_u0_dma_in_cnt_reg[2]/P0001  ;
  assign n5328 = \u4_u0_buf0_orig_m3_reg[1]/P0001  & ~\u4_u0_dma_in_cnt_reg[1]/P0001  ;
  assign n5329 = ~n5327 & ~n5328 ;
  assign n5330 = ~n5326 & n5329 ;
  assign n5331 = ~\u4_u0_buf0_orig_m3_reg[3]/P0001  & \u4_u0_dma_in_cnt_reg[3]/P0001  ;
  assign n5332 = ~\u4_u0_buf0_orig_m3_reg[2]/P0001  & \u4_u0_dma_in_cnt_reg[2]/P0001  ;
  assign n5333 = ~n5331 & ~n5332 ;
  assign n5334 = n5319 & n5333 ;
  assign n5335 = ~n5330 & n5334 ;
  assign n5336 = ~n5323 & ~n5335 ;
  assign n5337 = \u4_u0_buf0_orig_m3_reg[5]/P0001  & ~\u4_u0_dma_in_cnt_reg[5]/P0001  ;
  assign n5338 = \u4_u0_buf0_orig_m3_reg[6]/P0001  & ~\u4_u0_dma_in_cnt_reg[6]/P0001  ;
  assign n5339 = ~n5337 & ~n5338 ;
  assign n5340 = n5312 & n5339 ;
  assign n5341 = n5336 & n5340 ;
  assign n5342 = ~n5316 & ~n5341 ;
  assign n5343 = ~\u4_u0_buf0_orig_m3_reg[8]/P0001  & \u4_u0_dma_in_cnt_reg[8]/P0001  ;
  assign n5344 = ~\u4_u0_buf0_orig_m3_reg[9]/P0001  & \u4_u0_dma_in_cnt_reg[9]/P0001  ;
  assign n5345 = ~n5343 & ~n5344 ;
  assign n5346 = n5304 & n5345 ;
  assign n5347 = n5342 & n5346 ;
  assign n5348 = ~n5309 & ~n5347 ;
  assign n5349 = ~\u4_u1_buf0_orig_m3_reg[11]/P0001  & \u4_u1_dma_in_cnt_reg[11]/P0001  ;
  assign n5350 = \u4_u1_buf0_orig_m3_reg[11]/P0001  & ~\u4_u1_dma_in_cnt_reg[11]/P0001  ;
  assign n5351 = ~\u4_u1_buf0_orig_m3_reg[10]/P0001  & \u4_u1_dma_in_cnt_reg[10]/P0001  ;
  assign n5352 = ~n5350 & n5351 ;
  assign n5353 = ~n5349 & ~n5352 ;
  assign n5354 = \u4_u1_buf0_orig_m3_reg[9]/P0001  & ~\u4_u1_dma_in_cnt_reg[9]/P0001  ;
  assign n5355 = \u4_u1_buf0_orig_m3_reg[10]/P0001  & ~\u4_u1_dma_in_cnt_reg[10]/P0001  ;
  assign n5356 = ~n5354 & ~n5355 ;
  assign n5357 = ~n5350 & n5356 ;
  assign n5358 = n5353 & ~n5357 ;
  assign n5359 = \u4_u1_buf0_orig_m3_reg[8]/P0001  & ~\u4_u1_dma_in_cnt_reg[8]/P0001  ;
  assign n5360 = \u4_u1_buf0_orig_m3_reg[7]/P0001  & ~\u4_u1_dma_in_cnt_reg[7]/P0001  ;
  assign n5361 = ~n5359 & ~n5360 ;
  assign n5362 = ~\u4_u1_buf0_orig_m3_reg[7]/P0001  & \u4_u1_dma_in_cnt_reg[7]/P0001  ;
  assign n5363 = ~\u4_u1_buf0_orig_m3_reg[6]/P0001  & \u4_u1_dma_in_cnt_reg[6]/P0001  ;
  assign n5364 = ~n5362 & ~n5363 ;
  assign n5365 = n5361 & ~n5364 ;
  assign n5366 = ~\u4_u1_buf0_orig_m3_reg[5]/P0001  & \u4_u1_dma_in_cnt_reg[5]/P0001  ;
  assign n5367 = ~\u4_u1_buf0_orig_m3_reg[4]/P0001  & \u4_u1_dma_in_cnt_reg[4]/P0001  ;
  assign n5368 = ~n5366 & ~n5367 ;
  assign n5369 = \u4_u1_buf0_orig_m3_reg[3]/P0001  & ~\u4_u1_dma_in_cnt_reg[3]/P0001  ;
  assign n5370 = \u4_u1_buf0_orig_m3_reg[4]/P0001  & ~\u4_u1_dma_in_cnt_reg[4]/P0001  ;
  assign n5371 = ~n5369 & ~n5370 ;
  assign n5372 = n5368 & ~n5371 ;
  assign n5373 = ~\u4_u1_buf0_orig_m3_reg[1]/P0001  & \u4_u1_dma_in_cnt_reg[1]/P0001  ;
  assign n5374 = \u4_u1_buf0_orig_m3_reg[0]/P0001  & ~\u4_u1_dma_in_cnt_reg[0]/P0001  ;
  assign n5375 = ~n5373 & n5374 ;
  assign n5376 = \u4_u1_buf0_orig_m3_reg[2]/P0001  & ~\u4_u1_dma_in_cnt_reg[2]/P0001  ;
  assign n5377 = \u4_u1_buf0_orig_m3_reg[1]/P0001  & ~\u4_u1_dma_in_cnt_reg[1]/P0001  ;
  assign n5378 = ~n5376 & ~n5377 ;
  assign n5379 = ~n5375 & n5378 ;
  assign n5380 = ~\u4_u1_buf0_orig_m3_reg[3]/P0001  & \u4_u1_dma_in_cnt_reg[3]/P0001  ;
  assign n5381 = ~\u4_u1_buf0_orig_m3_reg[2]/P0001  & \u4_u1_dma_in_cnt_reg[2]/P0001  ;
  assign n5382 = ~n5380 & ~n5381 ;
  assign n5383 = n5368 & n5382 ;
  assign n5384 = ~n5379 & n5383 ;
  assign n5385 = ~n5372 & ~n5384 ;
  assign n5386 = \u4_u1_buf0_orig_m3_reg[5]/P0001  & ~\u4_u1_dma_in_cnt_reg[5]/P0001  ;
  assign n5387 = \u4_u1_buf0_orig_m3_reg[6]/P0001  & ~\u4_u1_dma_in_cnt_reg[6]/P0001  ;
  assign n5388 = ~n5386 & ~n5387 ;
  assign n5389 = n5361 & n5388 ;
  assign n5390 = n5385 & n5389 ;
  assign n5391 = ~n5365 & ~n5390 ;
  assign n5392 = ~\u4_u1_buf0_orig_m3_reg[8]/P0001  & \u4_u1_dma_in_cnt_reg[8]/P0001  ;
  assign n5393 = ~\u4_u1_buf0_orig_m3_reg[9]/P0001  & \u4_u1_dma_in_cnt_reg[9]/P0001  ;
  assign n5394 = ~n5392 & ~n5393 ;
  assign n5395 = n5353 & n5394 ;
  assign n5396 = n5391 & n5395 ;
  assign n5397 = ~n5358 & ~n5396 ;
  assign n5398 = ~n5116 & n5117 ;
  assign n5399 = ~n5013 & ~n5398 ;
  assign n5400 = \u1_u3_state_reg[2]/P0001  & ~\u1_u3_state_reg[4]/P0001  ;
  assign n5401 = n2372 & n5400 ;
  assign n5402 = ~\u1_u2_idma_done_reg/P0001  & n4918 ;
  assign n5403 = n5401 & n5402 ;
  assign n5404 = n3451 & n3458 ;
  assign n5405 = n5015 & n5404 ;
  assign n5406 = ~\u4_csr_reg[27]/NET0131  & n5017 ;
  assign n5407 = ~\u4_csr_reg[26]/NET0131  & ~n5406 ;
  assign n5408 = ~n2382 & ~n5407 ;
  assign n5409 = n3451 & n5408 ;
  assign n5410 = n3454 & ~n5409 ;
  assign n5411 = \u1_u3_state_reg[2]/P0001  & n5015 ;
  assign n5412 = ~n5410 & n5411 ;
  assign n5413 = ~n5405 & ~n5412 ;
  assign n5414 = ~n5403 & n5413 ;
  assign n5415 = ~n5399 & ~n5414 ;
  assign n5416 = ~n2382 & ~n3457 ;
  assign n5417 = n3451 & n5416 ;
  assign n5418 = n3454 & ~n5417 ;
  assign n5419 = \u1_u3_match_r_reg/P0001  & ~\u4_csr_reg[26]/NET0131  ;
  assign n5420 = ~n2383 & n5419 ;
  assign n5421 = ~n2379 & n5420 ;
  assign n5422 = ~\u1_u3_state_reg[4]/P0001  & ~n5421 ;
  assign n5423 = ~\u1_u3_state_reg[4]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n5424 = n5017 & n5423 ;
  assign n5425 = ~n5422 & ~n5424 ;
  assign n5426 = n5015 & n5425 ;
  assign n5427 = ~n5418 & n5426 ;
  assign n5428 = ~n4935 & n4936 ;
  assign n5429 = n4906 & n4919 ;
  assign n5430 = n4907 & n5429 ;
  assign n5431 = ~n5428 & n5430 ;
  assign n5432 = \u1_u3_state_reg[4]/P0001  & ~n4936 ;
  assign n5433 = n5431 & n5432 ;
  assign n5434 = ~n5427 & ~n5433 ;
  assign n5435 = ~n5399 & ~n5434 ;
  assign n5436 = ~n2382 & n3451 ;
  assign n5437 = \u1_u3_state_reg[1]/P0001  & ~n5021 ;
  assign n5438 = n5436 & ~n5437 ;
  assign n5439 = n3454 & n5015 ;
  assign n5440 = ~n5438 & n5439 ;
  assign n5441 = n5013 & n5440 ;
  assign n5442 = n5117 & n5440 ;
  assign n5443 = ~n5116 & n5442 ;
  assign n5444 = ~n5441 & ~n5443 ;
  assign n5445 = ~n2423 & ~n2424 ;
  assign n5446 = n2381 & n2384 ;
  assign n5447 = ~n3451 & n5446 ;
  assign n5448 = n5445 & ~n5447 ;
  assign n5449 = \u1_u3_int_upid_set_reg/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n5450 = ~\u4_u2_int_stat_reg[2]/P0001  & ~n5449 ;
  assign n5451 = rst_i_pad & ~\u4_u2_int_re_reg/P0001  ;
  assign n5452 = ~n5450 & n5451 ;
  assign n5453 = \u1_u3_int_upid_set_reg/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n5454 = ~\u4_u3_int_stat_reg[2]/P0001  & ~n5453 ;
  assign n5455 = rst_i_pad & ~\u4_u3_int_re_reg/P0001  ;
  assign n5456 = ~n5454 & n5455 ;
  assign n5457 = \u1_u3_int_upid_set_reg/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n5458 = ~\u4_u0_int_stat_reg[2]/P0001  & ~n5457 ;
  assign n5459 = rst_i_pad & ~\u4_u0_int_re_reg/P0001  ;
  assign n5460 = ~n5458 & n5459 ;
  assign n5461 = \u1_u3_int_upid_set_reg/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n5462 = ~\u4_u1_int_stat_reg[2]/P0001  & ~n5461 ;
  assign n5463 = rst_i_pad & ~\u4_u1_int_re_reg/P0001  ;
  assign n5464 = ~n5462 & n5463 ;
  assign n5465 = n3036 & n3614 ;
  assign n5466 = \u4_csr_reg[0]/P0001  & n3036 ;
  assign n5467 = ~n3617 & n5466 ;
  assign n5468 = ~n5465 & ~n5467 ;
  assign n5469 = \u1_u2_sizu_c_reg[0]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n5470 = ~n3833 & n5469 ;
  assign n5471 = \u1_u2_sizu_c_reg[0]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n5472 = n3033 & n5471 ;
  assign n5473 = ~n5470 & ~n5472 ;
  assign n5474 = ~n3967 & n5473 ;
  assign n5475 = n5468 & n5474 ;
  assign n5476 = \u4_csr_reg[10]/P0001  & n3036 ;
  assign n5477 = ~n3636 & n5476 ;
  assign n5478 = \u1_u2_sizu_c_reg[10]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n5479 = ~n3833 & n5478 ;
  assign n5480 = \u1_u2_sizu_c_reg[10]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n5481 = n3033 & n5480 ;
  assign n5482 = ~n5479 & ~n5481 ;
  assign n5483 = ~n3889 & n5482 ;
  assign n5484 = ~n5477 & n5483 ;
  assign n5485 = ~n3475 & n3611 ;
  assign n5486 = ~n3586 & n5485 ;
  assign n5487 = ~n3577 & n5486 ;
  assign n5488 = \u4_csr_reg[1]/P0001  & ~n3611 ;
  assign n5489 = \u4_csr_reg[1]/P0001  & n3565 ;
  assign n5490 = ~n3585 & n5489 ;
  assign n5491 = ~n5488 & ~n5490 ;
  assign n5492 = \u4_csr_reg[1]/P0001  & n3548 ;
  assign n5493 = n3574 & n5492 ;
  assign n5494 = ~n3531 & n5493 ;
  assign n5495 = ~n3530 & n5494 ;
  assign n5496 = n5491 & ~n5495 ;
  assign n5497 = ~n5487 & n5496 ;
  assign n5498 = n3036 & ~n5497 ;
  assign n5499 = \u1_u2_sizu_c_reg[1]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n5500 = ~n3833 & n5499 ;
  assign n5501 = \u1_u2_sizu_c_reg[1]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n5502 = n3033 & n5501 ;
  assign n5503 = ~n5500 & ~n5502 ;
  assign n5504 = ~n3954 & n5503 ;
  assign n5505 = ~n5498 & n5504 ;
  assign n5506 = \u4_csr_reg[2]/NET0131  & n3036 ;
  assign n5507 = ~n3617 & n5506 ;
  assign n5508 = n3036 & ~n3493 ;
  assign n5509 = n3617 & n5508 ;
  assign n5510 = ~n5507 & ~n5509 ;
  assign n5511 = \u1_u2_sizu_c_reg[2]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n5512 = ~n3833 & n5511 ;
  assign n5513 = \u1_u2_sizu_c_reg[2]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n5514 = n3033 & n5513 ;
  assign n5515 = ~n5512 & ~n5514 ;
  assign n5516 = ~n3941 & n5515 ;
  assign n5517 = n5510 & n5516 ;
  assign n5518 = \u4_csr_reg[3]/P0001  & n3036 ;
  assign n5519 = ~n3617 & n5518 ;
  assign n5520 = n3036 & ~n3511 ;
  assign n5521 = n3617 & n5520 ;
  assign n5522 = ~n5519 & ~n5521 ;
  assign n5523 = \u1_u2_sizu_c_reg[3]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n5524 = ~n3833 & n5523 ;
  assign n5525 = \u1_u2_sizu_c_reg[3]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n5526 = n3033 & n5525 ;
  assign n5527 = ~n5524 & ~n5526 ;
  assign n5528 = ~n3928 & n5527 ;
  assign n5529 = n5522 & n5528 ;
  assign n5530 = \u4_csr_reg[4]/NET0131  & n3036 ;
  assign n5531 = ~n3617 & n5530 ;
  assign n5532 = n3036 & ~n3503 ;
  assign n5533 = n3617 & n5532 ;
  assign n5534 = ~n5531 & ~n5533 ;
  assign n5535 = \u1_u2_sizu_c_reg[4]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n5536 = ~n3833 & n5535 ;
  assign n5537 = \u1_u2_sizu_c_reg[4]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n5538 = n3033 & n5537 ;
  assign n5539 = ~n5536 & ~n5538 ;
  assign n5540 = ~n3923 & n5539 ;
  assign n5541 = n5534 & n5540 ;
  assign n5542 = \u4_csr_reg[5]/NET0131  & n3036 ;
  assign n5543 = ~n3617 & n5542 ;
  assign n5544 = n3036 & ~n3525 ;
  assign n5545 = n3617 & n5544 ;
  assign n5546 = ~n5543 & ~n5545 ;
  assign n5547 = \u1_u2_sizu_c_reg[5]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n5548 = ~n3833 & n5547 ;
  assign n5549 = \u1_u2_sizu_c_reg[5]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n5550 = n3033 & n5549 ;
  assign n5551 = ~n5548 & ~n5550 ;
  assign n5552 = ~n3914 & n5551 ;
  assign n5553 = n5546 & n5552 ;
  assign n5554 = ~\u1_u2_idma_done_reg/P0001  & ~\u1_u3_state_reg[8]/P0001  ;
  assign n5555 = \u4_csr_reg[24]/P0001  & ~\u4_csr_reg[25]/P0001  ;
  assign n5556 = \u1_u2_idma_done_reg/P0001  & ~n5555 ;
  assign n5557 = n4918 & ~n5556 ;
  assign n5558 = n5401 & n5557 ;
  assign n5559 = ~n5554 & n5558 ;
  assign n5560 = n4949 & n4951 ;
  assign n5561 = n4947 & n5560 ;
  assign n5562 = ~n5559 & ~n5561 ;
  assign n5563 = \u1_u0_token_valid_str1_reg/P0001  & n4958 ;
  assign n5564 = ~\u1_u3_state_reg[8]/P0001  & ~n5563 ;
  assign n5565 = ~\u1_u3_rx_ack_to_reg/P0001  & n4962 ;
  assign n5566 = n4965 & n5565 ;
  assign n5567 = ~n5564 & n5566 ;
  assign n5568 = \u1_u3_state_reg[7]/P0001  & ~\u1_u3_state_reg[9]/P0001  ;
  assign n5569 = n4944 & n5568 ;
  assign n5570 = ~n5567 & ~n5569 ;
  assign n5571 = n5562 & n5570 ;
  assign n5572 = n5013 & ~n5571 ;
  assign n5573 = n5117 & ~n5571 ;
  assign n5574 = ~n5116 & n5573 ;
  assign n5575 = ~n5572 & ~n5574 ;
  assign n5576 = ~\u4_csr_reg[5]/NET0131  & ~\u4_csr_reg[6]/NET0131  ;
  assign n5577 = ~\u4_csr_reg[3]/P0001  & ~\u4_csr_reg[4]/NET0131  ;
  assign n5578 = n5576 & n5577 ;
  assign n5579 = ~\u4_csr_reg[1]/P0001  & ~\u4_csr_reg[2]/NET0131  ;
  assign n5580 = ~\u4_csr_reg[0]/P0001  & ~\u4_csr_reg[10]/P0001  ;
  assign n5581 = n5579 & n5580 ;
  assign n5582 = n5578 & n5581 ;
  assign n5583 = ~\u4_csr_reg[7]/P0001  & ~\u4_csr_reg[8]/P0001  ;
  assign n5584 = ~\u4_csr_reg[9]/NET0131  & n5583 ;
  assign n5585 = n5582 & n5584 ;
  assign n5586 = ~\u1_u3_state_reg[1]/P0001  & n5585 ;
  assign n5587 = n3458 & n5586 ;
  assign n5588 = n3451 & n5587 ;
  assign n5589 = n2376 & n5588 ;
  assign n5590 = n3455 & ~n5406 ;
  assign n5591 = ~\u1_u3_state_reg[1]/P0001  & ~\u4_csr_reg[26]/NET0131  ;
  assign n5592 = n2376 & n5591 ;
  assign n5593 = n5590 & n5592 ;
  assign n5594 = n3451 & n5593 ;
  assign n5595 = \u4_csr_reg[6]/NET0131  & ~n3840 ;
  assign n5596 = ~n3617 & n5595 ;
  assign n5597 = ~n3572 & ~n3840 ;
  assign n5598 = n3617 & n5597 ;
  assign n5599 = ~n5596 & ~n5598 ;
  assign n5600 = n3872 & ~n3875 ;
  assign n5601 = n5599 & n5600 ;
  assign n5602 = n3861 & ~n3864 ;
  assign n5603 = \u4_csr_reg[7]/P0001  & ~n3840 ;
  assign n5604 = ~n3617 & n5603 ;
  assign n5605 = ~n3538 & ~n3840 ;
  assign n5606 = n3617 & n5605 ;
  assign n5607 = ~n5604 & ~n5606 ;
  assign n5608 = n5602 & n5607 ;
  assign n5609 = ~n3831 & n3838 ;
  assign n5610 = \u4_csr_reg[8]/P0001  & ~n3840 ;
  assign n5611 = ~n3617 & n5610 ;
  assign n5612 = ~n3546 & ~n3840 ;
  assign n5613 = n3617 & n5612 ;
  assign n5614 = ~n5611 & ~n5613 ;
  assign n5615 = n5609 & n5614 ;
  assign n5616 = \u4_csr_reg[9]/NET0131  & ~n3840 ;
  assign n5617 = ~n3617 & n5616 ;
  assign n5618 = ~n3563 & ~n3840 ;
  assign n5619 = n3617 & n5618 ;
  assign n5620 = ~n5617 & ~n5619 ;
  assign n5621 = n3848 & ~n3852 ;
  assign n5622 = n5620 & n5621 ;
  assign n5623 = \u1_u3_state_reg[5]/P0001  & ~n4936 ;
  assign n5624 = ~n4912 & ~n5555 ;
  assign n5625 = n4911 & n5624 ;
  assign n5626 = ~n5623 & ~n5625 ;
  assign n5627 = n5431 & ~n5626 ;
  assign n5628 = n5013 & n5627 ;
  assign n5629 = n5117 & n5627 ;
  assign n5630 = ~n5116 & n5629 ;
  assign n5631 = ~n5628 & ~n5630 ;
  assign n5632 = ~\u1_u3_abort_reg/P0001  & n4968 ;
  assign n5633 = n4965 & n5632 ;
  assign n5634 = n5013 & n5633 ;
  assign n5635 = n5117 & n5633 ;
  assign n5636 = ~n5116 & n5635 ;
  assign n5637 = ~n5634 & ~n5636 ;
  assign n5638 = n4907 & ~n5625 ;
  assign n5639 = n5429 & n5638 ;
  assign n5640 = ~n5428 & n5639 ;
  assign n5641 = ~\u1_u3_state_reg[7]/P0001  & ~n4936 ;
  assign n5642 = n5013 & ~n5641 ;
  assign n5643 = n5117 & ~n5641 ;
  assign n5644 = ~n5116 & n5643 ;
  assign n5645 = ~n5642 & ~n5644 ;
  assign n5646 = n5640 & ~n5645 ;
  assign n5647 = ~\u1_u3_state_reg[6]/P0001  & \u1_u3_state_reg[8]/P0001  ;
  assign n5648 = n2370 & n5647 ;
  assign n5649 = n2375 & n5648 ;
  assign n5650 = n5013 & n5649 ;
  assign n5651 = n5117 & n5649 ;
  assign n5652 = ~n5116 & n5651 ;
  assign n5653 = ~n5650 & ~n5652 ;
  assign n5654 = n4916 & ~n5653 ;
  assign n5655 = n4918 & n5401 ;
  assign n5656 = ~\u1_u2_idma_done_reg/P0001  & \u1_u3_state_reg[3]/P0001  ;
  assign n5657 = ~n5556 & ~n5656 ;
  assign n5658 = n5655 & ~n5657 ;
  assign n5659 = \u1_u3_state_reg[3]/P0001  & ~n5563 ;
  assign n5660 = n5566 & n5659 ;
  assign n5661 = ~n5658 & ~n5660 ;
  assign n5662 = n5013 & ~n5661 ;
  assign n5663 = n5117 & ~n5661 ;
  assign n5664 = ~n5116 & n5663 ;
  assign n5665 = ~n5662 & ~n5664 ;
  assign n5666 = ~\u4_int_srcb_reg[2]/P0001  & ~\u4_nse_err_r_reg/P0001  ;
  assign n5667 = rst_i_pad & ~\u4_int_src_re_reg/P0001  ;
  assign n5668 = ~n5666 & n5667 ;
  assign n5669 = ~\u1_u3_adr_reg[8]/P0001  & n3546 ;
  assign n5670 = ~\u1_u3_adr_reg[11]/P0001  & n3601 ;
  assign n5671 = ~\u1_u3_adr_reg[12]/P0001  & n3594 ;
  assign n5672 = ~n5670 & ~n5671 ;
  assign n5673 = ~\u1_u3_adr_reg[10]/P0001  & n3555 ;
  assign n5674 = ~\u1_u3_adr_reg[9]/P0001  & n3563 ;
  assign n5675 = ~n5673 & ~n5674 ;
  assign n5676 = n5672 & n5675 ;
  assign n5677 = ~n5669 & n5676 ;
  assign n5678 = \u1_u3_adr_reg[9]/P0001  & ~n3563 ;
  assign n5679 = ~n5673 & n5678 ;
  assign n5680 = \u1_u3_adr_reg[11]/P0001  & ~n3601 ;
  assign n5681 = \u1_u3_adr_reg[10]/P0001  & ~n3555 ;
  assign n5682 = ~n5680 & ~n5681 ;
  assign n5683 = ~n5679 & n5682 ;
  assign n5684 = n5672 & ~n5683 ;
  assign n5685 = \u1_u3_adr_reg[13]/P0001  & ~n3609 ;
  assign n5686 = ~\u1_u3_adr_reg[13]/P0001  & n3609 ;
  assign n5687 = ~n5685 & ~n5686 ;
  assign n5688 = \u1_u3_adr_reg[12]/P0001  & ~n3594 ;
  assign n5689 = n5687 & ~n5688 ;
  assign n5690 = ~n5684 & n5689 ;
  assign n5691 = ~n5677 & n5690 ;
  assign n5692 = ~\u1_u3_adr_reg[6]/P0001  & n3572 ;
  assign n5693 = ~\u1_u3_adr_reg[7]/P0001  & n3538 ;
  assign n5694 = ~n5692 & ~n5693 ;
  assign n5695 = \u1_u3_adr_reg[6]/P0001  & ~n3572 ;
  assign n5696 = \u1_u3_adr_reg[5]/P0001  & ~n3525 ;
  assign n5697 = ~n5695 & ~n5696 ;
  assign n5698 = n5694 & ~n5697 ;
  assign n5699 = ~\u1_u3_adr_reg[5]/P0001  & n3525 ;
  assign n5700 = ~\u1_u3_adr_reg[4]/P0001  & n3503 ;
  assign n5701 = ~n5699 & ~n5700 ;
  assign n5702 = n5694 & n5701 ;
  assign n5703 = ~n5698 & ~n5702 ;
  assign n5704 = ~\u1_u3_adr_reg[1]/P0001  & n3475 ;
  assign n5705 = \u1_u3_adr_reg[0]/P0001  & ~n3483 ;
  assign n5706 = ~n5704 & n5705 ;
  assign n5707 = \u1_u3_adr_reg[2]/P0001  & ~n3493 ;
  assign n5708 = \u1_u3_adr_reg[1]/P0001  & ~n3475 ;
  assign n5709 = ~n5707 & ~n5708 ;
  assign n5710 = ~n5706 & n5709 ;
  assign n5711 = ~\u1_u3_adr_reg[3]/P0001  & n3511 ;
  assign n5712 = ~\u1_u3_adr_reg[2]/P0001  & n3493 ;
  assign n5713 = ~n5711 & ~n5712 ;
  assign n5714 = ~n5710 & n5713 ;
  assign n5715 = \u1_u3_adr_reg[4]/P0001  & ~n3503 ;
  assign n5716 = \u1_u3_adr_reg[3]/P0001  & ~n3511 ;
  assign n5717 = ~n5715 & ~n5716 ;
  assign n5718 = ~n5698 & n5717 ;
  assign n5719 = ~n5714 & n5718 ;
  assign n5720 = ~n5703 & ~n5719 ;
  assign n5721 = \u1_u3_adr_reg[8]/P0001  & ~n3546 ;
  assign n5722 = \u1_u3_adr_reg[7]/P0001  & ~n3538 ;
  assign n5723 = ~n5721 & ~n5722 ;
  assign n5724 = n5690 & n5723 ;
  assign n5725 = ~n5720 & n5724 ;
  assign n5726 = ~n5691 & ~n5725 ;
  assign n5727 = ~n5684 & ~n5688 ;
  assign n5728 = ~n5677 & n5727 ;
  assign n5729 = n5723 & n5727 ;
  assign n5730 = ~n5720 & n5729 ;
  assign n5731 = ~n5728 & ~n5730 ;
  assign n5732 = ~n5687 & n5731 ;
  assign n5733 = n5726 & ~n5732 ;
  assign n5734 = ~\u0_u0_state_reg[13]/NET0131  & ~\u0_u0_state_reg[14]/P0001  ;
  assign n5735 = ~\u0_u0_state_reg[0]/NET0131  & n5734 ;
  assign n5736 = ~\u0_u0_state_reg[8]/NET0131  & ~\u0_u0_state_reg[9]/P0001  ;
  assign n5737 = \u0_u0_state_reg[10]/P0001  & ~\u0_u0_state_reg[7]/NET0131  ;
  assign n5738 = n5736 & n5737 ;
  assign n5739 = n5735 & n5738 ;
  assign n5740 = ~\u0_u0_state_reg[4]/NET0131  & ~\u0_u0_state_reg[5]/P0001  ;
  assign n5741 = ~\u0_u0_state_reg[3]/P0001  & ~\u0_u0_state_reg[6]/NET0131  ;
  assign n5742 = n5740 & n5741 ;
  assign n5743 = ~\u0_u0_state_reg[1]/P0001  & ~\u0_u0_state_reg[2]/NET0131  ;
  assign n5744 = ~\u0_u0_state_reg[11]/NET0131  & ~\u0_u0_state_reg[12]/NET0131  ;
  assign n5745 = n5743 & n5744 ;
  assign n5746 = n5742 & n5745 ;
  assign n5747 = n5739 & n5746 ;
  assign n5748 = rst_i_pad & ~usb_vbus_pad_i_pad ;
  assign n5749 = ~\u0_u0_T2_gt_1_0_mS_reg/P0001  & ~\u0_u0_state_reg[11]/NET0131  ;
  assign n5750 = n5748 & ~n5749 ;
  assign n5751 = n5747 & n5750 ;
  assign n5752 = n5742 & n5743 ;
  assign n5753 = ~\u0_u0_state_reg[10]/P0001  & ~\u0_u0_state_reg[7]/NET0131  ;
  assign n5754 = ~\u0_u0_state_reg[8]/NET0131  & n5753 ;
  assign n5755 = ~\u0_u0_state_reg[0]/NET0131  & ~\u0_u0_state_reg[9]/P0001  ;
  assign n5756 = n5734 & n5755 ;
  assign n5757 = n5754 & n5756 ;
  assign n5758 = n5752 & n5757 ;
  assign n5759 = \LineState_r_reg[0]/P0001  & ~\LineState_r_reg[1]/P0001  ;
  assign n5760 = \u0_u0_ls_j_r_reg/P0001  & n5759 ;
  assign n5761 = ~\u0_u0_state_reg[11]/NET0131  & \u0_u0_state_reg[12]/NET0131  ;
  assign n5762 = n5760 & n5761 ;
  assign n5763 = n5758 & n5762 ;
  assign n5764 = \u0_u0_state_reg[11]/NET0131  & ~\u0_u0_state_reg[12]/NET0131  ;
  assign n5765 = ~\LineState_r_reg[0]/P0001  & ~\LineState_r_reg[1]/P0001  ;
  assign n5766 = \u0_u0_ls_se0_r_reg/P0001  & n5765 ;
  assign n5767 = ~\LineState_r_reg[0]/P0001  & \LineState_r_reg[1]/P0001  ;
  assign n5768 = \u0_u0_ls_k_r_reg/P0001  & n5767 ;
  assign n5769 = ~n5766 & ~n5768 ;
  assign n5770 = n5764 & n5769 ;
  assign n5771 = n5758 & n5770 ;
  assign n5772 = ~n5763 & ~n5771 ;
  assign n5773 = ~\u0_u0_chirp_cnt_is_6_reg/P0001  & n5748 ;
  assign n5774 = ~n5772 & n5773 ;
  assign n5775 = ~n5751 & ~n5774 ;
  assign n5776 = \u4_u3_csr0_reg[9]/P0001  & ~\u4_u3_dma_out_left_reg[7]/P0001  ;
  assign n5777 = \u4_u3_csr0_reg[10]/P0001  & ~\u4_u3_dma_out_left_reg[8]/P0001  ;
  assign n5778 = ~n5776 & ~n5777 ;
  assign n5779 = ~\u4_u3_csr0_reg[9]/P0001  & \u4_u3_dma_out_left_reg[7]/P0001  ;
  assign n5780 = ~\u4_u3_csr0_reg[8]/P0001  & \u4_u3_dma_out_left_reg[6]/P0001  ;
  assign n5781 = ~n5779 & ~n5780 ;
  assign n5782 = n5778 & ~n5781 ;
  assign n5783 = ~\u4_u3_csr0_reg[7]/P0001  & \u4_u3_dma_out_left_reg[5]/P0001  ;
  assign n5784 = ~\u4_u3_csr0_reg[6]/P0001  & \u4_u3_dma_out_left_reg[4]/P0001  ;
  assign n5785 = ~n5783 & ~n5784 ;
  assign n5786 = \u4_u3_csr0_reg[6]/P0001  & ~\u4_u3_dma_out_left_reg[4]/P0001  ;
  assign n5787 = \u4_u3_csr0_reg[5]/P0001  & ~\u4_u3_dma_out_left_reg[3]/P0001  ;
  assign n5788 = ~n5786 & ~n5787 ;
  assign n5789 = n5785 & ~n5788 ;
  assign n5790 = ~\u4_u3_csr0_reg[3]/NET0131  & \u4_u3_dma_out_left_reg[1]/P0001  ;
  assign n5791 = \u4_u3_csr0_reg[2]/P0001  & ~\u4_u3_dma_out_left_reg[0]/P0001  ;
  assign n5792 = ~n5790 & n5791 ;
  assign n5793 = \u4_u3_csr0_reg[4]/P0001  & ~\u4_u3_dma_out_left_reg[2]/P0001  ;
  assign n5794 = \u4_u3_csr0_reg[3]/NET0131  & ~\u4_u3_dma_out_left_reg[1]/P0001  ;
  assign n5795 = ~n5793 & ~n5794 ;
  assign n5796 = ~n5792 & n5795 ;
  assign n5797 = ~\u4_u3_csr0_reg[5]/P0001  & \u4_u3_dma_out_left_reg[3]/P0001  ;
  assign n5798 = ~\u4_u3_csr0_reg[4]/P0001  & \u4_u3_dma_out_left_reg[2]/P0001  ;
  assign n5799 = ~n5797 & ~n5798 ;
  assign n5800 = n5785 & n5799 ;
  assign n5801 = ~n5796 & n5800 ;
  assign n5802 = ~n5789 & ~n5801 ;
  assign n5803 = \u4_u3_csr0_reg[8]/P0001  & ~\u4_u3_dma_out_left_reg[6]/P0001  ;
  assign n5804 = \u4_u3_csr0_reg[7]/P0001  & ~\u4_u3_dma_out_left_reg[5]/P0001  ;
  assign n5805 = ~n5803 & ~n5804 ;
  assign n5806 = n5778 & n5805 ;
  assign n5807 = n5802 & n5806 ;
  assign n5808 = ~n5782 & ~n5807 ;
  assign n5809 = ~\u4_u3_csr0_reg[10]/P0001  & \u4_u3_dma_out_left_reg[8]/P0001  ;
  assign n5810 = ~\u4_u3_dma_out_left_reg[10]/P0001  & ~\u4_u3_dma_out_left_reg[11]/P0001  ;
  assign n5811 = ~\u4_u3_dma_out_left_reg[9]/P0001  & n5810 ;
  assign n5812 = ~n5809 & n5811 ;
  assign n5813 = n5808 & n5812 ;
  assign n5814 = \u4_u0_csr0_reg[9]/P0001  & ~\u4_u0_dma_out_left_reg[7]/P0001  ;
  assign n5815 = \u4_u0_csr0_reg[10]/P0001  & ~\u4_u0_dma_out_left_reg[8]/P0001  ;
  assign n5816 = ~n5814 & ~n5815 ;
  assign n5817 = ~\u4_u0_csr0_reg[9]/P0001  & \u4_u0_dma_out_left_reg[7]/P0001  ;
  assign n5818 = ~\u4_u0_csr0_reg[8]/P0001  & \u4_u0_dma_out_left_reg[6]/P0001  ;
  assign n5819 = ~n5817 & ~n5818 ;
  assign n5820 = n5816 & ~n5819 ;
  assign n5821 = ~\u4_u0_csr0_reg[7]/P0001  & \u4_u0_dma_out_left_reg[5]/P0001  ;
  assign n5822 = ~\u4_u0_csr0_reg[6]/P0001  & \u4_u0_dma_out_left_reg[4]/P0001  ;
  assign n5823 = ~n5821 & ~n5822 ;
  assign n5824 = \u4_u0_csr0_reg[6]/P0001  & ~\u4_u0_dma_out_left_reg[4]/P0001  ;
  assign n5825 = \u4_u0_csr0_reg[5]/P0001  & ~\u4_u0_dma_out_left_reg[3]/P0001  ;
  assign n5826 = ~n5824 & ~n5825 ;
  assign n5827 = n5823 & ~n5826 ;
  assign n5828 = ~\u4_u0_csr0_reg[3]/NET0131  & \u4_u0_dma_out_left_reg[1]/P0001  ;
  assign n5829 = \u4_u0_csr0_reg[2]/P0001  & ~\u4_u0_dma_out_left_reg[0]/P0001  ;
  assign n5830 = ~n5828 & n5829 ;
  assign n5831 = \u4_u0_csr0_reg[4]/P0001  & ~\u4_u0_dma_out_left_reg[2]/P0001  ;
  assign n5832 = \u4_u0_csr0_reg[3]/NET0131  & ~\u4_u0_dma_out_left_reg[1]/P0001  ;
  assign n5833 = ~n5831 & ~n5832 ;
  assign n5834 = ~n5830 & n5833 ;
  assign n5835 = ~\u4_u0_csr0_reg[5]/P0001  & \u4_u0_dma_out_left_reg[3]/P0001  ;
  assign n5836 = ~\u4_u0_csr0_reg[4]/P0001  & \u4_u0_dma_out_left_reg[2]/P0001  ;
  assign n5837 = ~n5835 & ~n5836 ;
  assign n5838 = n5823 & n5837 ;
  assign n5839 = ~n5834 & n5838 ;
  assign n5840 = ~n5827 & ~n5839 ;
  assign n5841 = \u4_u0_csr0_reg[8]/P0001  & ~\u4_u0_dma_out_left_reg[6]/P0001  ;
  assign n5842 = \u4_u0_csr0_reg[7]/P0001  & ~\u4_u0_dma_out_left_reg[5]/P0001  ;
  assign n5843 = ~n5841 & ~n5842 ;
  assign n5844 = n5816 & n5843 ;
  assign n5845 = n5840 & n5844 ;
  assign n5846 = ~n5820 & ~n5845 ;
  assign n5847 = ~\u4_u0_csr0_reg[10]/P0001  & \u4_u0_dma_out_left_reg[8]/P0001  ;
  assign n5848 = ~\u4_u0_dma_out_left_reg[10]/P0001  & ~\u4_u0_dma_out_left_reg[11]/P0001  ;
  assign n5849 = ~\u4_u0_dma_out_left_reg[9]/P0001  & n5848 ;
  assign n5850 = ~n5847 & n5849 ;
  assign n5851 = n5846 & n5850 ;
  assign n5852 = \u4_u1_csr0_reg[9]/P0001  & ~\u4_u1_dma_out_left_reg[7]/P0001  ;
  assign n5853 = \u4_u1_csr0_reg[10]/P0001  & ~\u4_u1_dma_out_left_reg[8]/P0001  ;
  assign n5854 = ~n5852 & ~n5853 ;
  assign n5855 = ~\u4_u1_csr0_reg[9]/P0001  & \u4_u1_dma_out_left_reg[7]/P0001  ;
  assign n5856 = ~\u4_u1_csr0_reg[8]/P0001  & \u4_u1_dma_out_left_reg[6]/P0001  ;
  assign n5857 = ~n5855 & ~n5856 ;
  assign n5858 = n5854 & ~n5857 ;
  assign n5859 = ~\u4_u1_csr0_reg[7]/P0001  & \u4_u1_dma_out_left_reg[5]/P0001  ;
  assign n5860 = ~\u4_u1_csr0_reg[6]/P0001  & \u4_u1_dma_out_left_reg[4]/P0001  ;
  assign n5861 = ~n5859 & ~n5860 ;
  assign n5862 = \u4_u1_csr0_reg[6]/P0001  & ~\u4_u1_dma_out_left_reg[4]/P0001  ;
  assign n5863 = \u4_u1_csr0_reg[5]/P0001  & ~\u4_u1_dma_out_left_reg[3]/P0001  ;
  assign n5864 = ~n5862 & ~n5863 ;
  assign n5865 = n5861 & ~n5864 ;
  assign n5866 = ~\u4_u1_csr0_reg[3]/NET0131  & \u4_u1_dma_out_left_reg[1]/P0001  ;
  assign n5867 = \u4_u1_csr0_reg[2]/P0001  & ~\u4_u1_dma_out_left_reg[0]/P0001  ;
  assign n5868 = ~n5866 & n5867 ;
  assign n5869 = \u4_u1_csr0_reg[4]/P0001  & ~\u4_u1_dma_out_left_reg[2]/P0001  ;
  assign n5870 = \u4_u1_csr0_reg[3]/NET0131  & ~\u4_u1_dma_out_left_reg[1]/P0001  ;
  assign n5871 = ~n5869 & ~n5870 ;
  assign n5872 = ~n5868 & n5871 ;
  assign n5873 = ~\u4_u1_csr0_reg[5]/P0001  & \u4_u1_dma_out_left_reg[3]/P0001  ;
  assign n5874 = ~\u4_u1_csr0_reg[4]/P0001  & \u4_u1_dma_out_left_reg[2]/P0001  ;
  assign n5875 = ~n5873 & ~n5874 ;
  assign n5876 = n5861 & n5875 ;
  assign n5877 = ~n5872 & n5876 ;
  assign n5878 = ~n5865 & ~n5877 ;
  assign n5879 = \u4_u1_csr0_reg[8]/P0001  & ~\u4_u1_dma_out_left_reg[6]/P0001  ;
  assign n5880 = \u4_u1_csr0_reg[7]/P0001  & ~\u4_u1_dma_out_left_reg[5]/P0001  ;
  assign n5881 = ~n5879 & ~n5880 ;
  assign n5882 = n5854 & n5881 ;
  assign n5883 = n5878 & n5882 ;
  assign n5884 = ~n5858 & ~n5883 ;
  assign n5885 = ~\u4_u1_csr0_reg[10]/P0001  & \u4_u1_dma_out_left_reg[8]/P0001  ;
  assign n5886 = ~\u4_u1_dma_out_left_reg[10]/P0001  & ~\u4_u1_dma_out_left_reg[11]/P0001  ;
  assign n5887 = ~\u4_u1_dma_out_left_reg[9]/P0001  & n5886 ;
  assign n5888 = ~n5885 & n5887 ;
  assign n5889 = n5884 & n5888 ;
  assign n5890 = \u4_u2_csr0_reg[9]/P0001  & ~\u4_u2_dma_out_left_reg[7]/P0001  ;
  assign n5891 = \u4_u2_csr0_reg[10]/P0001  & ~\u4_u2_dma_out_left_reg[8]/P0001  ;
  assign n5892 = ~n5890 & ~n5891 ;
  assign n5893 = ~\u4_u2_csr0_reg[9]/P0001  & \u4_u2_dma_out_left_reg[7]/P0001  ;
  assign n5894 = ~\u4_u2_csr0_reg[8]/P0001  & \u4_u2_dma_out_left_reg[6]/P0001  ;
  assign n5895 = ~n5893 & ~n5894 ;
  assign n5896 = n5892 & ~n5895 ;
  assign n5897 = ~\u4_u2_csr0_reg[7]/P0001  & \u4_u2_dma_out_left_reg[5]/P0001  ;
  assign n5898 = ~\u4_u2_csr0_reg[6]/P0001  & \u4_u2_dma_out_left_reg[4]/P0001  ;
  assign n5899 = ~n5897 & ~n5898 ;
  assign n5900 = \u4_u2_csr0_reg[6]/P0001  & ~\u4_u2_dma_out_left_reg[4]/P0001  ;
  assign n5901 = \u4_u2_csr0_reg[5]/P0001  & ~\u4_u2_dma_out_left_reg[3]/P0001  ;
  assign n5902 = ~n5900 & ~n5901 ;
  assign n5903 = n5899 & ~n5902 ;
  assign n5904 = ~\u4_u2_csr0_reg[3]/NET0131  & \u4_u2_dma_out_left_reg[1]/P0001  ;
  assign n5905 = \u4_u2_csr0_reg[2]/P0001  & ~\u4_u2_dma_out_left_reg[0]/P0001  ;
  assign n5906 = ~n5904 & n5905 ;
  assign n5907 = \u4_u2_csr0_reg[4]/P0001  & ~\u4_u2_dma_out_left_reg[2]/P0001  ;
  assign n5908 = \u4_u2_csr0_reg[3]/NET0131  & ~\u4_u2_dma_out_left_reg[1]/P0001  ;
  assign n5909 = ~n5907 & ~n5908 ;
  assign n5910 = ~n5906 & n5909 ;
  assign n5911 = ~\u4_u2_csr0_reg[5]/P0001  & \u4_u2_dma_out_left_reg[3]/P0001  ;
  assign n5912 = ~\u4_u2_csr0_reg[4]/P0001  & \u4_u2_dma_out_left_reg[2]/P0001  ;
  assign n5913 = ~n5911 & ~n5912 ;
  assign n5914 = n5899 & n5913 ;
  assign n5915 = ~n5910 & n5914 ;
  assign n5916 = ~n5903 & ~n5915 ;
  assign n5917 = \u4_u2_csr0_reg[8]/P0001  & ~\u4_u2_dma_out_left_reg[6]/P0001  ;
  assign n5918 = \u4_u2_csr0_reg[7]/P0001  & ~\u4_u2_dma_out_left_reg[5]/P0001  ;
  assign n5919 = ~n5917 & ~n5918 ;
  assign n5920 = n5892 & n5919 ;
  assign n5921 = n5916 & n5920 ;
  assign n5922 = ~n5896 & ~n5921 ;
  assign n5923 = ~\u4_u2_csr0_reg[10]/P0001  & \u4_u2_dma_out_left_reg[8]/P0001  ;
  assign n5924 = ~\u4_u2_dma_out_left_reg[10]/P0001  & ~\u4_u2_dma_out_left_reg[11]/P0001  ;
  assign n5925 = ~\u4_u2_dma_out_left_reg[9]/P0001  & n5924 ;
  assign n5926 = ~n5923 & n5925 ;
  assign n5927 = n5922 & n5926 ;
  assign n5928 = n5012 & ~n5015 ;
  assign n5929 = \u1_u3_match_r_reg/P0001  & \u1_u3_to_large_reg/P0001  ;
  assign n5930 = ~\u1_u3_buffer_overflow_reg/P0001  & ~n5929 ;
  assign n5931 = ~n5928 & n5930 ;
  assign n5932 = \u1_u0_token_valid_str1_reg/P0001  & n5930 ;
  assign n5933 = ~n5116 & n5932 ;
  assign n5934 = ~n5931 & ~n5933 ;
  assign n5935 = ~\u0_u0_T2_gt_1_0_mS_reg/P0001  & ~\u0_u0_state_reg[10]/P0001  ;
  assign n5936 = ~\u0_u0_state_reg[8]/NET0131  & \u0_u0_state_reg[9]/P0001  ;
  assign n5937 = n5753 & n5936 ;
  assign n5938 = n5735 & n5937 ;
  assign n5939 = n5746 & n5938 ;
  assign n5940 = ~n5935 & n5939 ;
  assign n5941 = ~\u0_u0_T2_gt_1_0_mS_reg/P0001  & n5747 ;
  assign n5942 = ~n5940 & ~n5941 ;
  assign n5943 = n5748 & ~n5942 ;
  assign n5944 = n5701 & n5716 ;
  assign n5945 = n5701 & n5713 ;
  assign n5946 = ~n5710 & n5945 ;
  assign n5947 = ~n5944 & ~n5946 ;
  assign n5948 = ~n5693 & n5695 ;
  assign n5949 = ~n5722 & ~n5948 ;
  assign n5950 = ~n5699 & n5715 ;
  assign n5951 = ~n5696 & ~n5950 ;
  assign n5952 = n5949 & n5951 ;
  assign n5953 = n5947 & n5952 ;
  assign n5954 = ~\u1_u3_adr_reg[6]/P0001  & n3538 ;
  assign n5955 = n3572 & n5954 ;
  assign n5956 = ~\u1_u3_adr_reg[6]/P0001  & ~\u1_u3_adr_reg[7]/P0001  ;
  assign n5957 = n3572 & n5956 ;
  assign n5958 = ~n5693 & ~n5957 ;
  assign n5959 = ~n5955 & n5958 ;
  assign n5960 = ~n5673 & ~n5686 ;
  assign n5961 = n5672 & n5960 ;
  assign n5962 = ~n5669 & ~n5674 ;
  assign n5963 = n5961 & n5962 ;
  assign n5964 = n5959 & n5963 ;
  assign n5965 = ~n5953 & n5964 ;
  assign n5966 = n5672 & ~n5682 ;
  assign n5967 = ~n5685 & ~n5688 ;
  assign n5968 = ~n5966 & n5967 ;
  assign n5969 = ~n5686 & ~n5968 ;
  assign n5970 = ~n5674 & n5721 ;
  assign n5971 = ~n5678 & ~n5970 ;
  assign n5972 = n5961 & ~n5971 ;
  assign n5973 = ~\u1_u3_adr_reg[14]/P0001  & ~n5972 ;
  assign n5974 = ~n5969 & n5973 ;
  assign n5975 = ~n5965 & n5974 ;
  assign n5976 = ~n5969 & ~n5972 ;
  assign n5977 = ~n5965 & n5976 ;
  assign n5978 = \u1_u3_adr_reg[14]/P0001  & ~n5977 ;
  assign n5979 = ~n5975 & ~n5978 ;
  assign n5980 = \u1_frame_no_same_reg/P0001  & \u1_mfm_cnt_reg[0]/P0001  ;
  assign n5981 = ~\u1_mfm_cnt_reg[1]/P0001  & ~n5980 ;
  assign n5982 = \u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_same_reg/P0001  ;
  assign n5983 = rst_i_pad & ~n5982 ;
  assign n5984 = \u1_mfm_cnt_reg[1]/P0001  & n5980 ;
  assign n5985 = n5983 & ~n5984 ;
  assign n5986 = ~n5981 & n5985 ;
  assign n5987 = \u1_u3_int_seqerr_set_reg/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n5988 = ~\u4_u2_int_stat_reg[5]/P0001  & ~n5987 ;
  assign n5989 = n5451 & ~n5988 ;
  assign n5990 = ~\u1_frame_no_same_reg/P0001  & ~\u1_mfm_cnt_reg[0]/P0001  ;
  assign n5991 = ~n5980 & ~n5990 ;
  assign n5992 = n5983 & n5991 ;
  assign n5993 = ~\u1_mfm_cnt_reg[2]/P0001  & ~n5984 ;
  assign n5994 = \u1_mfm_cnt_reg[1]/P0001  & \u1_mfm_cnt_reg[2]/P0001  ;
  assign n5995 = n5980 & n5994 ;
  assign n5996 = n5983 & ~n5995 ;
  assign n5997 = ~n5993 & n5996 ;
  assign n5998 = rst_i_pad & \u1_mfm_cnt_reg[3]/P0001  ;
  assign n5999 = ~n5982 & n5998 ;
  assign n6000 = ~n5995 & n5999 ;
  assign n6001 = rst_i_pad & ~\u1_mfm_cnt_reg[3]/P0001  ;
  assign n6002 = ~n5982 & n6001 ;
  assign n6003 = n5995 & n6002 ;
  assign n6004 = ~n6000 & ~n6003 ;
  assign n6005 = \u1_u3_int_seqerr_set_reg/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n6006 = ~\u4_u3_int_stat_reg[5]/P0001  & ~n6005 ;
  assign n6007 = n5455 & ~n6006 ;
  assign n6008 = \u1_u3_int_seqerr_set_reg/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n6009 = ~\u4_u0_int_stat_reg[5]/P0001  & ~n6008 ;
  assign n6010 = n5459 & ~n6009 ;
  assign n6011 = \u1_u3_int_seqerr_set_reg/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n6012 = ~\u4_u1_int_stat_reg[5]/P0001  & ~n6011 ;
  assign n6013 = n5463 & ~n6012 ;
  assign n6014 = \u1_u3_match_r_reg/P0001  & ~n2379 ;
  assign n6015 = ~\u1_u3_pid_IN_r_reg/P0001  & n2361 ;
  assign n6016 = ~\u1_u3_pid_IN_r_reg/P0001  & ~\u1_u3_pid_SETUP_r_reg/P0001  ;
  assign n6017 = ~\u4_csr_reg[27]/NET0131  & ~n6016 ;
  assign n6018 = ~\u1_u3_pid_OUT_r_reg/P0001  & ~\u1_u3_pid_PING_r_reg/P0001  ;
  assign n6019 = ~\u4_csr_reg[26]/NET0131  & n6018 ;
  assign n6020 = ~n6017 & n6019 ;
  assign n6021 = ~n6015 & ~n6020 ;
  assign n6022 = n6014 & ~n6021 ;
  assign n6023 = \u4_csr_reg[0]/P0001  & ~n3617 ;
  assign n6024 = ~n3614 & ~n6023 ;
  assign n6025 = \u4_csr_reg[10]/P0001  & ~n3636 ;
  assign n6026 = \u4_csr_reg[3]/P0001  & ~n3617 ;
  assign n6027 = ~n3691 & ~n6026 ;
  assign n6028 = \u4_csr_reg[4]/NET0131  & ~n3617 ;
  assign n6029 = ~n3704 & ~n6028 ;
  assign n6030 = \u4_csr_reg[5]/NET0131  & ~n3617 ;
  assign n6031 = ~n3720 & ~n6030 ;
  assign n6032 = \u4_csr_reg[6]/NET0131  & ~n3617 ;
  assign n6033 = ~n3733 & ~n6032 ;
  assign n6034 = \u4_csr_reg[7]/P0001  & ~n3617 ;
  assign n6035 = ~n3745 & ~n6034 ;
  assign n6036 = \u4_csr_reg[8]/P0001  & ~n3617 ;
  assign n6037 = ~n3758 & ~n6036 ;
  assign n6038 = \u4_csr_reg[9]/NET0131  & ~n3617 ;
  assign n6039 = ~n3771 & ~n6038 ;
  assign n6040 = \u1_u0_token_valid_str1_reg/P0001  & n2350 ;
  assign n6041 = ~n2378 & n6040 ;
  assign n6042 = ~n5012 & n6041 ;
  assign n6043 = \u1_u0_token_valid_str1_reg/P0001  & n6041 ;
  assign n6044 = ~n5116 & n6043 ;
  assign n6045 = ~n6042 & ~n6044 ;
  assign n6046 = \u1_u2_sizu_c_reg[8]/NET0131  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n6047 = \u1_u3_new_size_reg[8]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n6048 = ~n6046 & ~n6047 ;
  assign n6049 = \u1_u3_new_size_reg[9]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n6050 = \u1_u2_sizu_c_reg[9]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n6051 = ~n6049 & ~n6050 ;
  assign n6052 = n5959 & n5962 ;
  assign n6053 = ~n5953 & n6052 ;
  assign n6054 = ~n5673 & ~n5681 ;
  assign n6055 = n5971 & n6054 ;
  assign n6056 = ~n6053 & n6055 ;
  assign n6057 = ~n5971 & ~n6054 ;
  assign n6058 = n5962 & ~n6054 ;
  assign n6059 = n5959 & n6058 ;
  assign n6060 = ~n5953 & n6059 ;
  assign n6061 = ~n6057 & ~n6060 ;
  assign n6062 = ~n6056 & n6061 ;
  assign n6063 = ~n5671 & ~n5688 ;
  assign n6064 = ~n5670 & ~n5682 ;
  assign n6065 = ~n5670 & ~n5673 ;
  assign n6066 = ~n6064 & ~n6065 ;
  assign n6067 = n5971 & ~n6064 ;
  assign n6068 = ~n6053 & n6067 ;
  assign n6069 = ~n6066 & ~n6068 ;
  assign n6070 = ~n6063 & n6069 ;
  assign n6071 = n6063 & ~n6069 ;
  assign n6072 = ~n6070 & ~n6071 ;
  assign n6073 = ~n5720 & n5723 ;
  assign n6074 = ~n5674 & ~n5678 ;
  assign n6075 = ~n5669 & ~n6074 ;
  assign n6076 = ~n6073 & n6075 ;
  assign n6077 = n5669 & n6074 ;
  assign n6078 = n5723 & n6074 ;
  assign n6079 = ~n5720 & n6078 ;
  assign n6080 = ~n6077 & ~n6079 ;
  assign n6081 = ~n6076 & n6080 ;
  assign n6082 = \u1_u2_sizu_c_reg[10]/P0001  & n3555 ;
  assign n6083 = ~\u1_u2_sizu_c_reg[9]/P0001  & ~n3563 ;
  assign n6084 = \u1_u2_sizu_c_reg[9]/P0001  & n3563 ;
  assign n6085 = \u1_u2_sizu_c_reg[8]/NET0131  & n3546 ;
  assign n6086 = ~n6084 & ~n6085 ;
  assign n6087 = ~n6083 & ~n6086 ;
  assign n6088 = ~n6082 & ~n6087 ;
  assign n6089 = ~\u1_u2_sizu_c_reg[10]/P0001  & ~n3555 ;
  assign n6090 = \u1_u0_data_valid0_reg/P0001  & ~n6089 ;
  assign n6091 = ~n6088 & n6090 ;
  assign n6092 = \u1_u2_sizu_c_reg[7]/P0001  & n3538 ;
  assign n6093 = \u1_u2_sizu_c_reg[6]/P0001  & n3572 ;
  assign n6094 = ~n6092 & ~n6093 ;
  assign n6095 = ~\u1_u2_sizu_c_reg[5]/P0001  & ~n3525 ;
  assign n6096 = ~\u1_u2_sizu_c_reg[6]/P0001  & ~n3572 ;
  assign n6097 = ~n6095 & ~n6096 ;
  assign n6098 = n6094 & ~n6097 ;
  assign n6099 = ~\u1_u2_sizu_c_reg[3]/P0001  & ~n3511 ;
  assign n6100 = ~\u1_u2_sizu_c_reg[4]/P0001  & ~n3503 ;
  assign n6101 = ~n6099 & ~n6100 ;
  assign n6102 = \u1_u2_sizu_c_reg[2]/P0001  & n3493 ;
  assign n6103 = \u1_u2_sizu_c_reg[3]/P0001  & n3511 ;
  assign n6104 = ~n6102 & ~n6103 ;
  assign n6105 = n6101 & ~n6104 ;
  assign n6106 = \u1_u2_sizu_c_reg[0]/P0001  & n3483 ;
  assign n6107 = ~\u1_u2_sizu_c_reg[1]/P0001  & ~n6106 ;
  assign n6108 = ~\u1_u2_sizu_c_reg[2]/P0001  & ~n3493 ;
  assign n6109 = ~n6107 & ~n6108 ;
  assign n6110 = \u1_u2_sizu_c_reg[0]/P0001  & \u1_u2_sizu_c_reg[1]/P0001  ;
  assign n6111 = n3483 & n6110 ;
  assign n6112 = ~n3475 & ~n6111 ;
  assign n6113 = n6101 & ~n6112 ;
  assign n6114 = n6109 & n6113 ;
  assign n6115 = ~n6105 & ~n6114 ;
  assign n6116 = \u1_u2_sizu_c_reg[5]/P0001  & n3525 ;
  assign n6117 = \u1_u2_sizu_c_reg[4]/P0001  & n3503 ;
  assign n6118 = ~n6116 & ~n6117 ;
  assign n6119 = n6094 & n6118 ;
  assign n6120 = n6115 & n6119 ;
  assign n6121 = ~n6098 & ~n6120 ;
  assign n6122 = ~\u1_u2_sizu_c_reg[8]/NET0131  & ~n3546 ;
  assign n6123 = ~\u1_u2_sizu_c_reg[7]/P0001  & ~n3538 ;
  assign n6124 = ~n6122 & ~n6123 ;
  assign n6125 = ~n6083 & n6124 ;
  assign n6126 = n6090 & n6125 ;
  assign n6127 = n6121 & n6126 ;
  assign n6128 = ~n6091 & ~n6127 ;
  assign n6129 = n3610 & ~n6128 ;
  assign n6130 = n5744 & n5754 ;
  assign n6131 = n5742 & n5756 ;
  assign n6132 = n6130 & n6131 ;
  assign n6133 = \u0_u0_state_reg[1]/P0001  & ~\u0_u0_state_reg[2]/NET0131  ;
  assign n6134 = n6132 & n6133 ;
  assign n6135 = n5741 & n5744 ;
  assign n6136 = n5754 & n6135 ;
  assign n6137 = ~\u0_u0_state_reg[4]/NET0131  & \u0_u0_state_reg[5]/P0001  ;
  assign n6138 = n5743 & n6137 ;
  assign n6139 = n5756 & n6138 ;
  assign n6140 = n6136 & n6139 ;
  assign n6141 = ~n6134 & ~n6140 ;
  assign n6142 = n5743 & n5756 ;
  assign n6143 = n6136 & n6142 ;
  assign n6144 = \u0_u0_state_reg[4]/NET0131  & ~\u0_u0_state_reg[5]/P0001  ;
  assign n6145 = ~n6137 & ~n6144 ;
  assign n6146 = n6143 & ~n6145 ;
  assign n6147 = \u0_u0_T1_gt_3_0_mS_reg/P0001  & \u0_u0_mode_hs_reg/P0001  ;
  assign n6148 = ~\u0_u0_idle_long_reg/P0001  & ~\u0_u0_mode_hs_reg/P0001  ;
  assign n6149 = \u0_u0_T1_gt_2_5_uS_reg/P0001  & \u0_u0_T1_st_3_0_mS_reg/P0001  ;
  assign n6150 = n6148 & n6149 ;
  assign n6151 = ~n6147 & ~n6150 ;
  assign n6152 = ~n6146 & ~n6151 ;
  assign n6153 = ~n6141 & n6152 ;
  assign n6154 = n5736 & n5753 ;
  assign n6155 = \u0_u0_state_reg[0]/NET0131  & n5734 ;
  assign n6156 = n6154 & n6155 ;
  assign n6157 = n5746 & n6156 ;
  assign n6158 = ~n6146 & n6157 ;
  assign n6159 = n6141 & n6158 ;
  assign n6160 = n5765 & n6144 ;
  assign n6161 = n6143 & n6160 ;
  assign n6162 = ~n6134 & n6161 ;
  assign n6163 = ~\u0_u0_T2_wakeup_reg/P0001  & ~\u0_u0_state_reg[7]/NET0131  ;
  assign n6164 = n5743 & ~n6163 ;
  assign n6165 = n5756 & n6164 ;
  assign n6166 = n6136 & n6165 ;
  assign n6167 = n6137 & n6166 ;
  assign n6168 = ~n6162 & ~n6167 ;
  assign n6169 = ~n6159 & n6168 ;
  assign n6170 = ~n6153 & n6169 ;
  assign n6171 = n5740 & n5743 ;
  assign n6172 = n5756 & n6171 ;
  assign n6173 = \u0_u0_state_reg[3]/P0001  & ~\u0_u0_state_reg[6]/NET0131  ;
  assign n6174 = n5744 & n6173 ;
  assign n6175 = n5754 & n6174 ;
  assign n6176 = n6172 & n6175 ;
  assign n6177 = ~n6162 & n6176 ;
  assign n6178 = ~\u0_u0_state_reg[1]/P0001  & \u0_u0_state_reg[2]/NET0131  ;
  assign n6179 = n6132 & n6178 ;
  assign n6180 = ~n5939 & ~n6179 ;
  assign n6181 = ~n6177 & n6180 ;
  assign n6182 = ~n6170 & n6181 ;
  assign n6183 = ~n5939 & ~n6146 ;
  assign n6184 = ~n5939 & ~n6176 ;
  assign n6185 = ~n6179 & n6184 ;
  assign n6186 = ~n6183 & ~n6185 ;
  assign n6187 = \u0_u0_T2_gt_1_0_mS_reg/P0001  & ~n6140 ;
  assign n6188 = ~n6134 & n6187 ;
  assign n6189 = ~n6176 & ~n6188 ;
  assign n6190 = n6186 & ~n6189 ;
  assign n6191 = \u0_u0_T1_gt_2_5_uS_reg/P0001  & \u0_u0_ls_se0_r_reg/P0001  ;
  assign n6192 = n5765 & n6191 ;
  assign n6193 = n6176 & n6192 ;
  assign n6194 = \u0_u0_T2_gt_100_uS_reg/P0001  & \u0_u0_ls_j_r_reg/P0001  ;
  assign n6195 = n5759 & n6194 ;
  assign n6196 = \u0_u0_state_reg[9]/P0001  & ~n6195 ;
  assign n6197 = \u0_u0_T2_gt_100_uS_reg/P0001  & \u0_u0_ls_se0_r_reg/P0001  ;
  assign n6198 = n5765 & n6197 ;
  assign n6199 = ~n6196 & ~n6198 ;
  assign n6200 = n6179 & ~n6199 ;
  assign n6201 = ~n6193 & ~n6200 ;
  assign n6202 = \u0_u0_me_cnt_reg[6]/P0001  & \u0_u0_me_cnt_reg[7]/P0001  ;
  assign n6203 = ~\u0_u0_me_cnt_reg[2]/P0001  & \u0_u0_me_cnt_reg[3]/P0001  ;
  assign n6204 = n6202 & n6203 ;
  assign n6205 = ~\u0_u0_me_cnt_reg[4]/P0001  & ~\u0_u0_me_cnt_reg[5]/P0001  ;
  assign n6206 = ~\u0_u0_me_cnt_reg[0]/P0001  & ~\u0_u0_me_cnt_reg[1]/P0001  ;
  assign n6207 = n6205 & n6206 ;
  assign n6208 = n6204 & n6207 ;
  assign n6209 = n6201 & n6208 ;
  assign n6210 = ~n6190 & n6209 ;
  assign n6211 = ~n6182 & n6210 ;
  assign n6212 = \u1_hms_clk_reg/P0001  & \u1_sof_time_reg[0]/P0001  ;
  assign n6213 = \u1_sof_time_reg[6]/P0001  & \u1_sof_time_reg[8]/P0001  ;
  assign n6214 = \u1_sof_time_reg[7]/P0001  & n6213 ;
  assign n6215 = n6212 & n6214 ;
  assign n6216 = \u1_sof_time_reg[3]/P0001  & \u1_sof_time_reg[5]/P0001  ;
  assign n6217 = \u1_sof_time_reg[4]/P0001  & n6216 ;
  assign n6218 = \u1_sof_time_reg[1]/P0001  & \u1_sof_time_reg[2]/P0001  ;
  assign n6219 = \u1_sof_time_reg[10]/P0001  & \u1_sof_time_reg[9]/P0001  ;
  assign n6220 = n6218 & n6219 ;
  assign n6221 = n6217 & n6220 ;
  assign n6222 = n6215 & n6221 ;
  assign n6223 = ~\u1_clr_sof_time_reg/P0001  & \u1_sof_time_reg[11]/P0001  ;
  assign n6224 = ~n6222 & n6223 ;
  assign n6225 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_sof_time_reg[11]/P0001  ;
  assign n6226 = n6222 & n6225 ;
  assign n6227 = ~n6224 & ~n6226 ;
  assign n6228 = ~n5669 & n5675 ;
  assign n6229 = ~n5679 & ~n5681 ;
  assign n6230 = ~n5670 & ~n5680 ;
  assign n6231 = n6229 & n6230 ;
  assign n6232 = ~n6228 & n6231 ;
  assign n6233 = n5723 & n6231 ;
  assign n6234 = ~n5720 & n6233 ;
  assign n6235 = ~n6232 & ~n6234 ;
  assign n6236 = ~n6228 & n6229 ;
  assign n6237 = n5723 & n6229 ;
  assign n6238 = ~n5720 & n6237 ;
  assign n6239 = ~n6236 & ~n6238 ;
  assign n6240 = ~n6230 & n6239 ;
  assign n6241 = n6235 & ~n6240 ;
  assign n6242 = \u4_u3_csr0_reg[3]/NET0131  & ~\u4_u3_dma_in_cnt_reg[1]/P0001  ;
  assign n6243 = \u4_u3_csr0_reg[2]/P0001  & ~\u4_u3_dma_in_cnt_reg[0]/P0001  ;
  assign n6244 = ~n6242 & ~n6243 ;
  assign n6245 = ~\u4_u3_csr0_reg[4]/P0001  & \u4_u3_dma_in_cnt_reg[2]/P0001  ;
  assign n6246 = ~\u4_u3_csr0_reg[3]/NET0131  & \u4_u3_dma_in_cnt_reg[1]/P0001  ;
  assign n6247 = ~n6245 & ~n6246 ;
  assign n6248 = ~n6244 & n6247 ;
  assign n6249 = \u4_u3_csr0_reg[6]/P0001  & ~\u4_u3_dma_in_cnt_reg[4]/P0001  ;
  assign n6250 = \u4_u3_csr0_reg[7]/P0001  & ~\u4_u3_dma_in_cnt_reg[5]/P0001  ;
  assign n6251 = ~n6249 & ~n6250 ;
  assign n6252 = \u4_u3_csr0_reg[5]/P0001  & ~\u4_u3_dma_in_cnt_reg[3]/P0001  ;
  assign n6253 = \u4_u3_csr0_reg[4]/P0001  & ~\u4_u3_dma_in_cnt_reg[2]/P0001  ;
  assign n6254 = ~n6252 & ~n6253 ;
  assign n6255 = n6251 & n6254 ;
  assign n6256 = ~n6248 & n6255 ;
  assign n6257 = ~\u4_u3_csr0_reg[5]/P0001  & \u4_u3_dma_in_cnt_reg[3]/P0001  ;
  assign n6258 = ~\u4_u3_csr0_reg[6]/P0001  & \u4_u3_dma_in_cnt_reg[4]/P0001  ;
  assign n6259 = ~n6257 & ~n6258 ;
  assign n6260 = n6251 & ~n6259 ;
  assign n6261 = ~\u4_u3_csr0_reg[8]/P0001  & \u4_u3_dma_in_cnt_reg[6]/P0001  ;
  assign n6262 = ~\u4_u3_csr0_reg[7]/P0001  & \u4_u3_dma_in_cnt_reg[5]/P0001  ;
  assign n6263 = ~n6261 & ~n6262 ;
  assign n6264 = ~n6260 & n6263 ;
  assign n6265 = ~n6256 & n6264 ;
  assign n6266 = \u4_u3_csr0_reg[10]/P0001  & ~\u4_u3_dma_in_cnt_reg[8]/P0001  ;
  assign n6267 = \u4_u3_csr0_reg[9]/P0001  & ~\u4_u3_dma_in_cnt_reg[7]/P0001  ;
  assign n6268 = ~n6266 & ~n6267 ;
  assign n6269 = \u4_u3_csr0_reg[8]/P0001  & ~\u4_u3_dma_in_cnt_reg[6]/P0001  ;
  assign n6270 = n6268 & ~n6269 ;
  assign n6271 = ~n6265 & n6270 ;
  assign n6272 = \u4_u3_dma_in_cnt_reg[4]/P0001  & \u4_u3_dma_in_cnt_reg[6]/P0001  ;
  assign n6273 = \u4_u3_dma_in_cnt_reg[5]/P0001  & n6272 ;
  assign n6274 = \u4_u3_dma_in_cnt_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[1]/P0001  ;
  assign n6275 = \u4_u3_dma_in_cnt_reg[2]/P0001  & \u4_u3_dma_in_cnt_reg[3]/P0001  ;
  assign n6276 = n6274 & n6275 ;
  assign n6277 = n6273 & n6276 ;
  assign n6278 = \u4_u3_dma_in_cnt_reg[7]/P0001  & \u4_u3_dma_in_cnt_reg[8]/P0001  ;
  assign n6279 = n6277 & n6278 ;
  assign n6280 = \u4_u3_r5_reg/NET0131  & ~n6279 ;
  assign n6281 = ~\u1_u3_buf0_rl_reg/P0001  & ~\u1_u3_buf0_set_reg/P0001  ;
  assign n6282 = ~\u4_u3_set_r_reg/P0001  & n6281 ;
  assign n6283 = ~\u4_u3_csr0_reg[10]/P0001  & \u4_u3_dma_in_cnt_reg[8]/P0001  ;
  assign n6284 = \u4_u3_ep_match_r_reg/P0001  & ~n6283 ;
  assign n6285 = ~n6282 & n6284 ;
  assign n6286 = ~\u4_u3_csr0_reg[9]/P0001  & \u4_u3_dma_in_cnt_reg[7]/P0001  ;
  assign n6287 = ~n6266 & n6286 ;
  assign n6288 = n6285 & ~n6287 ;
  assign n6289 = ~n6280 & n6288 ;
  assign n6290 = ~n6271 & n6289 ;
  assign n6291 = \u4_u3_r5_reg/NET0131  & n6278 ;
  assign n6292 = n6277 & n6291 ;
  assign n6293 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[9]/P0001  ;
  assign n6294 = ~n6292 & n6293 ;
  assign n6295 = ~n6290 & n6294 ;
  assign n6296 = ~n6290 & ~n6292 ;
  assign n6297 = \u4_u3_csr1_reg[0]/P0001  & ~\u4_u3_dma_in_cnt_reg[9]/P0001  ;
  assign n6298 = ~n6296 & n6297 ;
  assign n6299 = ~n6295 & ~n6298 ;
  assign n6300 = \u4_u0_csr0_reg[3]/NET0131  & ~\u4_u0_dma_in_cnt_reg[1]/P0001  ;
  assign n6301 = \u4_u0_csr0_reg[2]/P0001  & ~\u4_u0_dma_in_cnt_reg[0]/P0001  ;
  assign n6302 = ~n6300 & ~n6301 ;
  assign n6303 = ~\u4_u0_csr0_reg[4]/P0001  & \u4_u0_dma_in_cnt_reg[2]/P0001  ;
  assign n6304 = ~\u4_u0_csr0_reg[3]/NET0131  & \u4_u0_dma_in_cnt_reg[1]/P0001  ;
  assign n6305 = ~n6303 & ~n6304 ;
  assign n6306 = ~n6302 & n6305 ;
  assign n6307 = \u4_u0_csr0_reg[6]/P0001  & ~\u4_u0_dma_in_cnt_reg[4]/P0001  ;
  assign n6308 = \u4_u0_csr0_reg[7]/P0001  & ~\u4_u0_dma_in_cnt_reg[5]/P0001  ;
  assign n6309 = ~n6307 & ~n6308 ;
  assign n6310 = \u4_u0_csr0_reg[5]/P0001  & ~\u4_u0_dma_in_cnt_reg[3]/P0001  ;
  assign n6311 = \u4_u0_csr0_reg[4]/P0001  & ~\u4_u0_dma_in_cnt_reg[2]/P0001  ;
  assign n6312 = ~n6310 & ~n6311 ;
  assign n6313 = n6309 & n6312 ;
  assign n6314 = ~n6306 & n6313 ;
  assign n6315 = ~\u4_u0_csr0_reg[5]/P0001  & \u4_u0_dma_in_cnt_reg[3]/P0001  ;
  assign n6316 = ~\u4_u0_csr0_reg[6]/P0001  & \u4_u0_dma_in_cnt_reg[4]/P0001  ;
  assign n6317 = ~n6315 & ~n6316 ;
  assign n6318 = n6309 & ~n6317 ;
  assign n6319 = ~\u4_u0_csr0_reg[8]/P0001  & \u4_u0_dma_in_cnt_reg[6]/P0001  ;
  assign n6320 = ~\u4_u0_csr0_reg[7]/P0001  & \u4_u0_dma_in_cnt_reg[5]/P0001  ;
  assign n6321 = ~n6319 & ~n6320 ;
  assign n6322 = ~n6318 & n6321 ;
  assign n6323 = ~n6314 & n6322 ;
  assign n6324 = \u4_u0_csr0_reg[10]/P0001  & ~\u4_u0_dma_in_cnt_reg[8]/P0001  ;
  assign n6325 = \u4_u0_csr0_reg[9]/P0001  & ~\u4_u0_dma_in_cnt_reg[7]/P0001  ;
  assign n6326 = ~n6324 & ~n6325 ;
  assign n6327 = \u4_u0_csr0_reg[8]/P0001  & ~\u4_u0_dma_in_cnt_reg[6]/P0001  ;
  assign n6328 = n6326 & ~n6327 ;
  assign n6329 = ~n6323 & n6328 ;
  assign n6330 = \u4_u0_dma_in_cnt_reg[4]/P0001  & \u4_u0_dma_in_cnt_reg[6]/P0001  ;
  assign n6331 = \u4_u0_dma_in_cnt_reg[5]/P0001  & n6330 ;
  assign n6332 = \u4_u0_dma_in_cnt_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[1]/P0001  ;
  assign n6333 = \u4_u0_dma_in_cnt_reg[2]/P0001  & \u4_u0_dma_in_cnt_reg[3]/P0001  ;
  assign n6334 = n6332 & n6333 ;
  assign n6335 = n6331 & n6334 ;
  assign n6336 = \u4_u0_dma_in_cnt_reg[7]/P0001  & \u4_u0_dma_in_cnt_reg[8]/P0001  ;
  assign n6337 = n6335 & n6336 ;
  assign n6338 = \u4_u0_r5_reg/NET0131  & ~n6337 ;
  assign n6339 = ~\u4_u0_set_r_reg/P0001  & n6281 ;
  assign n6340 = ~\u4_u0_csr0_reg[10]/P0001  & \u4_u0_dma_in_cnt_reg[8]/P0001  ;
  assign n6341 = \u4_u0_ep_match_r_reg/P0001  & ~n6340 ;
  assign n6342 = ~n6339 & n6341 ;
  assign n6343 = ~\u4_u0_csr0_reg[9]/P0001  & \u4_u0_dma_in_cnt_reg[7]/P0001  ;
  assign n6344 = ~n6324 & n6343 ;
  assign n6345 = n6342 & ~n6344 ;
  assign n6346 = ~n6338 & n6345 ;
  assign n6347 = ~n6329 & n6346 ;
  assign n6348 = \u4_u0_r5_reg/NET0131  & n6336 ;
  assign n6349 = n6335 & n6348 ;
  assign n6350 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[9]/P0001  ;
  assign n6351 = ~n6349 & n6350 ;
  assign n6352 = ~n6347 & n6351 ;
  assign n6353 = ~n6347 & ~n6349 ;
  assign n6354 = \u4_u0_csr1_reg[0]/P0001  & ~\u4_u0_dma_in_cnt_reg[9]/P0001  ;
  assign n6355 = ~n6353 & n6354 ;
  assign n6356 = ~n6352 & ~n6355 ;
  assign n6357 = \u4_u1_dma_in_cnt_reg[4]/P0001  & \u4_u1_dma_in_cnt_reg[6]/P0001  ;
  assign n6358 = \u4_u1_dma_in_cnt_reg[5]/P0001  & n6357 ;
  assign n6359 = \u4_u1_dma_in_cnt_reg[0]/P0001  & \u4_u1_dma_in_cnt_reg[1]/P0001  ;
  assign n6360 = \u4_u1_dma_in_cnt_reg[2]/P0001  & \u4_u1_dma_in_cnt_reg[3]/P0001  ;
  assign n6361 = n6359 & n6360 ;
  assign n6362 = n6358 & n6361 ;
  assign n6363 = \u4_u1_dma_in_cnt_reg[7]/P0001  & \u4_u1_dma_in_cnt_reg[8]/P0001  ;
  assign n6364 = \u4_u1_r5_reg/NET0131  & n6363 ;
  assign n6365 = n6362 & n6364 ;
  assign n6366 = n6362 & n6363 ;
  assign n6367 = \u4_u1_r5_reg/NET0131  & ~n6366 ;
  assign n6368 = ~\u4_u1_set_r_reg/P0001  & n6281 ;
  assign n6369 = \u4_u1_ep_match_r_reg/P0001  & ~n6368 ;
  assign n6370 = ~\u4_u1_csr0_reg[10]/P0001  & \u4_u1_dma_in_cnt_reg[8]/P0001  ;
  assign n6371 = \u4_u1_csr0_reg[10]/P0001  & ~\u4_u1_dma_in_cnt_reg[8]/P0001  ;
  assign n6372 = ~\u4_u1_csr0_reg[9]/P0001  & \u4_u1_dma_in_cnt_reg[7]/P0001  ;
  assign n6373 = ~n6371 & n6372 ;
  assign n6374 = ~n6370 & ~n6373 ;
  assign n6375 = n6369 & n6374 ;
  assign n6376 = ~n6367 & n6375 ;
  assign n6377 = ~n6365 & ~n6376 ;
  assign n6378 = ~\u4_u1_csr0_reg[8]/P0001  & \u4_u1_dma_in_cnt_reg[6]/P0001  ;
  assign n6379 = \u4_u1_csr0_reg[7]/P0001  & ~\u4_u1_dma_in_cnt_reg[5]/P0001  ;
  assign n6380 = ~n6378 & n6379 ;
  assign n6381 = \u4_u1_csr0_reg[6]/P0001  & ~\u4_u1_dma_in_cnt_reg[4]/P0001  ;
  assign n6382 = \u4_u1_csr0_reg[5]/P0001  & ~\u4_u1_dma_in_cnt_reg[3]/P0001  ;
  assign n6383 = ~n6381 & ~n6382 ;
  assign n6384 = ~\u4_u1_csr0_reg[5]/P0001  & \u4_u1_dma_in_cnt_reg[3]/P0001  ;
  assign n6385 = n6383 & n6384 ;
  assign n6386 = \u4_u1_csr0_reg[3]/NET0131  & ~\u4_u1_dma_in_cnt_reg[1]/P0001  ;
  assign n6387 = \u4_u1_csr0_reg[2]/P0001  & ~\u4_u1_dma_in_cnt_reg[0]/P0001  ;
  assign n6388 = ~n6386 & ~n6387 ;
  assign n6389 = ~\u4_u1_csr0_reg[4]/P0001  & \u4_u1_dma_in_cnt_reg[2]/P0001  ;
  assign n6390 = ~\u4_u1_csr0_reg[3]/NET0131  & \u4_u1_dma_in_cnt_reg[1]/P0001  ;
  assign n6391 = ~n6389 & ~n6390 ;
  assign n6392 = ~n6388 & n6391 ;
  assign n6393 = \u4_u1_csr0_reg[4]/P0001  & ~\u4_u1_dma_in_cnt_reg[2]/P0001  ;
  assign n6394 = n6383 & ~n6393 ;
  assign n6395 = ~n6392 & n6394 ;
  assign n6396 = ~n6385 & ~n6395 ;
  assign n6397 = ~\u4_u1_csr0_reg[7]/P0001  & \u4_u1_dma_in_cnt_reg[5]/P0001  ;
  assign n6398 = ~\u4_u1_csr0_reg[6]/P0001  & \u4_u1_dma_in_cnt_reg[4]/P0001  ;
  assign n6399 = ~n6397 & ~n6398 ;
  assign n6400 = ~n6378 & n6399 ;
  assign n6401 = n6396 & n6400 ;
  assign n6402 = ~n6380 & ~n6401 ;
  assign n6403 = \u4_u1_csr0_reg[9]/P0001  & ~\u4_u1_dma_in_cnt_reg[7]/P0001  ;
  assign n6404 = ~n6371 & ~n6403 ;
  assign n6405 = \u4_u1_csr0_reg[8]/P0001  & ~\u4_u1_dma_in_cnt_reg[6]/P0001  ;
  assign n6406 = n6404 & ~n6405 ;
  assign n6407 = ~n6365 & n6406 ;
  assign n6408 = n6402 & n6407 ;
  assign n6409 = ~n6377 & ~n6408 ;
  assign n6410 = \u4_u1_csr1_reg[0]/P0001  & \u4_u1_dma_in_cnt_reg[9]/P0001  ;
  assign n6411 = ~n6409 & n6410 ;
  assign n6412 = \u4_u1_csr1_reg[0]/P0001  & ~\u4_u1_dma_in_cnt_reg[9]/P0001  ;
  assign n6413 = n6409 & n6412 ;
  assign n6414 = ~n6411 & ~n6413 ;
  assign n6415 = ~\u4_u2_set_r_reg/P0001  & n6281 ;
  assign n6416 = \u4_u2_csr0_reg[10]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n6417 = ~\u4_u2_dma_in_cnt_reg[8]/P0001  & n6416 ;
  assign n6418 = ~n6415 & n6417 ;
  assign n6419 = ~\u4_u2_csr0_reg[10]/P0001  & \u4_u2_dma_in_cnt_reg[8]/P0001  ;
  assign n6420 = \u4_u2_ep_match_r_reg/P0001  & ~n6419 ;
  assign n6421 = ~n6415 & n6420 ;
  assign n6422 = ~\u4_u2_csr0_reg[9]/P0001  & \u4_u2_dma_in_cnt_reg[7]/P0001  ;
  assign n6423 = n6421 & ~n6422 ;
  assign n6424 = ~n6418 & ~n6423 ;
  assign n6425 = ~\u4_u2_csr0_reg[8]/P0001  & \u4_u2_dma_in_cnt_reg[6]/P0001  ;
  assign n6426 = \u4_u2_csr0_reg[7]/P0001  & ~\u4_u2_dma_in_cnt_reg[5]/P0001  ;
  assign n6427 = ~n6425 & n6426 ;
  assign n6428 = \u4_u2_csr0_reg[6]/P0001  & ~\u4_u2_dma_in_cnt_reg[4]/P0001  ;
  assign n6429 = \u4_u2_csr0_reg[5]/P0001  & ~\u4_u2_dma_in_cnt_reg[3]/P0001  ;
  assign n6430 = ~n6428 & ~n6429 ;
  assign n6431 = ~\u4_u2_csr0_reg[5]/P0001  & \u4_u2_dma_in_cnt_reg[3]/P0001  ;
  assign n6432 = n6430 & n6431 ;
  assign n6433 = \u4_u2_csr0_reg[3]/NET0131  & ~\u4_u2_dma_in_cnt_reg[1]/P0001  ;
  assign n6434 = \u4_u2_csr0_reg[2]/P0001  & ~\u4_u2_dma_in_cnt_reg[0]/P0001  ;
  assign n6435 = ~n6433 & ~n6434 ;
  assign n6436 = ~\u4_u2_csr0_reg[4]/P0001  & \u4_u2_dma_in_cnt_reg[2]/P0001  ;
  assign n6437 = ~\u4_u2_csr0_reg[3]/NET0131  & \u4_u2_dma_in_cnt_reg[1]/P0001  ;
  assign n6438 = ~n6436 & ~n6437 ;
  assign n6439 = ~n6435 & n6438 ;
  assign n6440 = \u4_u2_csr0_reg[4]/P0001  & ~\u4_u2_dma_in_cnt_reg[2]/P0001  ;
  assign n6441 = n6430 & ~n6440 ;
  assign n6442 = ~n6439 & n6441 ;
  assign n6443 = ~n6432 & ~n6442 ;
  assign n6444 = ~\u4_u2_csr0_reg[7]/P0001  & \u4_u2_dma_in_cnt_reg[5]/P0001  ;
  assign n6445 = ~\u4_u2_csr0_reg[6]/P0001  & \u4_u2_dma_in_cnt_reg[4]/P0001  ;
  assign n6446 = ~n6444 & ~n6445 ;
  assign n6447 = ~n6425 & n6446 ;
  assign n6448 = n6443 & n6447 ;
  assign n6449 = ~n6427 & ~n6448 ;
  assign n6450 = \u4_u2_csr0_reg[9]/P0001  & ~\u4_u2_dma_in_cnt_reg[7]/P0001  ;
  assign n6451 = \u4_u2_csr0_reg[8]/P0001  & ~\u4_u2_dma_in_cnt_reg[6]/P0001  ;
  assign n6452 = ~n6450 & ~n6451 ;
  assign n6453 = ~n6418 & n6452 ;
  assign n6454 = n6449 & n6453 ;
  assign n6455 = ~n6424 & ~n6454 ;
  assign n6456 = ~\u4_u2_r5_reg/NET0131  & ~n6455 ;
  assign n6457 = \u4_u2_dma_in_cnt_reg[9]/P0001  & ~\u4_u2_r5_reg/NET0131  ;
  assign n6458 = \u4_u2_dma_in_cnt_reg[4]/P0001  & \u4_u2_dma_in_cnt_reg[6]/P0001  ;
  assign n6459 = \u4_u2_dma_in_cnt_reg[5]/P0001  & n6458 ;
  assign n6460 = \u4_u2_dma_in_cnt_reg[0]/P0001  & \u4_u2_dma_in_cnt_reg[1]/P0001  ;
  assign n6461 = \u4_u2_dma_in_cnt_reg[2]/P0001  & \u4_u2_dma_in_cnt_reg[3]/P0001  ;
  assign n6462 = n6460 & n6461 ;
  assign n6463 = n6459 & n6462 ;
  assign n6464 = \u4_u2_dma_in_cnt_reg[7]/P0001  & \u4_u2_dma_in_cnt_reg[8]/P0001  ;
  assign n6465 = \u4_u2_dma_in_cnt_reg[9]/P0001  & n6464 ;
  assign n6466 = n6463 & n6465 ;
  assign n6467 = ~n6457 & ~n6466 ;
  assign n6468 = ~n6456 & ~n6467 ;
  assign n6469 = ~\u4_u2_dma_in_cnt_reg[9]/P0001  & ~\u4_u2_r5_reg/NET0131  ;
  assign n6470 = ~n6455 & n6469 ;
  assign n6471 = n6463 & n6464 ;
  assign n6472 = ~\u4_u2_dma_in_cnt_reg[9]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n6473 = ~n6471 & n6472 ;
  assign n6474 = \u4_u2_csr1_reg[0]/P0001  & ~n6473 ;
  assign n6475 = ~n6470 & n6474 ;
  assign n6476 = ~n6468 & n6475 ;
  assign n6477 = rst_i_pad & ~\u1_clr_sof_time_reg/P0001  ;
  assign n6478 = ~\u1_hms_clk_reg/P0001  & n6477 ;
  assign n6479 = \u1_hms_cnt_reg[0]/P0001  & \u1_hms_cnt_reg[1]/P0001  ;
  assign n6480 = ~\u1_hms_cnt_reg[0]/P0001  & ~\u1_hms_cnt_reg[1]/P0001  ;
  assign n6481 = ~n6479 & ~n6480 ;
  assign n6482 = n6478 & n6481 ;
  assign n6483 = \u1_hms_cnt_reg[2]/P0001  & n6479 ;
  assign n6484 = ~\u1_hms_cnt_reg[2]/P0001  & ~n6479 ;
  assign n6485 = ~n6483 & ~n6484 ;
  assign n6486 = n6478 & n6485 ;
  assign n6487 = ~\u1_hms_cnt_reg[3]/P0001  & ~n6483 ;
  assign n6488 = \u1_hms_cnt_reg[2]/P0001  & \u1_hms_cnt_reg[3]/P0001  ;
  assign n6489 = n6479 & n6488 ;
  assign n6490 = n6478 & ~n6489 ;
  assign n6491 = ~n6487 & n6490 ;
  assign n6492 = ~\u1_hms_clk_reg/P0001  & \u1_hms_cnt_reg[4]/P0001  ;
  assign n6493 = n6477 & n6492 ;
  assign n6494 = ~n6489 & n6493 ;
  assign n6495 = ~\u1_hms_clk_reg/P0001  & ~\u1_hms_cnt_reg[4]/P0001  ;
  assign n6496 = n6477 & n6495 ;
  assign n6497 = n6489 & n6496 ;
  assign n6498 = ~n6494 & ~n6497 ;
  assign n6499 = \u1_u0_token_valid_str1_reg/P0001  & ~n5116 ;
  assign n6500 = n5012 & ~n6499 ;
  assign n6501 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token0_reg[0]/NET0131  ;
  assign n6502 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[0]/P0001  ;
  assign n6503 = rst_i_pad & ~n6502 ;
  assign n6504 = ~n6501 & n6503 ;
  assign n6505 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token1_reg[2]/P0001  ;
  assign n6506 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[10]/P0001  ;
  assign n6507 = rst_i_pad & ~n6506 ;
  assign n6508 = ~n6505 & n6507 ;
  assign n6509 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token0_reg[1]/P0001  ;
  assign n6510 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[1]/P0001  ;
  assign n6511 = rst_i_pad & ~n6510 ;
  assign n6512 = ~n6509 & n6511 ;
  assign n6513 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token0_reg[3]/NET0131  ;
  assign n6514 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[3]/P0001  ;
  assign n6515 = rst_i_pad & ~n6514 ;
  assign n6516 = ~n6513 & n6515 ;
  assign n6517 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token0_reg[2]/NET0131  ;
  assign n6518 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[2]/P0001  ;
  assign n6519 = rst_i_pad & ~n6518 ;
  assign n6520 = ~n6517 & n6519 ;
  assign n6521 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token0_reg[4]/P0001  ;
  assign n6522 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[4]/P0001  ;
  assign n6523 = rst_i_pad & ~n6522 ;
  assign n6524 = ~n6521 & n6523 ;
  assign n6525 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token0_reg[5]/NET0131  ;
  assign n6526 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[5]/P0001  ;
  assign n6527 = rst_i_pad & ~n6526 ;
  assign n6528 = ~n6525 & n6527 ;
  assign n6529 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token0_reg[6]/P0001  ;
  assign n6530 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[6]/P0001  ;
  assign n6531 = rst_i_pad & ~n6530 ;
  assign n6532 = ~n6529 & n6531 ;
  assign n6533 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token0_reg[7]/P0001  ;
  assign n6534 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[7]/P0001  ;
  assign n6535 = rst_i_pad & ~n6534 ;
  assign n6536 = ~n6533 & n6535 ;
  assign n6537 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token1_reg[0]/P0001  ;
  assign n6538 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[8]/P0001  ;
  assign n6539 = rst_i_pad & ~n6538 ;
  assign n6540 = ~n6537 & n6539 ;
  assign n6541 = \u1_clr_sof_time_reg/P0001  & ~\u1_u0_token1_reg[1]/P0001  ;
  assign n6542 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_frame_no_r_reg[9]/P0001  ;
  assign n6543 = rst_i_pad & ~n6542 ;
  assign n6544 = ~n6541 & n6543 ;
  assign n6545 = \u1_u2_sizu_c_reg[4]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n6546 = \u1_u3_new_size_reg[4]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n6547 = ~n6545 & ~n6546 ;
  assign n6548 = \u1_u2_sizu_c_reg[5]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n6549 = \u1_u3_new_size_reg[5]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n6550 = ~n6548 & ~n6549 ;
  assign n6551 = \u1_u3_new_size_reg[6]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n6552 = \u1_u2_sizu_c_reg[6]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n6553 = ~n6551 & ~n6552 ;
  assign n6554 = \u1_u3_new_size_reg[7]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n6555 = \u1_u2_sizu_c_reg[7]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n6556 = ~n6554 & ~n6555 ;
  assign n6557 = ~n5692 & ~n5695 ;
  assign n6558 = ~n5944 & n5951 ;
  assign n6559 = ~n5946 & n6558 ;
  assign n6560 = n6557 & n6559 ;
  assign n6561 = ~n6557 & ~n6559 ;
  assign n6562 = ~n6560 & ~n6561 ;
  assign n6563 = ~n5669 & ~n5721 ;
  assign n6564 = ~n5959 & ~n6563 ;
  assign n6565 = n5952 & ~n6563 ;
  assign n6566 = n5947 & n6565 ;
  assign n6567 = ~n6564 & ~n6566 ;
  assign n6568 = n5959 & n6563 ;
  assign n6569 = ~n5953 & n6568 ;
  assign n6570 = n6567 & ~n6569 ;
  assign n6571 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[8]/P0001  ;
  assign n6572 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[7]/P0001  ;
  assign n6573 = n6277 & n6572 ;
  assign n6574 = ~n6571 & ~n6573 ;
  assign n6575 = n6280 & ~n6574 ;
  assign n6576 = ~\u4_u3_dma_in_cnt_reg[8]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n6577 = n6281 & n6576 ;
  assign n6578 = ~\u4_u3_dma_in_cnt_reg[8]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n6579 = \u4_u3_csr1_reg[0]/P0001  & ~\u4_u3_r5_reg/NET0131  ;
  assign n6580 = ~n6578 & n6579 ;
  assign n6581 = ~n6577 & n6580 ;
  assign n6582 = ~n6266 & ~n6283 ;
  assign n6583 = ~n6245 & ~n6257 ;
  assign n6584 = ~n6252 & ~n6583 ;
  assign n6585 = n6251 & n6584 ;
  assign n6586 = ~n6244 & ~n6246 ;
  assign n6587 = n6255 & ~n6586 ;
  assign n6588 = ~n6585 & ~n6587 ;
  assign n6589 = ~n6261 & ~n6286 ;
  assign n6590 = ~n6258 & ~n6262 ;
  assign n6591 = ~n6250 & ~n6590 ;
  assign n6592 = n6589 & ~n6591 ;
  assign n6593 = n6588 & n6592 ;
  assign n6594 = n6269 & ~n6286 ;
  assign n6595 = ~n6267 & ~n6594 ;
  assign n6596 = ~n6593 & n6595 ;
  assign n6597 = n6582 & ~n6596 ;
  assign n6598 = \u4_u3_ep_match_r_reg/P0001  & ~n6282 ;
  assign n6599 = ~n6582 & n6595 ;
  assign n6600 = ~n6593 & n6599 ;
  assign n6601 = n6598 & ~n6600 ;
  assign n6602 = ~n6597 & n6601 ;
  assign n6603 = n6581 & ~n6602 ;
  assign n6604 = ~n6575 & ~n6603 ;
  assign n6605 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[8]/P0001  ;
  assign n6606 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[7]/P0001  ;
  assign n6607 = n6335 & n6606 ;
  assign n6608 = ~n6605 & ~n6607 ;
  assign n6609 = n6338 & ~n6608 ;
  assign n6610 = ~\u4_u0_dma_in_cnt_reg[8]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n6611 = n6281 & n6610 ;
  assign n6612 = ~\u4_u0_dma_in_cnt_reg[8]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n6613 = \u4_u0_csr1_reg[0]/P0001  & ~\u4_u0_r5_reg/NET0131  ;
  assign n6614 = ~n6612 & n6613 ;
  assign n6615 = ~n6611 & n6614 ;
  assign n6616 = ~n6324 & ~n6340 ;
  assign n6617 = ~n6303 & ~n6315 ;
  assign n6618 = ~n6310 & ~n6617 ;
  assign n6619 = n6309 & n6618 ;
  assign n6620 = ~n6302 & ~n6304 ;
  assign n6621 = n6313 & ~n6620 ;
  assign n6622 = ~n6619 & ~n6621 ;
  assign n6623 = ~n6319 & ~n6343 ;
  assign n6624 = ~n6316 & ~n6320 ;
  assign n6625 = ~n6308 & ~n6624 ;
  assign n6626 = n6623 & ~n6625 ;
  assign n6627 = n6622 & n6626 ;
  assign n6628 = n6327 & ~n6343 ;
  assign n6629 = ~n6325 & ~n6628 ;
  assign n6630 = ~n6627 & n6629 ;
  assign n6631 = n6616 & ~n6630 ;
  assign n6632 = \u4_u0_ep_match_r_reg/P0001  & ~n6339 ;
  assign n6633 = ~n6616 & n6629 ;
  assign n6634 = ~n6627 & n6633 ;
  assign n6635 = n6632 & ~n6634 ;
  assign n6636 = ~n6631 & n6635 ;
  assign n6637 = n6615 & ~n6636 ;
  assign n6638 = ~n6609 & ~n6637 ;
  assign n6639 = ~\u4_u1_dma_in_cnt_reg[8]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n6640 = n6281 & n6639 ;
  assign n6641 = ~\u4_u1_dma_in_cnt_reg[8]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n6642 = \u4_u1_csr1_reg[0]/P0001  & ~\u4_u1_r5_reg/NET0131  ;
  assign n6643 = ~n6641 & n6642 ;
  assign n6644 = ~n6640 & n6643 ;
  assign n6645 = \u4_u1_dma_in_cnt_reg[7]/P0001  & n6362 ;
  assign n6646 = ~\u4_u1_dma_in_cnt_reg[8]/P0001  & ~n6645 ;
  assign n6647 = \u4_u1_csr1_reg[0]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n6648 = ~n6366 & n6647 ;
  assign n6649 = ~n6646 & n6648 ;
  assign n6650 = ~n6644 & ~n6649 ;
  assign n6651 = ~n6370 & ~n6371 ;
  assign n6652 = n6403 & n6651 ;
  assign n6653 = n6396 & n6399 ;
  assign n6654 = ~n6379 & ~n6405 ;
  assign n6655 = ~n6653 & n6654 ;
  assign n6656 = ~n6372 & ~n6378 ;
  assign n6657 = n6651 & n6656 ;
  assign n6658 = ~n6655 & n6657 ;
  assign n6659 = ~n6652 & ~n6658 ;
  assign n6660 = ~n6655 & n6656 ;
  assign n6661 = ~n6403 & ~n6651 ;
  assign n6662 = ~n6660 & n6661 ;
  assign n6663 = n6659 & ~n6662 ;
  assign n6664 = n6369 & ~n6649 ;
  assign n6665 = n6663 & n6664 ;
  assign n6666 = ~n6650 & ~n6665 ;
  assign n6667 = \u4_u2_ep_match_r_reg/P0001  & ~n6415 ;
  assign n6668 = \u4_u2_csr0_reg[10]/P0001  & ~\u4_u2_dma_in_cnt_reg[8]/P0001  ;
  assign n6669 = ~n6419 & ~n6668 ;
  assign n6670 = n6667 & n6669 ;
  assign n6671 = \u4_u2_ep_match_r_reg/P0001  & ~n6422 ;
  assign n6672 = ~n6415 & n6671 ;
  assign n6673 = ~n6670 & ~n6672 ;
  assign n6674 = n6452 & ~n6670 ;
  assign n6675 = n6449 & n6674 ;
  assign n6676 = ~n6673 & ~n6675 ;
  assign n6677 = \u4_u2_r5_reg/NET0131  & ~n6471 ;
  assign n6678 = \u4_u2_dma_in_cnt_reg[7]/P0001  & n6463 ;
  assign n6679 = ~\u4_u2_dma_in_cnt_reg[8]/P0001  & ~n6678 ;
  assign n6680 = n6677 & ~n6679 ;
  assign n6681 = ~n6422 & n6669 ;
  assign n6682 = ~n6680 & ~n6681 ;
  assign n6683 = n6452 & ~n6680 ;
  assign n6684 = n6449 & n6683 ;
  assign n6685 = ~n6682 & ~n6684 ;
  assign n6686 = n6676 & ~n6685 ;
  assign n6687 = ~\u4_u2_dma_in_cnt_reg[8]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n6688 = n6281 & n6687 ;
  assign n6689 = ~\u4_u2_dma_in_cnt_reg[8]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n6690 = ~\u4_u2_r5_reg/NET0131  & ~n6689 ;
  assign n6691 = ~n6688 & n6690 ;
  assign n6692 = ~n6680 & ~n6691 ;
  assign n6693 = \u4_u2_csr1_reg[0]/P0001  & ~n6692 ;
  assign n6694 = ~n6686 & n6693 ;
  assign n6695 = ~n6190 & n6201 ;
  assign n6696 = ~\u0_u0_me_ps2_reg[0]/P0001  & ~\u0_u0_me_ps2_reg[1]/P0001  ;
  assign n6697 = ~\u0_u0_me_ps2_reg[2]/P0001  & ~\u0_u0_me_ps2_reg[4]/P0001  ;
  assign n6698 = n6696 & n6697 ;
  assign n6699 = ~\u0_u0_me_ps2_reg[3]/P0001  & ~\u0_u0_me_ps2_reg[4]/P0001  ;
  assign n6700 = \u0_u0_me_ps2_reg[5]/P0001  & ~n6699 ;
  assign n6701 = ~n6698 & n6700 ;
  assign n6702 = ~\u0_u0_me_ps2_reg[6]/P0001  & ~\u0_u0_me_ps2_reg[7]/P0001  ;
  assign n6703 = ~n6701 & n6702 ;
  assign n6704 = n6695 & ~n6703 ;
  assign n6705 = ~n6182 & n6704 ;
  assign n6706 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & ~\u0_u0_me_ps_reg[0]/P0001  ;
  assign n6707 = n6695 & n6706 ;
  assign n6708 = ~n6182 & n6707 ;
  assign n6709 = \u0_u0_me_ps_reg[0]/P0001  & \u0_u0_me_ps_reg[1]/P0001  ;
  assign n6710 = \u0_u0_me_ps_reg[2]/P0001  & \u0_u0_me_ps_reg[3]/P0001  ;
  assign n6711 = n6709 & n6710 ;
  assign n6712 = \u0_u0_me_ps_reg[4]/P0001  & \u0_u0_me_ps_reg[5]/P0001  ;
  assign n6713 = n6711 & n6712 ;
  assign n6714 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & \u0_u0_me_ps_reg[5]/P0001  ;
  assign n6715 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & \u0_u0_me_ps_reg[4]/P0001  ;
  assign n6716 = n6711 & n6715 ;
  assign n6717 = ~n6714 & ~n6716 ;
  assign n6718 = ~n6713 & ~n6717 ;
  assign n6719 = n6695 & n6718 ;
  assign n6720 = ~n6182 & n6719 ;
  assign n6721 = ~\u0_u0_me_ps_reg[6]/P0001  & ~n6713 ;
  assign n6722 = \u0_u0_me_ps_reg[4]/P0001  & \u0_u0_me_ps_reg[6]/P0001  ;
  assign n6723 = \u0_u0_me_ps_reg[5]/P0001  & n6722 ;
  assign n6724 = n6711 & n6723 ;
  assign n6725 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & ~n6724 ;
  assign n6726 = ~n6721 & n6725 ;
  assign n6727 = n6695 & n6726 ;
  assign n6728 = ~n6182 & n6727 ;
  assign n6729 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & \u0_u0_me_ps_reg[7]/P0001  ;
  assign n6730 = ~n6724 & n6729 ;
  assign n6731 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & ~\u0_u0_me_ps_reg[7]/P0001  ;
  assign n6732 = n6724 & n6731 ;
  assign n6733 = ~n6730 & ~n6732 ;
  assign n6734 = n6695 & ~n6733 ;
  assign n6735 = ~n6182 & n6734 ;
  assign n6736 = ~\u4_u3_dma_out_cnt_reg[4]/P0001  & ~\u4_u3_dma_out_cnt_reg[6]/P0001  ;
  assign n6737 = ~\u4_u3_dma_out_cnt_reg[5]/P0001  & n6736 ;
  assign n6738 = ~\u4_u3_dma_in_cnt_reg[0]/P0001  & ~\u4_u3_dma_out_cnt_reg[1]/P0001  ;
  assign n6739 = ~\u4_u3_dma_out_cnt_reg[2]/P0001  & ~\u4_u3_dma_out_cnt_reg[3]/P0001  ;
  assign n6740 = n6738 & n6739 ;
  assign n6741 = n6737 & n6740 ;
  assign n6742 = ~\u4_u3_dma_out_cnt_reg[7]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n6743 = ~\u4_u3_dma_out_cnt_reg[8]/P0001  & n6742 ;
  assign n6744 = n6741 & n6743 ;
  assign n6745 = \u4_u3_csr1_reg[0]/P0001  & n6744 ;
  assign n6746 = ~\u4_u3_dma_out_cnt_reg[7]/P0001  & n6741 ;
  assign n6747 = \u4_u3_dma_out_cnt_reg[8]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n6748 = \u4_u3_csr1_reg[0]/P0001  & n6747 ;
  assign n6749 = ~n6746 & n6748 ;
  assign n6750 = ~n6745 & ~n6749 ;
  assign n6751 = ~\u4_u3_dma_out_cnt_reg[8]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n6752 = n6281 & n6751 ;
  assign n6753 = ~\u4_u3_dma_out_cnt_reg[8]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n6754 = n6579 & ~n6753 ;
  assign n6755 = ~n6752 & n6754 ;
  assign n6756 = n6750 & ~n6755 ;
  assign n6757 = \u4_u3_csr0_reg[9]/P0001  & \u4_u3_dma_out_cnt_reg[7]/P0001  ;
  assign n6758 = \u4_u3_csr0_reg[8]/P0001  & \u4_u3_dma_out_cnt_reg[6]/P0001  ;
  assign n6759 = ~n6757 & ~n6758 ;
  assign n6760 = ~\u4_u3_csr0_reg[8]/P0001  & ~\u4_u3_dma_out_cnt_reg[6]/P0001  ;
  assign n6761 = \u4_u3_csr0_reg[7]/P0001  & \u4_u3_dma_out_cnt_reg[5]/P0001  ;
  assign n6762 = ~n6760 & n6761 ;
  assign n6763 = \u4_u3_csr0_reg[6]/P0001  & \u4_u3_dma_out_cnt_reg[4]/P0001  ;
  assign n6764 = \u4_u3_csr0_reg[5]/P0001  & \u4_u3_dma_out_cnt_reg[3]/P0001  ;
  assign n6765 = ~n6763 & ~n6764 ;
  assign n6766 = ~\u4_u3_csr0_reg[5]/P0001  & ~\u4_u3_dma_out_cnt_reg[3]/P0001  ;
  assign n6767 = n6765 & n6766 ;
  assign n6768 = \u4_u3_csr0_reg[3]/NET0131  & \u4_u3_dma_out_cnt_reg[1]/P0001  ;
  assign n6769 = \u4_u3_csr0_reg[2]/P0001  & \u4_u3_dma_in_cnt_reg[0]/P0001  ;
  assign n6770 = ~n6768 & ~n6769 ;
  assign n6771 = ~\u4_u3_csr0_reg[4]/P0001  & ~\u4_u3_dma_out_cnt_reg[2]/P0001  ;
  assign n6772 = ~\u4_u3_csr0_reg[3]/NET0131  & ~\u4_u3_dma_out_cnt_reg[1]/P0001  ;
  assign n6773 = ~n6771 & ~n6772 ;
  assign n6774 = ~n6770 & n6773 ;
  assign n6775 = \u4_u3_csr0_reg[4]/P0001  & \u4_u3_dma_out_cnt_reg[2]/P0001  ;
  assign n6776 = n6765 & ~n6775 ;
  assign n6777 = ~n6774 & n6776 ;
  assign n6778 = ~n6767 & ~n6777 ;
  assign n6779 = ~\u4_u3_csr0_reg[7]/P0001  & ~\u4_u3_dma_out_cnt_reg[5]/P0001  ;
  assign n6780 = ~\u4_u3_csr0_reg[6]/P0001  & ~\u4_u3_dma_out_cnt_reg[4]/P0001  ;
  assign n6781 = ~n6779 & ~n6780 ;
  assign n6782 = ~n6760 & n6781 ;
  assign n6783 = n6778 & n6782 ;
  assign n6784 = ~n6762 & ~n6783 ;
  assign n6785 = n6759 & n6784 ;
  assign n6786 = \u4_u3_csr0_reg[10]/P0001  & \u4_u3_dma_out_cnt_reg[8]/P0001  ;
  assign n6787 = ~\u4_u3_csr0_reg[10]/P0001  & ~\u4_u3_dma_out_cnt_reg[8]/P0001  ;
  assign n6788 = ~n6786 & ~n6787 ;
  assign n6789 = ~\u4_u3_csr0_reg[9]/P0001  & ~\u4_u3_dma_out_cnt_reg[7]/P0001  ;
  assign n6790 = ~n6788 & ~n6789 ;
  assign n6791 = ~n6785 & n6790 ;
  assign n6792 = n6598 & ~n6791 ;
  assign n6793 = n6788 & n6789 ;
  assign n6794 = n6759 & n6788 ;
  assign n6795 = n6784 & n6794 ;
  assign n6796 = ~n6793 & ~n6795 ;
  assign n6797 = n6750 & n6796 ;
  assign n6798 = n6792 & n6797 ;
  assign n6799 = ~n6756 & ~n6798 ;
  assign n6800 = ~\u4_u0_dma_out_cnt_reg[4]/P0001  & ~\u4_u0_dma_out_cnt_reg[6]/P0001  ;
  assign n6801 = ~\u4_u0_dma_out_cnt_reg[5]/P0001  & n6800 ;
  assign n6802 = ~\u4_u0_dma_in_cnt_reg[0]/P0001  & ~\u4_u0_dma_out_cnt_reg[1]/P0001  ;
  assign n6803 = ~\u4_u0_dma_out_cnt_reg[2]/P0001  & ~\u4_u0_dma_out_cnt_reg[3]/P0001  ;
  assign n6804 = n6802 & n6803 ;
  assign n6805 = n6801 & n6804 ;
  assign n6806 = ~\u4_u0_dma_out_cnt_reg[7]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n6807 = ~\u4_u0_dma_out_cnt_reg[8]/P0001  & n6806 ;
  assign n6808 = n6805 & n6807 ;
  assign n6809 = \u4_u0_csr1_reg[0]/P0001  & n6808 ;
  assign n6810 = ~\u4_u0_dma_out_cnt_reg[7]/P0001  & n6805 ;
  assign n6811 = \u4_u0_dma_out_cnt_reg[8]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n6812 = \u4_u0_csr1_reg[0]/P0001  & n6811 ;
  assign n6813 = ~n6810 & n6812 ;
  assign n6814 = ~n6809 & ~n6813 ;
  assign n6815 = ~\u4_u0_dma_out_cnt_reg[8]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n6816 = n6281 & n6815 ;
  assign n6817 = ~\u4_u0_dma_out_cnt_reg[8]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n6818 = n6613 & ~n6817 ;
  assign n6819 = ~n6816 & n6818 ;
  assign n6820 = n6814 & ~n6819 ;
  assign n6821 = \u4_u0_csr0_reg[10]/P0001  & \u4_u0_dma_out_cnt_reg[8]/P0001  ;
  assign n6822 = ~\u4_u0_csr0_reg[10]/P0001  & ~\u4_u0_dma_out_cnt_reg[8]/P0001  ;
  assign n6823 = ~n6821 & ~n6822 ;
  assign n6824 = ~\u4_u0_csr0_reg[9]/P0001  & ~\u4_u0_dma_out_cnt_reg[7]/P0001  ;
  assign n6825 = n6823 & n6824 ;
  assign n6826 = ~\u4_u0_csr0_reg[8]/P0001  & ~\u4_u0_dma_out_cnt_reg[6]/P0001  ;
  assign n6827 = \u4_u0_csr0_reg[7]/P0001  & \u4_u0_dma_out_cnt_reg[5]/P0001  ;
  assign n6828 = ~n6826 & n6827 ;
  assign n6829 = \u4_u0_csr0_reg[6]/P0001  & \u4_u0_dma_out_cnt_reg[4]/P0001  ;
  assign n6830 = \u4_u0_csr0_reg[5]/P0001  & \u4_u0_dma_out_cnt_reg[3]/P0001  ;
  assign n6831 = ~n6829 & ~n6830 ;
  assign n6832 = ~\u4_u0_csr0_reg[5]/P0001  & ~\u4_u0_dma_out_cnt_reg[3]/P0001  ;
  assign n6833 = n6831 & n6832 ;
  assign n6834 = \u4_u0_csr0_reg[3]/NET0131  & \u4_u0_dma_out_cnt_reg[1]/P0001  ;
  assign n6835 = \u4_u0_csr0_reg[2]/P0001  & \u4_u0_dma_in_cnt_reg[0]/P0001  ;
  assign n6836 = ~n6834 & ~n6835 ;
  assign n6837 = ~\u4_u0_csr0_reg[4]/P0001  & ~\u4_u0_dma_out_cnt_reg[2]/P0001  ;
  assign n6838 = ~\u4_u0_csr0_reg[3]/NET0131  & ~\u4_u0_dma_out_cnt_reg[1]/P0001  ;
  assign n6839 = ~n6837 & ~n6838 ;
  assign n6840 = ~n6836 & n6839 ;
  assign n6841 = \u4_u0_csr0_reg[4]/P0001  & \u4_u0_dma_out_cnt_reg[2]/P0001  ;
  assign n6842 = n6831 & ~n6841 ;
  assign n6843 = ~n6840 & n6842 ;
  assign n6844 = ~n6833 & ~n6843 ;
  assign n6845 = ~\u4_u0_csr0_reg[7]/P0001  & ~\u4_u0_dma_out_cnt_reg[5]/P0001  ;
  assign n6846 = ~\u4_u0_csr0_reg[6]/P0001  & ~\u4_u0_dma_out_cnt_reg[4]/P0001  ;
  assign n6847 = ~n6845 & ~n6846 ;
  assign n6848 = ~n6826 & n6847 ;
  assign n6849 = n6844 & n6848 ;
  assign n6850 = ~n6828 & ~n6849 ;
  assign n6851 = \u4_u0_csr0_reg[9]/P0001  & \u4_u0_dma_out_cnt_reg[7]/P0001  ;
  assign n6852 = \u4_u0_csr0_reg[8]/P0001  & \u4_u0_dma_out_cnt_reg[6]/P0001  ;
  assign n6853 = ~n6851 & ~n6852 ;
  assign n6854 = n6823 & n6853 ;
  assign n6855 = n6850 & n6854 ;
  assign n6856 = ~n6825 & ~n6855 ;
  assign n6857 = n6850 & n6853 ;
  assign n6858 = ~n6823 & ~n6824 ;
  assign n6859 = ~n6857 & n6858 ;
  assign n6860 = n6856 & ~n6859 ;
  assign n6861 = n6632 & n6814 ;
  assign n6862 = n6860 & n6861 ;
  assign n6863 = ~n6820 & ~n6862 ;
  assign n6864 = ~\u4_u1_dma_out_cnt_reg[4]/P0001  & ~\u4_u1_dma_out_cnt_reg[6]/P0001  ;
  assign n6865 = ~\u4_u1_dma_out_cnt_reg[5]/P0001  & n6864 ;
  assign n6866 = ~\u4_u1_dma_in_cnt_reg[0]/P0001  & ~\u4_u1_dma_out_cnt_reg[1]/P0001  ;
  assign n6867 = ~\u4_u1_dma_out_cnt_reg[2]/P0001  & ~\u4_u1_dma_out_cnt_reg[3]/P0001  ;
  assign n6868 = n6866 & n6867 ;
  assign n6869 = n6865 & n6868 ;
  assign n6870 = ~\u4_u1_dma_out_cnt_reg[7]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n6871 = ~\u4_u1_dma_out_cnt_reg[8]/P0001  & n6870 ;
  assign n6872 = n6869 & n6871 ;
  assign n6873 = \u4_u1_csr1_reg[0]/P0001  & n6872 ;
  assign n6874 = ~\u4_u1_dma_out_cnt_reg[7]/P0001  & n6869 ;
  assign n6875 = \u4_u1_dma_out_cnt_reg[8]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n6876 = \u4_u1_csr1_reg[0]/P0001  & n6875 ;
  assign n6877 = ~n6874 & n6876 ;
  assign n6878 = ~n6873 & ~n6877 ;
  assign n6879 = ~\u4_u1_dma_out_cnt_reg[8]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n6880 = n6281 & n6879 ;
  assign n6881 = ~\u4_u1_dma_out_cnt_reg[8]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n6882 = n6642 & ~n6881 ;
  assign n6883 = ~n6880 & n6882 ;
  assign n6884 = n6878 & ~n6883 ;
  assign n6885 = \u4_u1_csr0_reg[10]/P0001  & \u4_u1_dma_out_cnt_reg[8]/P0001  ;
  assign n6886 = ~\u4_u1_csr0_reg[10]/P0001  & ~\u4_u1_dma_out_cnt_reg[8]/P0001  ;
  assign n6887 = ~n6885 & ~n6886 ;
  assign n6888 = ~\u4_u1_csr0_reg[9]/P0001  & ~\u4_u1_dma_out_cnt_reg[7]/P0001  ;
  assign n6889 = n6887 & n6888 ;
  assign n6890 = ~\u4_u1_csr0_reg[8]/P0001  & ~\u4_u1_dma_out_cnt_reg[6]/P0001  ;
  assign n6891 = \u4_u1_csr0_reg[7]/P0001  & \u4_u1_dma_out_cnt_reg[5]/P0001  ;
  assign n6892 = ~n6890 & n6891 ;
  assign n6893 = \u4_u1_csr0_reg[6]/P0001  & \u4_u1_dma_out_cnt_reg[4]/P0001  ;
  assign n6894 = \u4_u1_csr0_reg[5]/P0001  & \u4_u1_dma_out_cnt_reg[3]/P0001  ;
  assign n6895 = ~n6893 & ~n6894 ;
  assign n6896 = ~\u4_u1_csr0_reg[5]/P0001  & ~\u4_u1_dma_out_cnt_reg[3]/P0001  ;
  assign n6897 = n6895 & n6896 ;
  assign n6898 = \u4_u1_csr0_reg[3]/NET0131  & \u4_u1_dma_out_cnt_reg[1]/P0001  ;
  assign n6899 = \u4_u1_csr0_reg[2]/P0001  & \u4_u1_dma_in_cnt_reg[0]/P0001  ;
  assign n6900 = ~n6898 & ~n6899 ;
  assign n6901 = ~\u4_u1_csr0_reg[4]/P0001  & ~\u4_u1_dma_out_cnt_reg[2]/P0001  ;
  assign n6902 = ~\u4_u1_csr0_reg[3]/NET0131  & ~\u4_u1_dma_out_cnt_reg[1]/P0001  ;
  assign n6903 = ~n6901 & ~n6902 ;
  assign n6904 = ~n6900 & n6903 ;
  assign n6905 = \u4_u1_csr0_reg[4]/P0001  & \u4_u1_dma_out_cnt_reg[2]/P0001  ;
  assign n6906 = n6895 & ~n6905 ;
  assign n6907 = ~n6904 & n6906 ;
  assign n6908 = ~n6897 & ~n6907 ;
  assign n6909 = ~\u4_u1_csr0_reg[7]/P0001  & ~\u4_u1_dma_out_cnt_reg[5]/P0001  ;
  assign n6910 = ~\u4_u1_csr0_reg[6]/P0001  & ~\u4_u1_dma_out_cnt_reg[4]/P0001  ;
  assign n6911 = ~n6909 & ~n6910 ;
  assign n6912 = ~n6890 & n6911 ;
  assign n6913 = n6908 & n6912 ;
  assign n6914 = ~n6892 & ~n6913 ;
  assign n6915 = \u4_u1_csr0_reg[9]/P0001  & \u4_u1_dma_out_cnt_reg[7]/P0001  ;
  assign n6916 = \u4_u1_csr0_reg[8]/P0001  & \u4_u1_dma_out_cnt_reg[6]/P0001  ;
  assign n6917 = ~n6915 & ~n6916 ;
  assign n6918 = n6887 & n6917 ;
  assign n6919 = n6914 & n6918 ;
  assign n6920 = ~n6889 & ~n6919 ;
  assign n6921 = n6914 & n6917 ;
  assign n6922 = ~n6887 & ~n6888 ;
  assign n6923 = ~n6921 & n6922 ;
  assign n6924 = n6920 & ~n6923 ;
  assign n6925 = n6369 & n6878 ;
  assign n6926 = n6924 & n6925 ;
  assign n6927 = ~n6884 & ~n6926 ;
  assign n6928 = ~\u4_u2_dma_out_cnt_reg[4]/P0001  & ~\u4_u2_dma_out_cnt_reg[6]/P0001  ;
  assign n6929 = ~\u4_u2_dma_out_cnt_reg[5]/P0001  & n6928 ;
  assign n6930 = ~\u4_u2_dma_in_cnt_reg[0]/P0001  & ~\u4_u2_dma_out_cnt_reg[1]/P0001  ;
  assign n6931 = ~\u4_u2_dma_out_cnt_reg[2]/P0001  & ~\u4_u2_dma_out_cnt_reg[3]/P0001  ;
  assign n6932 = n6930 & n6931 ;
  assign n6933 = n6929 & n6932 ;
  assign n6934 = ~\u4_u2_dma_out_cnt_reg[7]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n6935 = ~\u4_u2_dma_out_cnt_reg[8]/P0001  & n6934 ;
  assign n6936 = n6933 & n6935 ;
  assign n6937 = \u4_u2_csr1_reg[0]/P0001  & n6936 ;
  assign n6938 = ~\u4_u2_dma_out_cnt_reg[7]/P0001  & n6933 ;
  assign n6939 = \u4_u2_dma_out_cnt_reg[8]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n6940 = \u4_u2_csr1_reg[0]/P0001  & n6939 ;
  assign n6941 = ~n6938 & n6940 ;
  assign n6942 = ~n6937 & ~n6941 ;
  assign n6943 = ~\u4_u2_dma_out_cnt_reg[8]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n6944 = n6281 & n6943 ;
  assign n6945 = ~\u4_u2_dma_out_cnt_reg[8]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n6946 = \u4_u2_csr1_reg[0]/P0001  & ~\u4_u2_r5_reg/NET0131  ;
  assign n6947 = ~n6945 & n6946 ;
  assign n6948 = ~n6944 & n6947 ;
  assign n6949 = n6942 & ~n6948 ;
  assign n6950 = \u4_u2_csr0_reg[9]/P0001  & \u4_u2_dma_out_cnt_reg[7]/P0001  ;
  assign n6951 = \u4_u2_csr0_reg[8]/P0001  & \u4_u2_dma_out_cnt_reg[6]/P0001  ;
  assign n6952 = ~n6950 & ~n6951 ;
  assign n6953 = ~\u4_u2_csr0_reg[8]/P0001  & ~\u4_u2_dma_out_cnt_reg[6]/P0001  ;
  assign n6954 = \u4_u2_csr0_reg[7]/P0001  & \u4_u2_dma_out_cnt_reg[5]/P0001  ;
  assign n6955 = ~n6953 & n6954 ;
  assign n6956 = \u4_u2_csr0_reg[6]/P0001  & \u4_u2_dma_out_cnt_reg[4]/P0001  ;
  assign n6957 = \u4_u2_csr0_reg[5]/P0001  & \u4_u2_dma_out_cnt_reg[3]/P0001  ;
  assign n6958 = ~n6956 & ~n6957 ;
  assign n6959 = ~\u4_u2_csr0_reg[5]/P0001  & ~\u4_u2_dma_out_cnt_reg[3]/P0001  ;
  assign n6960 = n6958 & n6959 ;
  assign n6961 = \u4_u2_csr0_reg[3]/NET0131  & \u4_u2_dma_out_cnt_reg[1]/P0001  ;
  assign n6962 = \u4_u2_csr0_reg[2]/P0001  & \u4_u2_dma_in_cnt_reg[0]/P0001  ;
  assign n6963 = ~n6961 & ~n6962 ;
  assign n6964 = ~\u4_u2_csr0_reg[4]/P0001  & ~\u4_u2_dma_out_cnt_reg[2]/P0001  ;
  assign n6965 = ~\u4_u2_csr0_reg[3]/NET0131  & ~\u4_u2_dma_out_cnt_reg[1]/P0001  ;
  assign n6966 = ~n6964 & ~n6965 ;
  assign n6967 = ~n6963 & n6966 ;
  assign n6968 = \u4_u2_csr0_reg[4]/P0001  & \u4_u2_dma_out_cnt_reg[2]/P0001  ;
  assign n6969 = n6958 & ~n6968 ;
  assign n6970 = ~n6967 & n6969 ;
  assign n6971 = ~n6960 & ~n6970 ;
  assign n6972 = ~\u4_u2_csr0_reg[7]/P0001  & ~\u4_u2_dma_out_cnt_reg[5]/P0001  ;
  assign n6973 = ~\u4_u2_csr0_reg[6]/P0001  & ~\u4_u2_dma_out_cnt_reg[4]/P0001  ;
  assign n6974 = ~n6972 & ~n6973 ;
  assign n6975 = ~n6953 & n6974 ;
  assign n6976 = n6971 & n6975 ;
  assign n6977 = ~n6955 & ~n6976 ;
  assign n6978 = n6952 & n6977 ;
  assign n6979 = \u4_u2_csr0_reg[10]/P0001  & \u4_u2_dma_out_cnt_reg[8]/P0001  ;
  assign n6980 = ~\u4_u2_csr0_reg[10]/P0001  & ~\u4_u2_dma_out_cnt_reg[8]/P0001  ;
  assign n6981 = ~n6979 & ~n6980 ;
  assign n6982 = ~\u4_u2_csr0_reg[9]/P0001  & ~\u4_u2_dma_out_cnt_reg[7]/P0001  ;
  assign n6983 = ~n6981 & ~n6982 ;
  assign n6984 = ~n6978 & n6983 ;
  assign n6985 = n6667 & ~n6984 ;
  assign n6986 = n6981 & n6982 ;
  assign n6987 = n6952 & n6981 ;
  assign n6988 = n6977 & n6987 ;
  assign n6989 = ~n6986 & ~n6988 ;
  assign n6990 = n6942 & n6989 ;
  assign n6991 = n6985 & n6990 ;
  assign n6992 = ~n6949 & ~n6991 ;
  assign n6993 = ~\u1_hms_clk_reg/P0001  & ~\u1_hms_cnt_reg[0]/P0001  ;
  assign n6994 = n6477 & n6993 ;
  assign n6995 = ~\u0_u0_me_cnt_reg[6]/P0001  & ~\u0_u0_me_cnt_reg[7]/P0001  ;
  assign n6996 = n6205 & n6995 ;
  assign n6997 = \u0_u0_me_cnt_reg[0]/P0001  & \u0_u0_me_cnt_reg[1]/P0001  ;
  assign n6998 = ~\u0_u0_me_cnt_reg[2]/P0001  & ~\u0_u0_me_cnt_reg[3]/P0001  ;
  assign n6999 = ~n6997 & n6998 ;
  assign n7000 = n6996 & n6999 ;
  assign n7001 = n6695 & ~n7000 ;
  assign n7002 = ~n6182 & n7001 ;
  assign n7003 = ~\u0_u0_me_cnt_reg[2]/P0001  & ~n6997 ;
  assign n7004 = \u0_u0_me_cnt_reg[3]/P0001  & ~n7003 ;
  assign n7005 = n6996 & ~n7004 ;
  assign n7006 = n6695 & ~n7005 ;
  assign n7007 = ~n6182 & n7006 ;
  assign n7008 = \u5_wb_ack_s1_reg/P0001  & ~\u5_wb_ack_s2_reg/P0001  ;
  assign n7009 = ~wb_ack_o_pad & n7008 ;
  assign n7010 = \u1_u2_rx_data_valid_r_reg/NET0131  & \u1_u2_sizu_c_reg[2]/P0001  ;
  assign n7011 = n6110 & n7010 ;
  assign n7012 = \u1_u2_sizu_c_reg[3]/P0001  & \u1_u2_sizu_c_reg[5]/P0001  ;
  assign n7013 = \u1_u2_sizu_c_reg[4]/P0001  & n7012 ;
  assign n7014 = n7011 & n7013 ;
  assign n7015 = \u1_u2_sizu_c_reg[6]/P0001  & \u1_u2_sizu_c_reg[7]/P0001  ;
  assign n7016 = n7014 & n7015 ;
  assign n7017 = ~\u1_u2_sizu_c_reg[8]/NET0131  & ~n7016 ;
  assign n7018 = rst_i_pad & ~\u1_u2_rx_dma_en_r_reg/P0001  ;
  assign n7019 = \u1_u2_sizu_c_reg[4]/P0001  & \u1_u2_sizu_c_reg[8]/NET0131  ;
  assign n7020 = n7012 & n7019 ;
  assign n7021 = n7011 & n7020 ;
  assign n7022 = n7015 & n7021 ;
  assign n7023 = n7018 & ~n7022 ;
  assign n7024 = ~n7017 & n7023 ;
  assign n7025 = \u0_u0_me_ps2_reg[0]/P0001  & \u0_u0_me_ps_2_5_us_reg/P0001  ;
  assign n7026 = ~\u0_u0_me_ps2_reg[0]/P0001  & ~\u0_u0_me_ps_2_5_us_reg/P0001  ;
  assign n7027 = ~n7025 & ~n7026 ;
  assign n7028 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & n7027 ;
  assign n7029 = n6695 & n7028 ;
  assign n7030 = ~n6182 & n7029 ;
  assign n7031 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & \u0_u0_me_ps2_reg[1]/P0001  ;
  assign n7032 = ~n7025 & n7031 ;
  assign n7033 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & ~\u0_u0_me_ps2_reg[1]/P0001  ;
  assign n7034 = n7025 & n7033 ;
  assign n7035 = ~n7032 & ~n7034 ;
  assign n7036 = n6695 & ~n7035 ;
  assign n7037 = ~n6182 & n7036 ;
  assign n7038 = \u0_u0_me_ps2_reg[1]/P0001  & \u0_u0_me_ps2_reg[2]/P0001  ;
  assign n7039 = n7025 & n7038 ;
  assign n7040 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & \u0_u0_me_ps2_reg[2]/P0001  ;
  assign n7041 = n7025 & n7031 ;
  assign n7042 = ~n7040 & ~n7041 ;
  assign n7043 = ~n7039 & ~n7042 ;
  assign n7044 = n6695 & n7043 ;
  assign n7045 = ~n6182 & n7044 ;
  assign n7046 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & \u0_u0_me_ps2_reg[3]/P0001  ;
  assign n7047 = ~n7039 & n7046 ;
  assign n7048 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & ~\u0_u0_me_ps2_reg[3]/P0001  ;
  assign n7049 = n7039 & n7048 ;
  assign n7050 = ~n7047 & ~n7049 ;
  assign n7051 = n6695 & ~n7050 ;
  assign n7052 = ~n6182 & n7051 ;
  assign n7053 = \u0_u0_me_ps2_reg[3]/P0001  & \u0_u0_me_ps2_reg[4]/P0001  ;
  assign n7054 = n7039 & n7053 ;
  assign n7055 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & \u0_u0_me_ps2_reg[4]/P0001  ;
  assign n7056 = n7039 & n7046 ;
  assign n7057 = ~n7055 & ~n7056 ;
  assign n7058 = ~n7054 & ~n7057 ;
  assign n7059 = n6695 & n7058 ;
  assign n7060 = ~n6182 & n7059 ;
  assign n7061 = \u0_u0_me_ps2_reg[3]/P0001  & \u0_u0_me_ps2_reg[5]/P0001  ;
  assign n7062 = \u0_u0_me_ps2_reg[4]/P0001  & n7061 ;
  assign n7063 = n7039 & n7062 ;
  assign n7064 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & \u0_u0_me_ps2_reg[5]/P0001  ;
  assign n7065 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & n7053 ;
  assign n7066 = n7039 & n7065 ;
  assign n7067 = ~n7064 & ~n7066 ;
  assign n7068 = ~n7063 & ~n7067 ;
  assign n7069 = n6695 & n7068 ;
  assign n7070 = ~n6182 & n7069 ;
  assign n7071 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & \u0_u0_me_ps2_reg[6]/P0001  ;
  assign n7072 = ~n7063 & n7071 ;
  assign n7073 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & ~\u0_u0_me_ps2_reg[6]/P0001  ;
  assign n7074 = n7063 & n7073 ;
  assign n7075 = ~n7072 & ~n7074 ;
  assign n7076 = n6695 & ~n7075 ;
  assign n7077 = ~n6182 & n7076 ;
  assign n7078 = \u0_u0_me_ps2_reg[6]/P0001  & \u0_u0_me_ps2_reg[7]/P0001  ;
  assign n7079 = n7063 & n7078 ;
  assign n7080 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & \u0_u0_me_ps2_reg[7]/P0001  ;
  assign n7081 = n7063 & n7071 ;
  assign n7082 = ~n7080 & ~n7081 ;
  assign n7083 = ~n7079 & ~n7082 ;
  assign n7084 = n6695 & n7083 ;
  assign n7085 = ~n6182 & n7084 ;
  assign n7086 = ~\u0_u0_me_ps_reg[0]/P0001  & ~\u0_u0_me_ps_reg[1]/P0001  ;
  assign n7087 = ~n6709 & ~n7086 ;
  assign n7088 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & n7087 ;
  assign n7089 = n6695 & n7088 ;
  assign n7090 = ~n6182 & n7089 ;
  assign n7091 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & \u0_u0_me_ps_reg[2]/P0001  ;
  assign n7092 = ~n6709 & n7091 ;
  assign n7093 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & ~\u0_u0_me_ps_reg[2]/P0001  ;
  assign n7094 = n6709 & n7093 ;
  assign n7095 = ~n7092 & ~n7094 ;
  assign n7096 = n6695 & ~n7095 ;
  assign n7097 = ~n6182 & n7096 ;
  assign n7098 = \u0_u0_me_ps_reg[2]/P0001  & n6709 ;
  assign n7099 = ~\u0_u0_me_ps_reg[3]/P0001  & ~n7098 ;
  assign n7100 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & ~n6711 ;
  assign n7101 = ~n7099 & n7100 ;
  assign n7102 = n6695 & n7101 ;
  assign n7103 = ~n6182 & n7102 ;
  assign n7104 = ~n6711 & n6715 ;
  assign n7105 = ~\u0_u0_me_ps_2_5_us_reg/P0001  & ~\u0_u0_me_ps_reg[4]/P0001  ;
  assign n7106 = n6711 & n7105 ;
  assign n7107 = ~n7104 & ~n7106 ;
  assign n7108 = n6695 & ~n7107 ;
  assign n7109 = ~n6182 & n7108 ;
  assign n7110 = n6212 & n6218 ;
  assign n7111 = n6217 & n7110 ;
  assign n7112 = \u1_sof_time_reg[6]/P0001  & n7111 ;
  assign n7113 = ~\u1_sof_time_reg[7]/P0001  & ~n7112 ;
  assign n7114 = \u1_sof_time_reg[6]/P0001  & \u1_sof_time_reg[7]/P0001  ;
  assign n7115 = n7111 & n7114 ;
  assign n7116 = ~\u1_clr_sof_time_reg/P0001  & ~n7115 ;
  assign n7117 = ~n7113 & n7116 ;
  assign n7118 = \u1_u3_pid_seq_err_reg/P0001  & \u1_u3_state_reg[4]/P0001  ;
  assign n7119 = n4907 & n5555 ;
  assign n7120 = n7118 & n7119 ;
  assign n7121 = n4936 & n7120 ;
  assign n7122 = n4935 & n7121 ;
  assign n7123 = ~\u1_frame_no_r_reg[8]/P0001  & ~\u1_u0_token1_reg[0]/P0001  ;
  assign n7124 = \u1_frame_no_r_reg[8]/P0001  & \u1_u0_token1_reg[0]/P0001  ;
  assign n7125 = ~n7123 & ~n7124 ;
  assign n7126 = \u1_u0_token_valid_str1_reg/P0001  & n2379 ;
  assign n7127 = ~n5097 & n7126 ;
  assign n7128 = n5114 & n7127 ;
  assign n7129 = ~\u1_frame_no_r_reg[7]/P0001  & ~\u1_u0_token0_reg[7]/P0001  ;
  assign n7130 = \u1_frame_no_r_reg[7]/P0001  & \u1_u0_token0_reg[7]/P0001  ;
  assign n7131 = ~n7129 & ~n7130 ;
  assign n7132 = ~\u1_frame_no_r_reg[9]/P0001  & \u1_u0_token1_reg[1]/P0001  ;
  assign n7133 = \u1_frame_no_r_reg[4]/P0001  & ~\u1_u0_token0_reg[4]/P0001  ;
  assign n7134 = ~n7132 & ~n7133 ;
  assign n7135 = ~n7131 & n7134 ;
  assign n7136 = ~\u1_frame_no_r_reg[6]/P0001  & \u1_u0_token0_reg[6]/P0001  ;
  assign n7137 = \u1_frame_no_r_reg[10]/P0001  & ~\u1_u0_token1_reg[2]/P0001  ;
  assign n7138 = ~n7136 & ~n7137 ;
  assign n7139 = ~\u1_frame_no_r_reg[10]/P0001  & \u1_u0_token1_reg[2]/P0001  ;
  assign n7140 = ~\u1_frame_no_r_reg[1]/P0001  & \u1_u0_token0_reg[1]/P0001  ;
  assign n7141 = ~n7139 & ~n7140 ;
  assign n7142 = n7138 & n7141 ;
  assign n7143 = \u1_frame_no_r_reg[2]/P0001  & ~\u1_u0_token0_reg[2]/NET0131  ;
  assign n7144 = \u1_frame_no_r_reg[1]/P0001  & ~\u1_u0_token0_reg[1]/P0001  ;
  assign n7145 = ~n7143 & ~n7144 ;
  assign n7146 = ~\u1_frame_no_r_reg[2]/P0001  & \u1_u0_token0_reg[2]/NET0131  ;
  assign n7147 = ~\u1_frame_no_r_reg[5]/P0001  & \u1_u0_token0_reg[5]/NET0131  ;
  assign n7148 = ~n7146 & ~n7147 ;
  assign n7149 = n7145 & n7148 ;
  assign n7150 = n7142 & n7149 ;
  assign n7151 = \u1_frame_no_r_reg[0]/P0001  & ~\u1_u0_token0_reg[0]/NET0131  ;
  assign n7152 = ~\u1_frame_no_r_reg[3]/P0001  & \u1_u0_token0_reg[3]/NET0131  ;
  assign n7153 = ~n7151 & ~n7152 ;
  assign n7154 = ~\u1_frame_no_r_reg[0]/P0001  & \u1_u0_token0_reg[0]/NET0131  ;
  assign n7155 = \u1_frame_no_r_reg[9]/P0001  & ~\u1_u0_token1_reg[1]/P0001  ;
  assign n7156 = ~n7154 & ~n7155 ;
  assign n7157 = n7153 & n7156 ;
  assign n7158 = \u1_frame_no_r_reg[6]/P0001  & ~\u1_u0_token0_reg[6]/P0001  ;
  assign n7159 = \u1_frame_no_r_reg[5]/P0001  & ~\u1_u0_token0_reg[5]/NET0131  ;
  assign n7160 = ~n7158 & ~n7159 ;
  assign n7161 = \u1_frame_no_r_reg[3]/P0001  & ~\u1_u0_token0_reg[3]/NET0131  ;
  assign n7162 = ~\u1_frame_no_r_reg[4]/P0001  & \u1_u0_token0_reg[4]/P0001  ;
  assign n7163 = ~n7161 & ~n7162 ;
  assign n7164 = n7160 & n7163 ;
  assign n7165 = n7157 & n7164 ;
  assign n7166 = n7150 & n7165 ;
  assign n7167 = n7135 & n7166 ;
  assign n7168 = n5079 & n7167 ;
  assign n7169 = n5063 & n7168 ;
  assign n7170 = n7128 & n7169 ;
  assign n7171 = ~n7125 & n7170 ;
  assign n7172 = \sram_data_i[0]_pad  & \wb_addr_i[17]_pad  ;
  assign n7173 = \u4_dout_reg[0]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n7174 = ~n7172 & ~n7173 ;
  assign n7175 = \sram_data_i[1]_pad  & \wb_addr_i[17]_pad  ;
  assign n7176 = \u4_dout_reg[1]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n7177 = ~n7175 & ~n7176 ;
  assign n7178 = \sram_data_i[2]_pad  & \wb_addr_i[17]_pad  ;
  assign n7179 = \u4_dout_reg[2]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n7180 = ~n7178 & ~n7179 ;
  assign n7181 = \sram_data_i[3]_pad  & \wb_addr_i[17]_pad  ;
  assign n7182 = \u4_dout_reg[3]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n7183 = ~n7181 & ~n7182 ;
  assign n7184 = ~n4459 & n4468 ;
  assign n7185 = ~n4454 & n7184 ;
  assign n7186 = ~n4462 & ~n4473 ;
  assign n7187 = ~n7185 & ~n7186 ;
  assign n7188 = n4468 & n7186 ;
  assign n7189 = ~n4459 & n7188 ;
  assign n7190 = ~n4454 & n7189 ;
  assign n7191 = ~n7187 & ~n7190 ;
  assign n7192 = n4542 & n4546 ;
  assign n7193 = ~n4460 & ~n4461 ;
  assign n7194 = ~n7192 & ~n7193 ;
  assign n7195 = n4546 & n7193 ;
  assign n7196 = n4542 & n7195 ;
  assign n7197 = ~n7194 & ~n7196 ;
  assign n7198 = ~\u0_rx_err_reg/P0001  & n4958 ;
  assign n7199 = \u1_u0_state_reg[1]/P0001  & ~\u1_u0_state_reg[3]/P0001  ;
  assign n7200 = n4909 & n7199 ;
  assign n7201 = ~n7198 & n7200 ;
  assign n7202 = \u0_rx_active_reg/P0001  & \u0_rx_valid_reg/P0001  ;
  assign n7203 = ~\u0_rx_err_reg/P0001  & n7202 ;
  assign n7204 = ~n2350 & ~n3447 ;
  assign n7205 = n7203 & ~n7204 ;
  assign n7206 = n7201 & n7205 ;
  assign n7207 = ~\u1_u0_state_reg[1]/P0001  & ~\u1_u0_state_reg[3]/P0001  ;
  assign n7208 = ~\u1_u0_state_reg[0]/P0001  & \u1_u0_state_reg[2]/P0001  ;
  assign n7209 = n7207 & n7208 ;
  assign n7210 = ~n7203 & n7209 ;
  assign n7211 = ~n4911 & ~n7210 ;
  assign n7212 = \u0_rx_active_reg/P0001  & \u1_u0_state_reg[2]/P0001  ;
  assign n7213 = ~n7211 & n7212 ;
  assign n7214 = ~n7206 & ~n7213 ;
  assign n7215 = rst_i_pad & ~n7214 ;
  assign n7216 = ~\u4_u3_r5_reg/NET0131  & ~n6287 ;
  assign n7217 = n6285 & n7216 ;
  assign n7218 = ~\u4_u3_dma_in_cnt_reg[10]/P0001  & ~n7217 ;
  assign n7219 = ~\u4_u3_dma_in_cnt_reg[10]/P0001  & n6270 ;
  assign n7220 = ~n6265 & n7219 ;
  assign n7221 = ~n7218 & ~n7220 ;
  assign n7222 = ~\u4_u3_dma_in_cnt_reg[10]/P0001  & ~\u4_u3_dma_in_cnt_reg[9]/P0001  ;
  assign n7223 = ~\u4_u3_r5_reg/NET0131  & ~n7222 ;
  assign n7224 = ~\u4_u3_r5_reg/NET0131  & ~n7223 ;
  assign n7225 = \u4_u3_dma_in_cnt_reg[7]/P0001  & \u4_u3_dma_in_cnt_reg[9]/P0001  ;
  assign n7226 = \u4_u3_dma_in_cnt_reg[8]/P0001  & n7225 ;
  assign n7227 = ~n7223 & n7226 ;
  assign n7228 = n6277 & n7227 ;
  assign n7229 = ~n7224 & ~n7228 ;
  assign n7230 = \u4_u3_dma_in_cnt_reg[11]/P0001  & ~n7229 ;
  assign n7231 = n7221 & n7230 ;
  assign n7232 = ~\u4_u3_dma_in_cnt_reg[11]/P0001  & ~n7221 ;
  assign n7233 = ~\u4_u3_dma_in_cnt_reg[11]/P0001  & n7229 ;
  assign n7234 = \u4_u3_csr1_reg[0]/P0001  & ~n7233 ;
  assign n7235 = ~n7232 & n7234 ;
  assign n7236 = ~n7231 & n7235 ;
  assign n7237 = ~\u4_u0_r5_reg/NET0131  & ~n6344 ;
  assign n7238 = n6342 & n7237 ;
  assign n7239 = ~\u4_u0_dma_in_cnt_reg[10]/P0001  & ~n7238 ;
  assign n7240 = ~\u4_u0_dma_in_cnt_reg[10]/P0001  & n6328 ;
  assign n7241 = ~n6323 & n7240 ;
  assign n7242 = ~n7239 & ~n7241 ;
  assign n7243 = ~\u4_u0_dma_in_cnt_reg[10]/P0001  & ~\u4_u0_dma_in_cnt_reg[9]/P0001  ;
  assign n7244 = ~\u4_u0_r5_reg/NET0131  & ~n7243 ;
  assign n7245 = ~\u4_u0_r5_reg/NET0131  & ~n7244 ;
  assign n7246 = \u4_u0_dma_in_cnt_reg[7]/P0001  & \u4_u0_dma_in_cnt_reg[9]/P0001  ;
  assign n7247 = \u4_u0_dma_in_cnt_reg[8]/P0001  & n7246 ;
  assign n7248 = ~n7244 & n7247 ;
  assign n7249 = n6335 & n7248 ;
  assign n7250 = ~n7245 & ~n7249 ;
  assign n7251 = \u4_u0_dma_in_cnt_reg[11]/P0001  & ~n7250 ;
  assign n7252 = n7242 & n7251 ;
  assign n7253 = ~\u4_u0_dma_in_cnt_reg[11]/P0001  & ~n7242 ;
  assign n7254 = ~\u4_u0_dma_in_cnt_reg[11]/P0001  & n7250 ;
  assign n7255 = \u4_u0_csr1_reg[0]/P0001  & ~n7254 ;
  assign n7256 = ~n7253 & n7255 ;
  assign n7257 = ~n7252 & n7256 ;
  assign n7258 = ~\u4_u1_r5_reg/NET0131  & ~n6370 ;
  assign n7259 = ~n6373 & n7258 ;
  assign n7260 = n6369 & n7259 ;
  assign n7261 = ~\u4_u1_dma_in_cnt_reg[10]/P0001  & ~n7260 ;
  assign n7262 = ~\u4_u1_dma_in_cnt_reg[10]/P0001  & n6406 ;
  assign n7263 = n6402 & n7262 ;
  assign n7264 = ~n7261 & ~n7263 ;
  assign n7265 = ~\u4_u1_dma_in_cnt_reg[10]/P0001  & ~\u4_u1_dma_in_cnt_reg[9]/P0001  ;
  assign n7266 = ~\u4_u1_r5_reg/NET0131  & ~n7265 ;
  assign n7267 = ~\u4_u1_r5_reg/NET0131  & ~n7266 ;
  assign n7268 = \u4_u1_dma_in_cnt_reg[7]/P0001  & \u4_u1_dma_in_cnt_reg[9]/P0001  ;
  assign n7269 = \u4_u1_dma_in_cnt_reg[8]/P0001  & n7268 ;
  assign n7270 = ~n7266 & n7269 ;
  assign n7271 = n6362 & n7270 ;
  assign n7272 = ~n7267 & ~n7271 ;
  assign n7273 = \u4_u1_dma_in_cnt_reg[11]/P0001  & ~n7272 ;
  assign n7274 = n7264 & n7273 ;
  assign n7275 = ~\u4_u1_dma_in_cnt_reg[10]/P0001  & ~\u4_u1_dma_in_cnt_reg[11]/P0001  ;
  assign n7276 = ~n7260 & n7275 ;
  assign n7277 = n6406 & n7275 ;
  assign n7278 = n6402 & n7277 ;
  assign n7279 = ~n7276 & ~n7278 ;
  assign n7280 = ~\u4_u1_dma_in_cnt_reg[11]/P0001  & n7272 ;
  assign n7281 = \u4_u1_csr1_reg[0]/P0001  & ~n7280 ;
  assign n7282 = n7279 & n7281 ;
  assign n7283 = ~n7274 & n7282 ;
  assign n7284 = ~\u4_u2_dma_in_cnt_reg[10]/P0001  & ~\u4_u2_dma_in_cnt_reg[9]/P0001  ;
  assign n7285 = ~\u4_u2_r5_reg/NET0131  & n7284 ;
  assign n7286 = n6455 & n7285 ;
  assign n7287 = \u4_u2_dma_in_cnt_reg[7]/P0001  & \u4_u2_dma_in_cnt_reg[9]/P0001  ;
  assign n7288 = \u4_u2_dma_in_cnt_reg[8]/P0001  & n7287 ;
  assign n7289 = n6463 & n7288 ;
  assign n7290 = \u4_u2_dma_in_cnt_reg[10]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n7291 = n7289 & n7290 ;
  assign n7292 = \u4_u2_csr1_reg[0]/P0001  & \u4_u2_dma_in_cnt_reg[11]/P0001  ;
  assign n7293 = ~n7291 & n7292 ;
  assign n7294 = ~n7286 & n7293 ;
  assign n7295 = \u4_u2_csr1_reg[0]/P0001  & ~\u4_u2_dma_in_cnt_reg[11]/P0001  ;
  assign n7296 = n7291 & n7295 ;
  assign n7297 = n7285 & n7295 ;
  assign n7298 = n6455 & n7297 ;
  assign n7299 = ~n7296 & ~n7298 ;
  assign n7300 = ~n7294 & n7299 ;
  assign n7301 = \u4_u3_dma_out_cnt_reg[9]/P0001  & ~n6787 ;
  assign n7302 = ~n6789 & n7301 ;
  assign n7303 = \u4_u3_dma_out_cnt_reg[9]/P0001  & n6786 ;
  assign n7304 = ~n7302 & ~n7303 ;
  assign n7305 = n6759 & ~n7303 ;
  assign n7306 = n6784 & n7305 ;
  assign n7307 = ~n7304 & ~n7306 ;
  assign n7308 = ~\u4_u3_dma_out_cnt_reg[4]/P0001  & ~\u4_u3_dma_out_cnt_reg[5]/P0001  ;
  assign n7309 = n6740 & n7308 ;
  assign n7310 = ~\u4_u3_dma_out_cnt_reg[8]/P0001  & ~\u4_u3_dma_out_cnt_reg[9]/P0001  ;
  assign n7311 = ~\u4_u3_dma_out_cnt_reg[6]/P0001  & ~\u4_u3_dma_out_cnt_reg[7]/P0001  ;
  assign n7312 = n7310 & n7311 ;
  assign n7313 = ~\u4_u3_dma_out_cnt_reg[10]/P0001  & n7312 ;
  assign n7314 = n7309 & n7313 ;
  assign n7315 = \u4_u3_r5_reg/NET0131  & ~n7314 ;
  assign n7316 = \u4_u3_dma_out_cnt_reg[10]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n7317 = ~n6282 & n7316 ;
  assign n7318 = ~n7315 & n7317 ;
  assign n7319 = n7307 & n7318 ;
  assign n7320 = ~\u4_u3_dma_out_cnt_reg[10]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n7321 = n7312 & n7320 ;
  assign n7322 = n7309 & n7321 ;
  assign n7323 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_out_cnt_reg[11]/P0001  ;
  assign n7324 = ~n7322 & n7323 ;
  assign n7325 = ~n7319 & n7324 ;
  assign n7326 = \u4_u3_csr1_reg[0]/P0001  & ~\u4_u3_dma_out_cnt_reg[11]/P0001  ;
  assign n7327 = n7322 & n7326 ;
  assign n7328 = n7318 & n7326 ;
  assign n7329 = n7307 & n7328 ;
  assign n7330 = ~n7327 & ~n7329 ;
  assign n7331 = ~n7325 & n7330 ;
  assign n7332 = ~n6787 & ~n6789 ;
  assign n7333 = ~n6786 & ~n7332 ;
  assign n7334 = n6759 & ~n6786 ;
  assign n7335 = n6784 & n7334 ;
  assign n7336 = ~n7333 & ~n7335 ;
  assign n7337 = ~\u4_u3_r5_reg/NET0131  & ~n7336 ;
  assign n7338 = ~\u4_u3_r5_reg/NET0131  & n6598 ;
  assign n7339 = ~\u4_u3_dma_out_cnt_reg[7]/P0001  & ~\u4_u3_dma_out_cnt_reg[8]/P0001  ;
  assign n7340 = \u4_u3_r5_reg/NET0131  & n7339 ;
  assign n7341 = n6741 & n7340 ;
  assign n7342 = ~n7338 & ~n7341 ;
  assign n7343 = \u4_u3_dma_out_cnt_reg[9]/P0001  & ~n7342 ;
  assign n7344 = ~n7337 & n7343 ;
  assign n7345 = ~\u4_u3_dma_out_cnt_reg[9]/P0001  & ~\u4_u3_r5_reg/NET0131  ;
  assign n7346 = ~n7336 & n7345 ;
  assign n7347 = ~\u4_u3_dma_out_cnt_reg[9]/P0001  & n7342 ;
  assign n7348 = \u4_u3_csr1_reg[0]/P0001  & ~n7347 ;
  assign n7349 = ~n7346 & n7348 ;
  assign n7350 = ~n7344 & n7349 ;
  assign n7351 = \u4_u0_dma_out_cnt_reg[9]/P0001  & ~n6822 ;
  assign n7352 = ~n6824 & n7351 ;
  assign n7353 = \u4_u0_dma_out_cnt_reg[9]/P0001  & n6821 ;
  assign n7354 = ~n7352 & ~n7353 ;
  assign n7355 = n6853 & ~n7353 ;
  assign n7356 = n6850 & n7355 ;
  assign n7357 = ~n7354 & ~n7356 ;
  assign n7358 = ~\u4_u0_dma_out_cnt_reg[4]/P0001  & ~\u4_u0_dma_out_cnt_reg[5]/P0001  ;
  assign n7359 = n6804 & n7358 ;
  assign n7360 = ~\u4_u0_dma_out_cnt_reg[8]/P0001  & ~\u4_u0_dma_out_cnt_reg[9]/P0001  ;
  assign n7361 = ~\u4_u0_dma_out_cnt_reg[6]/P0001  & ~\u4_u0_dma_out_cnt_reg[7]/P0001  ;
  assign n7362 = n7360 & n7361 ;
  assign n7363 = ~\u4_u0_dma_out_cnt_reg[10]/P0001  & n7362 ;
  assign n7364 = n7359 & n7363 ;
  assign n7365 = \u4_u0_r5_reg/NET0131  & ~n7364 ;
  assign n7366 = \u4_u0_dma_out_cnt_reg[10]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n7367 = ~n6339 & n7366 ;
  assign n7368 = ~n7365 & n7367 ;
  assign n7369 = n7357 & n7368 ;
  assign n7370 = ~\u4_u0_dma_out_cnt_reg[10]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n7371 = n7362 & n7370 ;
  assign n7372 = n7359 & n7371 ;
  assign n7373 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_out_cnt_reg[11]/P0001  ;
  assign n7374 = ~n7372 & n7373 ;
  assign n7375 = ~n7369 & n7374 ;
  assign n7376 = \u4_u0_csr1_reg[0]/P0001  & ~\u4_u0_dma_out_cnt_reg[11]/P0001  ;
  assign n7377 = n7372 & n7376 ;
  assign n7378 = n7368 & n7376 ;
  assign n7379 = n7357 & n7378 ;
  assign n7380 = ~n7377 & ~n7379 ;
  assign n7381 = ~n7375 & n7380 ;
  assign n7382 = ~n6822 & ~n6824 ;
  assign n7383 = ~n6821 & ~n7382 ;
  assign n7384 = ~n6821 & n6853 ;
  assign n7385 = n6850 & n7384 ;
  assign n7386 = ~n7383 & ~n7385 ;
  assign n7387 = ~\u4_u0_r5_reg/NET0131  & ~n7386 ;
  assign n7388 = ~\u4_u0_r5_reg/NET0131  & n6632 ;
  assign n7389 = ~\u4_u0_dma_out_cnt_reg[7]/P0001  & ~\u4_u0_dma_out_cnt_reg[8]/P0001  ;
  assign n7390 = \u4_u0_r5_reg/NET0131  & n7389 ;
  assign n7391 = n6805 & n7390 ;
  assign n7392 = ~n7388 & ~n7391 ;
  assign n7393 = \u4_u0_dma_out_cnt_reg[9]/P0001  & ~n7392 ;
  assign n7394 = ~n7387 & n7393 ;
  assign n7395 = ~\u4_u0_dma_out_cnt_reg[9]/P0001  & ~\u4_u0_r5_reg/NET0131  ;
  assign n7396 = ~n7386 & n7395 ;
  assign n7397 = ~\u4_u0_dma_out_cnt_reg[9]/P0001  & n7392 ;
  assign n7398 = \u4_u0_csr1_reg[0]/P0001  & ~n7397 ;
  assign n7399 = ~n7396 & n7398 ;
  assign n7400 = ~n7394 & n7399 ;
  assign n7401 = \u4_u1_dma_out_cnt_reg[9]/P0001  & ~n6886 ;
  assign n7402 = ~n6888 & n7401 ;
  assign n7403 = \u4_u1_dma_out_cnt_reg[9]/P0001  & n6885 ;
  assign n7404 = ~n7402 & ~n7403 ;
  assign n7405 = n6917 & ~n7403 ;
  assign n7406 = n6914 & n7405 ;
  assign n7407 = ~n7404 & ~n7406 ;
  assign n7408 = ~\u4_u1_dma_out_cnt_reg[4]/P0001  & ~\u4_u1_dma_out_cnt_reg[5]/P0001  ;
  assign n7409 = n6868 & n7408 ;
  assign n7410 = ~\u4_u1_dma_out_cnt_reg[8]/P0001  & ~\u4_u1_dma_out_cnt_reg[9]/P0001  ;
  assign n7411 = ~\u4_u1_dma_out_cnt_reg[6]/P0001  & ~\u4_u1_dma_out_cnt_reg[7]/P0001  ;
  assign n7412 = n7410 & n7411 ;
  assign n7413 = ~\u4_u1_dma_out_cnt_reg[10]/P0001  & n7412 ;
  assign n7414 = n7409 & n7413 ;
  assign n7415 = \u4_u1_r5_reg/NET0131  & ~n7414 ;
  assign n7416 = \u4_u1_dma_out_cnt_reg[10]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n7417 = ~n6368 & n7416 ;
  assign n7418 = ~n7415 & n7417 ;
  assign n7419 = n7407 & n7418 ;
  assign n7420 = ~\u4_u1_dma_out_cnt_reg[10]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n7421 = n7412 & n7420 ;
  assign n7422 = n7409 & n7421 ;
  assign n7423 = \u4_u1_csr1_reg[0]/P0001  & \u4_u1_dma_out_cnt_reg[11]/P0001  ;
  assign n7424 = ~n7422 & n7423 ;
  assign n7425 = ~n7419 & n7424 ;
  assign n7426 = \u4_u1_csr1_reg[0]/P0001  & ~\u4_u1_dma_out_cnt_reg[11]/P0001  ;
  assign n7427 = n7422 & n7426 ;
  assign n7428 = n7418 & n7426 ;
  assign n7429 = n7407 & n7428 ;
  assign n7430 = ~n7427 & ~n7429 ;
  assign n7431 = ~n7425 & n7430 ;
  assign n7432 = ~n6886 & ~n6888 ;
  assign n7433 = ~n6885 & ~n7432 ;
  assign n7434 = ~n6885 & n6917 ;
  assign n7435 = n6914 & n7434 ;
  assign n7436 = ~n7433 & ~n7435 ;
  assign n7437 = ~\u4_u1_r5_reg/NET0131  & ~n7436 ;
  assign n7438 = ~\u4_u1_r5_reg/NET0131  & n6369 ;
  assign n7439 = ~\u4_u1_dma_out_cnt_reg[7]/P0001  & ~\u4_u1_dma_out_cnt_reg[8]/P0001  ;
  assign n7440 = \u4_u1_r5_reg/NET0131  & n7439 ;
  assign n7441 = n6869 & n7440 ;
  assign n7442 = ~n7438 & ~n7441 ;
  assign n7443 = \u4_u1_dma_out_cnt_reg[9]/P0001  & ~n7442 ;
  assign n7444 = ~n7437 & n7443 ;
  assign n7445 = ~\u4_u1_dma_out_cnt_reg[9]/P0001  & ~\u4_u1_r5_reg/NET0131  ;
  assign n7446 = ~n7436 & n7445 ;
  assign n7447 = ~\u4_u1_dma_out_cnt_reg[9]/P0001  & n7442 ;
  assign n7448 = \u4_u1_csr1_reg[0]/P0001  & ~n7447 ;
  assign n7449 = ~n7446 & n7448 ;
  assign n7450 = ~n7444 & n7449 ;
  assign n7451 = \u4_u2_dma_out_cnt_reg[9]/P0001  & ~n6980 ;
  assign n7452 = ~n6982 & n7451 ;
  assign n7453 = \u4_u2_dma_out_cnt_reg[9]/P0001  & n6979 ;
  assign n7454 = ~n7452 & ~n7453 ;
  assign n7455 = n6952 & ~n7453 ;
  assign n7456 = n6977 & n7455 ;
  assign n7457 = ~n7454 & ~n7456 ;
  assign n7458 = ~\u4_u2_dma_out_cnt_reg[4]/P0001  & ~\u4_u2_dma_out_cnt_reg[5]/P0001  ;
  assign n7459 = n6932 & n7458 ;
  assign n7460 = ~\u4_u2_dma_out_cnt_reg[8]/P0001  & ~\u4_u2_dma_out_cnt_reg[9]/P0001  ;
  assign n7461 = ~\u4_u2_dma_out_cnt_reg[6]/P0001  & ~\u4_u2_dma_out_cnt_reg[7]/P0001  ;
  assign n7462 = n7460 & n7461 ;
  assign n7463 = ~\u4_u2_dma_out_cnt_reg[10]/P0001  & n7462 ;
  assign n7464 = n7459 & n7463 ;
  assign n7465 = \u4_u2_r5_reg/NET0131  & ~n7464 ;
  assign n7466 = \u4_u2_dma_out_cnt_reg[10]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n7467 = ~n6415 & n7466 ;
  assign n7468 = ~n7465 & n7467 ;
  assign n7469 = n7457 & n7468 ;
  assign n7470 = ~\u4_u2_dma_out_cnt_reg[10]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n7471 = n7462 & n7470 ;
  assign n7472 = n7459 & n7471 ;
  assign n7473 = \u4_u2_csr1_reg[0]/P0001  & \u4_u2_dma_out_cnt_reg[11]/P0001  ;
  assign n7474 = ~n7472 & n7473 ;
  assign n7475 = ~n7469 & n7474 ;
  assign n7476 = \u4_u2_csr1_reg[0]/P0001  & ~\u4_u2_dma_out_cnt_reg[11]/P0001  ;
  assign n7477 = n7472 & n7476 ;
  assign n7478 = n7468 & n7476 ;
  assign n7479 = n7457 & n7478 ;
  assign n7480 = ~n7477 & ~n7479 ;
  assign n7481 = ~n7475 & n7480 ;
  assign n7482 = ~n6980 & ~n6982 ;
  assign n7483 = ~n6979 & ~n7482 ;
  assign n7484 = n6952 & ~n6979 ;
  assign n7485 = n6977 & n7484 ;
  assign n7486 = ~n7483 & ~n7485 ;
  assign n7487 = ~\u4_u2_r5_reg/NET0131  & ~n7486 ;
  assign n7488 = ~\u4_u2_r5_reg/NET0131  & n6667 ;
  assign n7489 = ~\u4_u2_dma_out_cnt_reg[7]/P0001  & ~\u4_u2_dma_out_cnt_reg[8]/P0001  ;
  assign n7490 = \u4_u2_r5_reg/NET0131  & n7489 ;
  assign n7491 = n6933 & n7490 ;
  assign n7492 = ~n7488 & ~n7491 ;
  assign n7493 = \u4_u2_dma_out_cnt_reg[9]/P0001  & ~n7492 ;
  assign n7494 = ~n7487 & n7493 ;
  assign n7495 = ~\u4_u2_dma_out_cnt_reg[9]/P0001  & ~\u4_u2_r5_reg/NET0131  ;
  assign n7496 = ~n7486 & n7495 ;
  assign n7497 = ~\u4_u2_dma_out_cnt_reg[9]/P0001  & n7492 ;
  assign n7498 = \u4_u2_csr1_reg[0]/P0001  & ~n7497 ;
  assign n7499 = ~n7496 & n7498 ;
  assign n7500 = ~n7494 & n7499 ;
  assign n7501 = n6254 & ~n6586 ;
  assign n7502 = n6251 & n6270 ;
  assign n7503 = n7501 & n7502 ;
  assign n7504 = ~\u4_u3_dma_in_cnt_reg[9]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n7505 = ~n6283 & n7504 ;
  assign n7506 = ~n6282 & n7505 ;
  assign n7507 = ~n7503 & n7506 ;
  assign n7508 = ~\u4_u3_r5_reg/NET0131  & ~n7507 ;
  assign n7509 = n6251 & ~n6269 ;
  assign n7510 = n6584 & n7509 ;
  assign n7511 = ~n6250 & ~n6269 ;
  assign n7512 = ~n6590 & n7511 ;
  assign n7513 = n6589 & ~n7512 ;
  assign n7514 = ~n7510 & n7513 ;
  assign n7515 = ~\u4_u3_r5_reg/NET0131  & n6268 ;
  assign n7516 = ~n7514 & n7515 ;
  assign n7517 = \u4_u3_dma_in_cnt_reg[10]/P0001  & ~\u4_u3_r5_reg/NET0131  ;
  assign n7518 = \u4_u3_dma_in_cnt_reg[10]/P0001  & n7226 ;
  assign n7519 = n6277 & n7518 ;
  assign n7520 = ~n7517 & ~n7519 ;
  assign n7521 = ~n7516 & ~n7520 ;
  assign n7522 = ~n7508 & n7521 ;
  assign n7523 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[10]/P0001  ;
  assign n7524 = \u4_u3_csr1_reg[0]/P0001  & ~\u4_u3_r5_reg/NET0131  ;
  assign n7525 = \u4_u3_csr1_reg[0]/P0001  & n7226 ;
  assign n7526 = n6277 & n7525 ;
  assign n7527 = ~n7524 & ~n7526 ;
  assign n7528 = ~n7516 & ~n7527 ;
  assign n7529 = ~n7508 & n7528 ;
  assign n7530 = ~n7523 & ~n7529 ;
  assign n7531 = ~n7522 & ~n7530 ;
  assign n7532 = n6312 & ~n6620 ;
  assign n7533 = n6309 & n6328 ;
  assign n7534 = n7532 & n7533 ;
  assign n7535 = ~\u4_u0_dma_in_cnt_reg[9]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n7536 = ~n6340 & n7535 ;
  assign n7537 = ~n6339 & n7536 ;
  assign n7538 = ~n7534 & n7537 ;
  assign n7539 = ~\u4_u0_r5_reg/NET0131  & ~n7538 ;
  assign n7540 = n6309 & ~n6327 ;
  assign n7541 = n6618 & n7540 ;
  assign n7542 = ~n6308 & ~n6327 ;
  assign n7543 = ~n6624 & n7542 ;
  assign n7544 = n6623 & ~n7543 ;
  assign n7545 = ~n7541 & n7544 ;
  assign n7546 = ~\u4_u0_r5_reg/NET0131  & n6326 ;
  assign n7547 = ~n7545 & n7546 ;
  assign n7548 = \u4_u0_dma_in_cnt_reg[10]/P0001  & ~\u4_u0_r5_reg/NET0131  ;
  assign n7549 = \u4_u0_dma_in_cnt_reg[10]/P0001  & n7247 ;
  assign n7550 = n6335 & n7549 ;
  assign n7551 = ~n7548 & ~n7550 ;
  assign n7552 = ~n7547 & ~n7551 ;
  assign n7553 = ~n7539 & n7552 ;
  assign n7554 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[10]/P0001  ;
  assign n7555 = \u4_u0_csr1_reg[0]/P0001  & n7247 ;
  assign n7556 = n6335 & n7555 ;
  assign n7557 = ~n6613 & ~n7556 ;
  assign n7558 = ~n7547 & ~n7557 ;
  assign n7559 = ~n7539 & n7558 ;
  assign n7560 = ~n7554 & ~n7559 ;
  assign n7561 = ~n7553 & ~n7560 ;
  assign n7562 = \u4_u1_r5_reg/NET0131  & n7269 ;
  assign n7563 = n6362 & n7562 ;
  assign n7564 = ~n7438 & ~n7563 ;
  assign n7565 = ~\u4_u1_dma_in_cnt_reg[9]/P0001  & ~n6370 ;
  assign n7566 = ~n7564 & n7565 ;
  assign n7567 = ~n6404 & n7566 ;
  assign n7568 = n6656 & n7566 ;
  assign n7569 = ~n6655 & n7568 ;
  assign n7570 = ~n7567 & ~n7569 ;
  assign n7571 = \u4_u1_csr1_reg[0]/P0001  & \u4_u1_dma_in_cnt_reg[10]/P0001  ;
  assign n7572 = ~n7563 & n7571 ;
  assign n7573 = n7570 & n7572 ;
  assign n7574 = ~n7563 & n7570 ;
  assign n7575 = \u4_u1_csr1_reg[0]/P0001  & ~\u4_u1_dma_in_cnt_reg[10]/P0001  ;
  assign n7576 = ~n7574 & n7575 ;
  assign n7577 = ~n7573 & ~n7576 ;
  assign n7578 = ~\u4_u2_r5_reg/NET0131  & ~n6457 ;
  assign n7579 = ~n6457 & n7288 ;
  assign n7580 = n6463 & n7579 ;
  assign n7581 = ~n7578 & ~n7580 ;
  assign n7582 = \u4_u2_dma_in_cnt_reg[10]/P0001  & ~n7581 ;
  assign n7583 = ~n6456 & n7582 ;
  assign n7584 = ~\u4_u2_dma_in_cnt_reg[10]/P0001  & ~\u4_u2_r5_reg/NET0131  ;
  assign n7585 = ~n6455 & n7584 ;
  assign n7586 = ~\u4_u2_dma_in_cnt_reg[10]/P0001  & n7581 ;
  assign n7587 = \u4_u2_csr1_reg[0]/P0001  & ~n7586 ;
  assign n7588 = ~n7585 & n7587 ;
  assign n7589 = ~n7583 & n7588 ;
  assign n7590 = ~\u0_u0_me_cnt_100_ms_reg/P0001  & \u0_u0_me_ps2_0_5_ms_reg/P0001  ;
  assign n7591 = \u0_u0_me_cnt_reg[0]/P0001  & n7590 ;
  assign n7592 = ~\u0_u0_me_cnt_reg[1]/P0001  & ~n7591 ;
  assign n7593 = n6997 & n7590 ;
  assign n7594 = ~n7592 & ~n7593 ;
  assign n7595 = n6201 & n7594 ;
  assign n7596 = ~n6190 & n7595 ;
  assign n7597 = ~n6182 & n7596 ;
  assign n7598 = ~\u1_hms_clk_reg/P0001  & ~\u1_sof_time_reg[0]/P0001  ;
  assign n7599 = ~\u1_clr_sof_time_reg/P0001  & ~n6212 ;
  assign n7600 = ~n7598 & n7599 ;
  assign n7601 = ~\u0_u0_me_cnt_reg[0]/P0001  & ~n7590 ;
  assign n7602 = ~n7591 & ~n7601 ;
  assign n7603 = n6695 & n7602 ;
  assign n7604 = ~n6182 & n7603 ;
  assign n7605 = \u0_u0_me_cnt_reg[2]/P0001  & n7593 ;
  assign n7606 = ~\u0_u0_me_cnt_reg[2]/P0001  & ~n7593 ;
  assign n7607 = ~n7605 & ~n7606 ;
  assign n7608 = n6695 & n7607 ;
  assign n7609 = ~n6182 & n7608 ;
  assign n7610 = \u0_u0_me_cnt_reg[2]/P0001  & \u0_u0_me_cnt_reg[3]/P0001  ;
  assign n7611 = n7593 & n7610 ;
  assign n7612 = ~\u0_u0_me_cnt_reg[3]/P0001  & ~n7605 ;
  assign n7613 = ~n7611 & ~n7612 ;
  assign n7614 = n6695 & n7613 ;
  assign n7615 = ~n6182 & n7614 ;
  assign n7616 = \u0_u0_me_cnt_reg[2]/P0001  & \u0_u0_me_cnt_reg[4]/P0001  ;
  assign n7617 = \u0_u0_me_cnt_reg[3]/P0001  & n7616 ;
  assign n7618 = n7593 & n7617 ;
  assign n7619 = ~\u0_u0_me_cnt_reg[4]/P0001  & ~n7611 ;
  assign n7620 = ~n7618 & ~n7619 ;
  assign n7621 = n6201 & n7620 ;
  assign n7622 = ~n6190 & n7621 ;
  assign n7623 = ~n6182 & n7622 ;
  assign n7624 = \u0_u0_me_cnt_reg[5]/P0001  & n7618 ;
  assign n7625 = ~\u0_u0_me_cnt_reg[5]/P0001  & ~n7618 ;
  assign n7626 = ~n7624 & ~n7625 ;
  assign n7627 = n6695 & n7626 ;
  assign n7628 = ~n6182 & n7627 ;
  assign n7629 = \u0_u0_me_cnt_reg[5]/P0001  & \u0_u0_me_cnt_reg[6]/P0001  ;
  assign n7630 = n7618 & n7629 ;
  assign n7631 = n6201 & ~n7630 ;
  assign n7632 = ~n6190 & n7631 ;
  assign n7633 = ~\u0_u0_me_cnt_reg[6]/P0001  & ~n7624 ;
  assign n7634 = n7632 & ~n7633 ;
  assign n7635 = ~n6182 & n7634 ;
  assign n7636 = ~\u0_u0_me_cnt_reg[7]/P0001  & ~n7630 ;
  assign n7637 = n6201 & ~n7636 ;
  assign n7638 = ~n6190 & n7637 ;
  assign n7639 = \u0_u0_me_cnt_reg[5]/P0001  & \u0_u0_me_cnt_reg[7]/P0001  ;
  assign n7640 = \u0_u0_me_cnt_reg[6]/P0001  & n7639 ;
  assign n7641 = n7618 & n7640 ;
  assign n7642 = n7638 & ~n7641 ;
  assign n7643 = ~n6182 & n7642 ;
  assign n7644 = \u4_u2_dma_in_buf_sz1_reg/P0001  & n5171 ;
  assign n7645 = n5156 & n7644 ;
  assign n7646 = \u4_u0_dma_in_buf_sz1_reg/P0001  & n5140 ;
  assign n7647 = \u4_u1_dma_in_buf_sz1_reg/P0001  & n5175 ;
  assign n7648 = ~n7646 & ~n7647 ;
  assign n7649 = ~n7645 & n7648 ;
  assign n7650 = \u4_dma_in_buf_sz1_reg/P0001  & n5198 ;
  assign n7651 = \u4_u3_dma_in_buf_sz1_reg/P0001  & n5195 ;
  assign n7652 = ~n7650 & ~n7651 ;
  assign n7653 = n7649 & n7652 ;
  assign n7654 = \u1_sof_time_reg[9]/P0001  & n6218 ;
  assign n7655 = n6217 & n7654 ;
  assign n7656 = n6215 & n7655 ;
  assign n7657 = ~\u1_sof_time_reg[10]/P0001  & ~n7656 ;
  assign n7658 = ~\u1_clr_sof_time_reg/P0001  & ~n6222 ;
  assign n7659 = ~n7657 & n7658 ;
  assign n7660 = ~\u1_clr_sof_time_reg/P0001  & \u1_sof_time_reg[1]/P0001  ;
  assign n7661 = ~n6212 & n7660 ;
  assign n7662 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_sof_time_reg[1]/P0001  ;
  assign n7663 = n6212 & n7662 ;
  assign n7664 = ~n7661 & ~n7663 ;
  assign n7665 = \u1_sof_time_reg[1]/P0001  & n6212 ;
  assign n7666 = ~\u1_sof_time_reg[2]/P0001  & ~n7665 ;
  assign n7667 = ~\u1_clr_sof_time_reg/P0001  & ~n7110 ;
  assign n7668 = ~n7666 & n7667 ;
  assign n7669 = ~\u1_clr_sof_time_reg/P0001  & \u1_sof_time_reg[3]/P0001  ;
  assign n7670 = ~n7110 & n7669 ;
  assign n7671 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_sof_time_reg[3]/P0001  ;
  assign n7672 = n7110 & n7671 ;
  assign n7673 = ~n7670 & ~n7672 ;
  assign n7674 = \u1_sof_time_reg[3]/P0001  & n7110 ;
  assign n7675 = ~\u1_sof_time_reg[4]/P0001  & ~n7674 ;
  assign n7676 = \u1_sof_time_reg[3]/P0001  & \u1_sof_time_reg[4]/P0001  ;
  assign n7677 = n7110 & n7676 ;
  assign n7678 = ~\u1_clr_sof_time_reg/P0001  & ~n7677 ;
  assign n7679 = ~n7675 & n7678 ;
  assign n7680 = ~\u1_sof_time_reg[5]/P0001  & ~n7677 ;
  assign n7681 = ~\u1_clr_sof_time_reg/P0001  & ~n7111 ;
  assign n7682 = ~n7680 & n7681 ;
  assign n7683 = ~\u1_clr_sof_time_reg/P0001  & \u1_sof_time_reg[6]/P0001  ;
  assign n7684 = ~n7111 & n7683 ;
  assign n7685 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_sof_time_reg[6]/P0001  ;
  assign n7686 = n7111 & n7685 ;
  assign n7687 = ~n7684 & ~n7686 ;
  assign n7688 = n6217 & n6218 ;
  assign n7689 = n6215 & n7688 ;
  assign n7690 = ~\u1_clr_sof_time_reg/P0001  & \u1_sof_time_reg[8]/P0001  ;
  assign n7691 = ~\u1_clr_sof_time_reg/P0001  & n7114 ;
  assign n7692 = n7111 & n7691 ;
  assign n7693 = ~n7690 & ~n7692 ;
  assign n7694 = ~n7689 & ~n7693 ;
  assign n7695 = ~\u1_clr_sof_time_reg/P0001  & \u1_sof_time_reg[9]/P0001  ;
  assign n7696 = ~n7689 & n7695 ;
  assign n7697 = ~\u1_clr_sof_time_reg/P0001  & ~\u1_sof_time_reg[9]/P0001  ;
  assign n7698 = n6214 & n7697 ;
  assign n7699 = n7111 & n7698 ;
  assign n7700 = ~n7696 & ~n7699 ;
  assign n7701 = ~\u4_crc5_err_r_reg/P0001  & ~\u4_int_srcb_reg[0]/P0001  ;
  assign n7702 = n5667 & ~n7701 ;
  assign n7703 = ~\u1_u2_sizu_c_reg[10]/P0001  & \u4_csr_reg[10]/P0001  ;
  assign n7704 = \u1_u2_sizu_c_reg[9]/P0001  & ~\u4_csr_reg[9]/NET0131  ;
  assign n7705 = \u1_u2_sizu_c_reg[10]/P0001  & ~\u4_csr_reg[10]/P0001  ;
  assign n7706 = ~n7704 & ~n7705 ;
  assign n7707 = \u1_u2_sizu_c_reg[8]/NET0131  & ~\u4_csr_reg[8]/P0001  ;
  assign n7708 = \u1_u2_sizu_c_reg[7]/P0001  & ~\u4_csr_reg[7]/P0001  ;
  assign n7709 = ~n7707 & ~n7708 ;
  assign n7710 = ~\u1_u2_sizu_c_reg[9]/P0001  & \u4_csr_reg[9]/NET0131  ;
  assign n7711 = ~\u1_u2_sizu_c_reg[8]/NET0131  & \u4_csr_reg[8]/P0001  ;
  assign n7712 = ~n7710 & ~n7711 ;
  assign n7713 = ~n7709 & n7712 ;
  assign n7714 = n7706 & ~n7713 ;
  assign n7715 = ~n7703 & ~n7714 ;
  assign n7716 = ~\u1_u2_sizu_c_reg[4]/P0001  & \u4_csr_reg[4]/NET0131  ;
  assign n7717 = ~\u1_u2_sizu_c_reg[3]/P0001  & \u4_csr_reg[3]/P0001  ;
  assign n7718 = ~n7716 & ~n7717 ;
  assign n7719 = \u1_u2_sizu_c_reg[6]/P0001  & ~\u4_csr_reg[6]/NET0131  ;
  assign n7720 = \u1_u2_sizu_c_reg[5]/P0001  & ~\u4_csr_reg[5]/NET0131  ;
  assign n7721 = ~n7719 & ~n7720 ;
  assign n7722 = \u1_u2_sizu_c_reg[4]/P0001  & ~\u4_csr_reg[4]/NET0131  ;
  assign n7723 = n7721 & ~n7722 ;
  assign n7724 = ~n7718 & n7723 ;
  assign n7725 = ~\u1_u2_sizu_c_reg[7]/P0001  & \u4_csr_reg[7]/P0001  ;
  assign n7726 = ~n7711 & ~n7725 ;
  assign n7727 = n7706 & ~n7707 ;
  assign n7728 = ~n7726 & n7727 ;
  assign n7729 = ~n7703 & ~n7710 ;
  assign n7730 = ~n7705 & ~n7729 ;
  assign n7731 = ~\u1_u2_sizu_c_reg[6]/P0001  & \u4_csr_reg[6]/NET0131  ;
  assign n7732 = ~\u1_u2_sizu_c_reg[5]/P0001  & \u4_csr_reg[5]/NET0131  ;
  assign n7733 = ~n7731 & ~n7732 ;
  assign n7734 = ~n7719 & ~n7733 ;
  assign n7735 = ~n7730 & ~n7734 ;
  assign n7736 = ~n7728 & n7735 ;
  assign n7737 = ~n7724 & n7736 ;
  assign n7738 = ~n7715 & ~n7737 ;
  assign n7739 = ~\u4_csr_reg[16]/P0001  & n7738 ;
  assign n7740 = ~n7728 & ~n7730 ;
  assign n7741 = \u1_u2_sizu_c_reg[3]/P0001  & ~\u4_csr_reg[3]/P0001  ;
  assign n7742 = ~n7722 & ~n7741 ;
  assign n7743 = ~n7716 & ~n7732 ;
  assign n7744 = ~n7742 & n7743 ;
  assign n7745 = n7721 & ~n7744 ;
  assign n7746 = ~n7731 & ~n7745 ;
  assign n7747 = ~n7715 & ~n7746 ;
  assign n7748 = n7740 & ~n7747 ;
  assign n7749 = ~\u1_u2_sizu_c_reg[2]/P0001  & \u4_csr_reg[2]/NET0131  ;
  assign n7750 = ~\u1_u2_sizu_c_reg[0]/P0001  & \u4_csr_reg[0]/P0001  ;
  assign n7751 = ~\u1_u2_sizu_c_reg[1]/P0001  & \u4_csr_reg[1]/P0001  ;
  assign n7752 = ~n7750 & ~n7751 ;
  assign n7753 = \u1_u2_sizu_c_reg[2]/P0001  & ~\u4_csr_reg[2]/NET0131  ;
  assign n7754 = \u1_u2_sizu_c_reg[1]/P0001  & ~\u4_csr_reg[1]/P0001  ;
  assign n7755 = ~n7753 & ~n7754 ;
  assign n7756 = ~n7752 & n7755 ;
  assign n7757 = ~n7749 & ~n7756 ;
  assign n7758 = ~\u4_csr_reg[16]/P0001  & ~n7757 ;
  assign n7759 = ~n7748 & n7758 ;
  assign n7760 = ~n7739 & ~n7759 ;
  assign n7761 = \u1_u3_new_size_reg[2]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n7762 = \u1_u2_sizu_c_reg[2]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n7763 = ~n7761 & ~n7762 ;
  assign n7764 = \u1_u3_new_size_reg[3]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n7765 = \u1_u2_sizu_c_reg[3]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n7766 = ~n7764 & ~n7765 ;
  assign n7767 = ~n5700 & ~n5715 ;
  assign n7768 = ~n5716 & n7767 ;
  assign n7769 = ~n5714 & n7768 ;
  assign n7770 = ~n5711 & ~n7767 ;
  assign n7771 = ~n5710 & ~n5712 ;
  assign n7772 = ~n5716 & ~n7771 ;
  assign n7773 = n7770 & ~n7772 ;
  assign n7774 = ~n7769 & ~n7773 ;
  assign n7775 = ~n5714 & n5717 ;
  assign n7776 = ~n5696 & ~n5699 ;
  assign n7777 = ~n5700 & ~n7776 ;
  assign n7778 = ~n7775 & n7777 ;
  assign n7779 = n5700 & n7776 ;
  assign n7780 = n5717 & n7776 ;
  assign n7781 = ~n5714 & n7780 ;
  assign n7782 = ~n7779 & ~n7781 ;
  assign n7783 = ~n7778 & n7782 ;
  assign n7784 = ~n5693 & ~n5722 ;
  assign n7785 = ~n5692 & ~n5697 ;
  assign n7786 = ~n5692 & n5701 ;
  assign n7787 = ~n7785 & ~n7786 ;
  assign n7788 = n5717 & ~n7785 ;
  assign n7789 = ~n5714 & n7788 ;
  assign n7790 = ~n7787 & ~n7789 ;
  assign n7791 = ~n7784 & n7790 ;
  assign n7792 = n7784 & ~n7790 ;
  assign n7793 = ~n7791 & ~n7792 ;
  assign n7794 = ~n7708 & n7721 ;
  assign n7795 = n7727 & n7794 ;
  assign n7796 = n7742 & n7795 ;
  assign n7797 = ~\u4_csr_reg[17]/P0001  & ~n7796 ;
  assign n7798 = \u1_u2_sizu_c_reg[0]/P0001  & ~\u4_csr_reg[0]/P0001  ;
  assign n7799 = n7755 & ~n7798 ;
  assign n7800 = n7751 & ~n7753 ;
  assign n7801 = ~\u4_csr_reg[17]/P0001  & ~n7749 ;
  assign n7802 = ~n7800 & n7801 ;
  assign n7803 = ~n7799 & n7802 ;
  assign n7804 = ~n7797 & ~n7803 ;
  assign n7805 = ~n7738 & ~n7804 ;
  assign n7806 = \u1_u0_pid_reg[0]/NET0131  & \u1_u0_pid_reg[1]/NET0131  ;
  assign n7807 = n7203 & n7806 ;
  assign n7808 = n7200 & n7807 ;
  assign n7809 = rst_i_pad & n7808 ;
  assign n7810 = \u0_rx_active_reg/P0001  & \u1_u0_state_reg[3]/P0001  ;
  assign n7811 = rst_i_pad & n7810 ;
  assign n7812 = ~n7211 & n7811 ;
  assign n7813 = ~n7809 & ~n7812 ;
  assign n7814 = \u4_u2_buf0_orig_reg[27]/P0001  & ~\u4_u2_dma_in_cnt_reg[8]/P0001  ;
  assign n7815 = \u4_u2_buf0_orig_reg[26]/P0001  & ~\u4_u2_dma_in_cnt_reg[7]/P0001  ;
  assign n7816 = ~n7814 & ~n7815 ;
  assign n7817 = ~\u4_u2_buf0_orig_reg[25]/P0001  & \u4_u2_dma_in_cnt_reg[6]/P0001  ;
  assign n7818 = ~\u4_u2_buf0_orig_reg[26]/P0001  & \u4_u2_dma_in_cnt_reg[7]/P0001  ;
  assign n7819 = ~n7817 & ~n7818 ;
  assign n7820 = n7816 & ~n7819 ;
  assign n7821 = ~\u4_u2_buf0_orig_reg[23]/P0001  & \u4_u2_dma_in_cnt_reg[4]/P0001  ;
  assign n7822 = ~\u4_u2_buf0_orig_reg[24]/P0001  & \u4_u2_dma_in_cnt_reg[5]/P0001  ;
  assign n7823 = ~n7821 & ~n7822 ;
  assign n7824 = \u4_u2_buf0_orig_reg[23]/P0001  & ~\u4_u2_dma_in_cnt_reg[4]/P0001  ;
  assign n7825 = \u4_u2_buf0_orig_reg[22]/P0001  & ~\u4_u2_dma_in_cnt_reg[3]/P0001  ;
  assign n7826 = ~n7824 & ~n7825 ;
  assign n7827 = n7823 & ~n7826 ;
  assign n7828 = \u4_u2_buf0_orig_reg[19]/P0001  & ~\u4_u2_dma_in_cnt_reg[0]/P0001  ;
  assign n7829 = ~\u4_u2_buf0_orig_reg[20]/P0001  & \u4_u2_dma_in_cnt_reg[1]/P0001  ;
  assign n7830 = n7828 & ~n7829 ;
  assign n7831 = \u4_u2_buf0_orig_reg[21]/P0001  & ~\u4_u2_dma_in_cnt_reg[2]/P0001  ;
  assign n7832 = \u4_u2_buf0_orig_reg[20]/P0001  & ~\u4_u2_dma_in_cnt_reg[1]/P0001  ;
  assign n7833 = ~n7831 & ~n7832 ;
  assign n7834 = ~n7830 & n7833 ;
  assign n7835 = ~\u4_u2_buf0_orig_reg[21]/P0001  & \u4_u2_dma_in_cnt_reg[2]/P0001  ;
  assign n7836 = ~\u4_u2_buf0_orig_reg[22]/P0001  & \u4_u2_dma_in_cnt_reg[3]/P0001  ;
  assign n7837 = ~n7835 & ~n7836 ;
  assign n7838 = n7823 & n7837 ;
  assign n7839 = ~n7834 & n7838 ;
  assign n7840 = ~n7827 & ~n7839 ;
  assign n7841 = \u4_u2_buf0_orig_reg[25]/P0001  & ~\u4_u2_dma_in_cnt_reg[6]/P0001  ;
  assign n7842 = \u4_u2_buf0_orig_reg[24]/P0001  & ~\u4_u2_dma_in_cnt_reg[5]/P0001  ;
  assign n7843 = ~n7841 & ~n7842 ;
  assign n7844 = n7816 & n7843 ;
  assign n7845 = n7840 & n7844 ;
  assign n7846 = ~n7820 & ~n7845 ;
  assign n7847 = ~\u4_u2_buf0_orig_reg[30]/NET0131  & \u4_u2_dma_in_cnt_reg[11]/P0001  ;
  assign n7848 = \u4_u2_csr1_reg[11]/P0001  & ~\u4_u2_csr1_reg[12]/P0001  ;
  assign n7849 = \u4_u2_csr1_reg[0]/P0001  & n7848 ;
  assign n7850 = ~n7847 & n7849 ;
  assign n7851 = \u4_u2_buf0_orig_reg[30]/NET0131  & ~\u4_u2_dma_in_cnt_reg[11]/P0001  ;
  assign n7852 = ~\u4_u2_buf0_orig_reg[29]/NET0131  & \u4_u2_dma_in_cnt_reg[10]/P0001  ;
  assign n7853 = ~n7851 & n7852 ;
  assign n7854 = ~\u4_u2_buf0_orig_reg[27]/P0001  & \u4_u2_dma_in_cnt_reg[8]/P0001  ;
  assign n7855 = ~\u4_u2_buf0_orig_reg[28]/P0001  & \u4_u2_dma_in_cnt_reg[9]/P0001  ;
  assign n7856 = ~n7854 & ~n7855 ;
  assign n7857 = ~n7853 & n7856 ;
  assign n7858 = n7850 & n7857 ;
  assign n7859 = n7846 & n7858 ;
  assign n7860 = \u4_u2_buf0_orig_reg[28]/P0001  & ~\u4_u2_dma_in_cnt_reg[9]/P0001  ;
  assign n7861 = \u4_u2_buf0_orig_reg[29]/NET0131  & ~\u4_u2_dma_in_cnt_reg[10]/P0001  ;
  assign n7862 = ~n7851 & ~n7861 ;
  assign n7863 = ~n7860 & n7862 ;
  assign n7864 = n7850 & ~n7863 ;
  assign n7865 = ~n7853 & n7864 ;
  assign n7866 = ~\u4_u2_dma_out_cnt_reg[10]/P0001  & n7458 ;
  assign n7867 = ~\u4_u2_dma_out_cnt_reg[11]/P0001  & n6931 ;
  assign n7868 = n7866 & n7867 ;
  assign n7869 = n6930 & n7462 ;
  assign n7870 = n7868 & n7869 ;
  assign n7871 = \u4_u2_csr1_reg[0]/P0001  & n4355 ;
  assign n7872 = ~n7870 & n7871 ;
  assign n7873 = ~n7865 & ~n7872 ;
  assign n7874 = ~n7859 & n7873 ;
  assign n7875 = ~\u4_u2_r2_reg/P0001  & ~\u4_u2_r4_reg/P0001  ;
  assign n7876 = ~\u4_u2_r5_reg/NET0131  & n7875 ;
  assign n7877 = ~n7874 & n7876 ;
  assign n7878 = \u4_u3_buf0_orig_reg[26]/P0001  & ~\u4_u3_dma_in_cnt_reg[7]/P0001  ;
  assign n7879 = \u4_u3_buf0_orig_reg[27]/P0001  & ~\u4_u3_dma_in_cnt_reg[8]/P0001  ;
  assign n7880 = \u4_u3_buf0_orig_reg[28]/P0001  & ~\u4_u3_dma_in_cnt_reg[9]/P0001  ;
  assign n7881 = ~n7879 & ~n7880 ;
  assign n7882 = ~n7878 & n7881 ;
  assign n7883 = ~\u4_u3_buf0_orig_reg[25]/P0001  & \u4_u3_dma_in_cnt_reg[6]/P0001  ;
  assign n7884 = ~\u4_u3_buf0_orig_reg[26]/P0001  & \u4_u3_dma_in_cnt_reg[7]/P0001  ;
  assign n7885 = ~n7883 & ~n7884 ;
  assign n7886 = n7882 & ~n7885 ;
  assign n7887 = ~\u4_u3_buf0_orig_reg[24]/P0001  & \u4_u3_dma_in_cnt_reg[5]/P0001  ;
  assign n7888 = ~\u4_u3_buf0_orig_reg[23]/P0001  & \u4_u3_dma_in_cnt_reg[4]/P0001  ;
  assign n7889 = ~n7887 & ~n7888 ;
  assign n7890 = \u4_u3_buf0_orig_reg[23]/P0001  & ~\u4_u3_dma_in_cnt_reg[4]/P0001  ;
  assign n7891 = \u4_u3_buf0_orig_reg[22]/P0001  & ~\u4_u3_dma_in_cnt_reg[3]/P0001  ;
  assign n7892 = ~n7890 & ~n7891 ;
  assign n7893 = n7889 & ~n7892 ;
  assign n7894 = \u4_u3_buf0_orig_reg[19]/P0001  & ~\u4_u3_dma_in_cnt_reg[0]/P0001  ;
  assign n7895 = \u4_u3_dma_in_cnt_reg[1]/P0001  & ~n7894 ;
  assign n7896 = \u4_u3_buf0_orig_reg[20]/P0001  & ~n7895 ;
  assign n7897 = \u4_u3_buf0_orig_reg[21]/P0001  & ~\u4_u3_dma_in_cnt_reg[2]/P0001  ;
  assign n7898 = ~\u4_u3_dma_in_cnt_reg[1]/P0001  & n7894 ;
  assign n7899 = ~n7897 & ~n7898 ;
  assign n7900 = ~n7896 & n7899 ;
  assign n7901 = ~\u4_u3_buf0_orig_reg[22]/P0001  & \u4_u3_dma_in_cnt_reg[3]/P0001  ;
  assign n7902 = ~\u4_u3_buf0_orig_reg[21]/P0001  & \u4_u3_dma_in_cnt_reg[2]/P0001  ;
  assign n7903 = ~n7901 & ~n7902 ;
  assign n7904 = n7889 & n7903 ;
  assign n7905 = ~n7900 & n7904 ;
  assign n7906 = ~n7893 & ~n7905 ;
  assign n7907 = \u4_u3_buf0_orig_reg[25]/P0001  & ~\u4_u3_dma_in_cnt_reg[6]/P0001  ;
  assign n7908 = \u4_u3_buf0_orig_reg[24]/P0001  & ~\u4_u3_dma_in_cnt_reg[5]/P0001  ;
  assign n7909 = ~n7907 & ~n7908 ;
  assign n7910 = n7882 & n7909 ;
  assign n7911 = n7906 & n7910 ;
  assign n7912 = ~n7886 & ~n7911 ;
  assign n7913 = \u4_u3_buf0_orig_reg[30]/NET0131  & ~\u4_u3_dma_in_cnt_reg[11]/P0001  ;
  assign n7914 = ~\u4_u3_buf0_orig_reg[29]/NET0131  & \u4_u3_dma_in_cnt_reg[10]/P0001  ;
  assign n7915 = ~n7913 & n7914 ;
  assign n7916 = ~\u4_u3_buf0_orig_reg[30]/NET0131  & \u4_u3_dma_in_cnt_reg[11]/P0001  ;
  assign n7917 = \u4_u3_csr1_reg[11]/P0001  & ~\u4_u3_csr1_reg[12]/P0001  ;
  assign n7918 = \u4_u3_csr1_reg[0]/P0001  & n7917 ;
  assign n7919 = ~n7916 & n7918 ;
  assign n7920 = ~n7915 & n7919 ;
  assign n7921 = ~\u4_u3_buf0_orig_reg[28]/P0001  & \u4_u3_dma_in_cnt_reg[9]/P0001  ;
  assign n7922 = ~\u4_u3_buf0_orig_reg[27]/P0001  & \u4_u3_dma_in_cnt_reg[8]/P0001  ;
  assign n7923 = ~n7880 & n7922 ;
  assign n7924 = ~n7921 & ~n7923 ;
  assign n7925 = n7920 & n7924 ;
  assign n7926 = n7912 & n7925 ;
  assign n7927 = \u4_u3_buf0_orig_reg[29]/NET0131  & ~\u4_u3_dma_in_cnt_reg[10]/P0001  ;
  assign n7928 = ~n7913 & ~n7927 ;
  assign n7929 = ~n7915 & ~n7928 ;
  assign n7930 = n7919 & n7929 ;
  assign n7931 = ~\u4_u3_dma_out_cnt_reg[10]/P0001  & n7308 ;
  assign n7932 = ~\u4_u3_dma_out_cnt_reg[11]/P0001  & n6739 ;
  assign n7933 = n7931 & n7932 ;
  assign n7934 = n6738 & n7312 ;
  assign n7935 = n7933 & n7934 ;
  assign n7936 = \u4_u3_csr1_reg[0]/P0001  & n4366 ;
  assign n7937 = ~n7935 & n7936 ;
  assign n7938 = ~n7930 & ~n7937 ;
  assign n7939 = ~n7926 & n7938 ;
  assign n7940 = ~\u4_u3_r2_reg/P0001  & ~\u4_u3_r4_reg/P0001  ;
  assign n7941 = ~\u4_u3_r5_reg/NET0131  & n7940 ;
  assign n7942 = ~n7939 & n7941 ;
  assign n7943 = \u1_u2_sizu_c_reg[10]/P0001  & \u1_u2_sizu_c_reg[9]/P0001  ;
  assign n7944 = n7015 & n7943 ;
  assign n7945 = n7021 & n7944 ;
  assign n7946 = \u1_u2_sizu_c_reg[10]/P0001  & n7018 ;
  assign n7947 = \u1_u2_sizu_c_reg[9]/P0001  & n7018 ;
  assign n7948 = n7015 & n7947 ;
  assign n7949 = n7021 & n7948 ;
  assign n7950 = ~n7946 & ~n7949 ;
  assign n7951 = ~n7945 & ~n7950 ;
  assign n7952 = ~\u1_u2_word_done_r_reg/P0001  & \u1_u2_word_done_reg/NET0131  ;
  assign n7953 = \u5_state_reg[0]/P0001  & ~\u5_wb_req_s1_reg/P0001  ;
  assign n7954 = n2558 & n7953 ;
  assign n7955 = n2557 & n7954 ;
  assign n7956 = ~\u5_state_reg[3]/P0001  & ~\u5_state_reg[4]/P0001  ;
  assign n7957 = ~\u5_state_reg[0]/P0001  & ~\u5_state_reg[1]/P0001  ;
  assign n7958 = ~\u5_state_reg[2]/P0001  & \u5_state_reg[5]/NET0131  ;
  assign n7959 = n7957 & n7958 ;
  assign n7960 = n7956 & n7959 ;
  assign n7961 = rst_i_pad & ~n7960 ;
  assign n7962 = ~n7955 & n7961 ;
  assign n7963 = \u1_u2_rx_data_st_r_reg[2]/P0001  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n7964 = ~\u1_u2_dtmp_sel_r_reg/P0001  & n4033 ;
  assign n7965 = n7963 & n7964 ;
  assign n7966 = \u1_u2_rx_data_valid_r_reg/NET0131  & n4033 ;
  assign n7967 = \u1_u2_dtmp_r_reg[10]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7968 = ~n7966 & n7967 ;
  assign n7969 = ~n7965 & ~n7968 ;
  assign n7970 = \sram_data_i[10]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7971 = n7969 & ~n7970 ;
  assign n7972 = \u1_u2_rx_data_st_r_reg[3]/P0001  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n7973 = n7964 & n7972 ;
  assign n7974 = \u1_u2_dtmp_r_reg[11]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7975 = ~n7966 & n7974 ;
  assign n7976 = \sram_data_i[11]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7977 = ~n7975 & ~n7976 ;
  assign n7978 = ~n7973 & n7977 ;
  assign n7979 = \u1_u2_rx_data_st_r_reg[4]/P0001  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n7980 = n7964 & n7979 ;
  assign n7981 = \u1_u2_dtmp_r_reg[12]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7982 = ~n7966 & n7981 ;
  assign n7983 = \sram_data_i[12]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7984 = ~n7982 & ~n7983 ;
  assign n7985 = ~n7980 & n7984 ;
  assign n7986 = \u1_u2_rx_data_st_r_reg[5]/P0001  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n7987 = n7964 & n7986 ;
  assign n7988 = \u1_u2_dtmp_r_reg[13]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7989 = ~n7966 & n7988 ;
  assign n7990 = \sram_data_i[13]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7991 = ~n7989 & ~n7990 ;
  assign n7992 = ~n7987 & n7991 ;
  assign n7993 = \u1_u2_rx_data_st_r_reg[6]/P0001  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n7994 = n7964 & n7993 ;
  assign n7995 = \u1_u2_dtmp_r_reg[14]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7996 = ~n7966 & n7995 ;
  assign n7997 = ~n7994 & ~n7996 ;
  assign n7998 = \sram_data_i[14]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n7999 = n7997 & ~n7998 ;
  assign n8000 = \u1_u2_rx_data_st_r_reg[7]/P0001  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n8001 = n7964 & n8000 ;
  assign n8002 = \u1_u2_dtmp_r_reg[15]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8003 = ~n7966 & n8002 ;
  assign n8004 = ~n8001 & ~n8003 ;
  assign n8005 = \sram_data_i[15]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8006 = n8004 & ~n8005 ;
  assign n8007 = \u1_u2_rx_data_st_r_reg[0]/P0001  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n8008 = ~\u1_u2_dtmp_sel_r_reg/P0001  & n8007 ;
  assign n8009 = n4034 & n8008 ;
  assign n8010 = \u1_u2_rx_data_valid_r_reg/NET0131  & n4034 ;
  assign n8011 = \u1_u2_dtmp_r_reg[16]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8012 = ~n8010 & n8011 ;
  assign n8013 = ~n8009 & ~n8012 ;
  assign n8014 = \sram_data_i[16]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8015 = n8013 & ~n8014 ;
  assign n8016 = \u1_u2_rx_data_st_r_reg[1]/P0001  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n8017 = ~\u1_u2_dtmp_sel_r_reg/P0001  & n8016 ;
  assign n8018 = n4034 & n8017 ;
  assign n8019 = \u1_u2_dtmp_r_reg[17]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8020 = ~n8010 & n8019 ;
  assign n8021 = ~n8018 & ~n8020 ;
  assign n8022 = \sram_data_i[17]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8023 = n8021 & ~n8022 ;
  assign n8024 = ~\u1_u2_dtmp_sel_r_reg/P0001  & n7963 ;
  assign n8025 = n4034 & n8024 ;
  assign n8026 = \u1_u2_dtmp_r_reg[18]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8027 = ~n8010 & n8026 ;
  assign n8028 = ~n8025 & ~n8027 ;
  assign n8029 = \sram_data_i[18]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8030 = n8028 & ~n8029 ;
  assign n8031 = ~\u1_u2_dtmp_sel_r_reg/P0001  & \u1_u2_rx_data_valid_r_reg/NET0131  ;
  assign n8032 = n4034 & n8031 ;
  assign n8033 = \u1_u2_rx_data_st_r_reg[3]/P0001  & n8032 ;
  assign n8034 = \u1_u2_dtmp_r_reg[19]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8035 = ~n8010 & n8034 ;
  assign n8036 = \sram_data_i[19]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8037 = ~n8035 & ~n8036 ;
  assign n8038 = ~n8033 & n8037 ;
  assign n8039 = \u1_u2_rx_data_st_r_reg[4]/P0001  & n8032 ;
  assign n8040 = \u1_u2_dtmp_r_reg[20]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8041 = ~n8010 & n8040 ;
  assign n8042 = \sram_data_i[20]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8043 = ~n8041 & ~n8042 ;
  assign n8044 = ~n8039 & n8043 ;
  assign n8045 = \u1_u2_rx_data_st_r_reg[5]/P0001  & n8032 ;
  assign n8046 = \u1_u2_dtmp_r_reg[21]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8047 = ~n8010 & n8046 ;
  assign n8048 = \sram_data_i[21]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8049 = ~n8047 & ~n8048 ;
  assign n8050 = ~n8045 & n8049 ;
  assign n8051 = \u1_u2_rx_data_st_r_reg[6]/P0001  & n8032 ;
  assign n8052 = \u1_u2_dtmp_r_reg[22]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8053 = ~n8010 & n8052 ;
  assign n8054 = \sram_data_i[22]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8055 = ~n8053 & ~n8054 ;
  assign n8056 = ~n8051 & n8055 ;
  assign n8057 = \u1_u2_rx_data_st_r_reg[7]/P0001  & n8032 ;
  assign n8058 = \u1_u2_dtmp_r_reg[23]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8059 = ~n8010 & n8058 ;
  assign n8060 = \sram_data_i[23]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8061 = ~n8059 & ~n8060 ;
  assign n8062 = ~n8057 & n8061 ;
  assign n8063 = \u1_u2_adr_cb_reg[0]/NET0131  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8064 = n8007 & n8063 ;
  assign n8065 = \u1_u2_adr_cb_reg[1]/NET0131  & n8064 ;
  assign n8066 = \u1_u2_rx_data_valid_r_reg/NET0131  & n4018 ;
  assign n8067 = \u1_u2_dtmp_r_reg[24]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8068 = ~n8066 & n8067 ;
  assign n8069 = ~n8065 & ~n8068 ;
  assign n8070 = \sram_data_i[24]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8071 = n8069 & ~n8070 ;
  assign n8072 = n4018 & n8017 ;
  assign n8073 = \u1_u2_dtmp_r_reg[25]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8074 = ~n8066 & n8073 ;
  assign n8075 = \sram_data_i[25]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8076 = ~n8074 & ~n8075 ;
  assign n8077 = ~n8072 & n8076 ;
  assign n8078 = n4018 & n8024 ;
  assign n8079 = \u1_u2_dtmp_r_reg[26]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8080 = ~n8066 & n8079 ;
  assign n8081 = \sram_data_i[26]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8082 = ~n8080 & ~n8081 ;
  assign n8083 = ~n8078 & n8082 ;
  assign n8084 = n4018 & n8031 ;
  assign n8085 = \u1_u2_rx_data_st_r_reg[3]/P0001  & n8084 ;
  assign n8086 = \u1_u2_dtmp_r_reg[27]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8087 = ~n8066 & n8086 ;
  assign n8088 = \sram_data_i[27]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8089 = ~n8087 & ~n8088 ;
  assign n8090 = ~n8085 & n8089 ;
  assign n8091 = \u1_u2_rx_data_st_r_reg[4]/P0001  & n8084 ;
  assign n8092 = \u1_u2_dtmp_r_reg[28]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8093 = ~n8066 & n8092 ;
  assign n8094 = \sram_data_i[28]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8095 = ~n8093 & ~n8094 ;
  assign n8096 = ~n8091 & n8095 ;
  assign n8097 = \u1_u2_rx_data_st_r_reg[5]/P0001  & n8084 ;
  assign n8098 = \u1_u2_dtmp_r_reg[29]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8099 = ~n8066 & n8098 ;
  assign n8100 = \sram_data_i[29]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8101 = ~n8099 & ~n8100 ;
  assign n8102 = ~n8097 & n8101 ;
  assign n8103 = \u1_u2_rx_data_st_r_reg[6]/P0001  & n8084 ;
  assign n8104 = \u1_u2_dtmp_r_reg[30]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8105 = ~n8066 & n8104 ;
  assign n8106 = \sram_data_i[30]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8107 = ~n8105 & ~n8106 ;
  assign n8108 = ~n8103 & n8107 ;
  assign n8109 = \u1_u2_rx_data_st_r_reg[7]/P0001  & n8084 ;
  assign n8110 = \u1_u2_dtmp_r_reg[31]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8111 = ~n8066 & n8110 ;
  assign n8112 = \sram_data_i[31]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8113 = ~n8111 & ~n8112 ;
  assign n8114 = ~n8109 & n8113 ;
  assign n8115 = ~\u1_u2_adr_cb_reg[1]/NET0131  & n8064 ;
  assign n8116 = \u1_u2_dtmp_r_reg[8]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8117 = ~n7966 & n8116 ;
  assign n8118 = ~n8115 & ~n8117 ;
  assign n8119 = \sram_data_i[8]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8120 = n8118 & ~n8119 ;
  assign n8121 = n7964 & n8016 ;
  assign n8122 = \u1_u2_dtmp_r_reg[9]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8123 = ~n7966 & n8122 ;
  assign n8124 = ~n8121 & ~n8123 ;
  assign n8125 = \sram_data_i[9]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8126 = n8124 & ~n8125 ;
  assign n8127 = ~\u1_u2_adr_cb_reg[0]/NET0131  & ~\u1_u2_adr_cb_reg[1]/NET0131  ;
  assign n8128 = n8008 & n8127 ;
  assign n8129 = \u1_u2_rx_data_valid_r_reg/NET0131  & n8127 ;
  assign n8130 = \u1_u2_dtmp_r_reg[0]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8131 = ~n8129 & n8130 ;
  assign n8132 = ~n8128 & ~n8131 ;
  assign n8133 = \sram_data_i[0]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8134 = n8132 & ~n8133 ;
  assign n8135 = n8017 & n8127 ;
  assign n8136 = \u1_u2_dtmp_r_reg[1]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8137 = ~n8129 & n8136 ;
  assign n8138 = ~n8135 & ~n8137 ;
  assign n8139 = \sram_data_i[1]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8140 = n8138 & ~n8139 ;
  assign n8141 = n8024 & n8127 ;
  assign n8142 = \u1_u2_dtmp_r_reg[2]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8143 = ~n8129 & n8142 ;
  assign n8144 = ~n8141 & ~n8143 ;
  assign n8145 = \sram_data_i[2]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8146 = n8144 & ~n8145 ;
  assign n8147 = n8031 & n8127 ;
  assign n8148 = \u1_u2_rx_data_st_r_reg[3]/P0001  & n8147 ;
  assign n8149 = \u1_u2_dtmp_r_reg[3]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8150 = ~n8129 & n8149 ;
  assign n8151 = ~n8148 & ~n8150 ;
  assign n8152 = \sram_data_i[3]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8153 = n8151 & ~n8152 ;
  assign n8154 = \u1_u2_rx_data_st_r_reg[4]/P0001  & n8147 ;
  assign n8155 = \u1_u2_dtmp_r_reg[4]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8156 = ~n8129 & n8155 ;
  assign n8157 = ~n8154 & ~n8156 ;
  assign n8158 = \sram_data_i[4]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8159 = n8157 & ~n8158 ;
  assign n8160 = \u1_u2_rx_data_st_r_reg[5]/P0001  & n8147 ;
  assign n8161 = \u1_u2_dtmp_r_reg[5]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8162 = ~n8129 & n8161 ;
  assign n8163 = ~n8160 & ~n8162 ;
  assign n8164 = \sram_data_i[5]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8165 = n8163 & ~n8164 ;
  assign n8166 = \u1_u2_rx_data_st_r_reg[6]/P0001  & n8147 ;
  assign n8167 = \u1_u2_dtmp_r_reg[6]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8168 = ~n8129 & n8167 ;
  assign n8169 = ~n8166 & ~n8168 ;
  assign n8170 = \sram_data_i[6]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8171 = n8169 & ~n8170 ;
  assign n8172 = \u1_u2_rx_data_st_r_reg[7]/P0001  & n8147 ;
  assign n8173 = \u1_u2_dtmp_r_reg[7]/P0001  & ~\u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8174 = ~n8129 & n8173 ;
  assign n8175 = ~n8172 & ~n8174 ;
  assign n8176 = \sram_data_i[7]_pad  & \u1_u2_dtmp_sel_r_reg/P0001  ;
  assign n8177 = n8175 & ~n8176 ;
  assign n8178 = ~\u1_u3_abort_reg/P0001  & n4106 ;
  assign n8179 = n4103 & ~n8178 ;
  assign n8180 = ~\u1_u2_mack_r_reg/P0001  & ~n8179 ;
  assign n8181 = \u5_state_reg[0]/P0001  & n2558 ;
  assign n8182 = n2557 & n8181 ;
  assign n8183 = \u5_wb_req_s1_reg/P0001  & \wb_addr_i[17]_pad  ;
  assign n8184 = n8182 & n8183 ;
  assign n8185 = ~\u5_state_reg[0]/P0001  & ~\u5_state_reg[5]/NET0131  ;
  assign n8186 = n7956 & n8185 ;
  assign n8187 = \u5_state_reg[1]/P0001  & \u5_state_reg[2]/P0001  ;
  assign n8188 = ~n2558 & ~n8187 ;
  assign n8189 = n8186 & n8188 ;
  assign n8190 = ~\u2_wack_r_reg/P0001  & n8189 ;
  assign n8191 = ~n8184 & ~n8190 ;
  assign n8192 = ~\u1_u2_word_done_r_reg/P0001  & ~n8191 ;
  assign n8193 = ~n8180 & n8192 ;
  assign n8194 = rst_i_pad & ~\u2_wack_r_reg/P0001  ;
  assign n8195 = n8193 & n8194 ;
  assign n8196 = ~n4451 & ~n4456 ;
  assign n8197 = n4437 & ~n8196 ;
  assign n8198 = n4444 & ~n8196 ;
  assign n8199 = ~n4442 & n8198 ;
  assign n8200 = ~n8197 & ~n8199 ;
  assign n8201 = ~n4437 & n8196 ;
  assign n8202 = ~n4445 & n8201 ;
  assign n8203 = n8200 & ~n8202 ;
  assign n8204 = ~n4437 & ~n4456 ;
  assign n8205 = ~n4445 & n8204 ;
  assign n8206 = ~n4450 & ~n4455 ;
  assign n8207 = ~n4451 & ~n8206 ;
  assign n8208 = ~n8205 & n8207 ;
  assign n8209 = n4451 & n8206 ;
  assign n8210 = ~n4456 & n8206 ;
  assign n8211 = ~n4437 & n8210 ;
  assign n8212 = ~n4445 & n8211 ;
  assign n8213 = ~n8209 & ~n8212 ;
  assign n8214 = ~n8208 & n8213 ;
  assign n8215 = ~n4448 & ~n4466 ;
  assign n8216 = ~n4458 & n8215 ;
  assign n8217 = n4452 & n8215 ;
  assign n8218 = ~n4446 & n8217 ;
  assign n8219 = ~n8216 & ~n8218 ;
  assign n8220 = n4437 & n4452 ;
  assign n8221 = n4444 & n4452 ;
  assign n8222 = ~n4442 & n8221 ;
  assign n8223 = ~n8220 & ~n8222 ;
  assign n8224 = n4458 & ~n8215 ;
  assign n8225 = n8223 & n8224 ;
  assign n8226 = n8219 & ~n8225 ;
  assign n8227 = ~n4447 & ~n4465 ;
  assign n8228 = n4466 & n8227 ;
  assign n8229 = ~n4448 & n8227 ;
  assign n8230 = ~n4539 & n8229 ;
  assign n8231 = ~n4538 & n8230 ;
  assign n8232 = ~n8228 & ~n8231 ;
  assign n8233 = ~n4448 & ~n4539 ;
  assign n8234 = ~n4538 & n8233 ;
  assign n8235 = ~n4466 & ~n8227 ;
  assign n8236 = ~n8234 & n8235 ;
  assign n8237 = n8232 & ~n8236 ;
  assign n8238 = \u5_state_reg[2]/P0001  & ~\u5_wb_req_s1_reg/P0001  ;
  assign n8239 = rst_i_pad & n8238 ;
  assign n8240 = rst_i_pad & ~wb_we_i_pad ;
  assign n8241 = n8183 & n8240 ;
  assign n8242 = ~n8239 & ~n8241 ;
  assign n8243 = n8182 & ~n8242 ;
  assign n8244 = ~\u1_u2_word_done_r_reg/P0001  & \u2_wack_r_reg/P0001  ;
  assign n8245 = ~\u5_state_reg[1]/P0001  & \u5_state_reg[2]/P0001  ;
  assign n8246 = rst_i_pad & n8245 ;
  assign n8247 = n8186 & n8246 ;
  assign n8248 = ~n8244 & n8247 ;
  assign n8249 = ~\u1_u2_mack_r_reg/P0001  & n8247 ;
  assign n8250 = ~n8179 & n8249 ;
  assign n8251 = ~n8248 & ~n8250 ;
  assign n8252 = ~n8243 & n8251 ;
  assign n8253 = ~n6267 & ~n6286 ;
  assign n8254 = n6263 & n8253 ;
  assign n8255 = ~n6260 & n8254 ;
  assign n8256 = ~n6256 & n8255 ;
  assign n8257 = \u4_u3_dma_in_cnt_reg[7]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n8258 = ~n6277 & n8257 ;
  assign n8259 = ~\u4_u3_dma_in_cnt_reg[7]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n8260 = n6277 & n8259 ;
  assign n8261 = ~n8258 & ~n8260 ;
  assign n8262 = n6269 & n8253 ;
  assign n8263 = n8261 & ~n8262 ;
  assign n8264 = ~n8256 & n8263 ;
  assign n8265 = ~n6269 & ~n8253 ;
  assign n8266 = ~n6265 & n8265 ;
  assign n8267 = n6598 & ~n8266 ;
  assign n8268 = n8264 & n8267 ;
  assign n8269 = ~\u4_u3_dma_in_cnt_reg[7]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n8270 = n6281 & n8269 ;
  assign n8271 = ~\u4_u3_dma_in_cnt_reg[7]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n8272 = ~\u4_u3_r5_reg/NET0131  & ~n8271 ;
  assign n8273 = ~n8270 & n8272 ;
  assign n8274 = n8261 & ~n8273 ;
  assign n8275 = \u4_u3_csr1_reg[0]/P0001  & ~n8274 ;
  assign n8276 = ~n8268 & n8275 ;
  assign n8277 = ~n6325 & ~n6343 ;
  assign n8278 = ~n6327 & ~n8277 ;
  assign n8279 = ~n6323 & n8278 ;
  assign n8280 = n6632 & ~n8279 ;
  assign n8281 = n6321 & n8277 ;
  assign n8282 = ~n6318 & n8281 ;
  assign n8283 = ~n6314 & n8282 ;
  assign n8284 = \u4_u0_dma_in_cnt_reg[7]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n8285 = ~n6335 & n8284 ;
  assign n8286 = ~\u4_u0_dma_in_cnt_reg[7]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n8287 = n6335 & n8286 ;
  assign n8288 = ~n8285 & ~n8287 ;
  assign n8289 = n6327 & n8277 ;
  assign n8290 = n8288 & ~n8289 ;
  assign n8291 = ~n8283 & n8290 ;
  assign n8292 = n8280 & n8291 ;
  assign n8293 = ~\u4_u0_dma_in_cnt_reg[7]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n8294 = n6281 & n8293 ;
  assign n8295 = ~\u4_u0_dma_in_cnt_reg[7]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n8296 = ~\u4_u0_r5_reg/NET0131  & ~n8295 ;
  assign n8297 = ~n8294 & n8296 ;
  assign n8298 = n8288 & ~n8297 ;
  assign n8299 = \u4_u0_csr1_reg[0]/P0001  & ~n8298 ;
  assign n8300 = ~n8292 & n8299 ;
  assign n8301 = \u4_u1_dma_in_cnt_reg[7]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n8302 = ~n6362 & n8301 ;
  assign n8303 = ~\u4_u1_dma_in_cnt_reg[7]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n8304 = n6362 & n8303 ;
  assign n8305 = ~n8302 & ~n8304 ;
  assign n8306 = ~n6372 & ~n6403 ;
  assign n8307 = n6654 & ~n8306 ;
  assign n8308 = ~n6653 & n8307 ;
  assign n8309 = n6378 & ~n8306 ;
  assign n8310 = n6369 & ~n8309 ;
  assign n8311 = ~n8308 & n8310 ;
  assign n8312 = ~n6403 & n6656 ;
  assign n8313 = ~n6655 & n8312 ;
  assign n8314 = n8311 & ~n8313 ;
  assign n8315 = n8305 & n8314 ;
  assign n8316 = ~\u4_u1_dma_in_cnt_reg[7]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n8317 = n6281 & n8316 ;
  assign n8318 = ~\u4_u1_dma_in_cnt_reg[7]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n8319 = ~\u4_u1_r5_reg/NET0131  & ~n8318 ;
  assign n8320 = ~n8317 & n8319 ;
  assign n8321 = n8305 & ~n8320 ;
  assign n8322 = \u4_u1_csr1_reg[0]/P0001  & ~n8321 ;
  assign n8323 = ~n8315 & n8322 ;
  assign n8324 = n6443 & n6446 ;
  assign n8325 = ~n6426 & ~n6451 ;
  assign n8326 = ~n8324 & n8325 ;
  assign n8327 = ~n6422 & ~n6450 ;
  assign n8328 = ~n6425 & n8327 ;
  assign n8329 = ~n8326 & n8328 ;
  assign n8330 = ~n6451 & ~n8327 ;
  assign n8331 = ~n6426 & n8330 ;
  assign n8332 = ~n8324 & n8331 ;
  assign n8333 = \u4_u2_dma_in_cnt_reg[7]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n8334 = ~n6463 & n8333 ;
  assign n8335 = ~\u4_u2_dma_in_cnt_reg[7]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n8336 = n6463 & n8335 ;
  assign n8337 = ~n8334 & ~n8336 ;
  assign n8338 = n6425 & ~n8327 ;
  assign n8339 = n6667 & ~n8338 ;
  assign n8340 = n8337 & n8339 ;
  assign n8341 = ~n8332 & n8340 ;
  assign n8342 = ~n8329 & n8341 ;
  assign n8343 = ~\u4_u2_dma_in_cnt_reg[7]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n8344 = n6281 & n8343 ;
  assign n8345 = ~\u4_u2_dma_in_cnt_reg[7]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n8346 = ~\u4_u2_r5_reg/NET0131  & ~n8345 ;
  assign n8347 = ~n8344 & n8346 ;
  assign n8348 = n8337 & ~n8347 ;
  assign n8349 = \u4_u2_csr1_reg[0]/P0001  & ~n8348 ;
  assign n8350 = ~n8342 & n8349 ;
  assign n8351 = \u4_u3_csr1_reg[0]/P0001  & n6742 ;
  assign n8352 = n6741 & n8351 ;
  assign n8353 = \u4_u3_dma_out_cnt_reg[7]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n8354 = \u4_u3_csr1_reg[0]/P0001  & n8353 ;
  assign n8355 = ~n6741 & n8354 ;
  assign n8356 = ~n8352 & ~n8355 ;
  assign n8357 = ~\u4_u3_dma_out_cnt_reg[7]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n8358 = n6281 & n8357 ;
  assign n8359 = ~\u4_u3_dma_out_cnt_reg[7]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n8360 = n7524 & ~n8359 ;
  assign n8361 = ~n8358 & n8360 ;
  assign n8362 = n8356 & ~n8361 ;
  assign n8363 = n6759 & ~n6789 ;
  assign n8364 = n6784 & n8363 ;
  assign n8365 = n6778 & n6781 ;
  assign n8366 = ~n6758 & ~n6761 ;
  assign n8367 = ~n8365 & n8366 ;
  assign n8368 = ~n6757 & ~n6789 ;
  assign n8369 = ~n6760 & ~n8368 ;
  assign n8370 = ~n8367 & n8369 ;
  assign n8371 = ~n8364 & ~n8370 ;
  assign n8372 = n6598 & n8356 ;
  assign n8373 = n8371 & n8372 ;
  assign n8374 = ~n8362 & ~n8373 ;
  assign n8375 = \u4_u0_csr1_reg[0]/P0001  & n6806 ;
  assign n8376 = n6805 & n8375 ;
  assign n8377 = \u4_u0_dma_out_cnt_reg[7]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n8378 = \u4_u0_csr1_reg[0]/P0001  & n8377 ;
  assign n8379 = ~n6805 & n8378 ;
  assign n8380 = ~n8376 & ~n8379 ;
  assign n8381 = n6844 & n6847 ;
  assign n8382 = ~n6827 & ~n6852 ;
  assign n8383 = ~n8381 & n8382 ;
  assign n8384 = ~n6824 & ~n6851 ;
  assign n8385 = ~n6826 & ~n8384 ;
  assign n8386 = ~n8383 & n8385 ;
  assign n8387 = ~n6824 & n6853 ;
  assign n8388 = n6850 & n8387 ;
  assign n8389 = n6632 & ~n8388 ;
  assign n8390 = ~n8386 & n8389 ;
  assign n8391 = ~\u4_u0_dma_out_cnt_reg[7]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n8392 = n6281 & n8391 ;
  assign n8393 = ~\u4_u0_dma_out_cnt_reg[7]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n8394 = \u4_u0_csr1_reg[0]/P0001  & ~n8393 ;
  assign n8395 = ~n8392 & n8394 ;
  assign n8396 = ~\u4_u0_r5_reg/NET0131  & n8395 ;
  assign n8397 = ~n8390 & n8396 ;
  assign n8398 = n8380 & ~n8397 ;
  assign n8399 = \u4_u1_csr1_reg[0]/P0001  & n6870 ;
  assign n8400 = n6869 & n8399 ;
  assign n8401 = \u4_u1_dma_out_cnt_reg[7]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n8402 = \u4_u1_csr1_reg[0]/P0001  & n8401 ;
  assign n8403 = ~n6869 & n8402 ;
  assign n8404 = ~n8400 & ~n8403 ;
  assign n8405 = ~\u4_u1_dma_out_cnt_reg[7]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n8406 = n6281 & n8405 ;
  assign n8407 = ~\u4_u1_dma_out_cnt_reg[7]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n8408 = n6642 & ~n8407 ;
  assign n8409 = ~n8406 & n8408 ;
  assign n8410 = n8404 & ~n8409 ;
  assign n8411 = n6908 & n6911 ;
  assign n8412 = ~n6891 & ~n6916 ;
  assign n8413 = ~n8411 & n8412 ;
  assign n8414 = ~n6888 & ~n6915 ;
  assign n8415 = ~n6890 & ~n8414 ;
  assign n8416 = ~n8413 & n8415 ;
  assign n8417 = n6369 & ~n8416 ;
  assign n8418 = ~n6888 & n6917 ;
  assign n8419 = n6914 & n8418 ;
  assign n8420 = n8404 & ~n8419 ;
  assign n8421 = n8417 & n8420 ;
  assign n8422 = ~n8410 & ~n8421 ;
  assign n8423 = \u4_u2_csr1_reg[0]/P0001  & n6934 ;
  assign n8424 = n6933 & n8423 ;
  assign n8425 = \u4_u2_dma_out_cnt_reg[7]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n8426 = \u4_u2_csr1_reg[0]/P0001  & n8425 ;
  assign n8427 = ~n6933 & n8426 ;
  assign n8428 = ~n8424 & ~n8427 ;
  assign n8429 = n6971 & n6974 ;
  assign n8430 = ~n6951 & ~n6954 ;
  assign n8431 = ~n8429 & n8430 ;
  assign n8432 = ~n6950 & ~n6982 ;
  assign n8433 = ~n6953 & ~n8432 ;
  assign n8434 = ~n8431 & n8433 ;
  assign n8435 = n6952 & ~n6982 ;
  assign n8436 = n6977 & n8435 ;
  assign n8437 = n6667 & ~n8436 ;
  assign n8438 = ~n8434 & n8437 ;
  assign n8439 = ~\u4_u2_dma_out_cnt_reg[7]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n8440 = n6281 & n8439 ;
  assign n8441 = ~\u4_u2_dma_out_cnt_reg[7]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n8442 = \u4_u2_csr1_reg[0]/P0001  & ~n8441 ;
  assign n8443 = ~n8440 & n8442 ;
  assign n8444 = ~\u4_u2_r5_reg/NET0131  & n8443 ;
  assign n8445 = ~n8438 & n8444 ;
  assign n8446 = n8428 & ~n8445 ;
  assign n8447 = ~\u4_u3_r5_reg/NET0131  & ~n7307 ;
  assign n8448 = \u4_u3_ep_match_r_reg/P0001  & ~\u4_u3_r5_reg/NET0131  ;
  assign n8449 = ~n6282 & n8448 ;
  assign n8450 = \u4_u3_r5_reg/NET0131  & n7312 ;
  assign n8451 = n7309 & n8450 ;
  assign n8452 = ~n8449 & ~n8451 ;
  assign n8453 = \u4_u3_dma_out_cnt_reg[10]/P0001  & ~n8452 ;
  assign n8454 = ~n8447 & n8453 ;
  assign n8455 = ~\u4_u3_dma_out_cnt_reg[10]/P0001  & ~\u4_u3_r5_reg/NET0131  ;
  assign n8456 = ~n7307 & n8455 ;
  assign n8457 = ~\u4_u3_dma_out_cnt_reg[10]/P0001  & ~n8449 ;
  assign n8458 = ~n8451 & n8457 ;
  assign n8459 = \u4_u3_csr1_reg[0]/P0001  & ~n8458 ;
  assign n8460 = ~n8456 & n8459 ;
  assign n8461 = ~n8454 & n8460 ;
  assign n8462 = ~\u4_u0_r5_reg/NET0131  & ~n7357 ;
  assign n8463 = \u4_u0_ep_match_r_reg/P0001  & ~\u4_u0_r5_reg/NET0131  ;
  assign n8464 = ~n6339 & n8463 ;
  assign n8465 = \u4_u0_r5_reg/NET0131  & n7362 ;
  assign n8466 = n7359 & n8465 ;
  assign n8467 = ~n8464 & ~n8466 ;
  assign n8468 = \u4_u0_dma_out_cnt_reg[10]/P0001  & ~n8467 ;
  assign n8469 = ~n8462 & n8468 ;
  assign n8470 = ~\u4_u0_dma_out_cnt_reg[10]/P0001  & ~\u4_u0_r5_reg/NET0131  ;
  assign n8471 = ~n7357 & n8470 ;
  assign n8472 = ~\u4_u0_dma_out_cnt_reg[10]/P0001  & ~n8464 ;
  assign n8473 = ~n8466 & n8472 ;
  assign n8474 = \u4_u0_csr1_reg[0]/P0001  & ~n8473 ;
  assign n8475 = ~n8471 & n8474 ;
  assign n8476 = ~n8469 & n8475 ;
  assign n8477 = ~\u4_u1_r5_reg/NET0131  & ~n7407 ;
  assign n8478 = \u4_u1_ep_match_r_reg/P0001  & ~\u4_u1_r5_reg/NET0131  ;
  assign n8479 = ~n6368 & n8478 ;
  assign n8480 = \u4_u1_r5_reg/NET0131  & n7412 ;
  assign n8481 = n7409 & n8480 ;
  assign n8482 = ~n8479 & ~n8481 ;
  assign n8483 = \u4_u1_dma_out_cnt_reg[10]/P0001  & ~n8482 ;
  assign n8484 = ~n8477 & n8483 ;
  assign n8485 = ~\u4_u1_dma_out_cnt_reg[10]/P0001  & ~\u4_u1_r5_reg/NET0131  ;
  assign n8486 = ~n7407 & n8485 ;
  assign n8487 = ~\u4_u1_dma_out_cnt_reg[10]/P0001  & ~n8479 ;
  assign n8488 = ~n8481 & n8487 ;
  assign n8489 = \u4_u1_csr1_reg[0]/P0001  & ~n8488 ;
  assign n8490 = ~n8486 & n8489 ;
  assign n8491 = ~n8484 & n8490 ;
  assign n8492 = ~\u4_u2_r5_reg/NET0131  & ~n7457 ;
  assign n8493 = \u4_u2_ep_match_r_reg/P0001  & ~\u4_u2_r5_reg/NET0131  ;
  assign n8494 = ~n6415 & n8493 ;
  assign n8495 = \u4_u2_r5_reg/NET0131  & n7462 ;
  assign n8496 = n7459 & n8495 ;
  assign n8497 = ~n8494 & ~n8496 ;
  assign n8498 = \u4_u2_dma_out_cnt_reg[10]/P0001  & ~n8497 ;
  assign n8499 = ~n8492 & n8498 ;
  assign n8500 = ~\u4_u2_dma_out_cnt_reg[10]/P0001  & ~\u4_u2_r5_reg/NET0131  ;
  assign n8501 = ~n7457 & n8500 ;
  assign n8502 = ~\u4_u2_dma_out_cnt_reg[10]/P0001  & ~n8494 ;
  assign n8503 = ~n8496 & n8502 ;
  assign n8504 = \u4_u2_csr1_reg[0]/P0001  & ~n8503 ;
  assign n8505 = ~n8501 & n8504 ;
  assign n8506 = ~n8499 & n8505 ;
  assign n8507 = ~\u5_state_reg[2]/P0001  & n7957 ;
  assign n8508 = \u5_state_reg[3]/P0001  & n2556 ;
  assign n8509 = n8507 & n8508 ;
  assign n8510 = ~\u5_state_reg[4]/P0001  & ~n8509 ;
  assign n8511 = ~n8244 & n8510 ;
  assign n8512 = ~\u1_u2_mack_r_reg/P0001  & n8510 ;
  assign n8513 = ~n8179 & n8512 ;
  assign n8514 = ~n8511 & ~n8513 ;
  assign n8515 = ~n8189 & ~n8509 ;
  assign n8516 = rst_i_pad & ~n8515 ;
  assign n8517 = n8514 & n8516 ;
  assign n8518 = \u4_u3_dma_in_cnt_reg[4]/P0001  & \u4_u3_dma_in_cnt_reg[5]/P0001  ;
  assign n8519 = n6276 & n8518 ;
  assign n8520 = \u4_u3_r5_reg/NET0131  & ~n8519 ;
  assign n8521 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[5]/P0001  ;
  assign n8522 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[4]/P0001  ;
  assign n8523 = n6276 & n8522 ;
  assign n8524 = ~n8521 & ~n8523 ;
  assign n8525 = n8520 & ~n8524 ;
  assign n8526 = ~n6249 & ~n6259 ;
  assign n8527 = ~n6249 & n6254 ;
  assign n8528 = ~n6248 & n8527 ;
  assign n8529 = ~n8526 & ~n8528 ;
  assign n8530 = ~n6250 & ~n6262 ;
  assign n8531 = n6598 & n8530 ;
  assign n8532 = ~n8529 & n8531 ;
  assign n8533 = n6598 & ~n8530 ;
  assign n8534 = n8529 & n8533 ;
  assign n8535 = ~\u4_u3_dma_in_cnt_reg[5]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n8536 = n6281 & n8535 ;
  assign n8537 = ~\u4_u3_dma_in_cnt_reg[5]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n8538 = n7524 & ~n8537 ;
  assign n8539 = ~n8536 & n8538 ;
  assign n8540 = ~n8534 & n8539 ;
  assign n8541 = ~n8532 & n8540 ;
  assign n8542 = ~n8525 & ~n8541 ;
  assign n8543 = \u4_u0_dma_in_cnt_reg[4]/P0001  & \u4_u0_dma_in_cnt_reg[5]/P0001  ;
  assign n8544 = n6334 & n8543 ;
  assign n8545 = \u4_u0_r5_reg/NET0131  & ~n8544 ;
  assign n8546 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[5]/P0001  ;
  assign n8547 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[4]/P0001  ;
  assign n8548 = n6334 & n8547 ;
  assign n8549 = ~n8546 & ~n8548 ;
  assign n8550 = n8545 & ~n8549 ;
  assign n8551 = ~n6307 & ~n6317 ;
  assign n8552 = ~n6307 & n6312 ;
  assign n8553 = ~n6306 & n8552 ;
  assign n8554 = ~n8551 & ~n8553 ;
  assign n8555 = ~n6308 & ~n6320 ;
  assign n8556 = n6632 & n8555 ;
  assign n8557 = ~\u4_u0_dma_in_cnt_reg[5]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n8558 = n6281 & n8557 ;
  assign n8559 = ~\u4_u0_dma_in_cnt_reg[5]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n8560 = \u4_u0_csr1_reg[0]/P0001  & ~n8559 ;
  assign n8561 = ~n8558 & n8560 ;
  assign n8562 = ~n8556 & n8561 ;
  assign n8563 = ~n8554 & n8562 ;
  assign n8564 = n6632 & ~n8555 ;
  assign n8565 = n8561 & ~n8564 ;
  assign n8566 = n8554 & n8565 ;
  assign n8567 = ~n8563 & ~n8566 ;
  assign n8568 = ~\u4_u0_r5_reg/NET0131  & ~n8567 ;
  assign n8569 = ~n8550 & ~n8568 ;
  assign n8570 = \u4_u1_ep_match_r_reg/P0001  & ~n6398 ;
  assign n8571 = ~n6368 & n8570 ;
  assign n8572 = n6396 & n8571 ;
  assign n8573 = ~n6379 & ~n6397 ;
  assign n8574 = n6369 & n8573 ;
  assign n8575 = ~n8572 & ~n8574 ;
  assign n8576 = \u4_u1_dma_in_cnt_reg[4]/P0001  & n6361 ;
  assign n8577 = ~\u4_u1_dma_in_cnt_reg[5]/P0001  & ~n8576 ;
  assign n8578 = \u4_u1_dma_in_cnt_reg[4]/P0001  & \u4_u1_dma_in_cnt_reg[5]/P0001  ;
  assign n8579 = n6361 & n8578 ;
  assign n8580 = \u4_u1_r5_reg/NET0131  & ~n8579 ;
  assign n8581 = ~n8577 & n8580 ;
  assign n8582 = ~n6379 & n6399 ;
  assign n8583 = n6396 & n8582 ;
  assign n8584 = ~n8581 & ~n8583 ;
  assign n8585 = ~n8575 & n8584 ;
  assign n8586 = ~\u4_u1_dma_in_cnt_reg[5]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n8587 = n6281 & n8586 ;
  assign n8588 = ~\u4_u1_dma_in_cnt_reg[5]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n8589 = ~\u4_u1_r5_reg/NET0131  & ~n8588 ;
  assign n8590 = ~n8587 & n8589 ;
  assign n8591 = ~n8581 & ~n8590 ;
  assign n8592 = \u4_u1_csr1_reg[0]/P0001  & ~n8591 ;
  assign n8593 = ~n8585 & n8592 ;
  assign n8594 = ~n6426 & ~n6444 ;
  assign n8595 = n6667 & n8594 ;
  assign n8596 = \u4_u2_ep_match_r_reg/P0001  & ~n6445 ;
  assign n8597 = ~n6415 & n8596 ;
  assign n8598 = n6443 & n8597 ;
  assign n8599 = ~n8595 & ~n8598 ;
  assign n8600 = \u4_u2_dma_in_cnt_reg[4]/P0001  & n6462 ;
  assign n8601 = ~\u4_u2_dma_in_cnt_reg[5]/P0001  & ~n8600 ;
  assign n8602 = \u4_u2_dma_in_cnt_reg[4]/P0001  & \u4_u2_dma_in_cnt_reg[5]/P0001  ;
  assign n8603 = n6462 & n8602 ;
  assign n8604 = \u4_u2_r5_reg/NET0131  & ~n8603 ;
  assign n8605 = ~n8601 & n8604 ;
  assign n8606 = ~n6445 & n8594 ;
  assign n8607 = n6443 & n8606 ;
  assign n8608 = ~n8605 & ~n8607 ;
  assign n8609 = ~n8599 & n8608 ;
  assign n8610 = ~\u4_u2_dma_in_cnt_reg[5]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n8611 = n6281 & n8610 ;
  assign n8612 = ~\u4_u2_dma_in_cnt_reg[5]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n8613 = ~\u4_u2_r5_reg/NET0131  & ~n8612 ;
  assign n8614 = ~n8611 & n8613 ;
  assign n8615 = ~n8605 & ~n8614 ;
  assign n8616 = \u4_u2_csr1_reg[0]/P0001  & ~n8615 ;
  assign n8617 = ~n8609 & n8616 ;
  assign n8618 = \u5_state_reg[4]/P0001  & ~\u5_state_reg[5]/NET0131  ;
  assign n8619 = rst_i_pad & n8618 ;
  assign n8620 = ~\u5_state_reg[2]/P0001  & ~\u5_state_reg[3]/P0001  ;
  assign n8621 = n7957 & n8620 ;
  assign n8622 = n8619 & n8621 ;
  assign n8623 = \u1_u2_rx_data_valid_r_reg/NET0131  & \u1_u2_sizu_c_reg[0]/P0001  ;
  assign n8624 = \u1_u2_sizu_c_reg[1]/P0001  & n8623 ;
  assign n8625 = ~\u1_u2_sizu_c_reg[2]/P0001  & ~n8624 ;
  assign n8626 = ~n7011 & n7018 ;
  assign n8627 = ~n8625 & n8626 ;
  assign n8628 = \u1_u2_sizu_c_reg[3]/P0001  & n7018 ;
  assign n8629 = ~n7011 & n8628 ;
  assign n8630 = ~\u1_u2_sizu_c_reg[3]/P0001  & n7018 ;
  assign n8631 = \u1_u2_sizu_c_reg[1]/P0001  & \u1_u2_sizu_c_reg[2]/P0001  ;
  assign n8632 = n8623 & n8631 ;
  assign n8633 = n8630 & n8632 ;
  assign n8634 = ~n8629 & ~n8633 ;
  assign n8635 = \u1_u2_sizu_c_reg[3]/P0001  & n7011 ;
  assign n8636 = ~\u1_u2_sizu_c_reg[4]/P0001  & ~n8635 ;
  assign n8637 = \u1_u2_sizu_c_reg[3]/P0001  & \u1_u2_sizu_c_reg[4]/P0001  ;
  assign n8638 = n8632 & n8637 ;
  assign n8639 = n7018 & ~n8638 ;
  assign n8640 = ~n8636 & n8639 ;
  assign n8641 = ~\u1_u2_sizu_c_reg[5]/P0001  & ~n8638 ;
  assign n8642 = ~n7014 & n7018 ;
  assign n8643 = ~n8641 & n8642 ;
  assign n8644 = \u1_u2_sizu_c_reg[6]/P0001  & n7018 ;
  assign n8645 = ~n7014 & n8644 ;
  assign n8646 = ~\u1_u2_sizu_c_reg[6]/P0001  & n7018 ;
  assign n8647 = n7014 & n8646 ;
  assign n8648 = ~n8645 & ~n8647 ;
  assign n8649 = \u1_u2_sizu_c_reg[4]/P0001  & \u1_u2_sizu_c_reg[6]/P0001  ;
  assign n8650 = n7012 & n8649 ;
  assign n8651 = n7011 & n8650 ;
  assign n8652 = ~\u1_u2_sizu_c_reg[7]/P0001  & ~n8651 ;
  assign n8653 = ~n7016 & ~n8652 ;
  assign n8654 = n7018 & n8653 ;
  assign n8655 = ~n7022 & n7947 ;
  assign n8656 = ~\u1_u2_sizu_c_reg[9]/P0001  & n7018 ;
  assign n8657 = n7015 & n8656 ;
  assign n8658 = n7021 & n8657 ;
  assign n8659 = ~n8655 & ~n8658 ;
  assign n8660 = \u0_u0_state_reg[8]/NET0131  & ~\u0_u0_state_reg[9]/P0001  ;
  assign n8661 = n5753 & n8660 ;
  assign n8662 = n5735 & n8661 ;
  assign n8663 = n5746 & n8662 ;
  assign n8664 = ~n6133 & ~n6178 ;
  assign n8665 = n6132 & ~n8664 ;
  assign n8666 = n8663 & ~n8665 ;
  assign n8667 = n6178 & n6195 ;
  assign n8668 = \u0_u0_T1_gt_3_0_mS_reg/P0001  & ~\u0_u0_mode_hs_reg/P0001  ;
  assign n8669 = n6133 & n8668 ;
  assign n8670 = ~n6150 & n8669 ;
  assign n8671 = ~n8667 & ~n8670 ;
  assign n8672 = n6132 & ~n8671 ;
  assign n8673 = ~\u0_u0_idle_cnt1_clr_reg/P0001  & \u0_u0_idle_long_reg/P0001  ;
  assign n8674 = ~\u0_u0_T1_gt_5_0_mS_reg/P0001  & \u0_u0_ps_cnt_clr_reg/P0001  ;
  assign n8675 = ~\u0_u0_idle_cnt1_reg[4]/P0001  & ~n8674 ;
  assign n8676 = n8673 & ~n8675 ;
  assign n8677 = ~\u0_u0_idle_cnt1_next_reg[4]/P0001  & n8674 ;
  assign n8678 = n8676 & ~n8677 ;
  assign n8679 = ~n8672 & n8678 ;
  assign n8680 = ~n8666 & n8679 ;
  assign n8681 = \u4_u0_buf0_orig_reg[26]/P0001  & ~\u4_u0_dma_in_cnt_reg[7]/P0001  ;
  assign n8682 = \u4_u0_buf0_orig_reg[28]/P0001  & ~\u4_u0_dma_in_cnt_reg[9]/P0001  ;
  assign n8683 = \u4_u0_buf0_orig_reg[27]/P0001  & ~\u4_u0_dma_in_cnt_reg[8]/P0001  ;
  assign n8684 = ~n8682 & ~n8683 ;
  assign n8685 = ~n8681 & n8684 ;
  assign n8686 = ~\u4_u0_buf0_orig_reg[25]/P0001  & \u4_u0_dma_in_cnt_reg[6]/P0001  ;
  assign n8687 = ~\u4_u0_buf0_orig_reg[26]/P0001  & \u4_u0_dma_in_cnt_reg[7]/P0001  ;
  assign n8688 = ~n8686 & ~n8687 ;
  assign n8689 = n8685 & ~n8688 ;
  assign n8690 = ~\u4_u0_buf0_orig_reg[24]/P0001  & \u4_u0_dma_in_cnt_reg[5]/P0001  ;
  assign n8691 = ~\u4_u0_buf0_orig_reg[23]/P0001  & \u4_u0_dma_in_cnt_reg[4]/P0001  ;
  assign n8692 = ~n8690 & ~n8691 ;
  assign n8693 = \u4_u0_buf0_orig_reg[23]/P0001  & ~\u4_u0_dma_in_cnt_reg[4]/P0001  ;
  assign n8694 = \u4_u0_buf0_orig_reg[22]/P0001  & ~\u4_u0_dma_in_cnt_reg[3]/P0001  ;
  assign n8695 = ~n8693 & ~n8694 ;
  assign n8696 = n8692 & ~n8695 ;
  assign n8697 = \u4_u0_buf0_orig_reg[19]/P0001  & ~\u4_u0_dma_in_cnt_reg[0]/P0001  ;
  assign n8698 = \u4_u0_dma_in_cnt_reg[1]/P0001  & ~n8697 ;
  assign n8699 = \u4_u0_buf0_orig_reg[20]/P0001  & ~n8698 ;
  assign n8700 = \u4_u0_buf0_orig_reg[21]/P0001  & ~\u4_u0_dma_in_cnt_reg[2]/P0001  ;
  assign n8701 = ~\u4_u0_dma_in_cnt_reg[1]/P0001  & n8697 ;
  assign n8702 = ~n8700 & ~n8701 ;
  assign n8703 = ~n8699 & n8702 ;
  assign n8704 = ~\u4_u0_buf0_orig_reg[22]/P0001  & \u4_u0_dma_in_cnt_reg[3]/P0001  ;
  assign n8705 = ~\u4_u0_buf0_orig_reg[21]/P0001  & \u4_u0_dma_in_cnt_reg[2]/P0001  ;
  assign n8706 = ~n8704 & ~n8705 ;
  assign n8707 = n8692 & n8706 ;
  assign n8708 = ~n8703 & n8707 ;
  assign n8709 = ~n8696 & ~n8708 ;
  assign n8710 = \u4_u0_buf0_orig_reg[25]/P0001  & ~\u4_u0_dma_in_cnt_reg[6]/P0001  ;
  assign n8711 = \u4_u0_buf0_orig_reg[24]/P0001  & ~\u4_u0_dma_in_cnt_reg[5]/P0001  ;
  assign n8712 = ~n8710 & ~n8711 ;
  assign n8713 = n8685 & n8712 ;
  assign n8714 = n8709 & n8713 ;
  assign n8715 = ~n8689 & ~n8714 ;
  assign n8716 = \u4_u0_csr1_reg[11]/P0001  & ~\u4_u0_csr1_reg[12]/P0001  ;
  assign n8717 = ~\u4_u0_buf0_orig_reg[30]/NET0131  & \u4_u0_dma_in_cnt_reg[11]/P0001  ;
  assign n8718 = \u4_u0_csr1_reg[0]/P0001  & ~n8717 ;
  assign n8719 = n8716 & n8718 ;
  assign n8720 = ~\u4_u0_buf0_orig_reg[27]/P0001  & \u4_u0_dma_in_cnt_reg[8]/P0001  ;
  assign n8721 = ~n8682 & n8720 ;
  assign n8722 = ~\u4_u0_buf0_orig_reg[28]/P0001  & \u4_u0_dma_in_cnt_reg[9]/P0001  ;
  assign n8723 = ~\u4_u0_buf0_orig_reg[29]/NET0131  & \u4_u0_dma_in_cnt_reg[10]/P0001  ;
  assign n8724 = ~n8722 & ~n8723 ;
  assign n8725 = ~n8721 & n8724 ;
  assign n8726 = n8719 & n8725 ;
  assign n8727 = n8715 & n8726 ;
  assign n8728 = \u4_u0_buf0_orig_reg[30]/NET0131  & ~\u4_u0_dma_in_cnt_reg[11]/P0001  ;
  assign n8729 = \u4_u0_buf0_orig_reg[29]/NET0131  & ~\u4_u0_dma_in_cnt_reg[10]/P0001  ;
  assign n8730 = ~n8728 & ~n8729 ;
  assign n8731 = n8719 & ~n8730 ;
  assign n8732 = ~\u4_u0_dma_out_cnt_reg[10]/P0001  & ~\u4_u0_dma_out_cnt_reg[11]/P0001  ;
  assign n8733 = n6803 & n7358 ;
  assign n8734 = n8732 & n8733 ;
  assign n8735 = n6802 & n7362 ;
  assign n8736 = n8734 & n8735 ;
  assign n8737 = \u4_u0_csr1_reg[0]/P0001  & n4377 ;
  assign n8738 = ~n8736 & n8737 ;
  assign n8739 = ~n8731 & ~n8738 ;
  assign n8740 = ~n8727 & n8739 ;
  assign n8741 = ~\u4_u0_r2_reg/P0001  & ~\u4_u0_r4_reg/P0001  ;
  assign n8742 = ~\u4_u0_r5_reg/NET0131  & n8741 ;
  assign n8743 = ~n8740 & n8742 ;
  assign n8744 = \u4_u1_buf0_orig_reg[27]/P0001  & ~\u4_u1_dma_in_cnt_reg[8]/P0001  ;
  assign n8745 = \u4_u1_buf0_orig_reg[26]/P0001  & ~\u4_u1_dma_in_cnt_reg[7]/P0001  ;
  assign n8746 = ~n8744 & ~n8745 ;
  assign n8747 = ~\u4_u1_buf0_orig_reg[25]/P0001  & \u4_u1_dma_in_cnt_reg[6]/P0001  ;
  assign n8748 = ~\u4_u1_buf0_orig_reg[26]/P0001  & \u4_u1_dma_in_cnt_reg[7]/P0001  ;
  assign n8749 = ~n8747 & ~n8748 ;
  assign n8750 = n8746 & ~n8749 ;
  assign n8751 = ~\u4_u1_buf0_orig_reg[23]/P0001  & \u4_u1_dma_in_cnt_reg[4]/P0001  ;
  assign n8752 = ~\u4_u1_buf0_orig_reg[24]/P0001  & \u4_u1_dma_in_cnt_reg[5]/P0001  ;
  assign n8753 = ~n8751 & ~n8752 ;
  assign n8754 = \u4_u1_buf0_orig_reg[23]/P0001  & ~\u4_u1_dma_in_cnt_reg[4]/P0001  ;
  assign n8755 = \u4_u1_buf0_orig_reg[22]/P0001  & ~\u4_u1_dma_in_cnt_reg[3]/P0001  ;
  assign n8756 = ~n8754 & ~n8755 ;
  assign n8757 = n8753 & ~n8756 ;
  assign n8758 = \u4_u1_buf0_orig_reg[19]/P0001  & ~\u4_u1_dma_in_cnt_reg[0]/P0001  ;
  assign n8759 = ~\u4_u1_buf0_orig_reg[20]/P0001  & \u4_u1_dma_in_cnt_reg[1]/P0001  ;
  assign n8760 = n8758 & ~n8759 ;
  assign n8761 = \u4_u1_buf0_orig_reg[21]/P0001  & ~\u4_u1_dma_in_cnt_reg[2]/P0001  ;
  assign n8762 = \u4_u1_buf0_orig_reg[20]/P0001  & ~\u4_u1_dma_in_cnt_reg[1]/P0001  ;
  assign n8763 = ~n8761 & ~n8762 ;
  assign n8764 = ~n8760 & n8763 ;
  assign n8765 = ~\u4_u1_buf0_orig_reg[21]/P0001  & \u4_u1_dma_in_cnt_reg[2]/P0001  ;
  assign n8766 = ~\u4_u1_buf0_orig_reg[22]/P0001  & \u4_u1_dma_in_cnt_reg[3]/P0001  ;
  assign n8767 = ~n8765 & ~n8766 ;
  assign n8768 = n8753 & n8767 ;
  assign n8769 = ~n8764 & n8768 ;
  assign n8770 = ~n8757 & ~n8769 ;
  assign n8771 = \u4_u1_buf0_orig_reg[25]/P0001  & ~\u4_u1_dma_in_cnt_reg[6]/P0001  ;
  assign n8772 = \u4_u1_buf0_orig_reg[24]/P0001  & ~\u4_u1_dma_in_cnt_reg[5]/P0001  ;
  assign n8773 = ~n8771 & ~n8772 ;
  assign n8774 = n8746 & n8773 ;
  assign n8775 = n8770 & n8774 ;
  assign n8776 = ~n8750 & ~n8775 ;
  assign n8777 = ~\u4_u1_buf0_orig_reg[30]/NET0131  & \u4_u1_dma_in_cnt_reg[11]/P0001  ;
  assign n8778 = \u4_u1_csr1_reg[11]/P0001  & ~\u4_u1_csr1_reg[12]/P0001  ;
  assign n8779 = \u4_u1_csr1_reg[0]/P0001  & n8778 ;
  assign n8780 = ~n8777 & n8779 ;
  assign n8781 = \u4_u1_buf0_orig_reg[30]/NET0131  & ~\u4_u1_dma_in_cnt_reg[11]/P0001  ;
  assign n8782 = ~\u4_u1_buf0_orig_reg[29]/NET0131  & \u4_u1_dma_in_cnt_reg[10]/P0001  ;
  assign n8783 = ~n8781 & n8782 ;
  assign n8784 = ~\u4_u1_buf0_orig_reg[27]/P0001  & \u4_u1_dma_in_cnt_reg[8]/P0001  ;
  assign n8785 = ~\u4_u1_buf0_orig_reg[28]/P0001  & \u4_u1_dma_in_cnt_reg[9]/P0001  ;
  assign n8786 = ~n8784 & ~n8785 ;
  assign n8787 = ~n8783 & n8786 ;
  assign n8788 = n8780 & n8787 ;
  assign n8789 = n8776 & n8788 ;
  assign n8790 = \u4_u1_buf0_orig_reg[28]/P0001  & ~\u4_u1_dma_in_cnt_reg[9]/P0001  ;
  assign n8791 = \u4_u1_buf0_orig_reg[29]/NET0131  & ~\u4_u1_dma_in_cnt_reg[10]/P0001  ;
  assign n8792 = ~n8781 & ~n8791 ;
  assign n8793 = ~n8790 & n8792 ;
  assign n8794 = n8780 & ~n8793 ;
  assign n8795 = ~n8783 & n8794 ;
  assign n8796 = ~\u4_u1_dma_out_cnt_reg[10]/P0001  & ~\u4_u1_dma_out_cnt_reg[11]/P0001  ;
  assign n8797 = n6867 & n7408 ;
  assign n8798 = n8796 & n8797 ;
  assign n8799 = n6866 & n7412 ;
  assign n8800 = n8798 & n8799 ;
  assign n8801 = \u4_u1_csr1_reg[0]/P0001  & n4388 ;
  assign n8802 = ~n8800 & n8801 ;
  assign n8803 = ~n8795 & ~n8802 ;
  assign n8804 = ~n8789 & n8803 ;
  assign n8805 = ~\u4_u1_r2_reg/P0001  & ~\u4_u1_r4_reg/P0001  ;
  assign n8806 = ~\u4_u1_r5_reg/NET0131  & n8805 ;
  assign n8807 = ~n8804 & n8806 ;
  assign n8808 = n5080 & n7128 ;
  assign n8809 = ~\u1_u2_rx_data_valid_r_reg/NET0131  & ~\u1_u2_sizu_c_reg[0]/P0001  ;
  assign n8810 = n7018 & ~n8623 ;
  assign n8811 = ~n8809 & n8810 ;
  assign n8812 = ~\u1_u2_sizu_c_reg[1]/P0001  & ~n8623 ;
  assign n8813 = n7018 & ~n8624 ;
  assign n8814 = ~n8812 & n8813 ;
  assign n8815 = n2583 & n2584 ;
  assign n8816 = ~\wb_addr_i[2]_pad  & ~\wb_addr_i[3]_pad  ;
  assign n8817 = \u4_u0_csr0_reg[0]/P0001  & n8816 ;
  assign n8818 = \u4_u0_buf1_reg[0]/P0001  & n2731 ;
  assign n8819 = ~n8817 & ~n8818 ;
  assign n8820 = \wb_addr_i[2]_pad  & ~\wb_addr_i[3]_pad  ;
  assign n8821 = \u4_u0_int_stat_reg[0]/P0001  & n8820 ;
  assign n8822 = \u4_u0_buf0_reg[0]/P0001  & n2568 ;
  assign n8823 = ~n8821 & ~n8822 ;
  assign n8824 = n8819 & n8823 ;
  assign n8825 = n8815 & ~n8824 ;
  assign n8826 = n2563 & n2583 ;
  assign n8827 = \u4_u2_buf0_reg[0]/P0001  & n2568 ;
  assign n8828 = \u4_u2_csr0_reg[0]/P0001  & n8816 ;
  assign n8829 = ~n8827 & ~n8828 ;
  assign n8830 = \u4_u2_buf1_reg[0]/P0001  & n2731 ;
  assign n8831 = \u4_u2_int_stat_reg[0]/P0001  & n8820 ;
  assign n8832 = ~n8830 & ~n8831 ;
  assign n8833 = n8829 & n8832 ;
  assign n8834 = n8826 & ~n8833 ;
  assign n8835 = ~n8825 & ~n8834 ;
  assign n8836 = n2562 & n2563 ;
  assign n8837 = \u4_u3_csr0_reg[0]/P0001  & n8816 ;
  assign n8838 = \u4_u3_buf1_reg[0]/P0001  & n2731 ;
  assign n8839 = ~n8837 & ~n8838 ;
  assign n8840 = \u4_u3_int_stat_reg[0]/P0001  & n8820 ;
  assign n8841 = \u4_u3_buf0_reg[0]/P0001  & n2568 ;
  assign n8842 = ~n8840 & ~n8841 ;
  assign n8843 = n8839 & n8842 ;
  assign n8844 = n8836 & ~n8843 ;
  assign n8845 = n8835 & ~n8844 ;
  assign n8846 = \u4_funct_adr_reg[0]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8847 = n8820 & n8846 ;
  assign n8848 = \u0_u0_usb_suspend_reg/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8849 = n8816 & n8848 ;
  assign n8850 = ~n8847 & ~n8849 ;
  assign n8851 = \u4_int_srca_reg[0]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8852 = n2731 & n8851 ;
  assign n8853 = n8850 & ~n8852 ;
  assign n8854 = \u4_inta_msk_reg[0]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8855 = n2568 & n8854 ;
  assign n8856 = \u1_sof_time_reg[0]/P0001  & \wb_addr_i[4]_pad  ;
  assign n8857 = n8816 & n8856 ;
  assign n8858 = ~n8855 & ~n8857 ;
  assign n8859 = \u4_utmi_vend_stat_r_reg[0]/P0001  & \wb_addr_i[4]_pad  ;
  assign n8860 = n8820 & n8859 ;
  assign n8861 = n8858 & ~n8860 ;
  assign n8862 = n8853 & n8861 ;
  assign n8863 = ~\wb_addr_i[5]_pad  & ~\wb_addr_i[6]_pad  ;
  assign n8864 = n2561 & n8863 ;
  assign n8865 = ~n8862 & n8864 ;
  assign n8866 = n2562 & n2584 ;
  assign n8867 = \u4_u1_csr0_reg[0]/P0001  & n8816 ;
  assign n8868 = \u4_u1_buf1_reg[0]/P0001  & n2731 ;
  assign n8869 = ~n8867 & ~n8868 ;
  assign n8870 = \u4_u1_int_stat_reg[0]/P0001  & n8820 ;
  assign n8871 = \u4_u1_buf0_reg[0]/P0001  & n2568 ;
  assign n8872 = ~n8870 & ~n8871 ;
  assign n8873 = n8869 & n8872 ;
  assign n8874 = n8866 & ~n8873 ;
  assign n8875 = ~n8865 & ~n8874 ;
  assign n8876 = n8845 & n8875 ;
  assign n8877 = \u4_u0_csr0_reg[1]/P0001  & n8816 ;
  assign n8878 = \u4_u0_buf1_reg[1]/P0001  & n2731 ;
  assign n8879 = ~n8877 & ~n8878 ;
  assign n8880 = \u4_u0_int_stat_reg[1]/P0001  & n8820 ;
  assign n8881 = \u4_u0_buf0_reg[1]/P0001  & n2568 ;
  assign n8882 = ~n8880 & ~n8881 ;
  assign n8883 = n8879 & n8882 ;
  assign n8884 = n8815 & ~n8883 ;
  assign n8885 = \u4_u3_buf0_reg[1]/P0001  & n2568 ;
  assign n8886 = \u4_u3_csr0_reg[1]/P0001  & n8816 ;
  assign n8887 = ~n8885 & ~n8886 ;
  assign n8888 = \u4_u3_buf1_reg[1]/P0001  & n2731 ;
  assign n8889 = \u4_u3_int_stat_reg[1]/P0001  & n8820 ;
  assign n8890 = ~n8888 & ~n8889 ;
  assign n8891 = n8887 & n8890 ;
  assign n8892 = n8836 & ~n8891 ;
  assign n8893 = ~n8884 & ~n8892 ;
  assign n8894 = \u4_u2_csr0_reg[1]/P0001  & n8816 ;
  assign n8895 = \u4_u2_buf1_reg[1]/P0001  & n2731 ;
  assign n8896 = ~n8894 & ~n8895 ;
  assign n8897 = \u4_u2_int_stat_reg[1]/P0001  & n8820 ;
  assign n8898 = \u4_u2_buf0_reg[1]/P0001  & n2568 ;
  assign n8899 = ~n8897 & ~n8898 ;
  assign n8900 = n8896 & n8899 ;
  assign n8901 = n8826 & ~n8900 ;
  assign n8902 = n8893 & ~n8901 ;
  assign n8903 = \u4_funct_adr_reg[1]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8904 = n8820 & n8903 ;
  assign n8905 = \u0_u0_mode_hs_reg/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8906 = n8816 & n8905 ;
  assign n8907 = ~n8904 & ~n8906 ;
  assign n8908 = \u4_int_srca_reg[1]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8909 = n2731 & n8908 ;
  assign n8910 = n8907 & ~n8909 ;
  assign n8911 = \u4_inta_msk_reg[1]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8912 = n2568 & n8911 ;
  assign n8913 = \u1_sof_time_reg[1]/P0001  & \wb_addr_i[4]_pad  ;
  assign n8914 = n8816 & n8913 ;
  assign n8915 = ~n8912 & ~n8914 ;
  assign n8916 = \u4_utmi_vend_stat_r_reg[1]/P0001  & \wb_addr_i[4]_pad  ;
  assign n8917 = n8820 & n8916 ;
  assign n8918 = n8915 & ~n8917 ;
  assign n8919 = n8910 & n8918 ;
  assign n8920 = n8864 & ~n8919 ;
  assign n8921 = \u4_u1_csr0_reg[1]/P0001  & n8816 ;
  assign n8922 = \u4_u1_buf1_reg[1]/P0001  & n2731 ;
  assign n8923 = ~n8921 & ~n8922 ;
  assign n8924 = \u4_u1_int_stat_reg[1]/P0001  & n8820 ;
  assign n8925 = \u4_u1_buf0_reg[1]/P0001  & n2568 ;
  assign n8926 = ~n8924 & ~n8925 ;
  assign n8927 = n8923 & n8926 ;
  assign n8928 = n8866 & ~n8927 ;
  assign n8929 = ~n8920 & ~n8928 ;
  assign n8930 = n8902 & n8929 ;
  assign n8931 = \u4_u0_csr0_reg[2]/P0001  & n8816 ;
  assign n8932 = \u4_u0_buf1_reg[2]/P0001  & n2731 ;
  assign n8933 = ~n8931 & ~n8932 ;
  assign n8934 = \u4_u0_int_stat_reg[2]/P0001  & n8820 ;
  assign n8935 = \u4_u0_buf0_reg[2]/P0001  & n2568 ;
  assign n8936 = ~n8934 & ~n8935 ;
  assign n8937 = n8933 & n8936 ;
  assign n8938 = n8815 & ~n8937 ;
  assign n8939 = \u4_u3_buf0_reg[2]/P0001  & n2568 ;
  assign n8940 = \u4_u3_csr0_reg[2]/P0001  & n8816 ;
  assign n8941 = ~n8939 & ~n8940 ;
  assign n8942 = \u4_u3_buf1_reg[2]/P0001  & n2731 ;
  assign n8943 = \u4_u3_int_stat_reg[2]/P0001  & n8820 ;
  assign n8944 = ~n8942 & ~n8943 ;
  assign n8945 = n8941 & n8944 ;
  assign n8946 = n8836 & ~n8945 ;
  assign n8947 = ~n8938 & ~n8946 ;
  assign n8948 = \u4_u2_csr0_reg[2]/P0001  & n8816 ;
  assign n8949 = \u4_u2_buf1_reg[2]/P0001  & n2731 ;
  assign n8950 = ~n8948 & ~n8949 ;
  assign n8951 = \u4_u2_int_stat_reg[2]/P0001  & n8820 ;
  assign n8952 = \u4_u2_buf0_reg[2]/P0001  & n2568 ;
  assign n8953 = ~n8951 & ~n8952 ;
  assign n8954 = n8950 & n8953 ;
  assign n8955 = n8826 & ~n8954 ;
  assign n8956 = n8947 & ~n8955 ;
  assign n8957 = \u4_funct_adr_reg[2]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8958 = n8820 & n8957 ;
  assign n8959 = \u0_u0_usb_attached_reg/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8960 = n8816 & n8959 ;
  assign n8961 = ~n8958 & ~n8960 ;
  assign n8962 = \u4_int_srca_reg[2]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8963 = n2731 & n8962 ;
  assign n8964 = n8961 & ~n8963 ;
  assign n8965 = \u4_inta_msk_reg[2]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n8966 = n2568 & n8965 ;
  assign n8967 = \u1_sof_time_reg[2]/P0001  & \wb_addr_i[4]_pad  ;
  assign n8968 = n8816 & n8967 ;
  assign n8969 = ~n8966 & ~n8968 ;
  assign n8970 = \u4_utmi_vend_stat_r_reg[2]/P0001  & \wb_addr_i[4]_pad  ;
  assign n8971 = n8820 & n8970 ;
  assign n8972 = n8969 & ~n8971 ;
  assign n8973 = n8964 & n8972 ;
  assign n8974 = n8864 & ~n8973 ;
  assign n8975 = \u4_u1_csr0_reg[2]/P0001  & n8816 ;
  assign n8976 = \u4_u1_buf1_reg[2]/P0001  & n2731 ;
  assign n8977 = ~n8975 & ~n8976 ;
  assign n8978 = \u4_u1_int_stat_reg[2]/P0001  & n8820 ;
  assign n8979 = \u4_u1_buf0_reg[2]/P0001  & n2568 ;
  assign n8980 = ~n8978 & ~n8979 ;
  assign n8981 = n8977 & n8980 ;
  assign n8982 = n8866 & ~n8981 ;
  assign n8983 = ~n8974 & ~n8982 ;
  assign n8984 = n8956 & n8983 ;
  assign n8985 = \u4_u0_csr0_reg[3]/NET0131  & n8816 ;
  assign n8986 = \u4_u0_buf1_reg[3]/P0001  & n2731 ;
  assign n8987 = ~n8985 & ~n8986 ;
  assign n8988 = \u4_u0_int_stat_reg[3]/P0001  & n8820 ;
  assign n8989 = \u4_u0_buf0_reg[3]/P0001  & n2568 ;
  assign n8990 = ~n8988 & ~n8989 ;
  assign n8991 = n8987 & n8990 ;
  assign n8992 = n8815 & ~n8991 ;
  assign n8993 = \u4_u3_buf0_reg[3]/P0001  & n2568 ;
  assign n8994 = \u4_u3_csr0_reg[3]/NET0131  & n8816 ;
  assign n8995 = ~n8993 & ~n8994 ;
  assign n8996 = \u4_u3_buf1_reg[3]/P0001  & n2731 ;
  assign n8997 = \u4_u3_int_stat_reg[3]/P0001  & n8820 ;
  assign n8998 = ~n8996 & ~n8997 ;
  assign n8999 = n8995 & n8998 ;
  assign n9000 = n8836 & ~n8999 ;
  assign n9001 = ~n8992 & ~n9000 ;
  assign n9002 = \u4_u2_csr0_reg[3]/NET0131  & n8816 ;
  assign n9003 = \u4_u2_buf1_reg[3]/P0001  & n2731 ;
  assign n9004 = ~n9002 & ~n9003 ;
  assign n9005 = \u4_u2_int_stat_reg[3]/P0001  & n8820 ;
  assign n9006 = \u4_u2_buf0_reg[3]/P0001  & n2568 ;
  assign n9007 = ~n9005 & ~n9006 ;
  assign n9008 = n9004 & n9007 ;
  assign n9009 = n8826 & ~n9008 ;
  assign n9010 = n9001 & ~n9009 ;
  assign n9011 = \u4_funct_adr_reg[3]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n9012 = n8820 & n9011 ;
  assign n9013 = \u1_sof_time_reg[3]/P0001  & \wb_addr_i[4]_pad  ;
  assign n9014 = n8816 & n9013 ;
  assign n9015 = ~n9012 & ~n9014 ;
  assign n9016 = \u4_int_srca_reg[3]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n9017 = n2731 & n9016 ;
  assign n9018 = n9015 & ~n9017 ;
  assign n9019 = \u4_inta_msk_reg[3]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n9020 = n2568 & n9019 ;
  assign n9021 = \LineState_r_reg[0]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n9022 = n8816 & n9021 ;
  assign n9023 = ~n9020 & ~n9022 ;
  assign n9024 = \u4_utmi_vend_stat_r_reg[3]/P0001  & \wb_addr_i[4]_pad  ;
  assign n9025 = n8820 & n9024 ;
  assign n9026 = n9023 & ~n9025 ;
  assign n9027 = n9018 & n9026 ;
  assign n9028 = n8864 & ~n9027 ;
  assign n9029 = \u4_u1_csr0_reg[3]/NET0131  & n8816 ;
  assign n9030 = \u4_u1_buf1_reg[3]/P0001  & n2731 ;
  assign n9031 = ~n9029 & ~n9030 ;
  assign n9032 = \u4_u1_int_stat_reg[3]/P0001  & n8820 ;
  assign n9033 = \u4_u1_buf0_reg[3]/P0001  & n2568 ;
  assign n9034 = ~n9032 & ~n9033 ;
  assign n9035 = n9031 & n9034 ;
  assign n9036 = n8866 & ~n9035 ;
  assign n9037 = ~n9028 & ~n9036 ;
  assign n9038 = n9010 & n9037 ;
  assign n9039 = ~\u1_u0_pid_reg[2]/NET0131  & ~\u1_u3_this_dpid_reg[1]/P0001  ;
  assign n9040 = \u1_u0_pid_reg[2]/NET0131  & \u1_u3_this_dpid_reg[1]/P0001  ;
  assign n9041 = ~n9039 & ~n9040 ;
  assign n9042 = \u1_u0_pid_reg[0]/NET0131  & ~n9041 ;
  assign n9043 = ~\u1_u0_pid_reg[3]/NET0131  & ~\u1_u3_this_dpid_reg[0]/P0001  ;
  assign n9044 = \u1_u0_pid_reg[3]/NET0131  & \u1_u3_this_dpid_reg[0]/P0001  ;
  assign n9045 = ~n9043 & ~n9044 ;
  assign n9046 = \u1_u0_pid_reg[1]/NET0131  & ~n9045 ;
  assign n9047 = n9042 & n9046 ;
  assign n9048 = \u1_u2_sizu_c_reg[1]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n9049 = \u1_u3_new_size_reg[1]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n9050 = ~n9048 & ~n9049 ;
  assign n9051 = ~n5706 & ~n5708 ;
  assign n9052 = ~n5707 & ~n5712 ;
  assign n9053 = n9051 & n9052 ;
  assign n9054 = ~n9051 & ~n9052 ;
  assign n9055 = ~n9053 & ~n9054 ;
  assign n9056 = ~n5711 & ~n5716 ;
  assign n9057 = ~n7771 & ~n9056 ;
  assign n9058 = ~n5712 & n9056 ;
  assign n9059 = ~n5710 & n9058 ;
  assign n9060 = ~n9057 & ~n9059 ;
  assign n9061 = ~\u4_u3_buf0_orig_reg[28]/P0001  & \u4_u3_dma_out_cnt_reg[9]/P0001  ;
  assign n9062 = ~\u4_u3_buf0_orig_reg[27]/P0001  & \u4_u3_dma_out_cnt_reg[8]/P0001  ;
  assign n9063 = \u4_u3_buf0_orig_reg[27]/P0001  & ~\u4_u3_dma_out_cnt_reg[8]/P0001  ;
  assign n9064 = \u4_u3_buf0_orig_reg[26]/P0001  & ~\u4_u3_dma_out_cnt_reg[7]/P0001  ;
  assign n9065 = ~n9063 & ~n9064 ;
  assign n9066 = ~n9062 & ~n9065 ;
  assign n9067 = \u4_u3_buf0_orig_reg[25]/P0001  & ~\u4_u3_dma_out_cnt_reg[6]/P0001  ;
  assign n9068 = ~\u4_u3_buf0_orig_reg[24]/P0001  & \u4_u3_dma_out_cnt_reg[5]/P0001  ;
  assign n9069 = ~n9067 & n9068 ;
  assign n9070 = ~\u4_u3_buf0_orig_reg[23]/P0001  & \u4_u3_dma_out_cnt_reg[4]/P0001  ;
  assign n9071 = ~\u4_u3_buf0_orig_reg[22]/P0001  & \u4_u3_dma_out_cnt_reg[3]/P0001  ;
  assign n9072 = ~n9070 & ~n9071 ;
  assign n9073 = \u4_u3_buf0_orig_reg[22]/P0001  & ~\u4_u3_dma_out_cnt_reg[3]/P0001  ;
  assign n9074 = n9072 & n9073 ;
  assign n9075 = ~\u4_u3_buf0_orig_reg[20]/P0001  & \u4_u3_dma_out_cnt_reg[1]/P0001  ;
  assign n9076 = ~\u4_u3_buf0_orig_reg[19]/P0001  & \u4_u3_dma_in_cnt_reg[0]/P0001  ;
  assign n9077 = ~n9075 & ~n9076 ;
  assign n9078 = \u4_u3_buf0_orig_reg[21]/P0001  & ~\u4_u3_dma_out_cnt_reg[2]/P0001  ;
  assign n9079 = \u4_u3_buf0_orig_reg[20]/P0001  & ~\u4_u3_dma_out_cnt_reg[1]/P0001  ;
  assign n9080 = ~n9078 & ~n9079 ;
  assign n9081 = ~n9077 & n9080 ;
  assign n9082 = ~\u4_u3_buf0_orig_reg[21]/P0001  & \u4_u3_dma_out_cnt_reg[2]/P0001  ;
  assign n9083 = n9072 & ~n9082 ;
  assign n9084 = ~n9081 & n9083 ;
  assign n9085 = ~n9074 & ~n9084 ;
  assign n9086 = \u4_u3_buf0_orig_reg[24]/P0001  & ~\u4_u3_dma_out_cnt_reg[5]/P0001  ;
  assign n9087 = \u4_u3_buf0_orig_reg[23]/P0001  & ~\u4_u3_dma_out_cnt_reg[4]/P0001  ;
  assign n9088 = ~n9086 & ~n9087 ;
  assign n9089 = ~n9067 & n9088 ;
  assign n9090 = n9085 & n9089 ;
  assign n9091 = ~n9069 & ~n9090 ;
  assign n9092 = ~\u4_u3_buf0_orig_reg[26]/P0001  & \u4_u3_dma_out_cnt_reg[7]/P0001  ;
  assign n9093 = ~\u4_u3_buf0_orig_reg[25]/P0001  & \u4_u3_dma_out_cnt_reg[6]/P0001  ;
  assign n9094 = ~n9092 & ~n9093 ;
  assign n9095 = ~n9062 & n9094 ;
  assign n9096 = n9091 & n9095 ;
  assign n9097 = ~n9066 & ~n9096 ;
  assign n9098 = ~n9061 & ~n9097 ;
  assign n9099 = \u4_u3_buf0_orig_reg[29]/NET0131  & ~\u4_u3_dma_out_cnt_reg[10]/P0001  ;
  assign n9100 = ~\u4_u3_buf0_orig_reg[29]/NET0131  & \u4_u3_dma_out_cnt_reg[10]/P0001  ;
  assign n9101 = ~n9099 & ~n9100 ;
  assign n9102 = \u4_u3_buf0_orig_reg[28]/P0001  & ~\u4_u3_dma_out_cnt_reg[9]/P0001  ;
  assign n9103 = n9101 & ~n9102 ;
  assign n9104 = ~n9098 & n9103 ;
  assign n9105 = ~n9101 & n9102 ;
  assign n9106 = ~n9061 & ~n9101 ;
  assign n9107 = ~n9097 & n9106 ;
  assign n9108 = ~n9105 & ~n9107 ;
  assign n9109 = ~n9104 & n9108 ;
  assign n9110 = ~\u4_u0_buf0_orig_reg[28]/P0001  & \u4_u0_dma_out_cnt_reg[9]/P0001  ;
  assign n9111 = ~\u4_u0_buf0_orig_reg[27]/P0001  & \u4_u0_dma_out_cnt_reg[8]/P0001  ;
  assign n9112 = \u4_u0_buf0_orig_reg[27]/P0001  & ~\u4_u0_dma_out_cnt_reg[8]/P0001  ;
  assign n9113 = \u4_u0_buf0_orig_reg[26]/P0001  & ~\u4_u0_dma_out_cnt_reg[7]/P0001  ;
  assign n9114 = ~n9112 & ~n9113 ;
  assign n9115 = ~n9111 & ~n9114 ;
  assign n9116 = \u4_u0_buf0_orig_reg[25]/P0001  & ~\u4_u0_dma_out_cnt_reg[6]/P0001  ;
  assign n9117 = ~\u4_u0_buf0_orig_reg[24]/P0001  & \u4_u0_dma_out_cnt_reg[5]/P0001  ;
  assign n9118 = ~n9116 & n9117 ;
  assign n9119 = ~\u4_u0_buf0_orig_reg[23]/P0001  & \u4_u0_dma_out_cnt_reg[4]/P0001  ;
  assign n9120 = ~\u4_u0_buf0_orig_reg[22]/P0001  & \u4_u0_dma_out_cnt_reg[3]/P0001  ;
  assign n9121 = ~n9119 & ~n9120 ;
  assign n9122 = \u4_u0_buf0_orig_reg[22]/P0001  & ~\u4_u0_dma_out_cnt_reg[3]/P0001  ;
  assign n9123 = n9121 & n9122 ;
  assign n9124 = ~\u4_u0_buf0_orig_reg[20]/P0001  & \u4_u0_dma_out_cnt_reg[1]/P0001  ;
  assign n9125 = ~\u4_u0_buf0_orig_reg[19]/P0001  & \u4_u0_dma_in_cnt_reg[0]/P0001  ;
  assign n9126 = ~n9124 & ~n9125 ;
  assign n9127 = \u4_u0_buf0_orig_reg[21]/P0001  & ~\u4_u0_dma_out_cnt_reg[2]/P0001  ;
  assign n9128 = \u4_u0_buf0_orig_reg[20]/P0001  & ~\u4_u0_dma_out_cnt_reg[1]/P0001  ;
  assign n9129 = ~n9127 & ~n9128 ;
  assign n9130 = ~n9126 & n9129 ;
  assign n9131 = ~\u4_u0_buf0_orig_reg[21]/P0001  & \u4_u0_dma_out_cnt_reg[2]/P0001  ;
  assign n9132 = n9121 & ~n9131 ;
  assign n9133 = ~n9130 & n9132 ;
  assign n9134 = ~n9123 & ~n9133 ;
  assign n9135 = \u4_u0_buf0_orig_reg[24]/P0001  & ~\u4_u0_dma_out_cnt_reg[5]/P0001  ;
  assign n9136 = \u4_u0_buf0_orig_reg[23]/P0001  & ~\u4_u0_dma_out_cnt_reg[4]/P0001  ;
  assign n9137 = ~n9135 & ~n9136 ;
  assign n9138 = ~n9116 & n9137 ;
  assign n9139 = n9134 & n9138 ;
  assign n9140 = ~n9118 & ~n9139 ;
  assign n9141 = ~\u4_u0_buf0_orig_reg[26]/P0001  & \u4_u0_dma_out_cnt_reg[7]/P0001  ;
  assign n9142 = ~\u4_u0_buf0_orig_reg[25]/P0001  & \u4_u0_dma_out_cnt_reg[6]/P0001  ;
  assign n9143 = ~n9141 & ~n9142 ;
  assign n9144 = ~n9111 & n9143 ;
  assign n9145 = n9140 & n9144 ;
  assign n9146 = ~n9115 & ~n9145 ;
  assign n9147 = ~n9110 & ~n9146 ;
  assign n9148 = \u4_u0_buf0_orig_reg[29]/NET0131  & ~\u4_u0_dma_out_cnt_reg[10]/P0001  ;
  assign n9149 = ~\u4_u0_buf0_orig_reg[29]/NET0131  & \u4_u0_dma_out_cnt_reg[10]/P0001  ;
  assign n9150 = ~n9148 & ~n9149 ;
  assign n9151 = \u4_u0_buf0_orig_reg[28]/P0001  & ~\u4_u0_dma_out_cnt_reg[9]/P0001  ;
  assign n9152 = n9150 & ~n9151 ;
  assign n9153 = ~n9147 & n9152 ;
  assign n9154 = ~n9150 & n9151 ;
  assign n9155 = ~n9110 & ~n9150 ;
  assign n9156 = ~n9146 & n9155 ;
  assign n9157 = ~n9154 & ~n9156 ;
  assign n9158 = ~n9153 & n9157 ;
  assign n9159 = ~\u4_u1_buf0_orig_reg[28]/P0001  & \u4_u1_dma_out_cnt_reg[9]/P0001  ;
  assign n9160 = ~\u4_u1_buf0_orig_reg[27]/P0001  & \u4_u1_dma_out_cnt_reg[8]/P0001  ;
  assign n9161 = \u4_u1_buf0_orig_reg[27]/P0001  & ~\u4_u1_dma_out_cnt_reg[8]/P0001  ;
  assign n9162 = \u4_u1_buf0_orig_reg[26]/P0001  & ~\u4_u1_dma_out_cnt_reg[7]/P0001  ;
  assign n9163 = ~n9161 & ~n9162 ;
  assign n9164 = ~n9160 & ~n9163 ;
  assign n9165 = \u4_u1_buf0_orig_reg[25]/P0001  & ~\u4_u1_dma_out_cnt_reg[6]/P0001  ;
  assign n9166 = ~\u4_u1_buf0_orig_reg[24]/P0001  & \u4_u1_dma_out_cnt_reg[5]/P0001  ;
  assign n9167 = ~n9165 & n9166 ;
  assign n9168 = ~\u4_u1_buf0_orig_reg[23]/P0001  & \u4_u1_dma_out_cnt_reg[4]/P0001  ;
  assign n9169 = ~\u4_u1_buf0_orig_reg[22]/P0001  & \u4_u1_dma_out_cnt_reg[3]/P0001  ;
  assign n9170 = ~n9168 & ~n9169 ;
  assign n9171 = \u4_u1_buf0_orig_reg[22]/P0001  & ~\u4_u1_dma_out_cnt_reg[3]/P0001  ;
  assign n9172 = n9170 & n9171 ;
  assign n9173 = ~\u4_u1_buf0_orig_reg[20]/P0001  & \u4_u1_dma_out_cnt_reg[1]/P0001  ;
  assign n9174 = ~\u4_u1_buf0_orig_reg[19]/P0001  & \u4_u1_dma_in_cnt_reg[0]/P0001  ;
  assign n9175 = ~n9173 & ~n9174 ;
  assign n9176 = \u4_u1_buf0_orig_reg[21]/P0001  & ~\u4_u1_dma_out_cnt_reg[2]/P0001  ;
  assign n9177 = \u4_u1_buf0_orig_reg[20]/P0001  & ~\u4_u1_dma_out_cnt_reg[1]/P0001  ;
  assign n9178 = ~n9176 & ~n9177 ;
  assign n9179 = ~n9175 & n9178 ;
  assign n9180 = ~\u4_u1_buf0_orig_reg[21]/P0001  & \u4_u1_dma_out_cnt_reg[2]/P0001  ;
  assign n9181 = n9170 & ~n9180 ;
  assign n9182 = ~n9179 & n9181 ;
  assign n9183 = ~n9172 & ~n9182 ;
  assign n9184 = \u4_u1_buf0_orig_reg[24]/P0001  & ~\u4_u1_dma_out_cnt_reg[5]/P0001  ;
  assign n9185 = \u4_u1_buf0_orig_reg[23]/P0001  & ~\u4_u1_dma_out_cnt_reg[4]/P0001  ;
  assign n9186 = ~n9184 & ~n9185 ;
  assign n9187 = ~n9165 & n9186 ;
  assign n9188 = n9183 & n9187 ;
  assign n9189 = ~n9167 & ~n9188 ;
  assign n9190 = ~\u4_u1_buf0_orig_reg[26]/P0001  & \u4_u1_dma_out_cnt_reg[7]/P0001  ;
  assign n9191 = ~\u4_u1_buf0_orig_reg[25]/P0001  & \u4_u1_dma_out_cnt_reg[6]/P0001  ;
  assign n9192 = ~n9190 & ~n9191 ;
  assign n9193 = ~n9160 & n9192 ;
  assign n9194 = n9189 & n9193 ;
  assign n9195 = ~n9164 & ~n9194 ;
  assign n9196 = ~n9159 & ~n9195 ;
  assign n9197 = \u4_u1_buf0_orig_reg[29]/NET0131  & ~\u4_u1_dma_out_cnt_reg[10]/P0001  ;
  assign n9198 = ~\u4_u1_buf0_orig_reg[29]/NET0131  & \u4_u1_dma_out_cnt_reg[10]/P0001  ;
  assign n9199 = ~n9197 & ~n9198 ;
  assign n9200 = \u4_u1_buf0_orig_reg[28]/P0001  & ~\u4_u1_dma_out_cnt_reg[9]/P0001  ;
  assign n9201 = n9199 & ~n9200 ;
  assign n9202 = ~n9196 & n9201 ;
  assign n9203 = ~n9199 & n9200 ;
  assign n9204 = ~n9159 & ~n9199 ;
  assign n9205 = ~n9195 & n9204 ;
  assign n9206 = ~n9203 & ~n9205 ;
  assign n9207 = ~n9202 & n9206 ;
  assign n9208 = ~\u4_u2_buf0_orig_reg[28]/P0001  & \u4_u2_dma_out_cnt_reg[9]/P0001  ;
  assign n9209 = ~\u4_u2_buf0_orig_reg[27]/P0001  & \u4_u2_dma_out_cnt_reg[8]/P0001  ;
  assign n9210 = \u4_u2_buf0_orig_reg[27]/P0001  & ~\u4_u2_dma_out_cnt_reg[8]/P0001  ;
  assign n9211 = \u4_u2_buf0_orig_reg[26]/P0001  & ~\u4_u2_dma_out_cnt_reg[7]/P0001  ;
  assign n9212 = ~n9210 & ~n9211 ;
  assign n9213 = ~n9209 & ~n9212 ;
  assign n9214 = \u4_u2_buf0_orig_reg[25]/P0001  & ~\u4_u2_dma_out_cnt_reg[6]/P0001  ;
  assign n9215 = ~\u4_u2_buf0_orig_reg[24]/P0001  & \u4_u2_dma_out_cnt_reg[5]/P0001  ;
  assign n9216 = ~n9214 & n9215 ;
  assign n9217 = ~\u4_u2_buf0_orig_reg[23]/P0001  & \u4_u2_dma_out_cnt_reg[4]/P0001  ;
  assign n9218 = ~\u4_u2_buf0_orig_reg[22]/P0001  & \u4_u2_dma_out_cnt_reg[3]/P0001  ;
  assign n9219 = ~n9217 & ~n9218 ;
  assign n9220 = \u4_u2_buf0_orig_reg[22]/P0001  & ~\u4_u2_dma_out_cnt_reg[3]/P0001  ;
  assign n9221 = n9219 & n9220 ;
  assign n9222 = ~\u4_u2_buf0_orig_reg[20]/P0001  & \u4_u2_dma_out_cnt_reg[1]/P0001  ;
  assign n9223 = ~\u4_u2_buf0_orig_reg[19]/P0001  & \u4_u2_dma_in_cnt_reg[0]/P0001  ;
  assign n9224 = ~n9222 & ~n9223 ;
  assign n9225 = \u4_u2_buf0_orig_reg[21]/P0001  & ~\u4_u2_dma_out_cnt_reg[2]/P0001  ;
  assign n9226 = \u4_u2_buf0_orig_reg[20]/P0001  & ~\u4_u2_dma_out_cnt_reg[1]/P0001  ;
  assign n9227 = ~n9225 & ~n9226 ;
  assign n9228 = ~n9224 & n9227 ;
  assign n9229 = ~\u4_u2_buf0_orig_reg[21]/P0001  & \u4_u2_dma_out_cnt_reg[2]/P0001  ;
  assign n9230 = n9219 & ~n9229 ;
  assign n9231 = ~n9228 & n9230 ;
  assign n9232 = ~n9221 & ~n9231 ;
  assign n9233 = \u4_u2_buf0_orig_reg[24]/P0001  & ~\u4_u2_dma_out_cnt_reg[5]/P0001  ;
  assign n9234 = \u4_u2_buf0_orig_reg[23]/P0001  & ~\u4_u2_dma_out_cnt_reg[4]/P0001  ;
  assign n9235 = ~n9233 & ~n9234 ;
  assign n9236 = ~n9214 & n9235 ;
  assign n9237 = n9232 & n9236 ;
  assign n9238 = ~n9216 & ~n9237 ;
  assign n9239 = ~\u4_u2_buf0_orig_reg[26]/P0001  & \u4_u2_dma_out_cnt_reg[7]/P0001  ;
  assign n9240 = ~\u4_u2_buf0_orig_reg[25]/P0001  & \u4_u2_dma_out_cnt_reg[6]/P0001  ;
  assign n9241 = ~n9239 & ~n9240 ;
  assign n9242 = ~n9209 & n9241 ;
  assign n9243 = n9238 & n9242 ;
  assign n9244 = ~n9213 & ~n9243 ;
  assign n9245 = ~n9208 & ~n9244 ;
  assign n9246 = \u4_u2_buf0_orig_reg[29]/NET0131  & ~\u4_u2_dma_out_cnt_reg[10]/P0001  ;
  assign n9247 = ~\u4_u2_buf0_orig_reg[29]/NET0131  & \u4_u2_dma_out_cnt_reg[10]/P0001  ;
  assign n9248 = ~n9246 & ~n9247 ;
  assign n9249 = \u4_u2_buf0_orig_reg[28]/P0001  & ~\u4_u2_dma_out_cnt_reg[9]/P0001  ;
  assign n9250 = n9248 & ~n9249 ;
  assign n9251 = ~n9245 & n9250 ;
  assign n9252 = ~n9248 & n9249 ;
  assign n9253 = ~n9208 & ~n9248 ;
  assign n9254 = ~n9244 & n9253 ;
  assign n9255 = ~n9252 & ~n9254 ;
  assign n9256 = ~n9251 & n9255 ;
  assign n9257 = ~n6261 & ~n6269 ;
  assign n9258 = n6598 & n9257 ;
  assign n9259 = ~n6591 & n6598 ;
  assign n9260 = n6588 & n9259 ;
  assign n9261 = ~n9258 & ~n9260 ;
  assign n9262 = ~\u4_u3_dma_in_cnt_reg[6]/P0001  & ~n8519 ;
  assign n9263 = \u4_u3_r5_reg/NET0131  & ~n6277 ;
  assign n9264 = ~n9262 & n9263 ;
  assign n9265 = ~n6591 & n9257 ;
  assign n9266 = n6588 & n9265 ;
  assign n9267 = ~n9264 & ~n9266 ;
  assign n9268 = ~n9261 & n9267 ;
  assign n9269 = ~\u4_u3_dma_in_cnt_reg[6]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n9270 = n6281 & n9269 ;
  assign n9271 = ~\u4_u3_dma_in_cnt_reg[6]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n9272 = ~\u4_u3_r5_reg/NET0131  & ~n9271 ;
  assign n9273 = ~n9270 & n9272 ;
  assign n9274 = ~n9264 & ~n9273 ;
  assign n9275 = \u4_u3_csr1_reg[0]/P0001  & ~n9274 ;
  assign n9276 = ~n9268 & n9275 ;
  assign n9277 = ~\u4_u3_dma_out_cnt_reg[6]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n9278 = n7308 & n9277 ;
  assign n9279 = n6740 & n9278 ;
  assign n9280 = \u4_u3_csr1_reg[0]/P0001  & n9279 ;
  assign n9281 = \u4_u3_dma_out_cnt_reg[6]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n9282 = \u4_u3_csr1_reg[0]/P0001  & n9281 ;
  assign n9283 = ~n7309 & n9282 ;
  assign n9284 = ~n9280 & ~n9283 ;
  assign n9285 = ~n6758 & ~n6760 ;
  assign n9286 = n6761 & ~n9285 ;
  assign n9287 = n6781 & ~n9285 ;
  assign n9288 = n6778 & n9287 ;
  assign n9289 = ~n9286 & ~n9288 ;
  assign n9290 = ~n6761 & n9285 ;
  assign n9291 = ~n8365 & n9290 ;
  assign n9292 = n9289 & ~n9291 ;
  assign n9293 = n6598 & n9292 ;
  assign n9294 = ~\u4_u3_dma_out_cnt_reg[6]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n9295 = n6281 & n9294 ;
  assign n9296 = ~\u4_u3_dma_out_cnt_reg[6]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n9297 = \u4_u3_csr1_reg[0]/P0001  & ~n9296 ;
  assign n9298 = ~n9295 & n9297 ;
  assign n9299 = ~\u4_u3_r5_reg/NET0131  & n9298 ;
  assign n9300 = ~n9293 & n9299 ;
  assign n9301 = n9284 & ~n9300 ;
  assign n9302 = ~n6319 & ~n6327 ;
  assign n9303 = n6632 & n9302 ;
  assign n9304 = ~n6625 & n6632 ;
  assign n9305 = n6622 & n9304 ;
  assign n9306 = ~n9303 & ~n9305 ;
  assign n9307 = ~\u4_u0_dma_in_cnt_reg[6]/P0001  & ~n8544 ;
  assign n9308 = \u4_u0_r5_reg/NET0131  & ~n6335 ;
  assign n9309 = ~n9307 & n9308 ;
  assign n9310 = ~n6625 & n9302 ;
  assign n9311 = n6622 & n9310 ;
  assign n9312 = ~n9309 & ~n9311 ;
  assign n9313 = ~n9306 & n9312 ;
  assign n9314 = ~\u4_u0_dma_in_cnt_reg[6]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n9315 = n6281 & n9314 ;
  assign n9316 = ~\u4_u0_dma_in_cnt_reg[6]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n9317 = ~\u4_u0_r5_reg/NET0131  & ~n9316 ;
  assign n9318 = ~n9315 & n9317 ;
  assign n9319 = ~n9309 & ~n9318 ;
  assign n9320 = \u4_u0_csr1_reg[0]/P0001  & ~n9319 ;
  assign n9321 = ~n9313 & n9320 ;
  assign n9322 = ~\u4_u0_dma_out_cnt_reg[6]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n9323 = n7358 & n9322 ;
  assign n9324 = n6804 & n9323 ;
  assign n9325 = \u4_u0_csr1_reg[0]/P0001  & n9324 ;
  assign n9326 = \u4_u0_dma_out_cnt_reg[6]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n9327 = \u4_u0_csr1_reg[0]/P0001  & n9326 ;
  assign n9328 = ~n7359 & n9327 ;
  assign n9329 = ~n9325 & ~n9328 ;
  assign n9330 = ~n6826 & ~n6852 ;
  assign n9331 = n6827 & ~n9330 ;
  assign n9332 = n6847 & ~n9330 ;
  assign n9333 = n6844 & n9332 ;
  assign n9334 = ~n9331 & ~n9333 ;
  assign n9335 = ~n6827 & n9330 ;
  assign n9336 = ~n8381 & n9335 ;
  assign n9337 = n9334 & ~n9336 ;
  assign n9338 = n6632 & n9337 ;
  assign n9339 = ~\u4_u0_dma_out_cnt_reg[6]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n9340 = n6281 & n9339 ;
  assign n9341 = ~\u4_u0_dma_out_cnt_reg[6]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n9342 = \u4_u0_csr1_reg[0]/P0001  & ~n9341 ;
  assign n9343 = ~n9340 & n9342 ;
  assign n9344 = ~\u4_u0_r5_reg/NET0131  & n9343 ;
  assign n9345 = ~n9338 & n9344 ;
  assign n9346 = n9329 & ~n9345 ;
  assign n9347 = \u4_u1_r5_reg/NET0131  & ~n6362 ;
  assign n9348 = \u4_u1_csr1_reg[0]/P0001  & \u4_u1_dma_in_cnt_reg[6]/P0001  ;
  assign n9349 = \u4_u1_csr1_reg[0]/P0001  & n8578 ;
  assign n9350 = n6361 & n9349 ;
  assign n9351 = ~n9348 & ~n9350 ;
  assign n9352 = n9347 & ~n9351 ;
  assign n9353 = ~n6378 & ~n6405 ;
  assign n9354 = ~n6379 & ~n9353 ;
  assign n9355 = ~n6653 & n9354 ;
  assign n9356 = n6379 & n9353 ;
  assign n9357 = n6399 & n9353 ;
  assign n9358 = n6396 & n9357 ;
  assign n9359 = ~n9356 & ~n9358 ;
  assign n9360 = ~n9355 & n9359 ;
  assign n9361 = n6369 & n9360 ;
  assign n9362 = ~\u4_u1_dma_in_cnt_reg[6]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n9363 = n6281 & n9362 ;
  assign n9364 = ~\u4_u1_dma_in_cnt_reg[6]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n9365 = \u4_u1_csr1_reg[0]/P0001  & ~n9364 ;
  assign n9366 = ~n9363 & n9365 ;
  assign n9367 = ~\u4_u1_r5_reg/NET0131  & n9366 ;
  assign n9368 = ~n9361 & n9367 ;
  assign n9369 = ~n9352 & ~n9368 ;
  assign n9370 = ~\u4_u1_dma_out_cnt_reg[6]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n9371 = n7408 & n9370 ;
  assign n9372 = n6868 & n9371 ;
  assign n9373 = \u4_u1_csr1_reg[0]/P0001  & n9372 ;
  assign n9374 = \u4_u1_dma_out_cnt_reg[6]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n9375 = \u4_u1_csr1_reg[0]/P0001  & n9374 ;
  assign n9376 = ~n7409 & n9375 ;
  assign n9377 = ~n9373 & ~n9376 ;
  assign n9378 = ~n6890 & ~n6916 ;
  assign n9379 = n6891 & ~n9378 ;
  assign n9380 = n6911 & ~n9378 ;
  assign n9381 = n6908 & n9380 ;
  assign n9382 = ~n9379 & ~n9381 ;
  assign n9383 = ~n6891 & n9378 ;
  assign n9384 = ~n8411 & n9383 ;
  assign n9385 = n9382 & ~n9384 ;
  assign n9386 = n6369 & n9385 ;
  assign n9387 = ~\u4_u1_dma_out_cnt_reg[6]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n9388 = n6281 & n9387 ;
  assign n9389 = ~\u4_u1_dma_out_cnt_reg[6]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n9390 = \u4_u1_csr1_reg[0]/P0001  & ~n9389 ;
  assign n9391 = ~n9388 & n9390 ;
  assign n9392 = ~\u4_u1_r5_reg/NET0131  & n9391 ;
  assign n9393 = ~n9386 & n9392 ;
  assign n9394 = n9377 & ~n9393 ;
  assign n9395 = ~\u4_u2_dma_in_cnt_reg[6]/P0001  & ~n8603 ;
  assign n9396 = \u4_u2_csr1_reg[0]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n9397 = ~n6463 & n9396 ;
  assign n9398 = ~n9395 & n9397 ;
  assign n9399 = ~\u4_u2_dma_in_cnt_reg[6]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n9400 = n6281 & n9399 ;
  assign n9401 = ~\u4_u2_dma_in_cnt_reg[6]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n9402 = n6946 & ~n9401 ;
  assign n9403 = ~n9400 & n9402 ;
  assign n9404 = ~n9398 & ~n9403 ;
  assign n9405 = ~n6425 & ~n6451 ;
  assign n9406 = ~n6426 & ~n9405 ;
  assign n9407 = ~n8324 & n9406 ;
  assign n9408 = n6426 & n9405 ;
  assign n9409 = n6446 & n9405 ;
  assign n9410 = n6443 & n9409 ;
  assign n9411 = ~n9408 & ~n9410 ;
  assign n9412 = ~n9407 & n9411 ;
  assign n9413 = n6667 & ~n9398 ;
  assign n9414 = n9412 & n9413 ;
  assign n9415 = ~n9404 & ~n9414 ;
  assign n9416 = \u4_u2_dma_out_cnt_reg[6]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n9417 = ~n7459 & n9416 ;
  assign n9418 = ~\u4_u2_dma_out_cnt_reg[6]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n9419 = n7458 & n9418 ;
  assign n9420 = n6932 & n9419 ;
  assign n9421 = ~n9417 & ~n9420 ;
  assign n9422 = ~\u4_u2_dma_out_cnt_reg[6]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n9423 = n6281 & n9422 ;
  assign n9424 = ~\u4_u2_dma_out_cnt_reg[6]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n9425 = ~\u4_u2_r5_reg/NET0131  & ~n9424 ;
  assign n9426 = ~n9423 & n9425 ;
  assign n9427 = n9421 & ~n9426 ;
  assign n9428 = ~n6951 & ~n6953 ;
  assign n9429 = n6954 & ~n9428 ;
  assign n9430 = n6974 & ~n9428 ;
  assign n9431 = n6971 & n9430 ;
  assign n9432 = ~n9429 & ~n9431 ;
  assign n9433 = ~n6954 & n9428 ;
  assign n9434 = ~n8429 & n9433 ;
  assign n9435 = n9432 & ~n9434 ;
  assign n9436 = n6667 & n9421 ;
  assign n9437 = n9435 & n9436 ;
  assign n9438 = ~n9427 & ~n9437 ;
  assign n9439 = \u4_u2_csr1_reg[0]/P0001  & n9438 ;
  assign n9440 = ~n6249 & ~n6258 ;
  assign n9441 = n6584 & ~n9440 ;
  assign n9442 = n6598 & ~n9441 ;
  assign n9443 = ~n6584 & n9440 ;
  assign n9444 = ~n7501 & n9443 ;
  assign n9445 = n6254 & ~n9440 ;
  assign n9446 = ~n6586 & n9445 ;
  assign n9447 = \u4_u3_dma_in_cnt_reg[4]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n9448 = ~n6276 & n9447 ;
  assign n9449 = ~\u4_u3_dma_in_cnt_reg[4]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n9450 = n6276 & n9449 ;
  assign n9451 = ~n9448 & ~n9450 ;
  assign n9452 = ~n9446 & n9451 ;
  assign n9453 = ~n9444 & n9452 ;
  assign n9454 = n9442 & n9453 ;
  assign n9455 = ~\u4_u3_dma_in_cnt_reg[4]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n9456 = n6281 & n9455 ;
  assign n9457 = ~\u4_u3_dma_in_cnt_reg[4]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n9458 = ~\u4_u3_r5_reg/NET0131  & ~n9457 ;
  assign n9459 = ~n9456 & n9458 ;
  assign n9460 = n9451 & ~n9459 ;
  assign n9461 = \u4_u3_csr1_reg[0]/P0001  & ~n9460 ;
  assign n9462 = ~n9454 & n9461 ;
  assign n9463 = ~n6307 & ~n6316 ;
  assign n9464 = n6618 & ~n9463 ;
  assign n9465 = n6632 & ~n9464 ;
  assign n9466 = ~n6618 & n9463 ;
  assign n9467 = ~n7532 & n9466 ;
  assign n9468 = n6312 & ~n9463 ;
  assign n9469 = ~n6620 & n9468 ;
  assign n9470 = \u4_u0_dma_in_cnt_reg[4]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n9471 = ~n6334 & n9470 ;
  assign n9472 = ~\u4_u0_dma_in_cnt_reg[4]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n9473 = n6334 & n9472 ;
  assign n9474 = ~n9471 & ~n9473 ;
  assign n9475 = ~n9469 & n9474 ;
  assign n9476 = ~n9467 & n9475 ;
  assign n9477 = n9465 & n9476 ;
  assign n9478 = ~\u4_u0_dma_in_cnt_reg[4]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n9479 = n6281 & n9478 ;
  assign n9480 = ~\u4_u0_dma_in_cnt_reg[4]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n9481 = ~\u4_u0_r5_reg/NET0131  & ~n9480 ;
  assign n9482 = ~n9479 & n9481 ;
  assign n9483 = n9474 & ~n9482 ;
  assign n9484 = \u4_u0_csr1_reg[0]/P0001  & ~n9483 ;
  assign n9485 = ~n9477 & n9484 ;
  assign n9486 = \u4_u1_dma_in_cnt_reg[4]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n9487 = ~n6361 & n9486 ;
  assign n9488 = ~\u4_u1_dma_in_cnt_reg[4]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n9489 = n6361 & n9488 ;
  assign n9490 = ~n9487 & ~n9489 ;
  assign n9491 = ~n6381 & ~n6398 ;
  assign n9492 = ~n6382 & ~n6393 ;
  assign n9493 = ~n9491 & n9492 ;
  assign n9494 = ~n6392 & n9493 ;
  assign n9495 = n6384 & ~n9491 ;
  assign n9496 = n6369 & ~n9495 ;
  assign n9497 = ~n9494 & n9496 ;
  assign n9498 = ~n6392 & n9492 ;
  assign n9499 = ~n6384 & n9491 ;
  assign n9500 = ~n9498 & n9499 ;
  assign n9501 = n9497 & ~n9500 ;
  assign n9502 = n9490 & n9501 ;
  assign n9503 = ~\u4_u1_dma_in_cnt_reg[4]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n9504 = n6281 & n9503 ;
  assign n9505 = ~\u4_u1_dma_in_cnt_reg[4]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n9506 = ~\u4_u1_r5_reg/NET0131  & ~n9505 ;
  assign n9507 = ~n9504 & n9506 ;
  assign n9508 = n9490 & ~n9507 ;
  assign n9509 = \u4_u1_csr1_reg[0]/P0001  & ~n9508 ;
  assign n9510 = ~n9502 & n9509 ;
  assign n9511 = \u4_u2_dma_in_cnt_reg[4]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n9512 = ~n6462 & n9511 ;
  assign n9513 = ~\u4_u2_dma_in_cnt_reg[4]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n9514 = n6462 & n9513 ;
  assign n9515 = ~n9512 & ~n9514 ;
  assign n9516 = ~n6428 & ~n6445 ;
  assign n9517 = ~n6429 & ~n6440 ;
  assign n9518 = ~n9516 & n9517 ;
  assign n9519 = ~n6439 & n9518 ;
  assign n9520 = n6431 & ~n9516 ;
  assign n9521 = n6667 & ~n9520 ;
  assign n9522 = ~n9519 & n9521 ;
  assign n9523 = ~n6439 & n9517 ;
  assign n9524 = ~n6431 & n9516 ;
  assign n9525 = ~n9523 & n9524 ;
  assign n9526 = n9522 & ~n9525 ;
  assign n9527 = n9515 & n9526 ;
  assign n9528 = ~\u4_u2_dma_in_cnt_reg[4]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n9529 = n6281 & n9528 ;
  assign n9530 = ~\u4_u2_dma_in_cnt_reg[4]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n9531 = ~\u4_u2_r5_reg/NET0131  & ~n9530 ;
  assign n9532 = ~n9529 & n9531 ;
  assign n9533 = n9515 & ~n9532 ;
  assign n9534 = \u4_u2_csr1_reg[0]/P0001  & ~n9533 ;
  assign n9535 = ~n9527 & n9534 ;
  assign n9536 = ~n6764 & ~n6775 ;
  assign n9537 = ~n6774 & n9536 ;
  assign n9538 = ~n6763 & ~n6780 ;
  assign n9539 = ~n6766 & ~n9538 ;
  assign n9540 = ~n9537 & n9539 ;
  assign n9541 = n6598 & ~n9540 ;
  assign n9542 = n9536 & n9538 ;
  assign n9543 = ~n6774 & n9542 ;
  assign n9544 = \u4_u3_dma_out_cnt_reg[4]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n9545 = ~n6740 & n9544 ;
  assign n9546 = ~\u4_u3_dma_out_cnt_reg[4]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n9547 = n6740 & n9546 ;
  assign n9548 = ~n9545 & ~n9547 ;
  assign n9549 = n6766 & n9538 ;
  assign n9550 = n9548 & ~n9549 ;
  assign n9551 = ~n9543 & n9550 ;
  assign n9552 = n9541 & n9551 ;
  assign n9553 = ~\u4_u3_dma_out_cnt_reg[4]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n9554 = n6281 & n9553 ;
  assign n9555 = ~\u4_u3_dma_out_cnt_reg[4]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n9556 = ~\u4_u3_r5_reg/NET0131  & ~n9555 ;
  assign n9557 = ~n9554 & n9556 ;
  assign n9558 = n9548 & ~n9557 ;
  assign n9559 = \u4_u3_csr1_reg[0]/P0001  & ~n9558 ;
  assign n9560 = ~n9552 & n9559 ;
  assign n9561 = ~n6830 & ~n6841 ;
  assign n9562 = ~n6840 & n9561 ;
  assign n9563 = ~n6829 & ~n6846 ;
  assign n9564 = ~n6832 & ~n9563 ;
  assign n9565 = ~n9562 & n9564 ;
  assign n9566 = n6632 & ~n9565 ;
  assign n9567 = n9561 & n9563 ;
  assign n9568 = ~n6840 & n9567 ;
  assign n9569 = \u4_u0_dma_out_cnt_reg[4]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n9570 = ~n6804 & n9569 ;
  assign n9571 = ~\u4_u0_dma_out_cnt_reg[4]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n9572 = n6804 & n9571 ;
  assign n9573 = ~n9570 & ~n9572 ;
  assign n9574 = n6832 & n9563 ;
  assign n9575 = n9573 & ~n9574 ;
  assign n9576 = ~n9568 & n9575 ;
  assign n9577 = n9566 & n9576 ;
  assign n9578 = ~\u4_u0_dma_out_cnt_reg[4]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n9579 = n6281 & n9578 ;
  assign n9580 = ~\u4_u0_dma_out_cnt_reg[4]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n9581 = ~\u4_u0_r5_reg/NET0131  & ~n9580 ;
  assign n9582 = ~n9579 & n9581 ;
  assign n9583 = n9573 & ~n9582 ;
  assign n9584 = \u4_u0_csr1_reg[0]/P0001  & ~n9583 ;
  assign n9585 = ~n9577 & n9584 ;
  assign n9586 = ~n6894 & ~n6905 ;
  assign n9587 = ~n6904 & n9586 ;
  assign n9588 = ~n6893 & ~n6910 ;
  assign n9589 = ~n6896 & ~n9588 ;
  assign n9590 = ~n9587 & n9589 ;
  assign n9591 = n6369 & ~n9590 ;
  assign n9592 = n9586 & n9588 ;
  assign n9593 = ~n6904 & n9592 ;
  assign n9594 = \u4_u1_dma_out_cnt_reg[4]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n9595 = ~n6868 & n9594 ;
  assign n9596 = ~\u4_u1_dma_out_cnt_reg[4]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n9597 = n6868 & n9596 ;
  assign n9598 = ~n9595 & ~n9597 ;
  assign n9599 = n6896 & n9588 ;
  assign n9600 = n9598 & ~n9599 ;
  assign n9601 = ~n9593 & n9600 ;
  assign n9602 = n9591 & n9601 ;
  assign n9603 = ~\u4_u1_dma_out_cnt_reg[4]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n9604 = n6281 & n9603 ;
  assign n9605 = ~\u4_u1_dma_out_cnt_reg[4]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n9606 = ~\u4_u1_r5_reg/NET0131  & ~n9605 ;
  assign n9607 = ~n9604 & n9606 ;
  assign n9608 = n9598 & ~n9607 ;
  assign n9609 = \u4_u1_csr1_reg[0]/P0001  & ~n9608 ;
  assign n9610 = ~n9602 & n9609 ;
  assign n9611 = ~n6957 & ~n6968 ;
  assign n9612 = ~n6967 & n9611 ;
  assign n9613 = ~n6956 & ~n6973 ;
  assign n9614 = ~n6959 & ~n9613 ;
  assign n9615 = ~n9612 & n9614 ;
  assign n9616 = n6667 & ~n9615 ;
  assign n9617 = n9611 & n9613 ;
  assign n9618 = ~n6967 & n9617 ;
  assign n9619 = \u4_u2_dma_out_cnt_reg[4]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n9620 = ~n6932 & n9619 ;
  assign n9621 = ~\u4_u2_dma_out_cnt_reg[4]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n9622 = n6932 & n9621 ;
  assign n9623 = ~n9620 & ~n9622 ;
  assign n9624 = n6959 & n9613 ;
  assign n9625 = n9623 & ~n9624 ;
  assign n9626 = ~n9618 & n9625 ;
  assign n9627 = n9616 & n9626 ;
  assign n9628 = ~\u4_u2_dma_out_cnt_reg[4]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n9629 = n6281 & n9628 ;
  assign n9630 = ~\u4_u2_dma_out_cnt_reg[4]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n9631 = ~\u4_u2_r5_reg/NET0131  & ~n9630 ;
  assign n9632 = ~n9629 & n9631 ;
  assign n9633 = n9623 & ~n9632 ;
  assign n9634 = \u4_u2_csr1_reg[0]/P0001  & ~n9633 ;
  assign n9635 = ~n9627 & n9634 ;
  assign n9636 = \u4_u3_buf1_reg[0]/P0001  & ~n2734 ;
  assign n9637 = \u1_u3_idin_reg[0]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9638 = ~n2733 & n9637 ;
  assign n9639 = ~n9636 & ~n9638 ;
  assign n9640 = ~n2732 & ~n9639 ;
  assign n9641 = \wb_data_i[0]_pad  & n2731 ;
  assign n9642 = n2567 & n9641 ;
  assign n9643 = rst_i_pad & ~n9642 ;
  assign n9644 = ~n9640 & n9643 ;
  assign n9645 = \u4_u3_buf1_reg[12]/P0001  & ~n2734 ;
  assign n9646 = \u1_u3_idin_reg[12]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9647 = ~n2733 & n9646 ;
  assign n9648 = ~n9645 & ~n9647 ;
  assign n9649 = ~n2732 & ~n9648 ;
  assign n9650 = \wb_data_i[12]_pad  & n2731 ;
  assign n9651 = n2567 & n9650 ;
  assign n9652 = rst_i_pad & ~n9651 ;
  assign n9653 = ~n9649 & n9652 ;
  assign n9654 = \u4_u3_buf1_reg[16]/P0001  & ~n2734 ;
  assign n9655 = \u1_u3_idin_reg[16]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9656 = ~n2733 & n9655 ;
  assign n9657 = ~n9654 & ~n9656 ;
  assign n9658 = ~n2732 & ~n9657 ;
  assign n9659 = \wb_data_i[16]_pad  & n2731 ;
  assign n9660 = n2567 & n9659 ;
  assign n9661 = rst_i_pad & ~n9660 ;
  assign n9662 = ~n9658 & n9661 ;
  assign n9663 = \u4_u3_buf1_reg[17]/P0001  & ~n2734 ;
  assign n9664 = \u1_u3_idin_reg[17]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9665 = ~n2733 & n9664 ;
  assign n9666 = ~n9663 & ~n9665 ;
  assign n9667 = ~n2732 & ~n9666 ;
  assign n9668 = \wb_data_i[17]_pad  & n2731 ;
  assign n9669 = n2567 & n9668 ;
  assign n9670 = rst_i_pad & ~n9669 ;
  assign n9671 = ~n9667 & n9670 ;
  assign n9672 = \u4_u3_buf1_reg[18]/P0001  & ~n2734 ;
  assign n9673 = \u1_u3_idin_reg[18]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9674 = ~n2733 & n9673 ;
  assign n9675 = ~n9672 & ~n9674 ;
  assign n9676 = ~n2732 & ~n9675 ;
  assign n9677 = \wb_data_i[18]_pad  & n2731 ;
  assign n9678 = n2567 & n9677 ;
  assign n9679 = rst_i_pad & ~n9678 ;
  assign n9680 = ~n9676 & n9679 ;
  assign n9681 = \u4_u3_buf1_reg[19]/P0001  & ~n2734 ;
  assign n9682 = \u1_u3_idin_reg[19]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9683 = ~n2733 & n9682 ;
  assign n9684 = ~n9681 & ~n9683 ;
  assign n9685 = ~n2732 & ~n9684 ;
  assign n9686 = \wb_data_i[19]_pad  & n2731 ;
  assign n9687 = n2567 & n9686 ;
  assign n9688 = rst_i_pad & ~n9687 ;
  assign n9689 = ~n9685 & n9688 ;
  assign n9690 = \u4_u3_buf1_reg[1]/P0001  & ~n2734 ;
  assign n9691 = \u1_u3_idin_reg[1]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9692 = ~n2733 & n9691 ;
  assign n9693 = ~n9690 & ~n9692 ;
  assign n9694 = ~n2732 & ~n9693 ;
  assign n9695 = \wb_data_i[1]_pad  & n2731 ;
  assign n9696 = n2567 & n9695 ;
  assign n9697 = rst_i_pad & ~n9696 ;
  assign n9698 = ~n9694 & n9697 ;
  assign n9699 = \u4_u3_buf1_reg[20]/P0001  & ~n2734 ;
  assign n9700 = \u1_u3_idin_reg[20]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9701 = ~n2733 & n9700 ;
  assign n9702 = ~n9699 & ~n9701 ;
  assign n9703 = ~n2732 & ~n9702 ;
  assign n9704 = \wb_data_i[20]_pad  & n2731 ;
  assign n9705 = n2567 & n9704 ;
  assign n9706 = rst_i_pad & ~n9705 ;
  assign n9707 = ~n9703 & n9706 ;
  assign n9708 = \u4_u3_buf1_reg[21]/P0001  & ~n2734 ;
  assign n9709 = \u1_u3_idin_reg[21]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9710 = ~n2733 & n9709 ;
  assign n9711 = ~n9708 & ~n9710 ;
  assign n9712 = ~n2732 & ~n9711 ;
  assign n9713 = \wb_data_i[21]_pad  & n2731 ;
  assign n9714 = n2567 & n9713 ;
  assign n9715 = rst_i_pad & ~n9714 ;
  assign n9716 = ~n9712 & n9715 ;
  assign n9717 = \u4_u3_buf1_reg[22]/P0001  & ~n2734 ;
  assign n9718 = \u1_u3_idin_reg[22]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9719 = ~n2733 & n9718 ;
  assign n9720 = ~n9717 & ~n9719 ;
  assign n9721 = ~n2732 & ~n9720 ;
  assign n9722 = \wb_data_i[22]_pad  & n2731 ;
  assign n9723 = n2567 & n9722 ;
  assign n9724 = rst_i_pad & ~n9723 ;
  assign n9725 = ~n9721 & n9724 ;
  assign n9726 = \u4_u3_buf1_reg[23]/P0001  & ~n2734 ;
  assign n9727 = \u1_u3_idin_reg[23]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9728 = ~n2733 & n9727 ;
  assign n9729 = ~n9726 & ~n9728 ;
  assign n9730 = ~n2732 & ~n9729 ;
  assign n9731 = \wb_data_i[23]_pad  & n2731 ;
  assign n9732 = n2567 & n9731 ;
  assign n9733 = rst_i_pad & ~n9732 ;
  assign n9734 = ~n9730 & n9733 ;
  assign n9735 = \u4_u3_buf1_reg[24]/P0001  & ~n2734 ;
  assign n9736 = \u1_u3_idin_reg[24]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9737 = ~n2733 & n9736 ;
  assign n9738 = ~n9735 & ~n9737 ;
  assign n9739 = ~n2732 & ~n9738 ;
  assign n9740 = \wb_data_i[24]_pad  & n2731 ;
  assign n9741 = n2567 & n9740 ;
  assign n9742 = rst_i_pad & ~n9741 ;
  assign n9743 = ~n9739 & n9742 ;
  assign n9744 = \u4_u3_buf1_reg[25]/P0001  & ~n2734 ;
  assign n9745 = \u1_u3_idin_reg[25]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9746 = ~n2733 & n9745 ;
  assign n9747 = ~n9744 & ~n9746 ;
  assign n9748 = ~n2732 & ~n9747 ;
  assign n9749 = \wb_data_i[25]_pad  & n2731 ;
  assign n9750 = n2567 & n9749 ;
  assign n9751 = rst_i_pad & ~n9750 ;
  assign n9752 = ~n9748 & n9751 ;
  assign n9753 = \u4_u3_buf1_reg[26]/P0001  & ~n2734 ;
  assign n9754 = \u1_u3_idin_reg[26]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9755 = ~n2733 & n9754 ;
  assign n9756 = ~n9753 & ~n9755 ;
  assign n9757 = ~n2732 & ~n9756 ;
  assign n9758 = \wb_data_i[26]_pad  & n2731 ;
  assign n9759 = n2567 & n9758 ;
  assign n9760 = rst_i_pad & ~n9759 ;
  assign n9761 = ~n9757 & n9760 ;
  assign n9762 = \u4_u3_buf1_reg[27]/P0001  & ~n2734 ;
  assign n9763 = \u1_u3_idin_reg[27]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9764 = ~n2733 & n9763 ;
  assign n9765 = ~n9762 & ~n9764 ;
  assign n9766 = ~n2732 & ~n9765 ;
  assign n9767 = \wb_data_i[27]_pad  & n2731 ;
  assign n9768 = n2567 & n9767 ;
  assign n9769 = rst_i_pad & ~n9768 ;
  assign n9770 = ~n9766 & n9769 ;
  assign n9771 = \u4_u3_buf1_reg[28]/P0001  & ~n2734 ;
  assign n9772 = \u1_u3_idin_reg[28]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9773 = ~n2733 & n9772 ;
  assign n9774 = ~n9771 & ~n9773 ;
  assign n9775 = ~n2732 & ~n9774 ;
  assign n9776 = \wb_data_i[28]_pad  & n2731 ;
  assign n9777 = n2567 & n9776 ;
  assign n9778 = rst_i_pad & ~n9777 ;
  assign n9779 = ~n9775 & n9778 ;
  assign n9780 = \u4_u3_buf1_reg[29]/P0001  & ~n2734 ;
  assign n9781 = \u1_u3_idin_reg[29]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9782 = ~n2733 & n9781 ;
  assign n9783 = ~n9780 & ~n9782 ;
  assign n9784 = ~n2732 & ~n9783 ;
  assign n9785 = \wb_data_i[29]_pad  & n2731 ;
  assign n9786 = n2567 & n9785 ;
  assign n9787 = rst_i_pad & ~n9786 ;
  assign n9788 = ~n9784 & n9787 ;
  assign n9789 = \u4_u3_buf1_reg[2]/P0001  & ~n2734 ;
  assign n9790 = \u1_u3_idin_reg[2]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9791 = ~n2733 & n9790 ;
  assign n9792 = ~n9789 & ~n9791 ;
  assign n9793 = ~n2732 & ~n9792 ;
  assign n9794 = \wb_data_i[2]_pad  & n2731 ;
  assign n9795 = n2567 & n9794 ;
  assign n9796 = rst_i_pad & ~n9795 ;
  assign n9797 = ~n9793 & n9796 ;
  assign n9798 = \u4_u3_buf1_reg[30]/P0001  & ~n2734 ;
  assign n9799 = \u1_u3_idin_reg[30]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9800 = ~n2733 & n9799 ;
  assign n9801 = ~n9798 & ~n9800 ;
  assign n9802 = ~n2732 & ~n9801 ;
  assign n9803 = \wb_data_i[30]_pad  & n2731 ;
  assign n9804 = n2567 & n9803 ;
  assign n9805 = rst_i_pad & ~n9804 ;
  assign n9806 = ~n9802 & n9805 ;
  assign n9807 = \u4_u3_buf1_reg[31]/P0001  & ~n2734 ;
  assign n9808 = \u1_u3_idin_reg[31]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9809 = ~n2733 & n9808 ;
  assign n9810 = ~n9807 & ~n9809 ;
  assign n9811 = ~n2732 & ~n9810 ;
  assign n9812 = \wb_data_i[31]_pad  & n2731 ;
  assign n9813 = n2567 & n9812 ;
  assign n9814 = rst_i_pad & ~n9813 ;
  assign n9815 = ~n9811 & n9814 ;
  assign n9816 = \u4_u3_buf1_reg[3]/P0001  & ~n2734 ;
  assign n9817 = \u1_u3_idin_reg[3]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9818 = ~n2733 & n9817 ;
  assign n9819 = ~n9816 & ~n9818 ;
  assign n9820 = ~n2732 & ~n9819 ;
  assign n9821 = \wb_data_i[3]_pad  & n2731 ;
  assign n9822 = n2567 & n9821 ;
  assign n9823 = rst_i_pad & ~n9822 ;
  assign n9824 = ~n9820 & n9823 ;
  assign n9825 = \u4_u3_buf1_reg[8]/P0001  & ~n2734 ;
  assign n9826 = \u1_u3_idin_reg[8]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9827 = ~n2733 & n9826 ;
  assign n9828 = ~n9825 & ~n9827 ;
  assign n9829 = ~n2732 & ~n9828 ;
  assign n9830 = \wb_data_i[8]_pad  & n2731 ;
  assign n9831 = n2567 & n9830 ;
  assign n9832 = rst_i_pad & ~n9831 ;
  assign n9833 = ~n9829 & n9832 ;
  assign n9834 = \u4_u3_buf1_reg[9]/P0001  & ~n2734 ;
  assign n9835 = \u1_u3_idin_reg[9]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n9836 = ~n2733 & n9835 ;
  assign n9837 = ~n9834 & ~n9836 ;
  assign n9838 = ~n2732 & ~n9837 ;
  assign n9839 = \wb_data_i[9]_pad  & n2731 ;
  assign n9840 = n2567 & n9839 ;
  assign n9841 = rst_i_pad & ~n9840 ;
  assign n9842 = ~n9838 & n9841 ;
  assign n9843 = \wb_addr_i[17]_pad  & n2564 ;
  assign n9844 = ~\u5_state_reg[1]/P0001  & ~n9843 ;
  assign n9845 = n8182 & ~n9844 ;
  assign n9846 = rst_i_pad & n9845 ;
  assign n9847 = \u5_state_reg[1]/P0001  & ~n8244 ;
  assign n9848 = ~\u1_u2_mack_r_reg/P0001  & \u5_state_reg[1]/P0001  ;
  assign n9849 = ~n8179 & n9848 ;
  assign n9850 = ~n9847 & ~n9849 ;
  assign n9851 = ~\u5_state_reg[2]/P0001  & n8186 ;
  assign n9852 = rst_i_pad & n9851 ;
  assign n9853 = ~n9850 & n9852 ;
  assign n9854 = ~n9846 & ~n9853 ;
  assign n9855 = ~\u1_u2_wr_last_reg/P0001  & ~n8066 ;
  assign n9856 = \u1_u2_rx_data_done_r2_reg/P0001  & ~\u1_u3_abort_reg/P0001  ;
  assign n9857 = \u1_u2_state_reg[2]/NET0131  & ~n9856 ;
  assign n9858 = ~\u1_u2_state_reg[2]/NET0131  & ~\u1_u2_state_reg[3]/NET0131  ;
  assign n9859 = \u1_u2_state_reg[2]/NET0131  & \u1_u2_state_reg[3]/NET0131  ;
  assign n9860 = ~n9858 & ~n9859 ;
  assign n9861 = ~n9857 & n9860 ;
  assign n9862 = n4071 & n9861 ;
  assign n9863 = ~\u1_u2_rx_data_valid_r_reg/NET0131  & ~n8127 ;
  assign n9864 = n9862 & n9863 ;
  assign n9865 = \u4_u0_buf1_reg[0]/P0001  & ~n2755 ;
  assign n9866 = \u1_u3_idin_reg[0]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9867 = ~n2733 & n9866 ;
  assign n9868 = ~n9865 & ~n9867 ;
  assign n9869 = ~n2754 & ~n9868 ;
  assign n9870 = n2587 & n9641 ;
  assign n9871 = rst_i_pad & ~n9870 ;
  assign n9872 = ~n9869 & n9871 ;
  assign n9873 = \u4_u0_buf1_reg[12]/P0001  & ~n2755 ;
  assign n9874 = \u1_u3_idin_reg[12]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9875 = ~n2733 & n9874 ;
  assign n9876 = ~n9873 & ~n9875 ;
  assign n9877 = ~n2754 & ~n9876 ;
  assign n9878 = n2587 & n9650 ;
  assign n9879 = rst_i_pad & ~n9878 ;
  assign n9880 = ~n9877 & n9879 ;
  assign n9881 = \u4_u0_buf1_reg[16]/P0001  & ~n2755 ;
  assign n9882 = \u1_u3_idin_reg[16]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9883 = ~n2733 & n9882 ;
  assign n9884 = ~n9881 & ~n9883 ;
  assign n9885 = ~n2754 & ~n9884 ;
  assign n9886 = n2587 & n9659 ;
  assign n9887 = rst_i_pad & ~n9886 ;
  assign n9888 = ~n9885 & n9887 ;
  assign n9889 = \u4_u0_buf1_reg[17]/P0001  & ~n2755 ;
  assign n9890 = \u1_u3_idin_reg[17]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9891 = ~n2733 & n9890 ;
  assign n9892 = ~n9889 & ~n9891 ;
  assign n9893 = ~n2754 & ~n9892 ;
  assign n9894 = n2587 & n9668 ;
  assign n9895 = rst_i_pad & ~n9894 ;
  assign n9896 = ~n9893 & n9895 ;
  assign n9897 = \u4_u0_buf1_reg[18]/P0001  & ~n2755 ;
  assign n9898 = \u1_u3_idin_reg[18]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9899 = ~n2733 & n9898 ;
  assign n9900 = ~n9897 & ~n9899 ;
  assign n9901 = ~n2754 & ~n9900 ;
  assign n9902 = n2587 & n9677 ;
  assign n9903 = rst_i_pad & ~n9902 ;
  assign n9904 = ~n9901 & n9903 ;
  assign n9905 = \u4_u0_buf1_reg[19]/P0001  & ~n2755 ;
  assign n9906 = \u1_u3_idin_reg[19]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9907 = ~n2733 & n9906 ;
  assign n9908 = ~n9905 & ~n9907 ;
  assign n9909 = ~n2754 & ~n9908 ;
  assign n9910 = n2587 & n9686 ;
  assign n9911 = rst_i_pad & ~n9910 ;
  assign n9912 = ~n9909 & n9911 ;
  assign n9913 = \u4_u0_buf1_reg[1]/P0001  & ~n2755 ;
  assign n9914 = \u1_u3_idin_reg[1]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9915 = ~n2733 & n9914 ;
  assign n9916 = ~n9913 & ~n9915 ;
  assign n9917 = ~n2754 & ~n9916 ;
  assign n9918 = n2587 & n9695 ;
  assign n9919 = rst_i_pad & ~n9918 ;
  assign n9920 = ~n9917 & n9919 ;
  assign n9921 = \u4_u0_buf1_reg[20]/P0001  & ~n2755 ;
  assign n9922 = \u1_u3_idin_reg[20]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9923 = ~n2733 & n9922 ;
  assign n9924 = ~n9921 & ~n9923 ;
  assign n9925 = ~n2754 & ~n9924 ;
  assign n9926 = n2587 & n9704 ;
  assign n9927 = rst_i_pad & ~n9926 ;
  assign n9928 = ~n9925 & n9927 ;
  assign n9929 = \u4_u0_buf1_reg[21]/P0001  & ~n2755 ;
  assign n9930 = \u1_u3_idin_reg[21]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9931 = ~n2733 & n9930 ;
  assign n9932 = ~n9929 & ~n9931 ;
  assign n9933 = ~n2754 & ~n9932 ;
  assign n9934 = n2587 & n9713 ;
  assign n9935 = rst_i_pad & ~n9934 ;
  assign n9936 = ~n9933 & n9935 ;
  assign n9937 = \u4_u0_buf1_reg[22]/P0001  & ~n2755 ;
  assign n9938 = \u1_u3_idin_reg[22]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9939 = ~n2733 & n9938 ;
  assign n9940 = ~n9937 & ~n9939 ;
  assign n9941 = ~n2754 & ~n9940 ;
  assign n9942 = n2587 & n9722 ;
  assign n9943 = rst_i_pad & ~n9942 ;
  assign n9944 = ~n9941 & n9943 ;
  assign n9945 = \u4_u0_buf1_reg[23]/P0001  & ~n2755 ;
  assign n9946 = \u1_u3_idin_reg[23]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9947 = ~n2733 & n9946 ;
  assign n9948 = ~n9945 & ~n9947 ;
  assign n9949 = ~n2754 & ~n9948 ;
  assign n9950 = n2587 & n9731 ;
  assign n9951 = rst_i_pad & ~n9950 ;
  assign n9952 = ~n9949 & n9951 ;
  assign n9953 = \u4_u0_buf1_reg[24]/P0001  & ~n2755 ;
  assign n9954 = \u1_u3_idin_reg[24]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9955 = ~n2733 & n9954 ;
  assign n9956 = ~n9953 & ~n9955 ;
  assign n9957 = ~n2754 & ~n9956 ;
  assign n9958 = n2587 & n9740 ;
  assign n9959 = rst_i_pad & ~n9958 ;
  assign n9960 = ~n9957 & n9959 ;
  assign n9961 = \u4_u0_buf1_reg[25]/P0001  & ~n2755 ;
  assign n9962 = \u1_u3_idin_reg[25]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n9963 = ~n2733 & n9962 ;
  assign n9964 = ~n9961 & ~n9963 ;
  assign n9965 = ~n2754 & ~n9964 ;
  assign n9966 = n2587 & n9749 ;
  assign n9967 = rst_i_pad & ~n9966 ;
  assign n9968 = ~n9965 & n9967 ;
  assign n9969 = ~\u4_buf1_reg[27]/P0001  & \u4_csr_reg[10]/P0001  ;
  assign n9970 = ~\u4_buf1_reg[26]/NET0131  & \u4_csr_reg[9]/NET0131  ;
  assign n9971 = ~n9969 & ~n9970 ;
  assign n9972 = ~\u4_buf1_reg[28]/P0001  & ~\u4_buf1_reg[29]/P0001  ;
  assign n9973 = \u4_buf1_reg[27]/P0001  & ~\u4_csr_reg[10]/P0001  ;
  assign n9974 = ~\u4_buf1_reg[30]/P0001  & ~n9973 ;
  assign n9975 = n9972 & n9974 ;
  assign n9976 = ~n9971 & n9975 ;
  assign n9977 = ~\u4_buf1_reg[25]/NET0131  & \u4_csr_reg[8]/P0001  ;
  assign n9978 = ~\u4_buf1_reg[24]/NET0131  & \u4_csr_reg[7]/P0001  ;
  assign n9979 = ~n9977 & ~n9978 ;
  assign n9980 = \u4_buf1_reg[23]/NET0131  & ~\u4_csr_reg[6]/NET0131  ;
  assign n9981 = \u4_buf1_reg[24]/NET0131  & ~\u4_csr_reg[7]/P0001  ;
  assign n9982 = ~n9980 & ~n9981 ;
  assign n9983 = n9979 & ~n9982 ;
  assign n9984 = \u4_buf1_reg[22]/NET0131  & ~\u4_csr_reg[5]/NET0131  ;
  assign n9985 = \u4_buf1_reg[21]/NET0131  & ~\u4_csr_reg[4]/NET0131  ;
  assign n9986 = ~n9984 & ~n9985 ;
  assign n9987 = ~\u4_buf1_reg[21]/NET0131  & \u4_csr_reg[4]/NET0131  ;
  assign n9988 = ~\u4_buf1_reg[20]/NET0131  & \u4_csr_reg[3]/P0001  ;
  assign n9989 = ~n9987 & ~n9988 ;
  assign n9990 = n9986 & ~n9989 ;
  assign n9991 = \u4_buf1_reg[18]/P0001  & ~\u4_csr_reg[1]/P0001  ;
  assign n9992 = ~\u4_buf1_reg[17]/NET0131  & \u4_csr_reg[0]/P0001  ;
  assign n9993 = ~n9991 & n9992 ;
  assign n9994 = ~\u4_buf1_reg[18]/P0001  & \u4_csr_reg[1]/P0001  ;
  assign n9995 = ~\u4_buf1_reg[19]/NET0131  & \u4_csr_reg[2]/NET0131  ;
  assign n9996 = ~n9994 & ~n9995 ;
  assign n9997 = ~n9993 & n9996 ;
  assign n9998 = \u4_buf1_reg[20]/NET0131  & ~\u4_csr_reg[3]/P0001  ;
  assign n9999 = \u4_buf1_reg[19]/NET0131  & ~\u4_csr_reg[2]/NET0131  ;
  assign n10000 = ~n9998 & ~n9999 ;
  assign n10001 = n9986 & n10000 ;
  assign n10002 = ~n9997 & n10001 ;
  assign n10003 = ~n9990 & ~n10002 ;
  assign n10004 = ~\u4_buf1_reg[23]/NET0131  & \u4_csr_reg[6]/NET0131  ;
  assign n10005 = ~\u4_buf1_reg[22]/NET0131  & \u4_csr_reg[5]/NET0131  ;
  assign n10006 = ~n10004 & ~n10005 ;
  assign n10007 = n9979 & n10006 ;
  assign n10008 = n10003 & n10007 ;
  assign n10009 = ~n9983 & ~n10008 ;
  assign n10010 = \u4_buf1_reg[25]/NET0131  & ~\u4_csr_reg[8]/P0001  ;
  assign n10011 = \u4_buf1_reg[26]/NET0131  & ~\u4_csr_reg[9]/NET0131  ;
  assign n10012 = ~n10010 & ~n10011 ;
  assign n10013 = n9975 & n10012 ;
  assign n10014 = n10009 & n10013 ;
  assign n10015 = ~n9976 & ~n10014 ;
  assign n10016 = \u4_u0_buf1_reg[26]/P0001  & ~n2755 ;
  assign n10017 = \u1_u3_idin_reg[26]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10018 = ~n2733 & n10017 ;
  assign n10019 = ~n10016 & ~n10018 ;
  assign n10020 = ~n2754 & ~n10019 ;
  assign n10021 = n2587 & n9758 ;
  assign n10022 = rst_i_pad & ~n10021 ;
  assign n10023 = ~n10020 & n10022 ;
  assign n10024 = \u4_u0_buf1_reg[27]/P0001  & ~n2755 ;
  assign n10025 = \u1_u3_idin_reg[27]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10026 = ~n2733 & n10025 ;
  assign n10027 = ~n10024 & ~n10026 ;
  assign n10028 = ~n2754 & ~n10027 ;
  assign n10029 = n2587 & n9767 ;
  assign n10030 = rst_i_pad & ~n10029 ;
  assign n10031 = ~n10028 & n10030 ;
  assign n10032 = \u4_u0_buf1_reg[28]/P0001  & ~n2755 ;
  assign n10033 = \u1_u3_idin_reg[28]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10034 = ~n2733 & n10033 ;
  assign n10035 = ~n10032 & ~n10034 ;
  assign n10036 = ~n2754 & ~n10035 ;
  assign n10037 = n2587 & n9776 ;
  assign n10038 = rst_i_pad & ~n10037 ;
  assign n10039 = ~n10036 & n10038 ;
  assign n10040 = \u4_u0_buf1_reg[29]/P0001  & ~n2755 ;
  assign n10041 = \u1_u3_idin_reg[29]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10042 = ~n2733 & n10041 ;
  assign n10043 = ~n10040 & ~n10042 ;
  assign n10044 = ~n2754 & ~n10043 ;
  assign n10045 = n2587 & n9785 ;
  assign n10046 = rst_i_pad & ~n10045 ;
  assign n10047 = ~n10044 & n10046 ;
  assign n10048 = \u4_u0_buf1_reg[2]/P0001  & ~n2755 ;
  assign n10049 = \u1_u3_idin_reg[2]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10050 = ~n2733 & n10049 ;
  assign n10051 = ~n10048 & ~n10050 ;
  assign n10052 = ~n2754 & ~n10051 ;
  assign n10053 = n2587 & n9794 ;
  assign n10054 = rst_i_pad & ~n10053 ;
  assign n10055 = ~n10052 & n10054 ;
  assign n10056 = \u4_u0_buf1_reg[30]/P0001  & ~n2755 ;
  assign n10057 = \u1_u3_idin_reg[30]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10058 = ~n2733 & n10057 ;
  assign n10059 = ~n10056 & ~n10058 ;
  assign n10060 = ~n2754 & ~n10059 ;
  assign n10061 = n2587 & n9803 ;
  assign n10062 = rst_i_pad & ~n10061 ;
  assign n10063 = ~n10060 & n10062 ;
  assign n10064 = \u4_u0_buf1_reg[31]/P0001  & ~n2755 ;
  assign n10065 = \u1_u3_idin_reg[31]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10066 = ~n2733 & n10065 ;
  assign n10067 = ~n10064 & ~n10066 ;
  assign n10068 = ~n2754 & ~n10067 ;
  assign n10069 = n2587 & n9812 ;
  assign n10070 = rst_i_pad & ~n10069 ;
  assign n10071 = ~n10068 & n10070 ;
  assign n10072 = \u4_u0_buf1_reg[3]/P0001  & ~n2755 ;
  assign n10073 = \u1_u3_idin_reg[3]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10074 = ~n2733 & n10073 ;
  assign n10075 = ~n10072 & ~n10074 ;
  assign n10076 = ~n2754 & ~n10075 ;
  assign n10077 = n2587 & n9821 ;
  assign n10078 = rst_i_pad & ~n10077 ;
  assign n10079 = ~n10076 & n10078 ;
  assign n10080 = \u4_u0_buf1_reg[8]/P0001  & ~n2755 ;
  assign n10081 = \u1_u3_idin_reg[8]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10082 = ~n2733 & n10081 ;
  assign n10083 = ~n10080 & ~n10082 ;
  assign n10084 = ~n2754 & ~n10083 ;
  assign n10085 = n2587 & n9830 ;
  assign n10086 = rst_i_pad & ~n10085 ;
  assign n10087 = ~n10084 & n10086 ;
  assign n10088 = \u4_u0_buf1_reg[9]/P0001  & ~n2755 ;
  assign n10089 = \u1_u3_idin_reg[9]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10090 = ~n2733 & n10089 ;
  assign n10091 = ~n10088 & ~n10090 ;
  assign n10092 = ~n2754 & ~n10091 ;
  assign n10093 = n2587 & n9839 ;
  assign n10094 = rst_i_pad & ~n10093 ;
  assign n10095 = ~n10092 & n10094 ;
  assign n10096 = ~\u0_u0_idle_cnt1_next_reg[7]/P0001  & n8674 ;
  assign n10097 = ~\u0_u0_idle_cnt1_reg[7]/P0001  & ~n8674 ;
  assign n10098 = n8673 & ~n10097 ;
  assign n10099 = ~n10096 & n10098 ;
  assign n10100 = ~n8672 & n10099 ;
  assign n10101 = ~n8666 & n10100 ;
  assign n10102 = \u4_u1_buf1_reg[0]/P0001  & ~n2775 ;
  assign n10103 = \u1_u3_idin_reg[0]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10104 = ~n2733 & n10103 ;
  assign n10105 = ~n10102 & ~n10104 ;
  assign n10106 = ~n2774 & ~n10105 ;
  assign n10107 = n2620 & n9641 ;
  assign n10108 = rst_i_pad & ~n10107 ;
  assign n10109 = ~n10106 & n10108 ;
  assign n10110 = \u4_u1_buf1_reg[12]/P0001  & ~n2775 ;
  assign n10111 = \u1_u3_idin_reg[12]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10112 = ~n2733 & n10111 ;
  assign n10113 = ~n10110 & ~n10112 ;
  assign n10114 = ~n2774 & ~n10113 ;
  assign n10115 = n2620 & n9650 ;
  assign n10116 = rst_i_pad & ~n10115 ;
  assign n10117 = ~n10114 & n10116 ;
  assign n10118 = \u4_u1_buf1_reg[16]/P0001  & ~n2775 ;
  assign n10119 = \u1_u3_idin_reg[16]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10120 = ~n2733 & n10119 ;
  assign n10121 = ~n10118 & ~n10120 ;
  assign n10122 = ~n2774 & ~n10121 ;
  assign n10123 = n2620 & n9659 ;
  assign n10124 = rst_i_pad & ~n10123 ;
  assign n10125 = ~n10122 & n10124 ;
  assign n10126 = \u4_u1_buf1_reg[17]/P0001  & ~n2775 ;
  assign n10127 = \u1_u3_idin_reg[17]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10128 = ~n2733 & n10127 ;
  assign n10129 = ~n10126 & ~n10128 ;
  assign n10130 = ~n2774 & ~n10129 ;
  assign n10131 = n2620 & n9668 ;
  assign n10132 = rst_i_pad & ~n10131 ;
  assign n10133 = ~n10130 & n10132 ;
  assign n10134 = \u4_u1_buf1_reg[18]/P0001  & ~n2775 ;
  assign n10135 = \u1_u3_idin_reg[18]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10136 = ~n2733 & n10135 ;
  assign n10137 = ~n10134 & ~n10136 ;
  assign n10138 = ~n2774 & ~n10137 ;
  assign n10139 = n2620 & n9677 ;
  assign n10140 = rst_i_pad & ~n10139 ;
  assign n10141 = ~n10138 & n10140 ;
  assign n10142 = \u4_u1_buf1_reg[19]/P0001  & ~n2775 ;
  assign n10143 = \u1_u3_idin_reg[19]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10144 = ~n2733 & n10143 ;
  assign n10145 = ~n10142 & ~n10144 ;
  assign n10146 = ~n2774 & ~n10145 ;
  assign n10147 = n2620 & n9686 ;
  assign n10148 = rst_i_pad & ~n10147 ;
  assign n10149 = ~n10146 & n10148 ;
  assign n10150 = \u4_u1_buf1_reg[1]/P0001  & ~n2775 ;
  assign n10151 = \u1_u3_idin_reg[1]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10152 = ~n2733 & n10151 ;
  assign n10153 = ~n10150 & ~n10152 ;
  assign n10154 = ~n2774 & ~n10153 ;
  assign n10155 = n2620 & n9695 ;
  assign n10156 = rst_i_pad & ~n10155 ;
  assign n10157 = ~n10154 & n10156 ;
  assign n10158 = \u4_u1_buf1_reg[20]/P0001  & ~n2775 ;
  assign n10159 = \u1_u3_idin_reg[20]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10160 = ~n2733 & n10159 ;
  assign n10161 = ~n10158 & ~n10160 ;
  assign n10162 = ~n2774 & ~n10161 ;
  assign n10163 = n2620 & n9704 ;
  assign n10164 = rst_i_pad & ~n10163 ;
  assign n10165 = ~n10162 & n10164 ;
  assign n10166 = \u4_u1_buf1_reg[21]/P0001  & ~n2775 ;
  assign n10167 = \u1_u3_idin_reg[21]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10168 = ~n2733 & n10167 ;
  assign n10169 = ~n10166 & ~n10168 ;
  assign n10170 = ~n2774 & ~n10169 ;
  assign n10171 = n2620 & n9713 ;
  assign n10172 = rst_i_pad & ~n10171 ;
  assign n10173 = ~n10170 & n10172 ;
  assign n10174 = \u4_u1_buf1_reg[22]/P0001  & ~n2775 ;
  assign n10175 = \u1_u3_idin_reg[22]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10176 = ~n2733 & n10175 ;
  assign n10177 = ~n10174 & ~n10176 ;
  assign n10178 = ~n2774 & ~n10177 ;
  assign n10179 = n2620 & n9722 ;
  assign n10180 = rst_i_pad & ~n10179 ;
  assign n10181 = ~n10178 & n10180 ;
  assign n10182 = \u4_u1_buf1_reg[23]/P0001  & ~n2775 ;
  assign n10183 = \u1_u3_idin_reg[23]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10184 = ~n2733 & n10183 ;
  assign n10185 = ~n10182 & ~n10184 ;
  assign n10186 = ~n2774 & ~n10185 ;
  assign n10187 = n2620 & n9731 ;
  assign n10188 = rst_i_pad & ~n10187 ;
  assign n10189 = ~n10186 & n10188 ;
  assign n10190 = \u4_u1_buf1_reg[24]/P0001  & ~n2775 ;
  assign n10191 = \u1_u3_idin_reg[24]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10192 = ~n2733 & n10191 ;
  assign n10193 = ~n10190 & ~n10192 ;
  assign n10194 = ~n2774 & ~n10193 ;
  assign n10195 = n2620 & n9740 ;
  assign n10196 = rst_i_pad & ~n10195 ;
  assign n10197 = ~n10194 & n10196 ;
  assign n10198 = \u4_u1_buf1_reg[25]/P0001  & ~n2775 ;
  assign n10199 = \u1_u3_idin_reg[25]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10200 = ~n2733 & n10199 ;
  assign n10201 = ~n10198 & ~n10200 ;
  assign n10202 = ~n2774 & ~n10201 ;
  assign n10203 = n2620 & n9749 ;
  assign n10204 = rst_i_pad & ~n10203 ;
  assign n10205 = ~n10202 & n10204 ;
  assign n10206 = \u4_u1_buf1_reg[26]/P0001  & ~n2775 ;
  assign n10207 = \u1_u3_idin_reg[26]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10208 = ~n2733 & n10207 ;
  assign n10209 = ~n10206 & ~n10208 ;
  assign n10210 = ~n2774 & ~n10209 ;
  assign n10211 = n2620 & n9758 ;
  assign n10212 = rst_i_pad & ~n10211 ;
  assign n10213 = ~n10210 & n10212 ;
  assign n10214 = \u4_u1_buf1_reg[27]/P0001  & ~n2775 ;
  assign n10215 = \u1_u3_idin_reg[27]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10216 = ~n2733 & n10215 ;
  assign n10217 = ~n10214 & ~n10216 ;
  assign n10218 = ~n2774 & ~n10217 ;
  assign n10219 = n2620 & n9767 ;
  assign n10220 = rst_i_pad & ~n10219 ;
  assign n10221 = ~n10218 & n10220 ;
  assign n10222 = \u4_u1_buf1_reg[28]/P0001  & ~n2775 ;
  assign n10223 = \u1_u3_idin_reg[28]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10224 = ~n2733 & n10223 ;
  assign n10225 = ~n10222 & ~n10224 ;
  assign n10226 = ~n2774 & ~n10225 ;
  assign n10227 = n2620 & n9776 ;
  assign n10228 = rst_i_pad & ~n10227 ;
  assign n10229 = ~n10226 & n10228 ;
  assign n10230 = \u4_u1_buf1_reg[29]/P0001  & ~n2775 ;
  assign n10231 = \u1_u3_idin_reg[29]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10232 = ~n2733 & n10231 ;
  assign n10233 = ~n10230 & ~n10232 ;
  assign n10234 = ~n2774 & ~n10233 ;
  assign n10235 = n2620 & n9785 ;
  assign n10236 = rst_i_pad & ~n10235 ;
  assign n10237 = ~n10234 & n10236 ;
  assign n10238 = \u4_u1_buf1_reg[2]/P0001  & ~n2775 ;
  assign n10239 = \u1_u3_idin_reg[2]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10240 = ~n2733 & n10239 ;
  assign n10241 = ~n10238 & ~n10240 ;
  assign n10242 = ~n2774 & ~n10241 ;
  assign n10243 = n2620 & n9794 ;
  assign n10244 = rst_i_pad & ~n10243 ;
  assign n10245 = ~n10242 & n10244 ;
  assign n10246 = \u4_u1_buf1_reg[30]/P0001  & ~n2775 ;
  assign n10247 = \u1_u3_idin_reg[30]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10248 = ~n2733 & n10247 ;
  assign n10249 = ~n10246 & ~n10248 ;
  assign n10250 = ~n2774 & ~n10249 ;
  assign n10251 = n2620 & n9803 ;
  assign n10252 = rst_i_pad & ~n10251 ;
  assign n10253 = ~n10250 & n10252 ;
  assign n10254 = \u4_u1_buf1_reg[31]/P0001  & ~n2775 ;
  assign n10255 = \u1_u3_idin_reg[31]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10256 = ~n2733 & n10255 ;
  assign n10257 = ~n10254 & ~n10256 ;
  assign n10258 = ~n2774 & ~n10257 ;
  assign n10259 = n2620 & n9812 ;
  assign n10260 = rst_i_pad & ~n10259 ;
  assign n10261 = ~n10258 & n10260 ;
  assign n10262 = \u4_u1_buf1_reg[3]/P0001  & ~n2775 ;
  assign n10263 = \u1_u3_idin_reg[3]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10264 = ~n2733 & n10263 ;
  assign n10265 = ~n10262 & ~n10264 ;
  assign n10266 = ~n2774 & ~n10265 ;
  assign n10267 = n2620 & n9821 ;
  assign n10268 = rst_i_pad & ~n10267 ;
  assign n10269 = ~n10266 & n10268 ;
  assign n10270 = \u4_u1_buf1_reg[8]/P0001  & ~n2775 ;
  assign n10271 = \u1_u3_idin_reg[8]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10272 = ~n2733 & n10271 ;
  assign n10273 = ~n10270 & ~n10272 ;
  assign n10274 = ~n2774 & ~n10273 ;
  assign n10275 = n2620 & n9830 ;
  assign n10276 = rst_i_pad & ~n10275 ;
  assign n10277 = ~n10274 & n10276 ;
  assign n10278 = \u4_u1_buf1_reg[9]/P0001  & ~n2775 ;
  assign n10279 = \u1_u3_idin_reg[9]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10280 = ~n2733 & n10279 ;
  assign n10281 = ~n10278 & ~n10280 ;
  assign n10282 = ~n2774 & ~n10281 ;
  assign n10283 = n2620 & n9839 ;
  assign n10284 = rst_i_pad & ~n10283 ;
  assign n10285 = ~n10282 & n10284 ;
  assign n10286 = \u4_u2_buf1_reg[0]/P0001  & ~n2811 ;
  assign n10287 = \u1_u3_idin_reg[0]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10288 = ~n2733 & n10287 ;
  assign n10289 = ~n10286 & ~n10288 ;
  assign n10290 = ~n2810 & ~n10289 ;
  assign n10291 = n2635 & n9641 ;
  assign n10292 = rst_i_pad & ~n10291 ;
  assign n10293 = ~n10290 & n10292 ;
  assign n10294 = \u4_u2_buf1_reg[12]/P0001  & ~n2811 ;
  assign n10295 = \u1_u3_idin_reg[12]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10296 = ~n2733 & n10295 ;
  assign n10297 = ~n10294 & ~n10296 ;
  assign n10298 = ~n2810 & ~n10297 ;
  assign n10299 = n2635 & n9650 ;
  assign n10300 = rst_i_pad & ~n10299 ;
  assign n10301 = ~n10298 & n10300 ;
  assign n10302 = \u4_u2_buf1_reg[16]/P0001  & ~n2811 ;
  assign n10303 = \u1_u3_idin_reg[16]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10304 = ~n2733 & n10303 ;
  assign n10305 = ~n10302 & ~n10304 ;
  assign n10306 = ~n2810 & ~n10305 ;
  assign n10307 = n2635 & n9659 ;
  assign n10308 = rst_i_pad & ~n10307 ;
  assign n10309 = ~n10306 & n10308 ;
  assign n10310 = \u4_u2_buf1_reg[17]/P0001  & ~n2811 ;
  assign n10311 = \u1_u3_idin_reg[17]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10312 = ~n2733 & n10311 ;
  assign n10313 = ~n10310 & ~n10312 ;
  assign n10314 = ~n2810 & ~n10313 ;
  assign n10315 = n2635 & n9668 ;
  assign n10316 = rst_i_pad & ~n10315 ;
  assign n10317 = ~n10314 & n10316 ;
  assign n10318 = \u4_u2_buf1_reg[18]/P0001  & ~n2811 ;
  assign n10319 = \u1_u3_idin_reg[18]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10320 = ~n2733 & n10319 ;
  assign n10321 = ~n10318 & ~n10320 ;
  assign n10322 = ~n2810 & ~n10321 ;
  assign n10323 = n2635 & n9677 ;
  assign n10324 = rst_i_pad & ~n10323 ;
  assign n10325 = ~n10322 & n10324 ;
  assign n10326 = \u4_u2_buf1_reg[19]/P0001  & ~n2811 ;
  assign n10327 = \u1_u3_idin_reg[19]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10328 = ~n2733 & n10327 ;
  assign n10329 = ~n10326 & ~n10328 ;
  assign n10330 = ~n2810 & ~n10329 ;
  assign n10331 = n2635 & n9686 ;
  assign n10332 = rst_i_pad & ~n10331 ;
  assign n10333 = ~n10330 & n10332 ;
  assign n10334 = \u4_u2_buf1_reg[1]/P0001  & ~n2811 ;
  assign n10335 = \u1_u3_idin_reg[1]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10336 = ~n2733 & n10335 ;
  assign n10337 = ~n10334 & ~n10336 ;
  assign n10338 = ~n2810 & ~n10337 ;
  assign n10339 = n2635 & n9695 ;
  assign n10340 = rst_i_pad & ~n10339 ;
  assign n10341 = ~n10338 & n10340 ;
  assign n10342 = \u4_u2_buf1_reg[20]/P0001  & ~n2811 ;
  assign n10343 = \u1_u3_idin_reg[20]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10344 = ~n2733 & n10343 ;
  assign n10345 = ~n10342 & ~n10344 ;
  assign n10346 = ~n2810 & ~n10345 ;
  assign n10347 = n2635 & n9704 ;
  assign n10348 = rst_i_pad & ~n10347 ;
  assign n10349 = ~n10346 & n10348 ;
  assign n10350 = \u4_u2_buf1_reg[21]/P0001  & ~n2811 ;
  assign n10351 = \u1_u3_idin_reg[21]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10352 = ~n2733 & n10351 ;
  assign n10353 = ~n10350 & ~n10352 ;
  assign n10354 = ~n2810 & ~n10353 ;
  assign n10355 = n2635 & n9713 ;
  assign n10356 = rst_i_pad & ~n10355 ;
  assign n10357 = ~n10354 & n10356 ;
  assign n10358 = \u4_u2_buf1_reg[22]/P0001  & ~n2811 ;
  assign n10359 = \u1_u3_idin_reg[22]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10360 = ~n2733 & n10359 ;
  assign n10361 = ~n10358 & ~n10360 ;
  assign n10362 = ~n2810 & ~n10361 ;
  assign n10363 = n2635 & n9722 ;
  assign n10364 = rst_i_pad & ~n10363 ;
  assign n10365 = ~n10362 & n10364 ;
  assign n10366 = \u4_u2_buf1_reg[23]/P0001  & ~n2811 ;
  assign n10367 = \u1_u3_idin_reg[23]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10368 = ~n2733 & n10367 ;
  assign n10369 = ~n10366 & ~n10368 ;
  assign n10370 = ~n2810 & ~n10369 ;
  assign n10371 = n2635 & n9731 ;
  assign n10372 = rst_i_pad & ~n10371 ;
  assign n10373 = ~n10370 & n10372 ;
  assign n10374 = \u4_u2_buf1_reg[24]/P0001  & ~n2811 ;
  assign n10375 = \u1_u3_idin_reg[24]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10376 = ~n2733 & n10375 ;
  assign n10377 = ~n10374 & ~n10376 ;
  assign n10378 = ~n2810 & ~n10377 ;
  assign n10379 = n2635 & n9740 ;
  assign n10380 = rst_i_pad & ~n10379 ;
  assign n10381 = ~n10378 & n10380 ;
  assign n10382 = \u4_u2_buf1_reg[25]/P0001  & ~n2811 ;
  assign n10383 = \u1_u3_idin_reg[25]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10384 = ~n2733 & n10383 ;
  assign n10385 = ~n10382 & ~n10384 ;
  assign n10386 = ~n2810 & ~n10385 ;
  assign n10387 = n2635 & n9749 ;
  assign n10388 = rst_i_pad & ~n10387 ;
  assign n10389 = ~n10386 & n10388 ;
  assign n10390 = \u4_u2_buf1_reg[26]/P0001  & ~n2811 ;
  assign n10391 = \u1_u3_idin_reg[26]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10392 = ~n2733 & n10391 ;
  assign n10393 = ~n10390 & ~n10392 ;
  assign n10394 = ~n2810 & ~n10393 ;
  assign n10395 = n2635 & n9758 ;
  assign n10396 = rst_i_pad & ~n10395 ;
  assign n10397 = ~n10394 & n10396 ;
  assign n10398 = \u4_u2_buf1_reg[27]/P0001  & ~n2811 ;
  assign n10399 = \u1_u3_idin_reg[27]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10400 = ~n2733 & n10399 ;
  assign n10401 = ~n10398 & ~n10400 ;
  assign n10402 = ~n2810 & ~n10401 ;
  assign n10403 = n2635 & n9767 ;
  assign n10404 = rst_i_pad & ~n10403 ;
  assign n10405 = ~n10402 & n10404 ;
  assign n10406 = \u4_u2_buf1_reg[28]/P0001  & ~n2811 ;
  assign n10407 = \u1_u3_idin_reg[28]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10408 = ~n2733 & n10407 ;
  assign n10409 = ~n10406 & ~n10408 ;
  assign n10410 = ~n2810 & ~n10409 ;
  assign n10411 = n2635 & n9776 ;
  assign n10412 = rst_i_pad & ~n10411 ;
  assign n10413 = ~n10410 & n10412 ;
  assign n10414 = \u4_u2_buf1_reg[29]/P0001  & ~n2811 ;
  assign n10415 = \u1_u3_idin_reg[29]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10416 = ~n2733 & n10415 ;
  assign n10417 = ~n10414 & ~n10416 ;
  assign n10418 = ~n2810 & ~n10417 ;
  assign n10419 = n2635 & n9785 ;
  assign n10420 = rst_i_pad & ~n10419 ;
  assign n10421 = ~n10418 & n10420 ;
  assign n10422 = \u4_u2_buf1_reg[2]/P0001  & ~n2811 ;
  assign n10423 = \u1_u3_idin_reg[2]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10424 = ~n2733 & n10423 ;
  assign n10425 = ~n10422 & ~n10424 ;
  assign n10426 = ~n2810 & ~n10425 ;
  assign n10427 = n2635 & n9794 ;
  assign n10428 = rst_i_pad & ~n10427 ;
  assign n10429 = ~n10426 & n10428 ;
  assign n10430 = \u4_u2_buf1_reg[30]/P0001  & ~n2811 ;
  assign n10431 = \u1_u3_idin_reg[30]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10432 = ~n2733 & n10431 ;
  assign n10433 = ~n10430 & ~n10432 ;
  assign n10434 = ~n2810 & ~n10433 ;
  assign n10435 = n2635 & n9803 ;
  assign n10436 = rst_i_pad & ~n10435 ;
  assign n10437 = ~n10434 & n10436 ;
  assign n10438 = \u4_u2_buf1_reg[31]/P0001  & ~n2811 ;
  assign n10439 = \u1_u3_idin_reg[31]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10440 = ~n2733 & n10439 ;
  assign n10441 = ~n10438 & ~n10440 ;
  assign n10442 = ~n2810 & ~n10441 ;
  assign n10443 = n2635 & n9812 ;
  assign n10444 = rst_i_pad & ~n10443 ;
  assign n10445 = ~n10442 & n10444 ;
  assign n10446 = \u4_u2_buf1_reg[3]/P0001  & ~n2811 ;
  assign n10447 = \u1_u3_idin_reg[3]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10448 = ~n2733 & n10447 ;
  assign n10449 = ~n10446 & ~n10448 ;
  assign n10450 = ~n2810 & ~n10449 ;
  assign n10451 = n2635 & n9821 ;
  assign n10452 = rst_i_pad & ~n10451 ;
  assign n10453 = ~n10450 & n10452 ;
  assign n10454 = \u4_u2_buf1_reg[8]/P0001  & ~n2811 ;
  assign n10455 = \u1_u3_idin_reg[8]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10456 = ~n2733 & n10455 ;
  assign n10457 = ~n10454 & ~n10456 ;
  assign n10458 = ~n2810 & ~n10457 ;
  assign n10459 = n2635 & n9830 ;
  assign n10460 = rst_i_pad & ~n10459 ;
  assign n10461 = ~n10458 & n10460 ;
  assign n10462 = \u4_u2_buf1_reg[9]/P0001  & ~n2811 ;
  assign n10463 = \u1_u3_idin_reg[9]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10464 = ~n2733 & n10463 ;
  assign n10465 = ~n10462 & ~n10464 ;
  assign n10466 = ~n2810 & ~n10465 ;
  assign n10467 = n2635 & n9839 ;
  assign n10468 = rst_i_pad & ~n10467 ;
  assign n10469 = ~n10466 & n10468 ;
  assign n10470 = n7202 & n7207 ;
  assign n10471 = \u1_u0_state_reg[0]/P0001  & ~\u1_u0_state_reg[2]/P0001  ;
  assign n10472 = rst_i_pad & n10471 ;
  assign n10473 = n10470 & n10472 ;
  assign n10474 = ~n7198 & n7807 ;
  assign n10475 = n7200 & ~n10474 ;
  assign n10476 = ~n4958 & n7203 ;
  assign n10477 = ~n7204 & n10476 ;
  assign n10478 = \u0_rx_active_reg/P0001  & \u1_u0_state_reg[1]/P0001  ;
  assign n10479 = rst_i_pad & n10478 ;
  assign n10480 = ~n10477 & n10479 ;
  assign n10481 = n10475 & n10480 ;
  assign n10482 = ~n10473 & ~n10481 ;
  assign n10483 = \u0_rx_data_reg[6]/P0001  & ~\u0_rx_data_reg[7]/P0001  ;
  assign n10484 = ~\u0_rx_data_reg[6]/P0001  & \u0_rx_data_reg[7]/P0001  ;
  assign n10485 = ~n10483 & ~n10484 ;
  assign n10486 = \u1_u0_crc16_sum_reg[8]/P0001  & ~n10485 ;
  assign n10487 = ~\u1_u0_crc16_sum_reg[8]/P0001  & n10485 ;
  assign n10488 = ~n10486 & ~n10487 ;
  assign n10489 = \u0_rx_data_reg[2]/P0001  & ~\u0_rx_data_reg[3]/P0001  ;
  assign n10490 = ~\u0_rx_data_reg[2]/P0001  & \u0_rx_data_reg[3]/P0001  ;
  assign n10491 = ~n10489 & ~n10490 ;
  assign n10492 = \u0_rx_data_reg[0]/P0001  & ~\u0_rx_data_reg[1]/P0001  ;
  assign n10493 = ~\u0_rx_data_reg[0]/P0001  & \u0_rx_data_reg[1]/P0001  ;
  assign n10494 = ~n10492 & ~n10493 ;
  assign n10495 = ~n10491 & ~n10494 ;
  assign n10496 = n10491 & n10494 ;
  assign n10497 = ~n10495 & ~n10496 ;
  assign n10498 = \u0_rx_data_reg[4]/P0001  & ~\u0_rx_data_reg[5]/P0001  ;
  assign n10499 = ~\u0_rx_data_reg[4]/P0001  & \u0_rx_data_reg[5]/P0001  ;
  assign n10500 = ~n10498 & ~n10499 ;
  assign n10501 = ~\u1_u0_crc16_sum_reg[15]/P0001  & ~\u1_u0_crc16_sum_reg[7]/P0001  ;
  assign n10502 = \u1_u0_crc16_sum_reg[15]/P0001  & \u1_u0_crc16_sum_reg[7]/P0001  ;
  assign n10503 = ~n10501 & ~n10502 ;
  assign n10504 = n10500 & ~n10503 ;
  assign n10505 = ~n10497 & n10504 ;
  assign n10506 = ~n10500 & ~n10503 ;
  assign n10507 = n10497 & n10506 ;
  assign n10508 = ~n10505 & ~n10507 ;
  assign n10509 = ~n10500 & n10503 ;
  assign n10510 = ~n10497 & n10509 ;
  assign n10511 = n10500 & n10503 ;
  assign n10512 = n10497 & n10511 ;
  assign n10513 = ~n10510 & ~n10512 ;
  assign n10514 = n10508 & n10513 ;
  assign n10515 = ~n10488 & ~n10514 ;
  assign n10516 = n10488 & n10514 ;
  assign n10517 = ~n10515 & ~n10516 ;
  assign n10518 = n7200 & n7806 ;
  assign n10519 = ~n7198 & n10518 ;
  assign n10520 = ~n4911 & ~n10519 ;
  assign n10521 = n7203 & ~n10520 ;
  assign n10522 = \u1_u0_crc16_sum_reg[11]/P0001  & ~\u1_u0_crc16_sum_reg[12]/P0001  ;
  assign n10523 = ~\u1_u0_crc16_sum_reg[11]/P0001  & \u1_u0_crc16_sum_reg[12]/P0001  ;
  assign n10524 = ~n10522 & ~n10523 ;
  assign n10525 = \u1_u0_crc16_sum_reg[10]/P0001  & ~\u1_u0_crc16_sum_reg[9]/P0001  ;
  assign n10526 = ~\u1_u0_crc16_sum_reg[10]/P0001  & \u1_u0_crc16_sum_reg[9]/P0001  ;
  assign n10527 = ~n10525 & ~n10526 ;
  assign n10528 = \u1_u0_crc16_sum_reg[13]/P0001  & ~\u1_u0_crc16_sum_reg[14]/P0001  ;
  assign n10529 = ~\u1_u0_crc16_sum_reg[13]/P0001  & \u1_u0_crc16_sum_reg[14]/P0001  ;
  assign n10530 = ~n10528 & ~n10529 ;
  assign n10531 = n10527 & n10530 ;
  assign n10532 = ~n10527 & ~n10530 ;
  assign n10533 = ~n10531 & ~n10532 ;
  assign n10534 = n10524 & n10533 ;
  assign n10535 = ~n10524 & ~n10533 ;
  assign n10536 = ~n10534 & ~n10535 ;
  assign n10537 = n10521 & ~n10536 ;
  assign n10538 = ~n10517 & n10537 ;
  assign n10539 = n10521 & n10536 ;
  assign n10540 = ~n10497 & ~n10500 ;
  assign n10541 = n10497 & n10500 ;
  assign n10542 = ~n10540 & ~n10541 ;
  assign n10543 = \u1_u0_crc16_sum_reg[8]/P0001  & ~n10503 ;
  assign n10544 = ~\u1_u0_crc16_sum_reg[8]/P0001  & n10503 ;
  assign n10545 = ~n10543 & ~n10544 ;
  assign n10546 = ~n10485 & ~n10545 ;
  assign n10547 = n10485 & n10545 ;
  assign n10548 = ~n10546 & ~n10547 ;
  assign n10549 = n10542 & ~n10548 ;
  assign n10550 = ~n10542 & n10548 ;
  assign n10551 = ~n10549 & ~n10550 ;
  assign n10552 = n10539 & n10551 ;
  assign n10553 = \u0_rx_active_reg/P0001  & ~\u1_u0_rx_active_r_reg/P0001  ;
  assign n10554 = \u1_u0_crc16_sum_reg[15]/P0001  & ~n7203 ;
  assign n10555 = \u1_u0_crc16_sum_reg[15]/P0001  & ~n4911 ;
  assign n10556 = ~n10519 & n10555 ;
  assign n10557 = ~n10554 & ~n10556 ;
  assign n10558 = ~n10553 & n10557 ;
  assign n10559 = ~n10552 & n10558 ;
  assign n10560 = ~n10538 & n10559 ;
  assign n10561 = \u1_u0_crc16_sum_reg[12]/P0001  & \u1_u0_crc16_sum_reg[13]/P0001  ;
  assign n10562 = ~n4925 & ~n10561 ;
  assign n10563 = \u1_u0_crc16_sum_reg[14]/P0001  & ~\u1_u0_crc16_sum_reg[15]/P0001  ;
  assign n10564 = ~n4921 & ~n10563 ;
  assign n10565 = ~\u1_u0_crc16_sum_reg[9]/P0001  & ~n10564 ;
  assign n10566 = ~n10562 & n10565 ;
  assign n10567 = ~n10497 & n10566 ;
  assign n10568 = \u1_u0_crc16_sum_reg[9]/P0001  & ~n10564 ;
  assign n10569 = n10562 & n10568 ;
  assign n10570 = ~n10497 & n10569 ;
  assign n10571 = ~n10567 & ~n10570 ;
  assign n10572 = ~n10562 & n10568 ;
  assign n10573 = n10497 & n10572 ;
  assign n10574 = n10562 & n10565 ;
  assign n10575 = n10497 & n10574 ;
  assign n10576 = ~n10573 & ~n10575 ;
  assign n10577 = n10571 & n10576 ;
  assign n10578 = \u1_u0_crc16_sum_reg[9]/P0001  & n10564 ;
  assign n10579 = ~n10562 & n10578 ;
  assign n10580 = ~n10497 & n10579 ;
  assign n10581 = ~\u1_u0_crc16_sum_reg[9]/P0001  & n10564 ;
  assign n10582 = n10562 & n10581 ;
  assign n10583 = ~n10497 & n10582 ;
  assign n10584 = ~n10580 & ~n10583 ;
  assign n10585 = ~n10562 & n10581 ;
  assign n10586 = n10497 & n10585 ;
  assign n10587 = n10562 & n10578 ;
  assign n10588 = n10497 & n10587 ;
  assign n10589 = ~n10586 & ~n10588 ;
  assign n10590 = n10584 & n10589 ;
  assign n10591 = n10577 & n10590 ;
  assign n10592 = \u1_u0_crc16_sum_reg[10]/P0001  & \u1_u0_crc16_sum_reg[11]/P0001  ;
  assign n10593 = ~n4924 & ~n10592 ;
  assign n10594 = ~n10500 & ~n10593 ;
  assign n10595 = n10500 & n10593 ;
  assign n10596 = ~n10594 & ~n10595 ;
  assign n10597 = ~\u0_rx_data_reg[6]/P0001  & ~n10596 ;
  assign n10598 = \u0_rx_data_reg[6]/P0001  & n10596 ;
  assign n10599 = ~n10597 & ~n10598 ;
  assign n10600 = n10521 & n10599 ;
  assign n10601 = ~n10591 & n10600 ;
  assign n10602 = n10521 & ~n10599 ;
  assign n10603 = \u1_u0_crc16_sum_reg[9]/P0001  & ~n10497 ;
  assign n10604 = ~\u1_u0_crc16_sum_reg[9]/P0001  & n10497 ;
  assign n10605 = ~n10603 & ~n10604 ;
  assign n10606 = ~n10562 & ~n10564 ;
  assign n10607 = n10562 & n10564 ;
  assign n10608 = ~n10606 & ~n10607 ;
  assign n10609 = n10605 & ~n10608 ;
  assign n10610 = ~n10605 & n10608 ;
  assign n10611 = ~n10609 & ~n10610 ;
  assign n10612 = n10602 & n10611 ;
  assign n10613 = ~n10601 & ~n10612 ;
  assign n10614 = \u1_u0_crc16_sum_reg[1]/P0001  & ~n4911 ;
  assign n10615 = ~n10519 & n10614 ;
  assign n10616 = \u1_u0_crc16_sum_reg[1]/P0001  & ~n7203 ;
  assign n10617 = ~n10553 & ~n10616 ;
  assign n10618 = ~n10615 & n10617 ;
  assign n10619 = n10613 & n10618 ;
  assign n10620 = \u0_rx_active_reg/P0001  & ~\u1_u0_state_reg[0]/P0001  ;
  assign n10621 = ~n10477 & ~n10620 ;
  assign n10622 = n10475 & n10621 ;
  assign n10623 = n4911 & ~n10620 ;
  assign n10624 = n7203 & n7209 ;
  assign n10625 = rst_i_pad & ~n10624 ;
  assign n10626 = ~n10623 & n10625 ;
  assign n10627 = \u1_u0_state_reg[0]/P0001  & \u1_u0_state_reg[2]/P0001  ;
  assign n10628 = n7207 & ~n10627 ;
  assign n10629 = ~n4909 & ~n10620 ;
  assign n10630 = n10628 & n10629 ;
  assign n10631 = ~n7202 & n10630 ;
  assign n10632 = n10626 & ~n10631 ;
  assign n10633 = ~n10622 & n10632 ;
  assign n10634 = n8188 & n8244 ;
  assign n10635 = ~n8509 & ~n10634 ;
  assign n10636 = ~\u1_u2_mack_r_reg/P0001  & ~n8509 ;
  assign n10637 = ~n8179 & n10636 ;
  assign n10638 = ~n10635 & ~n10637 ;
  assign n10639 = ~n4435 & ~n4443 ;
  assign n10640 = n4442 & ~n10639 ;
  assign n10641 = ~n4442 & n10639 ;
  assign n10642 = ~n10640 & ~n10641 ;
  assign n10643 = ~n4435 & ~n4438 ;
  assign n10644 = ~n4441 & n10643 ;
  assign n10645 = ~n4433 & ~n4434 ;
  assign n10646 = ~n4443 & n10645 ;
  assign n10647 = ~n10644 & n10646 ;
  assign n10648 = ~n4443 & ~n10644 ;
  assign n10649 = ~n10645 & ~n10648 ;
  assign n10650 = ~n10647 & ~n10649 ;
  assign n10651 = \u4_int_srcb_reg[4]/P0001  & \u4_inta_msk_reg[4]/P0001  ;
  assign n10652 = \u4_int_srcb_reg[6]/P0001  & \u4_inta_msk_reg[6]/P0001  ;
  assign n10653 = ~n10651 & ~n10652 ;
  assign n10654 = \u4_int_srcb_reg[5]/P0001  & \u4_inta_msk_reg[5]/P0001  ;
  assign n10655 = \u4_int_srcb_reg[7]/P0001  & \u4_inta_msk_reg[7]/P0001  ;
  assign n10656 = ~n10654 & ~n10655 ;
  assign n10657 = n10653 & n10656 ;
  assign n10658 = ~\u4_u2_inta_reg/P0001  & ~\u4_u3_inta_reg/P0001  ;
  assign n10659 = ~\u4_u0_inta_reg/P0001  & ~\u4_u1_inta_reg/P0001  ;
  assign n10660 = n10658 & n10659 ;
  assign n10661 = \u4_int_srcb_reg[0]/P0001  & \u4_inta_msk_reg[0]/P0001  ;
  assign n10662 = \u4_int_srcb_reg[3]/P0001  & \u4_inta_msk_reg[3]/P0001  ;
  assign n10663 = ~n10661 & ~n10662 ;
  assign n10664 = n10660 & n10663 ;
  assign n10665 = n10657 & n10664 ;
  assign n10666 = \u4_int_srcb_reg[8]/P0001  & \u4_inta_msk_reg[8]/P0001  ;
  assign n10667 = \u4_int_srcb_reg[2]/P0001  & \u4_inta_msk_reg[2]/P0001  ;
  assign n10668 = ~n10666 & ~n10667 ;
  assign n10669 = \u4_int_srcb_reg[1]/P0001  & \u4_inta_msk_reg[1]/P0001  ;
  assign n10670 = n10668 & ~n10669 ;
  assign n10671 = n10665 & n10670 ;
  assign n10672 = \u4_int_srcb_reg[4]/P0001  & \u4_intb_msk_reg[4]/P0001  ;
  assign n10673 = \u4_int_srcb_reg[6]/P0001  & \u4_intb_msk_reg[6]/P0001  ;
  assign n10674 = ~n10672 & ~n10673 ;
  assign n10675 = \u4_int_srcb_reg[5]/P0001  & \u4_intb_msk_reg[5]/P0001  ;
  assign n10676 = \u4_int_srcb_reg[7]/P0001  & \u4_intb_msk_reg[7]/P0001  ;
  assign n10677 = ~n10675 & ~n10676 ;
  assign n10678 = n10674 & n10677 ;
  assign n10679 = ~\u4_u2_intb_reg/P0001  & ~\u4_u3_intb_reg/P0001  ;
  assign n10680 = ~\u4_u0_intb_reg/P0001  & ~\u4_u1_intb_reg/P0001  ;
  assign n10681 = n10679 & n10680 ;
  assign n10682 = \u4_int_srcb_reg[0]/P0001  & \u4_intb_msk_reg[0]/P0001  ;
  assign n10683 = \u4_int_srcb_reg[3]/P0001  & \u4_intb_msk_reg[3]/P0001  ;
  assign n10684 = ~n10682 & ~n10683 ;
  assign n10685 = n10681 & n10684 ;
  assign n10686 = n10678 & n10685 ;
  assign n10687 = \u4_int_srcb_reg[8]/P0001  & \u4_intb_msk_reg[8]/P0001  ;
  assign n10688 = \u4_int_srcb_reg[2]/P0001  & \u4_intb_msk_reg[2]/P0001  ;
  assign n10689 = ~n10687 & ~n10688 ;
  assign n10690 = \u4_int_srcb_reg[1]/P0001  & \u4_intb_msk_reg[1]/P0001  ;
  assign n10691 = n10689 & ~n10690 ;
  assign n10692 = n10686 & n10691 ;
  assign n10693 = ~\u4_u3_r5_reg/NET0131  & ~\u4_u3_set_r_reg/P0001  ;
  assign n10694 = n6281 & n10693 ;
  assign n10695 = \u4_u3_csr0_reg[2]/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n10696 = ~\u4_u3_r5_reg/NET0131  & ~n10695 ;
  assign n10697 = ~n10694 & ~n10696 ;
  assign n10698 = \u4_u3_csr1_reg[0]/P0001  & ~\u4_u3_dma_in_cnt_reg[0]/P0001  ;
  assign n10699 = n10697 & n10698 ;
  assign n10700 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[0]/P0001  ;
  assign n10701 = ~n10697 & n10700 ;
  assign n10702 = ~n10699 & ~n10701 ;
  assign n10703 = \u4_u0_csr0_reg[2]/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n10704 = ~\u4_u0_r5_reg/NET0131  & ~n10703 ;
  assign n10705 = ~\u4_u0_r5_reg/NET0131  & ~\u4_u0_set_r_reg/P0001  ;
  assign n10706 = n6281 & n10705 ;
  assign n10707 = ~n10704 & ~n10706 ;
  assign n10708 = \u4_u0_csr1_reg[0]/P0001  & ~\u4_u0_dma_in_cnt_reg[0]/P0001  ;
  assign n10709 = n10707 & n10708 ;
  assign n10710 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[0]/P0001  ;
  assign n10711 = ~n10707 & n10710 ;
  assign n10712 = ~n10709 & ~n10711 ;
  assign n10713 = \u4_u1_csr0_reg[2]/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n10714 = ~\u4_u1_r5_reg/NET0131  & ~n10713 ;
  assign n10715 = ~\u4_u1_r5_reg/NET0131  & ~\u4_u1_set_r_reg/P0001  ;
  assign n10716 = n6281 & n10715 ;
  assign n10717 = ~n10714 & ~n10716 ;
  assign n10718 = \u4_u1_csr1_reg[0]/P0001  & ~\u4_u1_dma_in_cnt_reg[0]/P0001  ;
  assign n10719 = n10717 & n10718 ;
  assign n10720 = \u4_u1_csr1_reg[0]/P0001  & \u4_u1_dma_in_cnt_reg[0]/P0001  ;
  assign n10721 = ~n10717 & n10720 ;
  assign n10722 = ~n10719 & ~n10721 ;
  assign n10723 = \u4_u2_csr0_reg[2]/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n10724 = ~\u4_u2_r5_reg/NET0131  & ~n10723 ;
  assign n10725 = ~\u4_u2_r5_reg/NET0131  & ~\u4_u2_set_r_reg/P0001  ;
  assign n10726 = n6281 & n10725 ;
  assign n10727 = ~n10724 & ~n10726 ;
  assign n10728 = \u4_u2_csr1_reg[0]/P0001  & ~\u4_u2_dma_in_cnt_reg[0]/P0001  ;
  assign n10729 = n10727 & n10728 ;
  assign n10730 = \u4_u2_csr1_reg[0]/P0001  & \u4_u2_dma_in_cnt_reg[0]/P0001  ;
  assign n10731 = ~n10727 & n10730 ;
  assign n10732 = ~n10729 & ~n10731 ;
  assign n10733 = ~n6768 & ~n6772 ;
  assign n10734 = n6769 & ~n10733 ;
  assign n10735 = n6598 & ~n10734 ;
  assign n10736 = \u4_u3_dma_in_cnt_reg[0]/P0001  & \u4_u3_dma_out_cnt_reg[1]/P0001  ;
  assign n10737 = ~n6738 & ~n10736 ;
  assign n10738 = \u4_u3_r5_reg/NET0131  & ~n10737 ;
  assign n10739 = ~n6769 & n10733 ;
  assign n10740 = ~n10738 & ~n10739 ;
  assign n10741 = n10735 & n10740 ;
  assign n10742 = ~\u4_u3_dma_out_cnt_reg[1]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n10743 = n6281 & n10742 ;
  assign n10744 = ~\u4_u3_dma_out_cnt_reg[1]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n10745 = ~\u4_u3_r5_reg/NET0131  & ~n10744 ;
  assign n10746 = ~n10743 & n10745 ;
  assign n10747 = ~n10738 & ~n10746 ;
  assign n10748 = \u4_u3_csr1_reg[0]/P0001  & ~n10747 ;
  assign n10749 = ~n10741 & n10748 ;
  assign n10750 = ~n6770 & ~n6772 ;
  assign n10751 = ~n6771 & ~n6775 ;
  assign n10752 = n10750 & ~n10751 ;
  assign n10753 = n6598 & ~n10752 ;
  assign n10754 = \u4_u3_dma_out_cnt_reg[2]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n10755 = ~n6738 & n10754 ;
  assign n10756 = ~\u4_u3_dma_out_cnt_reg[2]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n10757 = n6738 & n10756 ;
  assign n10758 = ~n10755 & ~n10757 ;
  assign n10759 = ~n10750 & n10751 ;
  assign n10760 = n10758 & ~n10759 ;
  assign n10761 = n10753 & n10760 ;
  assign n10762 = ~\u4_u3_dma_out_cnt_reg[2]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n10763 = n6281 & n10762 ;
  assign n10764 = ~\u4_u3_dma_out_cnt_reg[2]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n10765 = ~\u4_u3_r5_reg/NET0131  & ~n10764 ;
  assign n10766 = ~n10763 & n10765 ;
  assign n10767 = n10758 & ~n10766 ;
  assign n10768 = \u4_u3_csr1_reg[0]/P0001  & ~n10767 ;
  assign n10769 = ~n10761 & n10768 ;
  assign n10770 = \u4_u3_r5_reg/NET0131  & n6740 ;
  assign n10771 = ~\u4_u3_dma_out_cnt_reg[2]/P0001  & n6738 ;
  assign n10772 = \u4_u3_dma_out_cnt_reg[3]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n10773 = ~n10771 & n10772 ;
  assign n10774 = ~n10770 & ~n10773 ;
  assign n10775 = \u4_u3_csr1_reg[0]/P0001  & ~n10774 ;
  assign n10776 = ~n6774 & ~n6775 ;
  assign n10777 = ~n6764 & ~n6766 ;
  assign n10778 = ~n10776 & ~n10777 ;
  assign n10779 = ~n6775 & n10777 ;
  assign n10780 = ~n6774 & n10779 ;
  assign n10781 = n6598 & ~n10780 ;
  assign n10782 = ~n10778 & n10781 ;
  assign n10783 = ~\u4_u3_dma_out_cnt_reg[3]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n10784 = n6281 & n10783 ;
  assign n10785 = ~\u4_u3_dma_out_cnt_reg[3]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n10786 = \u4_u3_csr1_reg[0]/P0001  & ~n10785 ;
  assign n10787 = ~n10784 & n10786 ;
  assign n10788 = ~\u4_u3_r5_reg/NET0131  & n10787 ;
  assign n10789 = ~n10782 & n10788 ;
  assign n10790 = ~n10775 & ~n10789 ;
  assign n10791 = ~\u1_u2_mack_r_reg/P0001  & n4066 ;
  assign n10792 = \u1_u2_state_reg[4]/NET0131  & n10791 ;
  assign n10793 = \u1_u2_state_reg[4]/NET0131  & n4189 ;
  assign n10794 = ~n4103 & n10793 ;
  assign n10795 = ~n10792 & ~n10794 ;
  assign n10796 = \u1_u2_state_reg[4]/NET0131  & ~\u1_u2_wr_done_reg/P0001  ;
  assign n10797 = ~\u1_u2_wr_last_reg/P0001  & ~n10796 ;
  assign n10798 = ~\u1_u3_abort_reg/P0001  & ~n10797 ;
  assign n10799 = n4082 & n10798 ;
  assign n10800 = n10795 & ~n10799 ;
  assign n10801 = rst_i_pad & ~n10800 ;
  assign n10802 = ~n6834 & ~n6838 ;
  assign n10803 = n6835 & ~n10802 ;
  assign n10804 = n6632 & ~n10803 ;
  assign n10805 = \u4_u0_dma_in_cnt_reg[0]/P0001  & \u4_u0_dma_out_cnt_reg[1]/P0001  ;
  assign n10806 = ~n6802 & ~n10805 ;
  assign n10807 = \u4_u0_r5_reg/NET0131  & ~n10806 ;
  assign n10808 = ~n6835 & n10802 ;
  assign n10809 = ~n10807 & ~n10808 ;
  assign n10810 = n10804 & n10809 ;
  assign n10811 = ~\u4_u0_dma_out_cnt_reg[1]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n10812 = n6281 & n10811 ;
  assign n10813 = ~\u4_u0_dma_out_cnt_reg[1]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n10814 = ~\u4_u0_r5_reg/NET0131  & ~n10813 ;
  assign n10815 = ~n10812 & n10814 ;
  assign n10816 = ~n10807 & ~n10815 ;
  assign n10817 = \u4_u0_csr1_reg[0]/P0001  & ~n10816 ;
  assign n10818 = ~n10810 & n10817 ;
  assign n10819 = ~n6836 & ~n6838 ;
  assign n10820 = ~n6837 & ~n6841 ;
  assign n10821 = n10819 & ~n10820 ;
  assign n10822 = n6632 & ~n10821 ;
  assign n10823 = \u4_u0_dma_out_cnt_reg[2]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n10824 = ~n6802 & n10823 ;
  assign n10825 = ~\u4_u0_dma_out_cnt_reg[2]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n10826 = ~\u4_u0_dma_in_cnt_reg[0]/P0001  & ~\u4_u0_dma_out_cnt_reg[1]/P0001  ;
  assign n10827 = n10825 & n10826 ;
  assign n10828 = ~n10824 & ~n10827 ;
  assign n10829 = ~n10819 & n10820 ;
  assign n10830 = n10828 & ~n10829 ;
  assign n10831 = n10822 & n10830 ;
  assign n10832 = ~\u4_u0_dma_out_cnt_reg[2]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n10833 = n6281 & n10832 ;
  assign n10834 = ~\u4_u0_dma_out_cnt_reg[2]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n10835 = ~\u4_u0_r5_reg/NET0131  & ~n10834 ;
  assign n10836 = ~n10833 & n10835 ;
  assign n10837 = n10828 & ~n10836 ;
  assign n10838 = \u4_u0_csr1_reg[0]/P0001  & ~n10837 ;
  assign n10839 = ~n10831 & n10838 ;
  assign n10840 = \u4_u0_r5_reg/NET0131  & n6804 ;
  assign n10841 = \u4_u0_dma_out_cnt_reg[3]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n10842 = ~\u4_u0_dma_out_cnt_reg[2]/P0001  & n10826 ;
  assign n10843 = n10841 & ~n10842 ;
  assign n10844 = ~n10840 & ~n10843 ;
  assign n10845 = \u4_u0_csr1_reg[0]/P0001  & ~n10844 ;
  assign n10846 = ~n6840 & ~n6841 ;
  assign n10847 = ~n6830 & ~n6832 ;
  assign n10848 = ~n10846 & ~n10847 ;
  assign n10849 = ~n6841 & n10847 ;
  assign n10850 = ~n6840 & n10849 ;
  assign n10851 = n6632 & ~n10850 ;
  assign n10852 = ~n10848 & n10851 ;
  assign n10853 = ~\u4_u0_dma_out_cnt_reg[3]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n10854 = n6281 & n10853 ;
  assign n10855 = ~\u4_u0_dma_out_cnt_reg[3]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n10856 = n6613 & ~n10855 ;
  assign n10857 = ~n10854 & n10856 ;
  assign n10858 = ~n10852 & n10857 ;
  assign n10859 = ~n10845 & ~n10858 ;
  assign n10860 = ~n6898 & ~n6902 ;
  assign n10861 = n6899 & ~n10860 ;
  assign n10862 = n6369 & ~n10861 ;
  assign n10863 = \u4_u1_dma_in_cnt_reg[0]/P0001  & \u4_u1_dma_out_cnt_reg[1]/P0001  ;
  assign n10864 = ~n6866 & ~n10863 ;
  assign n10865 = \u4_u1_r5_reg/NET0131  & ~n10864 ;
  assign n10866 = ~n6899 & n10860 ;
  assign n10867 = ~n10865 & ~n10866 ;
  assign n10868 = n10862 & n10867 ;
  assign n10869 = ~\u4_u1_dma_out_cnt_reg[1]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n10870 = n6281 & n10869 ;
  assign n10871 = ~\u4_u1_dma_out_cnt_reg[1]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n10872 = ~\u4_u1_r5_reg/NET0131  & ~n10871 ;
  assign n10873 = ~n10870 & n10872 ;
  assign n10874 = ~n10865 & ~n10873 ;
  assign n10875 = \u4_u1_csr1_reg[0]/P0001  & ~n10874 ;
  assign n10876 = ~n10868 & n10875 ;
  assign n10877 = ~n6900 & ~n6902 ;
  assign n10878 = ~n6901 & ~n6905 ;
  assign n10879 = n10877 & ~n10878 ;
  assign n10880 = n6369 & ~n10879 ;
  assign n10881 = \u4_u1_dma_out_cnt_reg[2]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n10882 = ~n6866 & n10881 ;
  assign n10883 = ~\u4_u1_dma_out_cnt_reg[2]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n10884 = n6866 & n10883 ;
  assign n10885 = ~n10882 & ~n10884 ;
  assign n10886 = ~n10877 & n10878 ;
  assign n10887 = n10885 & ~n10886 ;
  assign n10888 = n10880 & n10887 ;
  assign n10889 = ~\u4_u1_dma_out_cnt_reg[2]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n10890 = n6281 & n10889 ;
  assign n10891 = ~\u4_u1_dma_out_cnt_reg[2]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n10892 = ~\u4_u1_r5_reg/NET0131  & ~n10891 ;
  assign n10893 = ~n10890 & n10892 ;
  assign n10894 = n10885 & ~n10893 ;
  assign n10895 = \u4_u1_csr1_reg[0]/P0001  & ~n10894 ;
  assign n10896 = ~n10888 & n10895 ;
  assign n10897 = \u4_u1_r5_reg/NET0131  & n6868 ;
  assign n10898 = ~\u4_u1_dma_out_cnt_reg[2]/P0001  & n6866 ;
  assign n10899 = \u4_u1_dma_out_cnt_reg[3]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n10900 = ~n10898 & n10899 ;
  assign n10901 = ~n10897 & ~n10900 ;
  assign n10902 = \u4_u1_csr1_reg[0]/P0001  & ~n10901 ;
  assign n10903 = ~n6904 & ~n6905 ;
  assign n10904 = ~n6894 & ~n6896 ;
  assign n10905 = ~n10903 & ~n10904 ;
  assign n10906 = ~n6905 & n10904 ;
  assign n10907 = ~n6904 & n10906 ;
  assign n10908 = n6369 & ~n10907 ;
  assign n10909 = ~n10905 & n10908 ;
  assign n10910 = ~\u4_u1_dma_out_cnt_reg[3]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n10911 = n6281 & n10910 ;
  assign n10912 = ~\u4_u1_dma_out_cnt_reg[3]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n10913 = ~\u4_u1_r5_reg/NET0131  & ~n10912 ;
  assign n10914 = ~n10911 & n10913 ;
  assign n10915 = \u4_u1_csr1_reg[0]/P0001  & n10914 ;
  assign n10916 = ~n10909 & n10915 ;
  assign n10917 = ~n10902 & ~n10916 ;
  assign n10918 = ~n6961 & ~n6965 ;
  assign n10919 = n6962 & ~n10918 ;
  assign n10920 = n6667 & ~n10919 ;
  assign n10921 = \u4_u2_dma_in_cnt_reg[0]/P0001  & \u4_u2_dma_out_cnt_reg[1]/P0001  ;
  assign n10922 = ~n6930 & ~n10921 ;
  assign n10923 = \u4_u2_r5_reg/NET0131  & ~n10922 ;
  assign n10924 = ~n6962 & n10918 ;
  assign n10925 = ~n10923 & ~n10924 ;
  assign n10926 = n10920 & n10925 ;
  assign n10927 = ~\u4_u2_dma_out_cnt_reg[1]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n10928 = n6281 & n10927 ;
  assign n10929 = ~\u4_u2_dma_out_cnt_reg[1]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n10930 = ~\u4_u2_r5_reg/NET0131  & ~n10929 ;
  assign n10931 = ~n10928 & n10930 ;
  assign n10932 = ~n10923 & ~n10931 ;
  assign n10933 = \u4_u2_csr1_reg[0]/P0001  & ~n10932 ;
  assign n10934 = ~n10926 & n10933 ;
  assign n10935 = ~n6963 & ~n6965 ;
  assign n10936 = ~n6964 & ~n6968 ;
  assign n10937 = n10935 & ~n10936 ;
  assign n10938 = n6667 & ~n10937 ;
  assign n10939 = \u4_u2_dma_out_cnt_reg[2]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n10940 = ~n6930 & n10939 ;
  assign n10941 = ~\u4_u2_dma_out_cnt_reg[2]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n10942 = n6930 & n10941 ;
  assign n10943 = ~n10940 & ~n10942 ;
  assign n10944 = ~n10935 & n10936 ;
  assign n10945 = n10943 & ~n10944 ;
  assign n10946 = n10938 & n10945 ;
  assign n10947 = ~\u4_u2_dma_out_cnt_reg[2]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n10948 = n6281 & n10947 ;
  assign n10949 = ~\u4_u2_dma_out_cnt_reg[2]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n10950 = ~\u4_u2_r5_reg/NET0131  & ~n10949 ;
  assign n10951 = ~n10948 & n10950 ;
  assign n10952 = n10943 & ~n10951 ;
  assign n10953 = \u4_u2_csr1_reg[0]/P0001  & ~n10952 ;
  assign n10954 = ~n10946 & n10953 ;
  assign n10955 = \u4_u2_r5_reg/NET0131  & n6932 ;
  assign n10956 = ~\u4_u2_dma_out_cnt_reg[2]/P0001  & n6930 ;
  assign n10957 = \u4_u2_dma_out_cnt_reg[3]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n10958 = ~n10956 & n10957 ;
  assign n10959 = ~n10955 & ~n10958 ;
  assign n10960 = \u4_u2_csr1_reg[0]/P0001  & ~n10959 ;
  assign n10961 = ~n6967 & ~n6968 ;
  assign n10962 = ~n6957 & ~n6959 ;
  assign n10963 = ~n10961 & ~n10962 ;
  assign n10964 = ~n6968 & n10962 ;
  assign n10965 = ~n6967 & n10964 ;
  assign n10966 = n6667 & ~n10965 ;
  assign n10967 = ~n10963 & n10966 ;
  assign n10968 = ~\u4_u2_dma_out_cnt_reg[3]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n10969 = n6281 & n10968 ;
  assign n10970 = ~\u4_u2_dma_out_cnt_reg[3]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n10971 = n6946 & ~n10970 ;
  assign n10972 = ~n10969 & n10971 ;
  assign n10973 = ~n10967 & n10972 ;
  assign n10974 = ~n10960 & ~n10973 ;
  assign n10975 = ~n6245 & ~n6253 ;
  assign n10976 = ~n6586 & ~n10975 ;
  assign n10977 = n6598 & ~n10976 ;
  assign n10978 = \u4_u3_dma_in_cnt_reg[2]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n10979 = ~n6274 & n10978 ;
  assign n10980 = ~\u4_u3_dma_in_cnt_reg[2]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n10981 = n6274 & n10980 ;
  assign n10982 = ~n10979 & ~n10981 ;
  assign n10983 = n6248 & ~n6253 ;
  assign n10984 = n10982 & ~n10983 ;
  assign n10985 = n10977 & n10984 ;
  assign n10986 = ~\u4_u3_dma_in_cnt_reg[2]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n10987 = n6281 & n10986 ;
  assign n10988 = ~\u4_u3_dma_in_cnt_reg[2]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n10989 = ~\u4_u3_r5_reg/NET0131  & ~n10988 ;
  assign n10990 = ~n10987 & n10989 ;
  assign n10991 = n10982 & ~n10990 ;
  assign n10992 = \u4_u3_csr1_reg[0]/P0001  & ~n10991 ;
  assign n10993 = ~n10985 & n10992 ;
  assign n10994 = \u4_u3_r5_reg/NET0131  & ~n6276 ;
  assign n10995 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[3]/P0001  ;
  assign n10996 = \u4_u3_csr1_reg[0]/P0001  & \u4_u3_dma_in_cnt_reg[2]/P0001  ;
  assign n10997 = n6274 & n10996 ;
  assign n10998 = ~n10995 & ~n10997 ;
  assign n10999 = n10994 & ~n10998 ;
  assign n11000 = ~n6248 & ~n6253 ;
  assign n11001 = ~n6252 & ~n6257 ;
  assign n11002 = ~n11000 & n11001 ;
  assign n11003 = ~n6253 & ~n11001 ;
  assign n11004 = ~n6248 & n11003 ;
  assign n11005 = n6598 & ~n11004 ;
  assign n11006 = ~n11002 & n11005 ;
  assign n11007 = ~\u4_u3_dma_in_cnt_reg[3]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n11008 = n6281 & n11007 ;
  assign n11009 = ~\u4_u3_dma_in_cnt_reg[3]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n11010 = \u4_u3_csr1_reg[0]/P0001  & ~n11009 ;
  assign n11011 = ~n11008 & n11010 ;
  assign n11012 = ~\u4_u3_r5_reg/NET0131  & n11011 ;
  assign n11013 = ~n11006 & n11012 ;
  assign n11014 = ~n10999 & ~n11013 ;
  assign n11015 = ~\u4_u3_dma_out_cnt_reg[5]/P0001  & n9546 ;
  assign n11016 = n6740 & n11015 ;
  assign n11017 = \u4_u3_csr1_reg[0]/P0001  & n11016 ;
  assign n11018 = ~\u4_u3_dma_out_cnt_reg[4]/P0001  & n6740 ;
  assign n11019 = \u4_u3_dma_out_cnt_reg[5]/P0001  & \u4_u3_r5_reg/NET0131  ;
  assign n11020 = \u4_u3_csr1_reg[0]/P0001  & n11019 ;
  assign n11021 = ~n11018 & n11020 ;
  assign n11022 = ~n11017 & ~n11021 ;
  assign n11023 = n6778 & ~n6780 ;
  assign n11024 = ~n6761 & ~n6779 ;
  assign n11025 = ~n11023 & n11024 ;
  assign n11026 = ~n6780 & ~n11024 ;
  assign n11027 = n6778 & n11026 ;
  assign n11028 = n6598 & ~n11027 ;
  assign n11029 = ~n11025 & n11028 ;
  assign n11030 = ~\u4_u3_dma_out_cnt_reg[5]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n11031 = n6281 & n11030 ;
  assign n11032 = ~\u4_u3_dma_out_cnt_reg[5]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n11033 = \u4_u3_csr1_reg[0]/P0001  & ~n11032 ;
  assign n11034 = ~n11031 & n11033 ;
  assign n11035 = ~\u4_u3_r5_reg/NET0131  & n11034 ;
  assign n11036 = ~n11029 & n11035 ;
  assign n11037 = n11022 & ~n11036 ;
  assign n11038 = ~n6303 & ~n6311 ;
  assign n11039 = ~n6620 & ~n11038 ;
  assign n11040 = n6632 & ~n11039 ;
  assign n11041 = \u4_u0_dma_in_cnt_reg[2]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n11042 = ~n6332 & n11041 ;
  assign n11043 = ~\u4_u0_dma_in_cnt_reg[2]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n11044 = n6332 & n11043 ;
  assign n11045 = ~n11042 & ~n11044 ;
  assign n11046 = n6306 & ~n6311 ;
  assign n11047 = n11045 & ~n11046 ;
  assign n11048 = n11040 & n11047 ;
  assign n11049 = ~\u4_u0_dma_in_cnt_reg[2]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n11050 = n6281 & n11049 ;
  assign n11051 = ~\u4_u0_dma_in_cnt_reg[2]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n11052 = ~\u4_u0_r5_reg/NET0131  & ~n11051 ;
  assign n11053 = ~n11050 & n11052 ;
  assign n11054 = n11045 & ~n11053 ;
  assign n11055 = \u4_u0_csr1_reg[0]/P0001  & ~n11054 ;
  assign n11056 = ~n11048 & n11055 ;
  assign n11057 = \u4_u0_r5_reg/NET0131  & ~n6334 ;
  assign n11058 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[3]/P0001  ;
  assign n11059 = \u4_u0_csr1_reg[0]/P0001  & \u4_u0_dma_in_cnt_reg[2]/P0001  ;
  assign n11060 = n6332 & n11059 ;
  assign n11061 = ~n11058 & ~n11060 ;
  assign n11062 = n11057 & ~n11061 ;
  assign n11063 = ~n6306 & ~n6311 ;
  assign n11064 = ~n6310 & ~n6315 ;
  assign n11065 = ~n11063 & n11064 ;
  assign n11066 = ~n6311 & ~n11064 ;
  assign n11067 = ~n6306 & n11066 ;
  assign n11068 = n6632 & ~n11067 ;
  assign n11069 = ~n11065 & n11068 ;
  assign n11070 = ~\u4_u0_dma_in_cnt_reg[3]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n11071 = n6281 & n11070 ;
  assign n11072 = ~\u4_u0_dma_in_cnt_reg[3]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n11073 = n6613 & ~n11072 ;
  assign n11074 = ~n11071 & n11073 ;
  assign n11075 = ~n11069 & n11074 ;
  assign n11076 = ~n11062 & ~n11075 ;
  assign n11077 = ~\u4_u0_dma_out_cnt_reg[5]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n11078 = ~\u4_u0_dma_out_cnt_reg[4]/P0001  & n11077 ;
  assign n11079 = n6804 & n11078 ;
  assign n11080 = \u4_u0_csr1_reg[0]/P0001  & n11079 ;
  assign n11081 = ~\u4_u0_dma_out_cnt_reg[4]/P0001  & n6804 ;
  assign n11082 = \u4_u0_dma_out_cnt_reg[5]/P0001  & \u4_u0_r5_reg/NET0131  ;
  assign n11083 = \u4_u0_csr1_reg[0]/P0001  & n11082 ;
  assign n11084 = ~n11081 & n11083 ;
  assign n11085 = ~n11080 & ~n11084 ;
  assign n11086 = n6844 & ~n6846 ;
  assign n11087 = ~n6827 & ~n6845 ;
  assign n11088 = ~n11086 & n11087 ;
  assign n11089 = ~n6846 & ~n11087 ;
  assign n11090 = n6844 & n11089 ;
  assign n11091 = n6632 & ~n11090 ;
  assign n11092 = ~n11088 & n11091 ;
  assign n11093 = ~\u4_u0_dma_out_cnt_reg[5]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n11094 = n6281 & n11093 ;
  assign n11095 = ~\u4_u0_dma_out_cnt_reg[5]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n11096 = n6613 & ~n11095 ;
  assign n11097 = ~n11094 & n11096 ;
  assign n11098 = ~n11092 & n11097 ;
  assign n11099 = n11085 & ~n11098 ;
  assign n11100 = ~n6388 & ~n6390 ;
  assign n11101 = ~n6389 & ~n6393 ;
  assign n11102 = ~n11100 & ~n11101 ;
  assign n11103 = n6369 & ~n11102 ;
  assign n11104 = \u4_u1_dma_in_cnt_reg[2]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n11105 = ~n6359 & n11104 ;
  assign n11106 = ~\u4_u1_dma_in_cnt_reg[2]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n11107 = n6359 & n11106 ;
  assign n11108 = ~n11105 & ~n11107 ;
  assign n11109 = n11100 & n11101 ;
  assign n11110 = n11108 & ~n11109 ;
  assign n11111 = n11103 & n11110 ;
  assign n11112 = ~\u4_u1_dma_in_cnt_reg[2]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n11113 = n6281 & n11112 ;
  assign n11114 = ~\u4_u1_dma_in_cnt_reg[2]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n11115 = ~\u4_u1_r5_reg/NET0131  & ~n11114 ;
  assign n11116 = ~n11113 & n11115 ;
  assign n11117 = n11108 & ~n11116 ;
  assign n11118 = \u4_u1_csr1_reg[0]/P0001  & ~n11117 ;
  assign n11119 = ~n11111 & n11118 ;
  assign n11120 = \u4_u1_r5_reg/NET0131  & ~n6361 ;
  assign n11121 = \u4_u1_csr1_reg[0]/P0001  & \u4_u1_dma_in_cnt_reg[3]/P0001  ;
  assign n11122 = \u4_u1_csr1_reg[0]/P0001  & \u4_u1_dma_in_cnt_reg[2]/P0001  ;
  assign n11123 = n6359 & n11122 ;
  assign n11124 = ~n11121 & ~n11123 ;
  assign n11125 = n11120 & ~n11124 ;
  assign n11126 = ~n6392 & ~n6393 ;
  assign n11127 = ~n6382 & ~n6384 ;
  assign n11128 = ~n11126 & n11127 ;
  assign n11129 = ~n6393 & ~n11127 ;
  assign n11130 = ~n6392 & n11129 ;
  assign n11131 = n6369 & ~n11130 ;
  assign n11132 = ~n11128 & n11131 ;
  assign n11133 = ~\u4_u1_dma_in_cnt_reg[3]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n11134 = n6281 & n11133 ;
  assign n11135 = ~\u4_u1_dma_in_cnt_reg[3]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n11136 = \u4_u1_csr1_reg[0]/P0001  & ~n11135 ;
  assign n11137 = ~n11134 & n11136 ;
  assign n11138 = ~\u4_u1_r5_reg/NET0131  & n11137 ;
  assign n11139 = ~n11132 & n11138 ;
  assign n11140 = ~n11125 & ~n11139 ;
  assign n11141 = ~\u4_u1_dma_out_cnt_reg[5]/P0001  & n9596 ;
  assign n11142 = n6868 & n11141 ;
  assign n11143 = \u4_u1_csr1_reg[0]/P0001  & n11142 ;
  assign n11144 = ~\u4_u1_dma_out_cnt_reg[4]/P0001  & n6868 ;
  assign n11145 = \u4_u1_dma_out_cnt_reg[5]/P0001  & \u4_u1_r5_reg/NET0131  ;
  assign n11146 = \u4_u1_csr1_reg[0]/P0001  & n11145 ;
  assign n11147 = ~n11144 & n11146 ;
  assign n11148 = ~n11143 & ~n11147 ;
  assign n11149 = n6908 & ~n6910 ;
  assign n11150 = ~n6891 & ~n6909 ;
  assign n11151 = ~n11149 & n11150 ;
  assign n11152 = ~n6910 & ~n11150 ;
  assign n11153 = n6908 & n11152 ;
  assign n11154 = n6369 & ~n11153 ;
  assign n11155 = ~n11151 & n11154 ;
  assign n11156 = ~\u4_u1_dma_out_cnt_reg[5]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n11157 = n6281 & n11156 ;
  assign n11158 = ~\u4_u1_dma_out_cnt_reg[5]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n11159 = \u4_u1_csr1_reg[0]/P0001  & ~n11158 ;
  assign n11160 = ~n11157 & n11159 ;
  assign n11161 = ~\u4_u1_r5_reg/NET0131  & n11160 ;
  assign n11162 = ~n11155 & n11161 ;
  assign n11163 = n11148 & ~n11162 ;
  assign n11164 = ~n6435 & ~n6437 ;
  assign n11165 = ~n6436 & ~n6440 ;
  assign n11166 = ~n11164 & ~n11165 ;
  assign n11167 = n6667 & ~n11166 ;
  assign n11168 = \u4_u2_dma_in_cnt_reg[2]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n11169 = ~n6460 & n11168 ;
  assign n11170 = ~\u4_u2_dma_in_cnt_reg[2]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n11171 = n6460 & n11170 ;
  assign n11172 = ~n11169 & ~n11171 ;
  assign n11173 = n11164 & n11165 ;
  assign n11174 = n11172 & ~n11173 ;
  assign n11175 = n11167 & n11174 ;
  assign n11176 = ~\u4_u2_dma_in_cnt_reg[2]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n11177 = n6281 & n11176 ;
  assign n11178 = ~\u4_u2_dma_in_cnt_reg[2]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n11179 = ~\u4_u2_r5_reg/NET0131  & ~n11178 ;
  assign n11180 = ~n11177 & n11179 ;
  assign n11181 = n11172 & ~n11180 ;
  assign n11182 = \u4_u2_csr1_reg[0]/P0001  & ~n11181 ;
  assign n11183 = ~n11175 & n11182 ;
  assign n11184 = \u4_u2_r5_reg/NET0131  & ~n6462 ;
  assign n11185 = \u4_u2_csr1_reg[0]/P0001  & \u4_u2_dma_in_cnt_reg[3]/P0001  ;
  assign n11186 = \u4_u2_csr1_reg[0]/P0001  & \u4_u2_dma_in_cnt_reg[2]/P0001  ;
  assign n11187 = n6460 & n11186 ;
  assign n11188 = ~n11185 & ~n11187 ;
  assign n11189 = n11184 & ~n11188 ;
  assign n11190 = ~n6439 & ~n6440 ;
  assign n11191 = ~n6429 & ~n6431 ;
  assign n11192 = ~n11190 & n11191 ;
  assign n11193 = ~n6440 & ~n11191 ;
  assign n11194 = ~n6439 & n11193 ;
  assign n11195 = n6667 & ~n11194 ;
  assign n11196 = ~n11192 & n11195 ;
  assign n11197 = ~\u4_u2_dma_in_cnt_reg[3]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n11198 = n6281 & n11197 ;
  assign n11199 = ~\u4_u2_dma_in_cnt_reg[3]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n11200 = n6946 & ~n11199 ;
  assign n11201 = ~n11198 & n11200 ;
  assign n11202 = ~n11196 & n11201 ;
  assign n11203 = ~n11189 & ~n11202 ;
  assign n11204 = ~\u4_u2_dma_out_cnt_reg[5]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n11205 = ~\u4_u2_dma_out_cnt_reg[4]/P0001  & n11204 ;
  assign n11206 = n6932 & n11205 ;
  assign n11207 = \u4_u2_csr1_reg[0]/P0001  & n11206 ;
  assign n11208 = ~\u4_u2_dma_out_cnt_reg[4]/P0001  & n6932 ;
  assign n11209 = \u4_u2_dma_out_cnt_reg[5]/P0001  & \u4_u2_r5_reg/NET0131  ;
  assign n11210 = \u4_u2_csr1_reg[0]/P0001  & n11209 ;
  assign n11211 = ~n11208 & n11210 ;
  assign n11212 = ~n11207 & ~n11211 ;
  assign n11213 = n6971 & ~n6973 ;
  assign n11214 = ~n6954 & ~n6972 ;
  assign n11215 = ~n11213 & n11214 ;
  assign n11216 = ~n6973 & ~n11214 ;
  assign n11217 = n6971 & n11216 ;
  assign n11218 = n6667 & ~n11217 ;
  assign n11219 = ~n11215 & n11218 ;
  assign n11220 = ~\u4_u2_dma_out_cnt_reg[5]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n11221 = n6281 & n11220 ;
  assign n11222 = ~\u4_u2_dma_out_cnt_reg[5]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n11223 = n6946 & ~n11222 ;
  assign n11224 = ~n11221 & n11223 ;
  assign n11225 = ~n11219 & n11224 ;
  assign n11226 = n11212 & ~n11225 ;
  assign n11227 = \u0_u0_idle_cnt1_reg[0]/P0001  & \u0_u0_idle_cnt1_reg[1]/P0001  ;
  assign n11228 = ~\u0_u0_idle_cnt1_reg[2]/P0001  & ~n11227 ;
  assign n11229 = \u0_u0_idle_cnt1_reg[3]/P0001  & ~n11228 ;
  assign n11230 = ~\u0_u0_idle_cnt1_reg[4]/P0001  & ~\u0_u0_idle_cnt1_reg[5]/P0001  ;
  assign n11231 = ~\u0_u0_idle_cnt1_reg[6]/P0001  & ~\u0_u0_idle_cnt1_reg[7]/P0001  ;
  assign n11232 = n11230 & n11231 ;
  assign n11233 = ~n11229 & n11232 ;
  assign n11234 = ~n8672 & ~n11233 ;
  assign n11235 = ~n8666 & n11234 ;
  assign n11236 = ~n6242 & ~n6246 ;
  assign n11237 = ~n6243 & ~n11236 ;
  assign n11238 = n6598 & ~n11237 ;
  assign n11239 = ~\u4_u3_dma_in_cnt_reg[0]/P0001  & ~\u4_u3_dma_in_cnt_reg[1]/P0001  ;
  assign n11240 = \u4_u3_r5_reg/NET0131  & ~n6274 ;
  assign n11241 = ~n11239 & n11240 ;
  assign n11242 = n6243 & n11236 ;
  assign n11243 = ~n11241 & ~n11242 ;
  assign n11244 = n11238 & n11243 ;
  assign n11245 = ~\u4_u3_dma_in_cnt_reg[1]/P0001  & ~\u4_u3_set_r_reg/P0001  ;
  assign n11246 = n6281 & n11245 ;
  assign n11247 = ~\u4_u3_dma_in_cnt_reg[1]/P0001  & ~\u4_u3_ep_match_r_reg/P0001  ;
  assign n11248 = ~\u4_u3_r5_reg/NET0131  & ~n11247 ;
  assign n11249 = ~n11246 & n11248 ;
  assign n11250 = ~n11241 & ~n11249 ;
  assign n11251 = \u4_u3_csr1_reg[0]/P0001  & ~n11250 ;
  assign n11252 = ~n11244 & n11251 ;
  assign n11253 = ~n6300 & ~n6304 ;
  assign n11254 = ~n6301 & ~n11253 ;
  assign n11255 = n6632 & ~n11254 ;
  assign n11256 = ~\u4_u0_dma_in_cnt_reg[0]/P0001  & ~\u4_u0_dma_in_cnt_reg[1]/P0001  ;
  assign n11257 = \u4_u0_r5_reg/NET0131  & ~n6332 ;
  assign n11258 = ~n11256 & n11257 ;
  assign n11259 = n6301 & n11253 ;
  assign n11260 = ~n11258 & ~n11259 ;
  assign n11261 = n11255 & n11260 ;
  assign n11262 = ~\u4_u0_dma_in_cnt_reg[1]/P0001  & ~\u4_u0_set_r_reg/P0001  ;
  assign n11263 = n6281 & n11262 ;
  assign n11264 = ~\u4_u0_dma_in_cnt_reg[1]/P0001  & ~\u4_u0_ep_match_r_reg/P0001  ;
  assign n11265 = ~\u4_u0_r5_reg/NET0131  & ~n11264 ;
  assign n11266 = ~n11263 & n11265 ;
  assign n11267 = ~n11258 & ~n11266 ;
  assign n11268 = \u4_u0_csr1_reg[0]/P0001  & ~n11267 ;
  assign n11269 = ~n11261 & n11268 ;
  assign n11270 = ~n6386 & ~n6390 ;
  assign n11271 = ~n6387 & ~n11270 ;
  assign n11272 = n6369 & ~n11271 ;
  assign n11273 = ~\u4_u1_dma_in_cnt_reg[0]/P0001  & ~\u4_u1_dma_in_cnt_reg[1]/P0001  ;
  assign n11274 = \u4_u1_r5_reg/NET0131  & ~n6359 ;
  assign n11275 = ~n11273 & n11274 ;
  assign n11276 = n6387 & n11270 ;
  assign n11277 = ~n11275 & ~n11276 ;
  assign n11278 = n11272 & n11277 ;
  assign n11279 = ~\u4_u1_dma_in_cnt_reg[1]/P0001  & ~\u4_u1_set_r_reg/P0001  ;
  assign n11280 = n6281 & n11279 ;
  assign n11281 = ~\u4_u1_dma_in_cnt_reg[1]/P0001  & ~\u4_u1_ep_match_r_reg/P0001  ;
  assign n11282 = ~\u4_u1_r5_reg/NET0131  & ~n11281 ;
  assign n11283 = ~n11280 & n11282 ;
  assign n11284 = ~n11275 & ~n11283 ;
  assign n11285 = \u4_u1_csr1_reg[0]/P0001  & ~n11284 ;
  assign n11286 = ~n11278 & n11285 ;
  assign n11287 = ~n6433 & ~n6437 ;
  assign n11288 = ~n6434 & ~n11287 ;
  assign n11289 = n6667 & ~n11288 ;
  assign n11290 = ~\u4_u2_dma_in_cnt_reg[0]/P0001  & ~\u4_u2_dma_in_cnt_reg[1]/P0001  ;
  assign n11291 = \u4_u2_r5_reg/NET0131  & ~n6460 ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11293 = n6434 & n11287 ;
  assign n11294 = ~n11292 & ~n11293 ;
  assign n11295 = n11289 & n11294 ;
  assign n11296 = ~\u4_u2_dma_in_cnt_reg[1]/P0001  & ~\u4_u2_set_r_reg/P0001  ;
  assign n11297 = n6281 & n11296 ;
  assign n11298 = ~\u4_u2_dma_in_cnt_reg[1]/P0001  & ~\u4_u2_ep_match_r_reg/P0001  ;
  assign n11299 = ~\u4_u2_r5_reg/NET0131  & ~n11298 ;
  assign n11300 = ~n11297 & n11299 ;
  assign n11301 = ~n11292 & ~n11300 ;
  assign n11302 = \u4_u2_csr1_reg[0]/P0001  & ~n11301 ;
  assign n11303 = ~n11295 & n11302 ;
  assign n11304 = \u4_u2_int_stat_reg[0]/P0001  & n5451 ;
  assign n11305 = \u1_u3_rx_ack_to_reg/P0001  & n4962 ;
  assign n11306 = n4965 & n11305 ;
  assign n11307 = ~\u1_u3_state_reg[2]/P0001  & \u1_u3_tx_data_to_reg/P0001  ;
  assign n11308 = n2372 & n11307 ;
  assign n11309 = n4919 & n11308 ;
  assign n11310 = ~n11306 & ~n11309 ;
  assign n11311 = \u4_u2_ep_match_r_reg/P0001  & n5451 ;
  assign n11312 = ~n11310 & n11311 ;
  assign n11313 = ~n11304 & ~n11312 ;
  assign n11314 = \wb_data_i[0]_pad  & n2568 ;
  assign n11315 = n2567 & n11314 ;
  assign n11316 = rst_i_pad & ~n11315 ;
  assign n11317 = ~\u4_u3_buf0_reg[0]/P0001  & ~n2574 ;
  assign n11318 = ~\u1_u3_idin_reg[0]/P0001  & n2574 ;
  assign n11319 = ~n11317 & ~n11318 ;
  assign n11320 = ~n2573 & ~n11319 ;
  assign n11321 = ~\u4_u3_buf0_orig_reg[0]/P0001  & n2573 ;
  assign n11322 = ~n11320 & ~n11321 ;
  assign n11323 = ~n2572 & n11322 ;
  assign n11324 = n11316 & ~n11323 ;
  assign n11325 = \wb_data_i[12]_pad  & n2568 ;
  assign n11326 = n2567 & n11325 ;
  assign n11327 = rst_i_pad & ~n11326 ;
  assign n11328 = ~\u4_u3_buf0_reg[12]/P0001  & ~n2574 ;
  assign n11329 = ~\u1_u3_idin_reg[12]/P0001  & n2574 ;
  assign n11330 = ~n11328 & ~n11329 ;
  assign n11331 = ~n2573 & ~n11330 ;
  assign n11332 = ~\u4_u3_buf0_orig_reg[12]/P0001  & n2573 ;
  assign n11333 = ~n11331 & ~n11332 ;
  assign n11334 = ~n2572 & n11333 ;
  assign n11335 = n11327 & ~n11334 ;
  assign n11336 = \wb_data_i[16]_pad  & n2568 ;
  assign n11337 = n2567 & n11336 ;
  assign n11338 = rst_i_pad & ~n11337 ;
  assign n11339 = ~\u4_u3_buf0_reg[16]/P0001  & ~n2574 ;
  assign n11340 = ~\u1_u3_idin_reg[16]/P0001  & n2574 ;
  assign n11341 = ~n11339 & ~n11340 ;
  assign n11342 = ~n2573 & ~n11341 ;
  assign n11343 = ~\u4_u3_buf0_orig_reg[16]/P0001  & n2573 ;
  assign n11344 = ~n11342 & ~n11343 ;
  assign n11345 = ~n2572 & n11344 ;
  assign n11346 = n11338 & ~n11345 ;
  assign n11347 = \wb_data_i[17]_pad  & n2568 ;
  assign n11348 = n2567 & n11347 ;
  assign n11349 = rst_i_pad & ~n11348 ;
  assign n11350 = ~\u4_u3_buf0_reg[17]/P0001  & ~n2574 ;
  assign n11351 = ~\u1_u3_idin_reg[17]/P0001  & n2574 ;
  assign n11352 = ~n11350 & ~n11351 ;
  assign n11353 = ~n2573 & ~n11352 ;
  assign n11354 = ~\u4_u3_buf0_orig_reg[17]/P0001  & n2573 ;
  assign n11355 = ~n11353 & ~n11354 ;
  assign n11356 = ~n2572 & n11355 ;
  assign n11357 = n11349 & ~n11356 ;
  assign n11358 = \wb_data_i[18]_pad  & n2568 ;
  assign n11359 = n2567 & n11358 ;
  assign n11360 = rst_i_pad & ~n11359 ;
  assign n11361 = ~\u4_u3_buf0_reg[18]/P0001  & ~n2574 ;
  assign n11362 = ~\u1_u3_idin_reg[18]/P0001  & n2574 ;
  assign n11363 = ~n11361 & ~n11362 ;
  assign n11364 = ~n2573 & ~n11363 ;
  assign n11365 = ~\u4_u3_buf0_orig_reg[18]/P0001  & n2573 ;
  assign n11366 = ~n11364 & ~n11365 ;
  assign n11367 = ~n2572 & n11366 ;
  assign n11368 = n11360 & ~n11367 ;
  assign n11369 = \wb_data_i[19]_pad  & n2568 ;
  assign n11370 = n2567 & n11369 ;
  assign n11371 = rst_i_pad & ~n11370 ;
  assign n11372 = ~\u4_u3_buf0_reg[19]/P0001  & ~n2574 ;
  assign n11373 = ~\u1_u3_idin_reg[19]/P0001  & n2574 ;
  assign n11374 = ~n11372 & ~n11373 ;
  assign n11375 = ~n2573 & ~n11374 ;
  assign n11376 = ~\u4_u3_buf0_orig_reg[19]/P0001  & n2573 ;
  assign n11377 = ~n11375 & ~n11376 ;
  assign n11378 = ~n2572 & n11377 ;
  assign n11379 = n11371 & ~n11378 ;
  assign n11380 = \wb_data_i[1]_pad  & n2568 ;
  assign n11381 = n2567 & n11380 ;
  assign n11382 = rst_i_pad & ~n11381 ;
  assign n11383 = ~\u4_u3_buf0_reg[1]/P0001  & ~n2574 ;
  assign n11384 = ~\u1_u3_idin_reg[1]/P0001  & n2574 ;
  assign n11385 = ~n11383 & ~n11384 ;
  assign n11386 = ~n2573 & ~n11385 ;
  assign n11387 = ~\u4_u3_buf0_orig_reg[1]/P0001  & n2573 ;
  assign n11388 = ~n11386 & ~n11387 ;
  assign n11389 = ~n2572 & n11388 ;
  assign n11390 = n11382 & ~n11389 ;
  assign n11391 = \wb_data_i[20]_pad  & n2568 ;
  assign n11392 = n2567 & n11391 ;
  assign n11393 = rst_i_pad & ~n11392 ;
  assign n11394 = ~\u4_u3_buf0_reg[20]/P0001  & ~n2574 ;
  assign n11395 = ~\u1_u3_idin_reg[20]/P0001  & n2574 ;
  assign n11396 = ~n11394 & ~n11395 ;
  assign n11397 = ~n2573 & ~n11396 ;
  assign n11398 = ~\u4_u3_buf0_orig_reg[20]/P0001  & n2573 ;
  assign n11399 = ~n11397 & ~n11398 ;
  assign n11400 = ~n2572 & n11399 ;
  assign n11401 = n11393 & ~n11400 ;
  assign n11402 = \wb_data_i[21]_pad  & n2568 ;
  assign n11403 = n2567 & n11402 ;
  assign n11404 = rst_i_pad & ~n11403 ;
  assign n11405 = ~\u4_u3_buf0_reg[21]/P0001  & ~n2574 ;
  assign n11406 = ~\u1_u3_idin_reg[21]/P0001  & n2574 ;
  assign n11407 = ~n11405 & ~n11406 ;
  assign n11408 = ~n2573 & ~n11407 ;
  assign n11409 = ~\u4_u3_buf0_orig_reg[21]/P0001  & n2573 ;
  assign n11410 = ~n11408 & ~n11409 ;
  assign n11411 = ~n2572 & n11410 ;
  assign n11412 = n11404 & ~n11411 ;
  assign n11413 = \wb_data_i[22]_pad  & n2568 ;
  assign n11414 = n2567 & n11413 ;
  assign n11415 = rst_i_pad & ~n11414 ;
  assign n11416 = ~\u4_u3_buf0_reg[22]/P0001  & ~n2574 ;
  assign n11417 = ~\u1_u3_idin_reg[22]/P0001  & n2574 ;
  assign n11418 = ~n11416 & ~n11417 ;
  assign n11419 = ~n2573 & ~n11418 ;
  assign n11420 = ~\u4_u3_buf0_orig_reg[22]/P0001  & n2573 ;
  assign n11421 = ~n11419 & ~n11420 ;
  assign n11422 = ~n2572 & n11421 ;
  assign n11423 = n11415 & ~n11422 ;
  assign n11424 = \wb_data_i[23]_pad  & n2568 ;
  assign n11425 = n2567 & n11424 ;
  assign n11426 = rst_i_pad & ~n11425 ;
  assign n11427 = ~\u4_u3_buf0_reg[23]/P0001  & ~n2574 ;
  assign n11428 = ~\u1_u3_idin_reg[23]/P0001  & n2574 ;
  assign n11429 = ~n11427 & ~n11428 ;
  assign n11430 = ~n2573 & ~n11429 ;
  assign n11431 = ~\u4_u3_buf0_orig_reg[23]/P0001  & n2573 ;
  assign n11432 = ~n11430 & ~n11431 ;
  assign n11433 = ~n2572 & n11432 ;
  assign n11434 = n11426 & ~n11433 ;
  assign n11435 = \wb_data_i[24]_pad  & n2568 ;
  assign n11436 = n2567 & n11435 ;
  assign n11437 = rst_i_pad & ~n11436 ;
  assign n11438 = ~\u4_u3_buf0_reg[24]/P0001  & ~n2574 ;
  assign n11439 = ~\u1_u3_idin_reg[24]/P0001  & n2574 ;
  assign n11440 = ~n11438 & ~n11439 ;
  assign n11441 = ~n2573 & ~n11440 ;
  assign n11442 = ~\u4_u3_buf0_orig_reg[24]/P0001  & n2573 ;
  assign n11443 = ~n11441 & ~n11442 ;
  assign n11444 = ~n2572 & n11443 ;
  assign n11445 = n11437 & ~n11444 ;
  assign n11446 = \wb_data_i[25]_pad  & n2568 ;
  assign n11447 = n2567 & n11446 ;
  assign n11448 = rst_i_pad & ~n11447 ;
  assign n11449 = ~\u4_u3_buf0_reg[25]/P0001  & ~n2574 ;
  assign n11450 = ~\u1_u3_idin_reg[25]/P0001  & n2574 ;
  assign n11451 = ~n11449 & ~n11450 ;
  assign n11452 = ~n2573 & ~n11451 ;
  assign n11453 = ~\u4_u3_buf0_orig_reg[25]/P0001  & n2573 ;
  assign n11454 = ~n11452 & ~n11453 ;
  assign n11455 = ~n2572 & n11454 ;
  assign n11456 = n11448 & ~n11455 ;
  assign n11457 = \wb_data_i[26]_pad  & n2568 ;
  assign n11458 = n2567 & n11457 ;
  assign n11459 = rst_i_pad & ~n11458 ;
  assign n11460 = ~\u4_u3_buf0_reg[26]/P0001  & ~n2574 ;
  assign n11461 = ~\u1_u3_idin_reg[26]/P0001  & n2574 ;
  assign n11462 = ~n11460 & ~n11461 ;
  assign n11463 = ~n2573 & ~n11462 ;
  assign n11464 = ~\u4_u3_buf0_orig_reg[26]/P0001  & n2573 ;
  assign n11465 = ~n11463 & ~n11464 ;
  assign n11466 = ~n2572 & n11465 ;
  assign n11467 = n11459 & ~n11466 ;
  assign n11468 = \wb_data_i[27]_pad  & n2568 ;
  assign n11469 = n2567 & n11468 ;
  assign n11470 = rst_i_pad & ~n11469 ;
  assign n11471 = ~\u4_u3_buf0_reg[27]/P0001  & ~n2574 ;
  assign n11472 = ~\u1_u3_idin_reg[27]/P0001  & n2574 ;
  assign n11473 = ~n11471 & ~n11472 ;
  assign n11474 = ~n2573 & ~n11473 ;
  assign n11475 = ~\u4_u3_buf0_orig_reg[27]/P0001  & n2573 ;
  assign n11476 = ~n11474 & ~n11475 ;
  assign n11477 = ~n2572 & n11476 ;
  assign n11478 = n11470 & ~n11477 ;
  assign n11479 = \wb_data_i[28]_pad  & n2568 ;
  assign n11480 = n2567 & n11479 ;
  assign n11481 = rst_i_pad & ~n11480 ;
  assign n11482 = ~\u4_u3_buf0_reg[28]/P0001  & ~n2574 ;
  assign n11483 = ~\u1_u3_idin_reg[28]/P0001  & n2574 ;
  assign n11484 = ~n11482 & ~n11483 ;
  assign n11485 = ~n2573 & ~n11484 ;
  assign n11486 = ~\u4_u3_buf0_orig_reg[28]/P0001  & n2573 ;
  assign n11487 = ~n11485 & ~n11486 ;
  assign n11488 = ~n2572 & n11487 ;
  assign n11489 = n11481 & ~n11488 ;
  assign n11490 = \wb_data_i[29]_pad  & n2568 ;
  assign n11491 = n2567 & n11490 ;
  assign n11492 = rst_i_pad & ~n11491 ;
  assign n11493 = ~\u4_u3_buf0_reg[29]/P0001  & ~n2574 ;
  assign n11494 = ~\u1_u3_idin_reg[29]/P0001  & n2574 ;
  assign n11495 = ~n11493 & ~n11494 ;
  assign n11496 = ~n2573 & ~n11495 ;
  assign n11497 = ~\u4_u3_buf0_orig_reg[29]/NET0131  & n2573 ;
  assign n11498 = ~n11496 & ~n11497 ;
  assign n11499 = ~n2572 & n11498 ;
  assign n11500 = n11492 & ~n11499 ;
  assign n11501 = \wb_data_i[2]_pad  & n2568 ;
  assign n11502 = n2567 & n11501 ;
  assign n11503 = rst_i_pad & ~n11502 ;
  assign n11504 = ~\u4_u3_buf0_reg[2]/P0001  & ~n2574 ;
  assign n11505 = ~\u1_u3_idin_reg[2]/P0001  & n2574 ;
  assign n11506 = ~n11504 & ~n11505 ;
  assign n11507 = ~n2573 & ~n11506 ;
  assign n11508 = ~\u4_u3_buf0_orig_reg[2]/P0001  & n2573 ;
  assign n11509 = ~n11507 & ~n11508 ;
  assign n11510 = ~n2572 & n11509 ;
  assign n11511 = n11503 & ~n11510 ;
  assign n11512 = \wb_data_i[30]_pad  & n2568 ;
  assign n11513 = n2567 & n11512 ;
  assign n11514 = rst_i_pad & ~n11513 ;
  assign n11515 = ~\u4_u3_buf0_reg[30]/P0001  & ~n2574 ;
  assign n11516 = ~\u1_u3_idin_reg[30]/P0001  & n2574 ;
  assign n11517 = ~n11515 & ~n11516 ;
  assign n11518 = ~n2573 & ~n11517 ;
  assign n11519 = ~\u4_u3_buf0_orig_reg[30]/NET0131  & n2573 ;
  assign n11520 = ~n11518 & ~n11519 ;
  assign n11521 = ~n2572 & n11520 ;
  assign n11522 = n11514 & ~n11521 ;
  assign n11523 = \wb_data_i[31]_pad  & n2568 ;
  assign n11524 = n2567 & n11523 ;
  assign n11525 = rst_i_pad & ~n11524 ;
  assign n11526 = ~\u4_u3_buf0_reg[31]/P0001  & ~n2574 ;
  assign n11527 = ~\u1_u3_idin_reg[31]/P0001  & n2574 ;
  assign n11528 = ~n11526 & ~n11527 ;
  assign n11529 = ~n2573 & ~n11528 ;
  assign n11530 = ~\u4_u3_buf0_orig_reg[31]/P0001  & n2573 ;
  assign n11531 = ~n11529 & ~n11530 ;
  assign n11532 = ~n2572 & n11531 ;
  assign n11533 = n11525 & ~n11532 ;
  assign n11534 = \wb_data_i[3]_pad  & n2568 ;
  assign n11535 = n2567 & n11534 ;
  assign n11536 = rst_i_pad & ~n11535 ;
  assign n11537 = ~\u4_u3_buf0_reg[3]/P0001  & ~n2574 ;
  assign n11538 = ~\u1_u3_idin_reg[3]/P0001  & n2574 ;
  assign n11539 = ~n11537 & ~n11538 ;
  assign n11540 = ~n2573 & ~n11539 ;
  assign n11541 = ~\u4_u3_buf0_orig_reg[3]/P0001  & n2573 ;
  assign n11542 = ~n11540 & ~n11541 ;
  assign n11543 = ~n2572 & n11542 ;
  assign n11544 = n11536 & ~n11543 ;
  assign n11545 = \wb_data_i[8]_pad  & n2568 ;
  assign n11546 = n2567 & n11545 ;
  assign n11547 = rst_i_pad & ~n11546 ;
  assign n11548 = ~\u4_u3_buf0_reg[8]/P0001  & ~n2574 ;
  assign n11549 = ~\u1_u3_idin_reg[8]/P0001  & n2574 ;
  assign n11550 = ~n11548 & ~n11549 ;
  assign n11551 = ~n2573 & ~n11550 ;
  assign n11552 = ~\u4_u3_buf0_orig_reg[8]/P0001  & n2573 ;
  assign n11553 = ~n11551 & ~n11552 ;
  assign n11554 = ~n2572 & n11553 ;
  assign n11555 = n11547 & ~n11554 ;
  assign n11556 = \wb_data_i[9]_pad  & n2568 ;
  assign n11557 = n2567 & n11556 ;
  assign n11558 = rst_i_pad & ~n11557 ;
  assign n11559 = ~\u4_u3_buf0_reg[9]/P0001  & ~n2574 ;
  assign n11560 = ~\u1_u3_idin_reg[9]/P0001  & n2574 ;
  assign n11561 = ~n11559 & ~n11560 ;
  assign n11562 = ~n2573 & ~n11561 ;
  assign n11563 = ~\u4_u3_buf0_orig_reg[9]/P0001  & n2573 ;
  assign n11564 = ~n11562 & ~n11563 ;
  assign n11565 = ~n2572 & n11564 ;
  assign n11566 = n11558 & ~n11565 ;
  assign n11567 = \u4_u3_int_stat_reg[0]/P0001  & n5455 ;
  assign n11568 = \u4_u3_ep_match_r_reg/P0001  & n5455 ;
  assign n11569 = ~n11310 & n11568 ;
  assign n11570 = ~n11567 & ~n11569 ;
  assign n11571 = n4061 & n4074 ;
  assign n11572 = n4070 & n11571 ;
  assign n11573 = n9856 & n11572 ;
  assign n11574 = ~\u1_u2_wr_done_reg/P0001  & ~\u1_u2_wr_last_reg/P0001  ;
  assign n11575 = ~\u1_u3_abort_reg/P0001  & n11574 ;
  assign n11576 = n4082 & n11575 ;
  assign n11577 = ~n11573 & ~n11576 ;
  assign n11578 = rst_i_pad & ~n11577 ;
  assign n11579 = n2587 & n11314 ;
  assign n11580 = rst_i_pad & ~n11579 ;
  assign n11581 = ~\u4_u0_buf0_reg[0]/P0001  & ~n2592 ;
  assign n11582 = ~\u1_u3_idin_reg[0]/P0001  & n2592 ;
  assign n11583 = ~n11581 & ~n11582 ;
  assign n11584 = ~n2591 & ~n11583 ;
  assign n11585 = ~\u4_u0_buf0_orig_reg[0]/P0001  & n2591 ;
  assign n11586 = ~n11584 & ~n11585 ;
  assign n11587 = ~n2590 & n11586 ;
  assign n11588 = n11580 & ~n11587 ;
  assign n11589 = n2587 & n11325 ;
  assign n11590 = rst_i_pad & ~n11589 ;
  assign n11591 = ~\u4_u0_buf0_reg[12]/P0001  & ~n2592 ;
  assign n11592 = ~\u1_u3_idin_reg[12]/P0001  & n2592 ;
  assign n11593 = ~n11591 & ~n11592 ;
  assign n11594 = ~n2591 & ~n11593 ;
  assign n11595 = ~\u4_u0_buf0_orig_reg[12]/P0001  & n2591 ;
  assign n11596 = ~n11594 & ~n11595 ;
  assign n11597 = ~n2590 & n11596 ;
  assign n11598 = n11590 & ~n11597 ;
  assign n11599 = n2587 & n11336 ;
  assign n11600 = rst_i_pad & ~n11599 ;
  assign n11601 = ~\u4_u0_buf0_reg[16]/P0001  & ~n2592 ;
  assign n11602 = ~\u1_u3_idin_reg[16]/P0001  & n2592 ;
  assign n11603 = ~n11601 & ~n11602 ;
  assign n11604 = ~n2591 & ~n11603 ;
  assign n11605 = ~\u4_u0_buf0_orig_reg[16]/P0001  & n2591 ;
  assign n11606 = ~n11604 & ~n11605 ;
  assign n11607 = ~n2590 & n11606 ;
  assign n11608 = n11600 & ~n11607 ;
  assign n11609 = n2587 & n11347 ;
  assign n11610 = rst_i_pad & ~n11609 ;
  assign n11611 = ~\u4_u0_buf0_reg[17]/P0001  & ~n2592 ;
  assign n11612 = ~\u1_u3_idin_reg[17]/P0001  & n2592 ;
  assign n11613 = ~n11611 & ~n11612 ;
  assign n11614 = ~n2591 & ~n11613 ;
  assign n11615 = ~\u4_u0_buf0_orig_reg[17]/P0001  & n2591 ;
  assign n11616 = ~n11614 & ~n11615 ;
  assign n11617 = ~n2590 & n11616 ;
  assign n11618 = n11610 & ~n11617 ;
  assign n11619 = n2587 & n11358 ;
  assign n11620 = rst_i_pad & ~n11619 ;
  assign n11621 = ~\u4_u0_buf0_reg[18]/P0001  & ~n2592 ;
  assign n11622 = ~\u1_u3_idin_reg[18]/P0001  & n2592 ;
  assign n11623 = ~n11621 & ~n11622 ;
  assign n11624 = ~n2591 & ~n11623 ;
  assign n11625 = ~\u4_u0_buf0_orig_reg[18]/P0001  & n2591 ;
  assign n11626 = ~n11624 & ~n11625 ;
  assign n11627 = ~n2590 & n11626 ;
  assign n11628 = n11620 & ~n11627 ;
  assign n11629 = n2587 & n11369 ;
  assign n11630 = rst_i_pad & ~n11629 ;
  assign n11631 = ~\u4_u0_buf0_reg[19]/P0001  & ~n2592 ;
  assign n11632 = ~\u1_u3_idin_reg[19]/P0001  & n2592 ;
  assign n11633 = ~n11631 & ~n11632 ;
  assign n11634 = ~n2591 & ~n11633 ;
  assign n11635 = ~\u4_u0_buf0_orig_reg[19]/P0001  & n2591 ;
  assign n11636 = ~n11634 & ~n11635 ;
  assign n11637 = ~n2590 & n11636 ;
  assign n11638 = n11630 & ~n11637 ;
  assign n11639 = n2587 & n11380 ;
  assign n11640 = rst_i_pad & ~n11639 ;
  assign n11641 = ~\u4_u0_buf0_reg[1]/P0001  & ~n2592 ;
  assign n11642 = ~\u1_u3_idin_reg[1]/P0001  & n2592 ;
  assign n11643 = ~n11641 & ~n11642 ;
  assign n11644 = ~n2591 & ~n11643 ;
  assign n11645 = ~\u4_u0_buf0_orig_reg[1]/P0001  & n2591 ;
  assign n11646 = ~n11644 & ~n11645 ;
  assign n11647 = ~n2590 & n11646 ;
  assign n11648 = n11640 & ~n11647 ;
  assign n11649 = n2587 & n11391 ;
  assign n11650 = rst_i_pad & ~n11649 ;
  assign n11651 = ~\u4_u0_buf0_reg[20]/P0001  & ~n2592 ;
  assign n11652 = ~\u1_u3_idin_reg[20]/P0001  & n2592 ;
  assign n11653 = ~n11651 & ~n11652 ;
  assign n11654 = ~n2591 & ~n11653 ;
  assign n11655 = ~\u4_u0_buf0_orig_reg[20]/P0001  & n2591 ;
  assign n11656 = ~n11654 & ~n11655 ;
  assign n11657 = ~n2590 & n11656 ;
  assign n11658 = n11650 & ~n11657 ;
  assign n11659 = n2587 & n11402 ;
  assign n11660 = rst_i_pad & ~n11659 ;
  assign n11661 = ~\u4_u0_buf0_reg[21]/P0001  & ~n2592 ;
  assign n11662 = ~\u1_u3_idin_reg[21]/P0001  & n2592 ;
  assign n11663 = ~n11661 & ~n11662 ;
  assign n11664 = ~n2591 & ~n11663 ;
  assign n11665 = ~\u4_u0_buf0_orig_reg[21]/P0001  & n2591 ;
  assign n11666 = ~n11664 & ~n11665 ;
  assign n11667 = ~n2590 & n11666 ;
  assign n11668 = n11660 & ~n11667 ;
  assign n11669 = n2587 & n11413 ;
  assign n11670 = rst_i_pad & ~n11669 ;
  assign n11671 = ~\u4_u0_buf0_reg[22]/P0001  & ~n2592 ;
  assign n11672 = ~\u1_u3_idin_reg[22]/P0001  & n2592 ;
  assign n11673 = ~n11671 & ~n11672 ;
  assign n11674 = ~n2591 & ~n11673 ;
  assign n11675 = ~\u4_u0_buf0_orig_reg[22]/P0001  & n2591 ;
  assign n11676 = ~n11674 & ~n11675 ;
  assign n11677 = ~n2590 & n11676 ;
  assign n11678 = n11670 & ~n11677 ;
  assign n11679 = n2587 & n11424 ;
  assign n11680 = rst_i_pad & ~n11679 ;
  assign n11681 = ~\u4_u0_buf0_reg[23]/P0001  & ~n2592 ;
  assign n11682 = ~\u1_u3_idin_reg[23]/P0001  & n2592 ;
  assign n11683 = ~n11681 & ~n11682 ;
  assign n11684 = ~n2591 & ~n11683 ;
  assign n11685 = ~\u4_u0_buf0_orig_reg[23]/P0001  & n2591 ;
  assign n11686 = ~n11684 & ~n11685 ;
  assign n11687 = ~n2590 & n11686 ;
  assign n11688 = n11680 & ~n11687 ;
  assign n11689 = n2587 & n11435 ;
  assign n11690 = rst_i_pad & ~n11689 ;
  assign n11691 = ~\u4_u0_buf0_reg[24]/P0001  & ~n2592 ;
  assign n11692 = ~\u1_u3_idin_reg[24]/P0001  & n2592 ;
  assign n11693 = ~n11691 & ~n11692 ;
  assign n11694 = ~n2591 & ~n11693 ;
  assign n11695 = ~\u4_u0_buf0_orig_reg[24]/P0001  & n2591 ;
  assign n11696 = ~n11694 & ~n11695 ;
  assign n11697 = ~n2590 & n11696 ;
  assign n11698 = n11690 & ~n11697 ;
  assign n11699 = n2587 & n11446 ;
  assign n11700 = rst_i_pad & ~n11699 ;
  assign n11701 = ~\u4_u0_buf0_reg[25]/P0001  & ~n2592 ;
  assign n11702 = ~\u1_u3_idin_reg[25]/P0001  & n2592 ;
  assign n11703 = ~n11701 & ~n11702 ;
  assign n11704 = ~n2591 & ~n11703 ;
  assign n11705 = ~\u4_u0_buf0_orig_reg[25]/P0001  & n2591 ;
  assign n11706 = ~n11704 & ~n11705 ;
  assign n11707 = ~n2590 & n11706 ;
  assign n11708 = n11700 & ~n11707 ;
  assign n11709 = n2587 & n11457 ;
  assign n11710 = rst_i_pad & ~n11709 ;
  assign n11711 = ~\u4_u0_buf0_reg[26]/P0001  & ~n2592 ;
  assign n11712 = ~\u1_u3_idin_reg[26]/P0001  & n2592 ;
  assign n11713 = ~n11711 & ~n11712 ;
  assign n11714 = ~n2591 & ~n11713 ;
  assign n11715 = ~\u4_u0_buf0_orig_reg[26]/P0001  & n2591 ;
  assign n11716 = ~n11714 & ~n11715 ;
  assign n11717 = ~n2590 & n11716 ;
  assign n11718 = n11710 & ~n11717 ;
  assign n11719 = n2587 & n11468 ;
  assign n11720 = rst_i_pad & ~n11719 ;
  assign n11721 = ~\u4_u0_buf0_reg[27]/P0001  & ~n2592 ;
  assign n11722 = ~\u1_u3_idin_reg[27]/P0001  & n2592 ;
  assign n11723 = ~n11721 & ~n11722 ;
  assign n11724 = ~n2591 & ~n11723 ;
  assign n11725 = ~\u4_u0_buf0_orig_reg[27]/P0001  & n2591 ;
  assign n11726 = ~n11724 & ~n11725 ;
  assign n11727 = ~n2590 & n11726 ;
  assign n11728 = n11720 & ~n11727 ;
  assign n11729 = n2587 & n11479 ;
  assign n11730 = rst_i_pad & ~n11729 ;
  assign n11731 = ~\u4_u0_buf0_reg[28]/P0001  & ~n2592 ;
  assign n11732 = ~\u1_u3_idin_reg[28]/P0001  & n2592 ;
  assign n11733 = ~n11731 & ~n11732 ;
  assign n11734 = ~n2591 & ~n11733 ;
  assign n11735 = ~\u4_u0_buf0_orig_reg[28]/P0001  & n2591 ;
  assign n11736 = ~n11734 & ~n11735 ;
  assign n11737 = ~n2590 & n11736 ;
  assign n11738 = n11730 & ~n11737 ;
  assign n11739 = n2587 & n11490 ;
  assign n11740 = rst_i_pad & ~n11739 ;
  assign n11741 = ~\u4_u0_buf0_reg[29]/P0001  & ~n2592 ;
  assign n11742 = ~\u1_u3_idin_reg[29]/P0001  & n2592 ;
  assign n11743 = ~n11741 & ~n11742 ;
  assign n11744 = ~n2591 & ~n11743 ;
  assign n11745 = ~\u4_u0_buf0_orig_reg[29]/NET0131  & n2591 ;
  assign n11746 = ~n11744 & ~n11745 ;
  assign n11747 = ~n2590 & n11746 ;
  assign n11748 = n11740 & ~n11747 ;
  assign n11749 = n2587 & n11501 ;
  assign n11750 = rst_i_pad & ~n11749 ;
  assign n11751 = ~\u4_u0_buf0_reg[2]/P0001  & ~n2592 ;
  assign n11752 = ~\u1_u3_idin_reg[2]/P0001  & n2592 ;
  assign n11753 = ~n11751 & ~n11752 ;
  assign n11754 = ~n2591 & ~n11753 ;
  assign n11755 = ~\u4_u0_buf0_orig_reg[2]/P0001  & n2591 ;
  assign n11756 = ~n11754 & ~n11755 ;
  assign n11757 = ~n2590 & n11756 ;
  assign n11758 = n11750 & ~n11757 ;
  assign n11759 = n2587 & n11512 ;
  assign n11760 = rst_i_pad & ~n11759 ;
  assign n11761 = ~\u4_u0_buf0_reg[30]/P0001  & ~n2592 ;
  assign n11762 = ~\u1_u3_idin_reg[30]/P0001  & n2592 ;
  assign n11763 = ~n11761 & ~n11762 ;
  assign n11764 = ~n2591 & ~n11763 ;
  assign n11765 = ~\u4_u0_buf0_orig_reg[30]/NET0131  & n2591 ;
  assign n11766 = ~n11764 & ~n11765 ;
  assign n11767 = ~n2590 & n11766 ;
  assign n11768 = n11760 & ~n11767 ;
  assign n11769 = n2587 & n11523 ;
  assign n11770 = rst_i_pad & ~n11769 ;
  assign n11771 = ~\u4_u0_buf0_reg[31]/P0001  & ~n2592 ;
  assign n11772 = ~\u1_u3_idin_reg[31]/P0001  & n2592 ;
  assign n11773 = ~n11771 & ~n11772 ;
  assign n11774 = ~n2591 & ~n11773 ;
  assign n11775 = ~\u4_u0_buf0_orig_reg[31]/P0001  & n2591 ;
  assign n11776 = ~n11774 & ~n11775 ;
  assign n11777 = ~n2590 & n11776 ;
  assign n11778 = n11770 & ~n11777 ;
  assign n11779 = n2587 & n11534 ;
  assign n11780 = rst_i_pad & ~n11779 ;
  assign n11781 = ~\u4_u0_buf0_reg[3]/P0001  & ~n2592 ;
  assign n11782 = ~\u1_u3_idin_reg[3]/P0001  & n2592 ;
  assign n11783 = ~n11781 & ~n11782 ;
  assign n11784 = ~n2591 & ~n11783 ;
  assign n11785 = ~\u4_u0_buf0_orig_reg[3]/P0001  & n2591 ;
  assign n11786 = ~n11784 & ~n11785 ;
  assign n11787 = ~n2590 & n11786 ;
  assign n11788 = n11780 & ~n11787 ;
  assign n11789 = n2587 & n11545 ;
  assign n11790 = rst_i_pad & ~n11789 ;
  assign n11791 = ~\u4_u0_buf0_reg[8]/P0001  & ~n2592 ;
  assign n11792 = ~\u1_u3_idin_reg[8]/P0001  & n2592 ;
  assign n11793 = ~n11791 & ~n11792 ;
  assign n11794 = ~n2591 & ~n11793 ;
  assign n11795 = ~\u4_u0_buf0_orig_reg[8]/P0001  & n2591 ;
  assign n11796 = ~n11794 & ~n11795 ;
  assign n11797 = ~n2590 & n11796 ;
  assign n11798 = n11790 & ~n11797 ;
  assign n11799 = n2587 & n11556 ;
  assign n11800 = rst_i_pad & ~n11799 ;
  assign n11801 = ~\u4_u0_buf0_reg[9]/P0001  & ~n2592 ;
  assign n11802 = ~\u1_u3_idin_reg[9]/P0001  & n2592 ;
  assign n11803 = ~n11801 & ~n11802 ;
  assign n11804 = ~n2591 & ~n11803 ;
  assign n11805 = ~\u4_u0_buf0_orig_reg[9]/P0001  & n2591 ;
  assign n11806 = ~n11804 & ~n11805 ;
  assign n11807 = ~n2590 & n11806 ;
  assign n11808 = n11800 & ~n11807 ;
  assign n11809 = ~\u0_u0_idle_cnt1_next_reg[3]/P0001  & n8674 ;
  assign n11810 = ~\u0_u0_idle_cnt1_reg[3]/P0001  & ~n8674 ;
  assign n11811 = n8673 & ~n11810 ;
  assign n11812 = ~n11809 & n11811 ;
  assign n11813 = ~n8672 & n11812 ;
  assign n11814 = ~n8666 & n11813 ;
  assign n11815 = \u4_u0_int_stat_reg[0]/P0001  & n5459 ;
  assign n11816 = \u4_u0_ep_match_r_reg/P0001  & n5459 ;
  assign n11817 = ~n11310 & n11816 ;
  assign n11818 = ~n11815 & ~n11817 ;
  assign n11819 = n2620 & n11314 ;
  assign n11820 = rst_i_pad & ~n11819 ;
  assign n11821 = ~\u4_u1_buf0_reg[0]/P0001  & ~n2625 ;
  assign n11822 = ~\u1_u3_idin_reg[0]/P0001  & n2625 ;
  assign n11823 = ~n11821 & ~n11822 ;
  assign n11824 = ~n2624 & ~n11823 ;
  assign n11825 = ~\u4_u1_buf0_orig_reg[0]/P0001  & n2624 ;
  assign n11826 = ~n11824 & ~n11825 ;
  assign n11827 = ~n2623 & n11826 ;
  assign n11828 = n11820 & ~n11827 ;
  assign n11829 = n2620 & n11325 ;
  assign n11830 = rst_i_pad & ~n11829 ;
  assign n11831 = ~\u4_u1_buf0_reg[12]/P0001  & ~n2625 ;
  assign n11832 = ~\u1_u3_idin_reg[12]/P0001  & n2625 ;
  assign n11833 = ~n11831 & ~n11832 ;
  assign n11834 = ~n2624 & ~n11833 ;
  assign n11835 = ~\u4_u1_buf0_orig_reg[12]/P0001  & n2624 ;
  assign n11836 = ~n11834 & ~n11835 ;
  assign n11837 = ~n2623 & n11836 ;
  assign n11838 = n11830 & ~n11837 ;
  assign n11839 = n2620 & n11336 ;
  assign n11840 = rst_i_pad & ~n11839 ;
  assign n11841 = ~\u4_u1_buf0_reg[16]/P0001  & ~n2625 ;
  assign n11842 = ~\u1_u3_idin_reg[16]/P0001  & n2625 ;
  assign n11843 = ~n11841 & ~n11842 ;
  assign n11844 = ~n2624 & ~n11843 ;
  assign n11845 = ~\u4_u1_buf0_orig_reg[16]/P0001  & n2624 ;
  assign n11846 = ~n11844 & ~n11845 ;
  assign n11847 = ~n2623 & n11846 ;
  assign n11848 = n11840 & ~n11847 ;
  assign n11849 = n2620 & n11347 ;
  assign n11850 = rst_i_pad & ~n11849 ;
  assign n11851 = ~\u4_u1_buf0_reg[17]/P0001  & ~n2625 ;
  assign n11852 = ~\u1_u3_idin_reg[17]/P0001  & n2625 ;
  assign n11853 = ~n11851 & ~n11852 ;
  assign n11854 = ~n2624 & ~n11853 ;
  assign n11855 = ~\u4_u1_buf0_orig_reg[17]/P0001  & n2624 ;
  assign n11856 = ~n11854 & ~n11855 ;
  assign n11857 = ~n2623 & n11856 ;
  assign n11858 = n11850 & ~n11857 ;
  assign n11859 = n2620 & n11358 ;
  assign n11860 = rst_i_pad & ~n11859 ;
  assign n11861 = ~\u4_u1_buf0_reg[18]/P0001  & ~n2625 ;
  assign n11862 = ~\u1_u3_idin_reg[18]/P0001  & n2625 ;
  assign n11863 = ~n11861 & ~n11862 ;
  assign n11864 = ~n2624 & ~n11863 ;
  assign n11865 = ~\u4_u1_buf0_orig_reg[18]/P0001  & n2624 ;
  assign n11866 = ~n11864 & ~n11865 ;
  assign n11867 = ~n2623 & n11866 ;
  assign n11868 = n11860 & ~n11867 ;
  assign n11869 = n2620 & n11369 ;
  assign n11870 = rst_i_pad & ~n11869 ;
  assign n11871 = ~\u4_u1_buf0_reg[19]/P0001  & ~n2625 ;
  assign n11872 = ~\u1_u3_idin_reg[19]/P0001  & n2625 ;
  assign n11873 = ~n11871 & ~n11872 ;
  assign n11874 = ~n2624 & ~n11873 ;
  assign n11875 = ~\u4_u1_buf0_orig_reg[19]/P0001  & n2624 ;
  assign n11876 = ~n11874 & ~n11875 ;
  assign n11877 = ~n2623 & n11876 ;
  assign n11878 = n11870 & ~n11877 ;
  assign n11879 = n2620 & n11380 ;
  assign n11880 = rst_i_pad & ~n11879 ;
  assign n11881 = ~\u4_u1_buf0_reg[1]/P0001  & ~n2625 ;
  assign n11882 = ~\u1_u3_idin_reg[1]/P0001  & n2625 ;
  assign n11883 = ~n11881 & ~n11882 ;
  assign n11884 = ~n2624 & ~n11883 ;
  assign n11885 = ~\u4_u1_buf0_orig_reg[1]/P0001  & n2624 ;
  assign n11886 = ~n11884 & ~n11885 ;
  assign n11887 = ~n2623 & n11886 ;
  assign n11888 = n11880 & ~n11887 ;
  assign n11889 = n2620 & n11391 ;
  assign n11890 = rst_i_pad & ~n11889 ;
  assign n11891 = ~\u4_u1_buf0_reg[20]/P0001  & ~n2625 ;
  assign n11892 = ~\u1_u3_idin_reg[20]/P0001  & n2625 ;
  assign n11893 = ~n11891 & ~n11892 ;
  assign n11894 = ~n2624 & ~n11893 ;
  assign n11895 = ~\u4_u1_buf0_orig_reg[20]/P0001  & n2624 ;
  assign n11896 = ~n11894 & ~n11895 ;
  assign n11897 = ~n2623 & n11896 ;
  assign n11898 = n11890 & ~n11897 ;
  assign n11899 = n2620 & n11402 ;
  assign n11900 = rst_i_pad & ~n11899 ;
  assign n11901 = ~\u4_u1_buf0_reg[21]/P0001  & ~n2625 ;
  assign n11902 = ~\u1_u3_idin_reg[21]/P0001  & n2625 ;
  assign n11903 = ~n11901 & ~n11902 ;
  assign n11904 = ~n2624 & ~n11903 ;
  assign n11905 = ~\u4_u1_buf0_orig_reg[21]/P0001  & n2624 ;
  assign n11906 = ~n11904 & ~n11905 ;
  assign n11907 = ~n2623 & n11906 ;
  assign n11908 = n11900 & ~n11907 ;
  assign n11909 = n2620 & n11413 ;
  assign n11910 = rst_i_pad & ~n11909 ;
  assign n11911 = ~\u4_u1_buf0_reg[22]/P0001  & ~n2625 ;
  assign n11912 = ~\u1_u3_idin_reg[22]/P0001  & n2625 ;
  assign n11913 = ~n11911 & ~n11912 ;
  assign n11914 = ~n2624 & ~n11913 ;
  assign n11915 = ~\u4_u1_buf0_orig_reg[22]/P0001  & n2624 ;
  assign n11916 = ~n11914 & ~n11915 ;
  assign n11917 = ~n2623 & n11916 ;
  assign n11918 = n11910 & ~n11917 ;
  assign n11919 = n2620 & n11424 ;
  assign n11920 = rst_i_pad & ~n11919 ;
  assign n11921 = ~\u4_u1_buf0_reg[23]/P0001  & ~n2625 ;
  assign n11922 = ~\u1_u3_idin_reg[23]/P0001  & n2625 ;
  assign n11923 = ~n11921 & ~n11922 ;
  assign n11924 = ~n2624 & ~n11923 ;
  assign n11925 = ~\u4_u1_buf0_orig_reg[23]/P0001  & n2624 ;
  assign n11926 = ~n11924 & ~n11925 ;
  assign n11927 = ~n2623 & n11926 ;
  assign n11928 = n11920 & ~n11927 ;
  assign n11929 = n2620 & n11435 ;
  assign n11930 = rst_i_pad & ~n11929 ;
  assign n11931 = ~\u4_u1_buf0_reg[24]/P0001  & ~n2625 ;
  assign n11932 = ~\u1_u3_idin_reg[24]/P0001  & n2625 ;
  assign n11933 = ~n11931 & ~n11932 ;
  assign n11934 = ~n2624 & ~n11933 ;
  assign n11935 = ~\u4_u1_buf0_orig_reg[24]/P0001  & n2624 ;
  assign n11936 = ~n11934 & ~n11935 ;
  assign n11937 = ~n2623 & n11936 ;
  assign n11938 = n11930 & ~n11937 ;
  assign n11939 = n2620 & n11446 ;
  assign n11940 = rst_i_pad & ~n11939 ;
  assign n11941 = ~\u4_u1_buf0_reg[25]/P0001  & ~n2625 ;
  assign n11942 = ~\u1_u3_idin_reg[25]/P0001  & n2625 ;
  assign n11943 = ~n11941 & ~n11942 ;
  assign n11944 = ~n2624 & ~n11943 ;
  assign n11945 = ~\u4_u1_buf0_orig_reg[25]/P0001  & n2624 ;
  assign n11946 = ~n11944 & ~n11945 ;
  assign n11947 = ~n2623 & n11946 ;
  assign n11948 = n11940 & ~n11947 ;
  assign n11949 = n2620 & n11457 ;
  assign n11950 = rst_i_pad & ~n11949 ;
  assign n11951 = ~\u4_u1_buf0_reg[26]/P0001  & ~n2625 ;
  assign n11952 = ~\u1_u3_idin_reg[26]/P0001  & n2625 ;
  assign n11953 = ~n11951 & ~n11952 ;
  assign n11954 = ~n2624 & ~n11953 ;
  assign n11955 = ~\u4_u1_buf0_orig_reg[26]/P0001  & n2624 ;
  assign n11956 = ~n11954 & ~n11955 ;
  assign n11957 = ~n2623 & n11956 ;
  assign n11958 = n11950 & ~n11957 ;
  assign n11959 = n2620 & n11468 ;
  assign n11960 = rst_i_pad & ~n11959 ;
  assign n11961 = ~\u4_u1_buf0_reg[27]/P0001  & ~n2625 ;
  assign n11962 = ~\u1_u3_idin_reg[27]/P0001  & n2625 ;
  assign n11963 = ~n11961 & ~n11962 ;
  assign n11964 = ~n2624 & ~n11963 ;
  assign n11965 = ~\u4_u1_buf0_orig_reg[27]/P0001  & n2624 ;
  assign n11966 = ~n11964 & ~n11965 ;
  assign n11967 = ~n2623 & n11966 ;
  assign n11968 = n11960 & ~n11967 ;
  assign n11969 = n2620 & n11479 ;
  assign n11970 = rst_i_pad & ~n11969 ;
  assign n11971 = ~\u4_u1_buf0_reg[28]/P0001  & ~n2625 ;
  assign n11972 = ~\u1_u3_idin_reg[28]/P0001  & n2625 ;
  assign n11973 = ~n11971 & ~n11972 ;
  assign n11974 = ~n2624 & ~n11973 ;
  assign n11975 = ~\u4_u1_buf0_orig_reg[28]/P0001  & n2624 ;
  assign n11976 = ~n11974 & ~n11975 ;
  assign n11977 = ~n2623 & n11976 ;
  assign n11978 = n11970 & ~n11977 ;
  assign n11979 = n2620 & n11490 ;
  assign n11980 = rst_i_pad & ~n11979 ;
  assign n11981 = ~\u4_u1_buf0_reg[29]/P0001  & ~n2625 ;
  assign n11982 = ~\u1_u3_idin_reg[29]/P0001  & n2625 ;
  assign n11983 = ~n11981 & ~n11982 ;
  assign n11984 = ~n2624 & ~n11983 ;
  assign n11985 = ~\u4_u1_buf0_orig_reg[29]/NET0131  & n2624 ;
  assign n11986 = ~n11984 & ~n11985 ;
  assign n11987 = ~n2623 & n11986 ;
  assign n11988 = n11980 & ~n11987 ;
  assign n11989 = n2620 & n11501 ;
  assign n11990 = rst_i_pad & ~n11989 ;
  assign n11991 = ~\u4_u1_buf0_reg[2]/P0001  & ~n2625 ;
  assign n11992 = ~\u1_u3_idin_reg[2]/P0001  & n2625 ;
  assign n11993 = ~n11991 & ~n11992 ;
  assign n11994 = ~n2624 & ~n11993 ;
  assign n11995 = ~\u4_u1_buf0_orig_reg[2]/P0001  & n2624 ;
  assign n11996 = ~n11994 & ~n11995 ;
  assign n11997 = ~n2623 & n11996 ;
  assign n11998 = n11990 & ~n11997 ;
  assign n11999 = n2620 & n11512 ;
  assign n12000 = rst_i_pad & ~n11999 ;
  assign n12001 = ~\u4_u1_buf0_reg[30]/P0001  & ~n2625 ;
  assign n12002 = ~\u1_u3_idin_reg[30]/P0001  & n2625 ;
  assign n12003 = ~n12001 & ~n12002 ;
  assign n12004 = ~n2624 & ~n12003 ;
  assign n12005 = ~\u4_u1_buf0_orig_reg[30]/NET0131  & n2624 ;
  assign n12006 = ~n12004 & ~n12005 ;
  assign n12007 = ~n2623 & n12006 ;
  assign n12008 = n12000 & ~n12007 ;
  assign n12009 = n2620 & n11523 ;
  assign n12010 = rst_i_pad & ~n12009 ;
  assign n12011 = ~\u4_u1_buf0_reg[31]/P0001  & ~n2625 ;
  assign n12012 = ~\u1_u3_idin_reg[31]/P0001  & n2625 ;
  assign n12013 = ~n12011 & ~n12012 ;
  assign n12014 = ~n2624 & ~n12013 ;
  assign n12015 = ~\u4_u1_buf0_orig_reg[31]/P0001  & n2624 ;
  assign n12016 = ~n12014 & ~n12015 ;
  assign n12017 = ~n2623 & n12016 ;
  assign n12018 = n12010 & ~n12017 ;
  assign n12019 = n2620 & n11534 ;
  assign n12020 = rst_i_pad & ~n12019 ;
  assign n12021 = ~\u4_u1_buf0_reg[3]/P0001  & ~n2625 ;
  assign n12022 = ~\u1_u3_idin_reg[3]/P0001  & n2625 ;
  assign n12023 = ~n12021 & ~n12022 ;
  assign n12024 = ~n2624 & ~n12023 ;
  assign n12025 = ~\u4_u1_buf0_orig_reg[3]/P0001  & n2624 ;
  assign n12026 = ~n12024 & ~n12025 ;
  assign n12027 = ~n2623 & n12026 ;
  assign n12028 = n12020 & ~n12027 ;
  assign n12029 = n2620 & n11545 ;
  assign n12030 = rst_i_pad & ~n12029 ;
  assign n12031 = ~\u4_u1_buf0_reg[8]/P0001  & ~n2625 ;
  assign n12032 = ~\u1_u3_idin_reg[8]/P0001  & n2625 ;
  assign n12033 = ~n12031 & ~n12032 ;
  assign n12034 = ~n2624 & ~n12033 ;
  assign n12035 = ~\u4_u1_buf0_orig_reg[8]/P0001  & n2624 ;
  assign n12036 = ~n12034 & ~n12035 ;
  assign n12037 = ~n2623 & n12036 ;
  assign n12038 = n12030 & ~n12037 ;
  assign n12039 = n2620 & n11556 ;
  assign n12040 = rst_i_pad & ~n12039 ;
  assign n12041 = ~\u4_u1_buf0_reg[9]/P0001  & ~n2625 ;
  assign n12042 = ~\u1_u3_idin_reg[9]/P0001  & n2625 ;
  assign n12043 = ~n12041 & ~n12042 ;
  assign n12044 = ~n2624 & ~n12043 ;
  assign n12045 = ~\u4_u1_buf0_orig_reg[9]/P0001  & n2624 ;
  assign n12046 = ~n12044 & ~n12045 ;
  assign n12047 = ~n2623 & n12046 ;
  assign n12048 = n12040 & ~n12047 ;
  assign n12049 = \u4_u1_int_stat_reg[0]/P0001  & n5463 ;
  assign n12050 = \u4_u1_ep_match_r_reg/P0001  & n5463 ;
  assign n12051 = ~n11310 & n12050 ;
  assign n12052 = ~n12049 & ~n12051 ;
  assign n12053 = n2635 & n11314 ;
  assign n12054 = rst_i_pad & ~n12053 ;
  assign n12055 = ~\u4_u2_buf0_reg[0]/P0001  & ~n2640 ;
  assign n12056 = ~\u1_u3_idin_reg[0]/P0001  & n2640 ;
  assign n12057 = ~n12055 & ~n12056 ;
  assign n12058 = ~n2639 & ~n12057 ;
  assign n12059 = ~\u4_u2_buf0_orig_reg[0]/P0001  & n2639 ;
  assign n12060 = ~n12058 & ~n12059 ;
  assign n12061 = ~n2638 & n12060 ;
  assign n12062 = n12054 & ~n12061 ;
  assign n12063 = n2635 & n11325 ;
  assign n12064 = rst_i_pad & ~n12063 ;
  assign n12065 = ~\u4_u2_buf0_reg[12]/P0001  & ~n2640 ;
  assign n12066 = ~\u1_u3_idin_reg[12]/P0001  & n2640 ;
  assign n12067 = ~n12065 & ~n12066 ;
  assign n12068 = ~n2639 & ~n12067 ;
  assign n12069 = ~\u4_u2_buf0_orig_reg[12]/P0001  & n2639 ;
  assign n12070 = ~n12068 & ~n12069 ;
  assign n12071 = ~n2638 & n12070 ;
  assign n12072 = n12064 & ~n12071 ;
  assign n12073 = n2635 & n11336 ;
  assign n12074 = rst_i_pad & ~n12073 ;
  assign n12075 = ~\u4_u2_buf0_reg[16]/P0001  & ~n2640 ;
  assign n12076 = ~\u1_u3_idin_reg[16]/P0001  & n2640 ;
  assign n12077 = ~n12075 & ~n12076 ;
  assign n12078 = ~n2639 & ~n12077 ;
  assign n12079 = ~\u4_u2_buf0_orig_reg[16]/P0001  & n2639 ;
  assign n12080 = ~n12078 & ~n12079 ;
  assign n12081 = ~n2638 & n12080 ;
  assign n12082 = n12074 & ~n12081 ;
  assign n12083 = n2635 & n11347 ;
  assign n12084 = rst_i_pad & ~n12083 ;
  assign n12085 = ~\u4_u2_buf0_reg[17]/P0001  & ~n2640 ;
  assign n12086 = ~\u1_u3_idin_reg[17]/P0001  & n2640 ;
  assign n12087 = ~n12085 & ~n12086 ;
  assign n12088 = ~n2639 & ~n12087 ;
  assign n12089 = ~\u4_u2_buf0_orig_reg[17]/P0001  & n2639 ;
  assign n12090 = ~n12088 & ~n12089 ;
  assign n12091 = ~n2638 & n12090 ;
  assign n12092 = n12084 & ~n12091 ;
  assign n12093 = n2635 & n11358 ;
  assign n12094 = rst_i_pad & ~n12093 ;
  assign n12095 = ~\u4_u2_buf0_reg[18]/P0001  & ~n2640 ;
  assign n12096 = ~\u1_u3_idin_reg[18]/P0001  & n2640 ;
  assign n12097 = ~n12095 & ~n12096 ;
  assign n12098 = ~n2639 & ~n12097 ;
  assign n12099 = ~\u4_u2_buf0_orig_reg[18]/P0001  & n2639 ;
  assign n12100 = ~n12098 & ~n12099 ;
  assign n12101 = ~n2638 & n12100 ;
  assign n12102 = n12094 & ~n12101 ;
  assign n12103 = n2635 & n11369 ;
  assign n12104 = rst_i_pad & ~n12103 ;
  assign n12105 = ~\u4_u2_buf0_reg[19]/P0001  & ~n2640 ;
  assign n12106 = ~\u1_u3_idin_reg[19]/P0001  & n2640 ;
  assign n12107 = ~n12105 & ~n12106 ;
  assign n12108 = ~n2639 & ~n12107 ;
  assign n12109 = ~\u4_u2_buf0_orig_reg[19]/P0001  & n2639 ;
  assign n12110 = ~n12108 & ~n12109 ;
  assign n12111 = ~n2638 & n12110 ;
  assign n12112 = n12104 & ~n12111 ;
  assign n12113 = n2635 & n11380 ;
  assign n12114 = rst_i_pad & ~n12113 ;
  assign n12115 = ~\u4_u2_buf0_reg[1]/P0001  & ~n2640 ;
  assign n12116 = ~\u1_u3_idin_reg[1]/P0001  & n2640 ;
  assign n12117 = ~n12115 & ~n12116 ;
  assign n12118 = ~n2639 & ~n12117 ;
  assign n12119 = ~\u4_u2_buf0_orig_reg[1]/P0001  & n2639 ;
  assign n12120 = ~n12118 & ~n12119 ;
  assign n12121 = ~n2638 & n12120 ;
  assign n12122 = n12114 & ~n12121 ;
  assign n12123 = n2635 & n11391 ;
  assign n12124 = rst_i_pad & ~n12123 ;
  assign n12125 = ~\u4_u2_buf0_reg[20]/P0001  & ~n2640 ;
  assign n12126 = ~\u1_u3_idin_reg[20]/P0001  & n2640 ;
  assign n12127 = ~n12125 & ~n12126 ;
  assign n12128 = ~n2639 & ~n12127 ;
  assign n12129 = ~\u4_u2_buf0_orig_reg[20]/P0001  & n2639 ;
  assign n12130 = ~n12128 & ~n12129 ;
  assign n12131 = ~n2638 & n12130 ;
  assign n12132 = n12124 & ~n12131 ;
  assign n12133 = n2635 & n11402 ;
  assign n12134 = rst_i_pad & ~n12133 ;
  assign n12135 = ~\u4_u2_buf0_reg[21]/P0001  & ~n2640 ;
  assign n12136 = ~\u1_u3_idin_reg[21]/P0001  & n2640 ;
  assign n12137 = ~n12135 & ~n12136 ;
  assign n12138 = ~n2639 & ~n12137 ;
  assign n12139 = ~\u4_u2_buf0_orig_reg[21]/P0001  & n2639 ;
  assign n12140 = ~n12138 & ~n12139 ;
  assign n12141 = ~n2638 & n12140 ;
  assign n12142 = n12134 & ~n12141 ;
  assign n12143 = n2635 & n11413 ;
  assign n12144 = rst_i_pad & ~n12143 ;
  assign n12145 = ~\u4_u2_buf0_reg[22]/P0001  & ~n2640 ;
  assign n12146 = ~\u1_u3_idin_reg[22]/P0001  & n2640 ;
  assign n12147 = ~n12145 & ~n12146 ;
  assign n12148 = ~n2639 & ~n12147 ;
  assign n12149 = ~\u4_u2_buf0_orig_reg[22]/P0001  & n2639 ;
  assign n12150 = ~n12148 & ~n12149 ;
  assign n12151 = ~n2638 & n12150 ;
  assign n12152 = n12144 & ~n12151 ;
  assign n12153 = n2635 & n11424 ;
  assign n12154 = rst_i_pad & ~n12153 ;
  assign n12155 = ~\u4_u2_buf0_reg[23]/P0001  & ~n2640 ;
  assign n12156 = ~\u1_u3_idin_reg[23]/P0001  & n2640 ;
  assign n12157 = ~n12155 & ~n12156 ;
  assign n12158 = ~n2639 & ~n12157 ;
  assign n12159 = ~\u4_u2_buf0_orig_reg[23]/P0001  & n2639 ;
  assign n12160 = ~n12158 & ~n12159 ;
  assign n12161 = ~n2638 & n12160 ;
  assign n12162 = n12154 & ~n12161 ;
  assign n12163 = n2635 & n11435 ;
  assign n12164 = rst_i_pad & ~n12163 ;
  assign n12165 = ~\u4_u2_buf0_reg[24]/P0001  & ~n2640 ;
  assign n12166 = ~\u1_u3_idin_reg[24]/P0001  & n2640 ;
  assign n12167 = ~n12165 & ~n12166 ;
  assign n12168 = ~n2639 & ~n12167 ;
  assign n12169 = ~\u4_u2_buf0_orig_reg[24]/P0001  & n2639 ;
  assign n12170 = ~n12168 & ~n12169 ;
  assign n12171 = ~n2638 & n12170 ;
  assign n12172 = n12164 & ~n12171 ;
  assign n12173 = n2635 & n11446 ;
  assign n12174 = rst_i_pad & ~n12173 ;
  assign n12175 = ~\u4_u2_buf0_reg[25]/P0001  & ~n2640 ;
  assign n12176 = ~\u1_u3_idin_reg[25]/P0001  & n2640 ;
  assign n12177 = ~n12175 & ~n12176 ;
  assign n12178 = ~n2639 & ~n12177 ;
  assign n12179 = ~\u4_u2_buf0_orig_reg[25]/P0001  & n2639 ;
  assign n12180 = ~n12178 & ~n12179 ;
  assign n12181 = ~n2638 & n12180 ;
  assign n12182 = n12174 & ~n12181 ;
  assign n12183 = n2635 & n11457 ;
  assign n12184 = rst_i_pad & ~n12183 ;
  assign n12185 = ~\u4_u2_buf0_reg[26]/P0001  & ~n2640 ;
  assign n12186 = ~\u1_u3_idin_reg[26]/P0001  & n2640 ;
  assign n12187 = ~n12185 & ~n12186 ;
  assign n12188 = ~n2639 & ~n12187 ;
  assign n12189 = ~\u4_u2_buf0_orig_reg[26]/P0001  & n2639 ;
  assign n12190 = ~n12188 & ~n12189 ;
  assign n12191 = ~n2638 & n12190 ;
  assign n12192 = n12184 & ~n12191 ;
  assign n12193 = n2635 & n11468 ;
  assign n12194 = rst_i_pad & ~n12193 ;
  assign n12195 = ~\u4_u2_buf0_reg[27]/P0001  & ~n2640 ;
  assign n12196 = ~\u1_u3_idin_reg[27]/P0001  & n2640 ;
  assign n12197 = ~n12195 & ~n12196 ;
  assign n12198 = ~n2639 & ~n12197 ;
  assign n12199 = ~\u4_u2_buf0_orig_reg[27]/P0001  & n2639 ;
  assign n12200 = ~n12198 & ~n12199 ;
  assign n12201 = ~n2638 & n12200 ;
  assign n12202 = n12194 & ~n12201 ;
  assign n12203 = n2635 & n11479 ;
  assign n12204 = rst_i_pad & ~n12203 ;
  assign n12205 = ~\u4_u2_buf0_reg[28]/P0001  & ~n2640 ;
  assign n12206 = ~\u1_u3_idin_reg[28]/P0001  & n2640 ;
  assign n12207 = ~n12205 & ~n12206 ;
  assign n12208 = ~n2639 & ~n12207 ;
  assign n12209 = ~\u4_u2_buf0_orig_reg[28]/P0001  & n2639 ;
  assign n12210 = ~n12208 & ~n12209 ;
  assign n12211 = ~n2638 & n12210 ;
  assign n12212 = n12204 & ~n12211 ;
  assign n12213 = n2635 & n11490 ;
  assign n12214 = rst_i_pad & ~n12213 ;
  assign n12215 = ~\u4_u2_buf0_reg[29]/P0001  & ~n2640 ;
  assign n12216 = ~\u1_u3_idin_reg[29]/P0001  & n2640 ;
  assign n12217 = ~n12215 & ~n12216 ;
  assign n12218 = ~n2639 & ~n12217 ;
  assign n12219 = ~\u4_u2_buf0_orig_reg[29]/NET0131  & n2639 ;
  assign n12220 = ~n12218 & ~n12219 ;
  assign n12221 = ~n2638 & n12220 ;
  assign n12222 = n12214 & ~n12221 ;
  assign n12223 = n2635 & n11501 ;
  assign n12224 = rst_i_pad & ~n12223 ;
  assign n12225 = ~\u4_u2_buf0_reg[2]/P0001  & ~n2640 ;
  assign n12226 = ~\u1_u3_idin_reg[2]/P0001  & n2640 ;
  assign n12227 = ~n12225 & ~n12226 ;
  assign n12228 = ~n2639 & ~n12227 ;
  assign n12229 = ~\u4_u2_buf0_orig_reg[2]/P0001  & n2639 ;
  assign n12230 = ~n12228 & ~n12229 ;
  assign n12231 = ~n2638 & n12230 ;
  assign n12232 = n12224 & ~n12231 ;
  assign n12233 = n2635 & n11512 ;
  assign n12234 = rst_i_pad & ~n12233 ;
  assign n12235 = ~\u4_u2_buf0_reg[30]/P0001  & ~n2640 ;
  assign n12236 = ~\u1_u3_idin_reg[30]/P0001  & n2640 ;
  assign n12237 = ~n12235 & ~n12236 ;
  assign n12238 = ~n2639 & ~n12237 ;
  assign n12239 = ~\u4_u2_buf0_orig_reg[30]/NET0131  & n2639 ;
  assign n12240 = ~n12238 & ~n12239 ;
  assign n12241 = ~n2638 & n12240 ;
  assign n12242 = n12234 & ~n12241 ;
  assign n12243 = n2635 & n11523 ;
  assign n12244 = rst_i_pad & ~n12243 ;
  assign n12245 = ~\u4_u2_buf0_reg[31]/P0001  & ~n2640 ;
  assign n12246 = ~\u1_u3_idin_reg[31]/P0001  & n2640 ;
  assign n12247 = ~n12245 & ~n12246 ;
  assign n12248 = ~n2639 & ~n12247 ;
  assign n12249 = ~\u4_u2_buf0_orig_reg[31]/P0001  & n2639 ;
  assign n12250 = ~n12248 & ~n12249 ;
  assign n12251 = ~n2638 & n12250 ;
  assign n12252 = n12244 & ~n12251 ;
  assign n12253 = n2635 & n11534 ;
  assign n12254 = rst_i_pad & ~n12253 ;
  assign n12255 = ~\u4_u2_buf0_reg[3]/P0001  & ~n2640 ;
  assign n12256 = ~\u1_u3_idin_reg[3]/P0001  & n2640 ;
  assign n12257 = ~n12255 & ~n12256 ;
  assign n12258 = ~n2639 & ~n12257 ;
  assign n12259 = ~\u4_u2_buf0_orig_reg[3]/P0001  & n2639 ;
  assign n12260 = ~n12258 & ~n12259 ;
  assign n12261 = ~n2638 & n12260 ;
  assign n12262 = n12254 & ~n12261 ;
  assign n12263 = n2635 & n11545 ;
  assign n12264 = rst_i_pad & ~n12263 ;
  assign n12265 = ~\u4_u2_buf0_reg[8]/P0001  & ~n2640 ;
  assign n12266 = ~\u1_u3_idin_reg[8]/P0001  & n2640 ;
  assign n12267 = ~n12265 & ~n12266 ;
  assign n12268 = ~n2639 & ~n12267 ;
  assign n12269 = ~\u4_u2_buf0_orig_reg[8]/P0001  & n2639 ;
  assign n12270 = ~n12268 & ~n12269 ;
  assign n12271 = ~n2638 & n12270 ;
  assign n12272 = n12264 & ~n12271 ;
  assign n12273 = n2635 & n11556 ;
  assign n12274 = rst_i_pad & ~n12273 ;
  assign n12275 = ~\u4_u2_buf0_reg[9]/P0001  & ~n2640 ;
  assign n12276 = ~\u1_u3_idin_reg[9]/P0001  & n2640 ;
  assign n12277 = ~n12275 & ~n12276 ;
  assign n12278 = ~n2639 & ~n12277 ;
  assign n12279 = ~\u4_u2_buf0_orig_reg[9]/P0001  & n2639 ;
  assign n12280 = ~n12278 & ~n12279 ;
  assign n12281 = ~n2638 & n12280 ;
  assign n12282 = n12274 & ~n12281 ;
  assign n12283 = ~\u4_attach_r1_reg/P0001  & \u4_attach_r_reg/P0001  ;
  assign n12284 = ~\u4_int_srcb_reg[5]/P0001  & ~n12283 ;
  assign n12285 = n5667 & ~n12284 ;
  assign n12286 = \u4_attach_r1_reg/P0001  & ~\u4_attach_r_reg/P0001  ;
  assign n12287 = ~\u4_int_srcb_reg[6]/P0001  & ~n12286 ;
  assign n12288 = n5667 & ~n12287 ;
  assign n12289 = \u0_u0_mode_hs_reg/P0001  & \u4_csr_reg[11]/P0001  ;
  assign n12290 = \u4_csr_reg[29]/P0001  & n12289 ;
  assign n12291 = \u0_u0_mode_hs_reg/P0001  & \u4_csr_reg[12]/P0001  ;
  assign n12292 = \u4_csr_reg[24]/P0001  & \u4_csr_reg[27]/NET0131  ;
  assign n12293 = n12291 & n12292 ;
  assign n12294 = n12290 & n12293 ;
  assign n12295 = ~n2358 & ~n12294 ;
  assign n12296 = ~\u4_csr_reg[28]/P0001  & n12289 ;
  assign n12297 = n12293 & ~n12296 ;
  assign n12298 = ~n2358 & ~n12297 ;
  assign n12299 = ~n12295 & ~n12298 ;
  assign n12300 = ~\u1_u3_setup_token_reg/P0001  & \u4_csr_reg[28]/P0001  ;
  assign n12301 = ~n3036 & n12300 ;
  assign n12302 = n12299 & ~n12301 ;
  assign n12303 = \u4_csr_reg[12]/P0001  & ~\u4_csr_reg[29]/P0001  ;
  assign n12304 = n12289 & n12303 ;
  assign n12305 = n12292 & n12304 ;
  assign n12306 = n12295 & ~n12305 ;
  assign n12307 = ~n12297 & ~n12306 ;
  assign n12308 = n5007 & n7806 ;
  assign n12309 = ~n2358 & n12308 ;
  assign n12310 = ~n12305 & n12309 ;
  assign n12311 = ~n12294 & n12309 ;
  assign n12312 = ~n12310 & ~n12311 ;
  assign n12313 = n12307 & ~n12312 ;
  assign n12314 = n12297 & n12308 ;
  assign n12315 = ~\u4_csr_reg[25]/P0001  & n12291 ;
  assign n12316 = ~n12290 & n12315 ;
  assign n12317 = \u4_csr_reg[24]/P0001  & ~n12316 ;
  assign n12318 = ~\u4_csr_reg[24]/P0001  & ~\u4_csr_reg[26]/NET0131  ;
  assign n12319 = \u4_csr_reg[27]/NET0131  & ~n12318 ;
  assign n12320 = ~\u4_csr_reg[28]/P0001  & ~n12319 ;
  assign n12321 = ~n12317 & n12320 ;
  assign n12322 = ~n12314 & ~n12321 ;
  assign n12323 = n12306 & ~n12322 ;
  assign n12324 = ~n12313 & ~n12323 ;
  assign n12325 = ~n12302 & n12324 ;
  assign n12326 = ~n9208 & ~n9249 ;
  assign n12327 = n9244 & ~n12326 ;
  assign n12328 = ~n9244 & n12326 ;
  assign n12329 = ~n12327 & ~n12328 ;
  assign n12330 = ~n9061 & ~n9102 ;
  assign n12331 = n9097 & ~n12330 ;
  assign n12332 = ~n9097 & n12330 ;
  assign n12333 = ~n12331 & ~n12332 ;
  assign n12334 = ~\u0_u0_state_reg[6]/NET0131  & ~\u0_u0_state_reg[7]/NET0131  ;
  assign n12335 = ~\u0_u0_state_reg[8]/NET0131  & n12334 ;
  assign n12336 = n5740 & n12335 ;
  assign n12337 = ~\u0_u0_state_reg[0]/NET0131  & ~\u0_u0_state_reg[2]/NET0131  ;
  assign n12338 = ~\u0_u0_state_reg[1]/P0001  & ~\u0_u0_state_reg[3]/P0001  ;
  assign n12339 = n12337 & n12338 ;
  assign n12340 = n12336 & n12339 ;
  assign n12341 = ~\u0_u0_state_reg[10]/P0001  & n5744 ;
  assign n12342 = \u0_u0_state_reg[13]/NET0131  & ~\u0_u0_state_reg[9]/P0001  ;
  assign n12343 = ~\u0_u0_state_reg[14]/P0001  & ~\u0_u0_state_reg[4]/NET0131  ;
  assign n12344 = n12342 & n12343 ;
  assign n12345 = n12341 & n12344 ;
  assign n12346 = n12340 & n12345 ;
  assign n12347 = \u0_u0_T2_wakeup_reg/P0001  & ~\u0_u0_state_reg[1]/P0001  ;
  assign n12348 = \u0_u0_state_reg[5]/P0001  & n12347 ;
  assign n12349 = \u0_u0_state_reg[1]/P0001  & ~\u0_u0_state_reg[5]/P0001  ;
  assign n12350 = n6147 & n12349 ;
  assign n12351 = ~TermSel_pad_o_pad & ~n12350 ;
  assign n12352 = ~n12348 & n12351 ;
  assign n12353 = \u0_u0_mode_hs_reg/P0001  & \u0_u0_state_reg[4]/NET0131  ;
  assign n12354 = n5765 & n12353 ;
  assign n12355 = ~n12352 & ~n12354 ;
  assign n12356 = ~n12346 & n12355 ;
  assign n12357 = ~\u0_u0_state_reg[10]/P0001  & ~\u0_u0_state_reg[13]/NET0131  ;
  assign n12358 = \u0_u0_state_reg[0]/NET0131  & ~\u0_u0_state_reg[7]/NET0131  ;
  assign n12359 = n5736 & n12358 ;
  assign n12360 = ~\u0_u0_state_reg[14]/P0001  & n12359 ;
  assign n12361 = ~\u0_u0_state_reg[1]/P0001  & ~\u0_u0_state_reg[5]/P0001  ;
  assign n12362 = ~\u0_u0_state_reg[2]/NET0131  & n12361 ;
  assign n12363 = n5742 & n12362 ;
  assign n12364 = n12360 & n12363 ;
  assign n12365 = n5744 & n12364 ;
  assign n12366 = ~\u0_u0_state_reg[3]/P0001  & n12337 ;
  assign n12367 = \u0_u0_state_reg[14]/P0001  & \u0_u0_state_reg[9]/P0001  ;
  assign n12368 = ~\u0_u0_state_reg[14]/P0001  & ~\u0_u0_state_reg[9]/P0001  ;
  assign n12369 = ~n12367 & ~n12368 ;
  assign n12370 = n12361 & n12369 ;
  assign n12371 = n12366 & n12370 ;
  assign n12372 = n5744 & n12336 ;
  assign n12373 = n12371 & n12372 ;
  assign n12374 = ~n12365 & ~n12373 ;
  assign n12375 = n12357 & ~n12374 ;
  assign n12376 = ~n12356 & ~n12375 ;
  assign n12377 = ~n9110 & ~n9151 ;
  assign n12378 = n9146 & ~n12377 ;
  assign n12379 = ~n9146 & n12377 ;
  assign n12380 = ~n12378 & ~n12379 ;
  assign n12381 = ~n9159 & ~n9200 ;
  assign n12382 = n9195 & ~n12381 ;
  assign n12383 = ~n9195 & n12381 ;
  assign n12384 = ~n12382 & ~n12383 ;
  assign n12385 = \sram_data_i[22]_pad  & \wb_addr_i[17]_pad  ;
  assign n12386 = \u4_dout_reg[22]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n12387 = ~n12385 & ~n12386 ;
  assign n12388 = \sram_data_i[23]_pad  & \wb_addr_i[17]_pad  ;
  assign n12389 = \u4_dout_reg[23]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n12390 = ~n12388 & ~n12389 ;
  assign n12391 = \sram_data_i[4]_pad  & \wb_addr_i[17]_pad  ;
  assign n12392 = \u4_dout_reg[4]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n12393 = ~n12391 & ~n12392 ;
  assign n12394 = \sram_data_i[7]_pad  & \wb_addr_i[17]_pad  ;
  assign n12395 = \u4_dout_reg[7]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n12396 = ~n12394 & ~n12395 ;
  assign n12397 = \u1_u2_sizu_c_reg[0]/P0001  & \u1_u3_out_to_small_r_reg/P0001  ;
  assign n12398 = \u1_u3_new_size_reg[0]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n12399 = ~n12397 & ~n12398 ;
  assign n12400 = n9238 & n9241 ;
  assign n12401 = ~n9209 & ~n9210 ;
  assign n12402 = ~n9211 & ~n12401 ;
  assign n12403 = ~n12400 & n12402 ;
  assign n12404 = n9211 & n12401 ;
  assign n12405 = n9241 & n12401 ;
  assign n12406 = n9238 & n12405 ;
  assign n12407 = ~n12404 & ~n12406 ;
  assign n12408 = ~n12403 & n12407 ;
  assign n12409 = \u4_u3_buf0_orig_reg[19]/P0001  & \u4_u3_buf0_orig_reg[20]/P0001  ;
  assign n12410 = ~\u4_u3_buf0_orig_reg[21]/P0001  & ~\u4_u3_buf0_orig_reg[22]/P0001  ;
  assign n12411 = ~n12409 & n12410 ;
  assign n12412 = ~\u4_u3_buf0_orig_reg[23]/P0001  & ~\u4_u3_buf0_orig_reg[24]/P0001  ;
  assign n12413 = ~\u4_u3_buf0_orig_reg[25]/P0001  & ~\u4_u3_buf0_orig_reg[26]/P0001  ;
  assign n12414 = n12412 & n12413 ;
  assign n12415 = n12411 & n12414 ;
  assign n12416 = ~\u4_u3_buf0_orig_reg[27]/P0001  & ~\u4_u3_buf0_orig_reg[28]/P0001  ;
  assign n12417 = ~\u4_u3_buf0_orig_reg[29]/NET0131  & n12416 ;
  assign n12418 = \u4_u3_buf0_orig_reg[30]/NET0131  & n12417 ;
  assign n12419 = n12415 & n12418 ;
  assign n12420 = n12415 & n12417 ;
  assign n12421 = ~\u4_u3_buf0_orig_reg[30]/NET0131  & ~n12420 ;
  assign n12422 = ~n12419 & ~n12421 ;
  assign n12423 = ~n5704 & ~n5708 ;
  assign n12424 = ~n5705 & ~n12423 ;
  assign n12425 = n5705 & n12423 ;
  assign n12426 = ~n12424 & ~n12425 ;
  assign n12427 = n9091 & n9094 ;
  assign n12428 = ~n9062 & ~n9063 ;
  assign n12429 = ~n9064 & ~n12428 ;
  assign n12430 = ~n12427 & n12429 ;
  assign n12431 = n9064 & n12428 ;
  assign n12432 = n9094 & n12428 ;
  assign n12433 = n9091 & n12432 ;
  assign n12434 = ~n12431 & ~n12433 ;
  assign n12435 = ~n12430 & n12434 ;
  assign n12436 = ~\u4_u0_buf0_orig_reg[23]/P0001  & ~\u4_u0_buf0_orig_reg[24]/P0001  ;
  assign n12437 = ~\u4_u0_buf0_orig_reg[25]/P0001  & ~\u4_u0_buf0_orig_reg[26]/P0001  ;
  assign n12438 = n12436 & n12437 ;
  assign n12439 = \u4_u0_buf0_orig_reg[19]/P0001  & \u4_u0_buf0_orig_reg[20]/P0001  ;
  assign n12440 = ~\u4_u0_buf0_orig_reg[21]/P0001  & ~\u4_u0_buf0_orig_reg[22]/P0001  ;
  assign n12441 = ~n12439 & n12440 ;
  assign n12442 = ~\u4_u0_buf0_orig_reg[27]/P0001  & ~\u4_u0_buf0_orig_reg[29]/NET0131  ;
  assign n12443 = ~\u4_u0_buf0_orig_reg[28]/P0001  & n12442 ;
  assign n12444 = n12441 & n12443 ;
  assign n12445 = n12438 & n12444 ;
  assign n12446 = \u4_u0_buf0_orig_reg[30]/NET0131  & ~n12445 ;
  assign n12447 = ~\u4_u0_buf0_orig_reg[27]/P0001  & ~\u4_u0_buf0_orig_reg[28]/P0001  ;
  assign n12448 = ~\u4_u0_buf0_orig_reg[29]/NET0131  & ~\u4_u0_buf0_orig_reg[30]/NET0131  ;
  assign n12449 = n12447 & n12448 ;
  assign n12450 = n12438 & n12449 ;
  assign n12451 = n12441 & n12450 ;
  assign n12452 = ~n12446 & ~n12451 ;
  assign n12453 = n9140 & n9143 ;
  assign n12454 = ~n9111 & ~n9112 ;
  assign n12455 = ~n9113 & ~n12454 ;
  assign n12456 = ~n12453 & n12455 ;
  assign n12457 = n9113 & n12454 ;
  assign n12458 = n9143 & n12454 ;
  assign n12459 = n9140 & n12458 ;
  assign n12460 = ~n12457 & ~n12459 ;
  assign n12461 = ~n12456 & n12460 ;
  assign n12462 = \u4_u1_buf0_orig_reg[19]/P0001  & \u4_u1_buf0_orig_reg[20]/P0001  ;
  assign n12463 = ~\u4_u1_buf0_orig_reg[21]/P0001  & ~\u4_u1_buf0_orig_reg[22]/P0001  ;
  assign n12464 = ~n12462 & n12463 ;
  assign n12465 = ~\u4_u1_buf0_orig_reg[23]/P0001  & ~\u4_u1_buf0_orig_reg[24]/P0001  ;
  assign n12466 = ~\u4_u1_buf0_orig_reg[25]/P0001  & ~\u4_u1_buf0_orig_reg[26]/P0001  ;
  assign n12467 = n12465 & n12466 ;
  assign n12468 = n12464 & n12467 ;
  assign n12469 = ~\u4_u1_buf0_orig_reg[27]/P0001  & ~\u4_u1_buf0_orig_reg[28]/P0001  ;
  assign n12470 = ~\u4_u1_buf0_orig_reg[29]/NET0131  & n12469 ;
  assign n12471 = \u4_u1_buf0_orig_reg[30]/NET0131  & n12470 ;
  assign n12472 = n12468 & n12471 ;
  assign n12473 = n12468 & n12470 ;
  assign n12474 = ~\u4_u1_buf0_orig_reg[30]/NET0131  & ~n12473 ;
  assign n12475 = ~n12472 & ~n12474 ;
  assign n12476 = n9189 & n9192 ;
  assign n12477 = ~n9160 & ~n9161 ;
  assign n12478 = ~n9162 & ~n12477 ;
  assign n12479 = ~n12476 & n12478 ;
  assign n12480 = n9162 & n12477 ;
  assign n12481 = n9192 & n12477 ;
  assign n12482 = n9189 & n12481 ;
  assign n12483 = ~n12480 & ~n12482 ;
  assign n12484 = ~n12479 & n12483 ;
  assign n12485 = \u4_u2_buf0_orig_reg[19]/P0001  & \u4_u2_buf0_orig_reg[20]/P0001  ;
  assign n12486 = ~\u4_u2_buf0_orig_reg[21]/P0001  & ~\u4_u2_buf0_orig_reg[22]/P0001  ;
  assign n12487 = ~n12485 & n12486 ;
  assign n12488 = ~\u4_u2_buf0_orig_reg[23]/P0001  & ~\u4_u2_buf0_orig_reg[24]/P0001  ;
  assign n12489 = ~\u4_u2_buf0_orig_reg[25]/P0001  & ~\u4_u2_buf0_orig_reg[26]/P0001  ;
  assign n12490 = n12488 & n12489 ;
  assign n12491 = n12487 & n12490 ;
  assign n12492 = ~\u4_u2_buf0_orig_reg[27]/P0001  & ~\u4_u2_buf0_orig_reg[28]/P0001  ;
  assign n12493 = ~\u4_u2_buf0_orig_reg[29]/NET0131  & n12492 ;
  assign n12494 = \u4_u2_buf0_orig_reg[30]/NET0131  & n12493 ;
  assign n12495 = n12491 & n12494 ;
  assign n12496 = n12491 & n12493 ;
  assign n12497 = ~\u4_u2_buf0_orig_reg[30]/NET0131  & ~n12496 ;
  assign n12498 = ~n12495 & ~n12497 ;
  assign n12499 = \u1_u0_rxv2_reg/P0001  & ~n4936 ;
  assign n12500 = rst_i_pad & n12499 ;
  assign n12501 = ~\u0_rx_err_reg/P0001  & \u1_u0_rxv1_reg/P0001  ;
  assign n12502 = n7202 & n12501 ;
  assign n12503 = rst_i_pad & n12502 ;
  assign n12504 = ~n10520 & n12503 ;
  assign n12505 = ~n12500 & ~n12504 ;
  assign n12506 = \u1_u3_buffer_done_reg/P0001  & \u1_u3_state_reg[8]/P0001  ;
  assign n12507 = ~\u1_u3_buf0_not_aloc_reg/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n12508 = n12506 & n12507 ;
  assign n12509 = ~\u4_u2_int_stat_reg[3]/P0001  & ~n12508 ;
  assign n12510 = ~\u4_u2_int_stat_reg[3]/P0001  & ~n2793 ;
  assign n12511 = ~n2794 & n12510 ;
  assign n12512 = ~n12509 & ~n12511 ;
  assign n12513 = n5451 & n12512 ;
  assign n12514 = ~\u1_u3_buf0_not_aloc_reg/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n12515 = n12506 & n12514 ;
  assign n12516 = ~\u4_u3_int_stat_reg[3]/P0001  & ~n12515 ;
  assign n12517 = ~\u4_u3_int_stat_reg[3]/P0001  & ~n2793 ;
  assign n12518 = ~n2794 & n12517 ;
  assign n12519 = ~n12516 & ~n12518 ;
  assign n12520 = n5455 & n12519 ;
  assign n12521 = ~\u0_u0_state_reg[13]/NET0131  & \u0_u0_state_reg[9]/P0001  ;
  assign n12522 = ~n12342 & ~n12521 ;
  assign n12523 = n12343 & ~n12522 ;
  assign n12524 = n12341 & n12523 ;
  assign n12525 = n12340 & n12524 ;
  assign n12526 = XcvSelect_pad_o_pad & ~n12354 ;
  assign n12527 = ~n12525 & n12526 ;
  assign n12528 = ~\u0_u0_state_reg[13]/NET0131  & \u0_u0_state_reg[14]/P0001  ;
  assign n12529 = ~\u0_u0_state_reg[10]/P0001  & ~\u0_u0_state_reg[9]/P0001  ;
  assign n12530 = n5744 & n12529 ;
  assign n12531 = n12339 & n12530 ;
  assign n12532 = n12336 & n12531 ;
  assign n12533 = n12528 & n12532 ;
  assign n12534 = \u0_u0_state_reg[1]/P0001  & n6147 ;
  assign n12535 = ~n6157 & ~n12534 ;
  assign n12536 = ~n12533 & n12535 ;
  assign n12537 = ~n12527 & n12536 ;
  assign n12538 = susp_o_pad & ~\u4_suspend_r1_reg/P0001  ;
  assign n12539 = ~\u4_int_srcb_reg[3]/P0001  & ~n12538 ;
  assign n12540 = n5667 & ~n12539 ;
  assign n12541 = ~susp_o_pad & \u4_suspend_r1_reg/P0001  ;
  assign n12542 = ~\u4_int_srcb_reg[4]/P0001  & ~n12541 ;
  assign n12543 = n5667 & ~n12542 ;
  assign n12544 = ~\u0_u0_idle_cnt1_next_reg[0]/P0001  & n8674 ;
  assign n12545 = ~\u0_u0_idle_cnt1_reg[0]/P0001  & ~n8674 ;
  assign n12546 = n8673 & ~n12545 ;
  assign n12547 = ~n12544 & n12546 ;
  assign n12548 = ~n8672 & n12547 ;
  assign n12549 = ~n8666 & n12548 ;
  assign n12550 = ~\u0_u0_idle_cnt1_next_reg[1]/P0001  & n8674 ;
  assign n12551 = ~\u0_u0_idle_cnt1_reg[1]/P0001  & ~n8674 ;
  assign n12552 = n8673 & ~n12551 ;
  assign n12553 = ~n12550 & n12552 ;
  assign n12554 = ~n8672 & n12553 ;
  assign n12555 = ~n8666 & n12554 ;
  assign n12556 = ~\u0_u0_idle_cnt1_next_reg[2]/P0001  & n8674 ;
  assign n12557 = ~\u0_u0_idle_cnt1_reg[2]/P0001  & ~n8674 ;
  assign n12558 = n8673 & ~n12557 ;
  assign n12559 = ~n12556 & n12558 ;
  assign n12560 = ~n8672 & n12559 ;
  assign n12561 = ~n8666 & n12560 ;
  assign n12562 = ~\u0_u0_idle_cnt1_next_reg[5]/P0001  & n8674 ;
  assign n12563 = ~\u0_u0_idle_cnt1_reg[5]/P0001  & ~n8674 ;
  assign n12564 = n8673 & ~n12563 ;
  assign n12565 = ~n12562 & n12564 ;
  assign n12566 = ~n8672 & n12565 ;
  assign n12567 = ~n8666 & n12566 ;
  assign n12568 = ~\u0_u0_idle_cnt1_next_reg[6]/P0001  & n8674 ;
  assign n12569 = ~\u0_u0_idle_cnt1_reg[6]/P0001  & ~n8674 ;
  assign n12570 = n8673 & ~n12569 ;
  assign n12571 = ~n12568 & n12570 ;
  assign n12572 = ~n8672 & n12571 ;
  assign n12573 = ~n8666 & n12572 ;
  assign n12574 = ~\u0_u0_idle_cnt1_reg[0]/P0001  & ~\u0_u0_idle_cnt1_reg[1]/P0001  ;
  assign n12575 = ~\u0_u0_idle_cnt1_reg[2]/P0001  & ~\u0_u0_idle_cnt1_reg[3]/P0001  ;
  assign n12576 = n12574 & n12575 ;
  assign n12577 = \u0_u0_idle_cnt1_reg[4]/P0001  & \u0_u0_idle_cnt1_reg[6]/P0001  ;
  assign n12578 = ~n12576 & n12577 ;
  assign n12579 = \u0_u0_idle_cnt1_reg[5]/P0001  & \u0_u0_idle_cnt1_reg[6]/P0001  ;
  assign n12580 = ~\u0_u0_idle_cnt1_reg[7]/P0001  & ~n12579 ;
  assign n12581 = ~n12578 & n12580 ;
  assign n12582 = ~n8672 & ~n12581 ;
  assign n12583 = ~n8666 & n12582 ;
  assign n12584 = ~\u1_u3_buf0_not_aloc_reg/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n12585 = n12506 & n12584 ;
  assign n12586 = ~\u4_u0_int_stat_reg[3]/P0001  & ~n12585 ;
  assign n12587 = ~\u4_u0_int_stat_reg[3]/P0001  & ~n2793 ;
  assign n12588 = ~n2794 & n12587 ;
  assign n12589 = ~n12586 & ~n12588 ;
  assign n12590 = n5459 & n12589 ;
  assign n12591 = ~n2358 & ~n12290 ;
  assign n12592 = n12297 & n12591 ;
  assign n12593 = n12305 & n12308 ;
  assign n12594 = n12592 & n12593 ;
  assign n12595 = \u4_csr_reg[24]/P0001  & ~\u4_csr_reg[27]/NET0131  ;
  assign n12596 = ~\u4_csr_reg[25]/P0001  & \u4_csr_reg[28]/P0001  ;
  assign n12597 = n12595 & n12596 ;
  assign n12598 = n12304 & n12597 ;
  assign n12599 = ~n12592 & n12598 ;
  assign n12600 = n12295 & n12599 ;
  assign n12601 = ~\u1_u3_setup_token_reg/P0001  & \u4_csr_reg[29]/P0001  ;
  assign n12602 = n3036 & n12601 ;
  assign n12603 = n12299 & ~n12602 ;
  assign n12604 = ~n12600 & ~n12603 ;
  assign n12605 = ~n12594 & n12604 ;
  assign n12606 = \u0_u0_idle_long_reg/P0001  & ~\u0_u0_ps_cnt_clr_reg/P0001  ;
  assign n12607 = ~\u0_u0_ps_cnt_reg[0]/P0001  & n12606 ;
  assign n12608 = ~n8672 & n12607 ;
  assign n12609 = ~n8666 & n12608 ;
  assign n12610 = \u0_u0_ps_cnt_reg[0]/P0001  & ~\u0_u0_ps_cnt_reg[1]/P0001  ;
  assign n12611 = ~\u0_u0_ps_cnt_reg[0]/P0001  & \u0_u0_ps_cnt_reg[1]/P0001  ;
  assign n12612 = ~n12610 & ~n12611 ;
  assign n12613 = n12606 & ~n12612 ;
  assign n12614 = ~n8672 & n12613 ;
  assign n12615 = ~n8666 & n12614 ;
  assign n12616 = \u0_u0_ps_cnt_reg[0]/P0001  & \u0_u0_ps_cnt_reg[1]/P0001  ;
  assign n12617 = ~\u0_u0_ps_cnt_reg[2]/P0001  & ~n12616 ;
  assign n12618 = \u0_u0_ps_cnt_reg[2]/P0001  & n12616 ;
  assign n12619 = ~n12617 & ~n12618 ;
  assign n12620 = n12606 & n12619 ;
  assign n12621 = ~n8672 & n12620 ;
  assign n12622 = ~n8666 & n12621 ;
  assign n12623 = ~\u0_u0_ps_cnt_reg[3]/P0001  & ~n12618 ;
  assign n12624 = \u0_u0_ps_cnt_reg[2]/P0001  & \u0_u0_ps_cnt_reg[3]/P0001  ;
  assign n12625 = n12616 & n12624 ;
  assign n12626 = n12606 & ~n12625 ;
  assign n12627 = ~n12623 & n12626 ;
  assign n12628 = ~n8672 & n12627 ;
  assign n12629 = ~n8666 & n12628 ;
  assign n12630 = \u1_u3_rx_ack_to_cnt_reg[0]/P0001  & \u1_u3_rx_ack_to_cnt_reg[1]/P0001  ;
  assign n12631 = \u1_u3_rx_ack_to_cnt_reg[2]/P0001  & \u1_u3_rx_ack_to_cnt_reg[3]/P0001  ;
  assign n12632 = n12630 & n12631 ;
  assign n12633 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & \u1_u3_rx_ack_to_cnt_reg[4]/P0001  ;
  assign n12634 = ~n12632 & n12633 ;
  assign n12635 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & ~\u1_u3_rx_ack_to_cnt_reg[4]/P0001  ;
  assign n12636 = n12632 & n12635 ;
  assign n12637 = ~n12634 & ~n12636 ;
  assign n12638 = n6133 & ~n6150 ;
  assign n12639 = ~\u0_u0_T1_gt_3_0_mS_reg/P0001  & \u0_u0_state_reg[1]/P0001  ;
  assign n12640 = n12638 & n12639 ;
  assign n12641 = n6132 & n12640 ;
  assign n12642 = ~\u0_u0_state_reg[0]/NET0131  & ~\u0_u0_state_reg[8]/NET0131  ;
  assign n12643 = n5753 & n12642 ;
  assign n12644 = n5746 & n12643 ;
  assign n12645 = \u0_u0_state_reg[13]/NET0131  & ~\u0_u0_state_reg[14]/P0001  ;
  assign n12646 = ~n12528 & ~n12645 ;
  assign n12647 = ~\u0_u0_state_reg[9]/P0001  & ~n12646 ;
  assign n12648 = \u0_u0_state_reg[13]/NET0131  & ~\u0_u0_state_reg[1]/P0001  ;
  assign n12649 = ~n5766 & n12648 ;
  assign n12650 = n12647 & ~n12649 ;
  assign n12651 = n12644 & n12650 ;
  assign n12652 = ~n12641 & ~n12651 ;
  assign n12653 = n6130 & n6172 ;
  assign n12654 = ~\u0_u0_T2_gt_100_uS_reg/P0001  & ~\u0_u0_state_reg[1]/P0001  ;
  assign n12655 = ~\u0_u0_state_reg[3]/P0001  & \u0_u0_state_reg[6]/NET0131  ;
  assign n12656 = ~n12654 & n12655 ;
  assign n12657 = n12653 & n12656 ;
  assign n12658 = ~\u0_u0_me_cnt_100_ms_reg/P0001  & ~\u0_u0_state_reg[1]/P0001  ;
  assign n12659 = n8663 & ~n12658 ;
  assign n12660 = ~n12657 & ~n12659 ;
  assign n12661 = n12652 & n12660 ;
  assign n12662 = n5748 & ~n12661 ;
  assign n12663 = \u1_u3_tx_data_to_cnt_reg[0]/P0001  & \u1_u3_tx_data_to_cnt_reg[1]/P0001  ;
  assign n12664 = \u1_u3_tx_data_to_cnt_reg[2]/P0001  & \u1_u3_tx_data_to_cnt_reg[3]/P0001  ;
  assign n12665 = n12663 & n12664 ;
  assign n12666 = ~\u0_rx_active_reg/P0001  & \u1_u3_tx_data_to_cnt_reg[4]/P0001  ;
  assign n12667 = ~n12665 & n12666 ;
  assign n12668 = ~\u0_rx_active_reg/P0001  & ~\u1_u3_tx_data_to_cnt_reg[4]/P0001  ;
  assign n12669 = n12665 & n12668 ;
  assign n12670 = ~n12667 & ~n12669 ;
  assign n12671 = ~\u1_u3_buf0_not_aloc_reg/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n12672 = n12506 & n12671 ;
  assign n12673 = ~\u4_u1_int_stat_reg[3]/P0001  & ~n12672 ;
  assign n12674 = ~\u4_u1_int_stat_reg[3]/P0001  & ~n2793 ;
  assign n12675 = ~n2794 & n12674 ;
  assign n12676 = ~n12673 & ~n12675 ;
  assign n12677 = n5463 & n12676 ;
  assign n12678 = \u1_u0_crc16_sum_reg[8]/P0001  & ~\u1_u0_crc16_sum_reg[9]/P0001  ;
  assign n12679 = ~n10485 & n12678 ;
  assign n12680 = n4929 & ~n10483 ;
  assign n12681 = ~n10484 & n12680 ;
  assign n12682 = ~n12679 & ~n12681 ;
  assign n12683 = ~\u1_u0_crc16_sum_reg[8]/P0001  & \u1_u0_crc16_sum_reg[9]/P0001  ;
  assign n12684 = ~n10485 & n12683 ;
  assign n12685 = \u1_u0_crc16_sum_reg[8]/P0001  & \u1_u0_crc16_sum_reg[9]/P0001  ;
  assign n12686 = n10485 & n12685 ;
  assign n12687 = ~n12684 & ~n12686 ;
  assign n12688 = n12682 & n12687 ;
  assign n12689 = ~n10593 & ~n10608 ;
  assign n12690 = ~n12688 & n12689 ;
  assign n12691 = n10593 & ~n10608 ;
  assign n12692 = n12688 & n12691 ;
  assign n12693 = ~n12690 & ~n12692 ;
  assign n12694 = n10593 & n10608 ;
  assign n12695 = ~n12688 & n12694 ;
  assign n12696 = ~n10593 & n10608 ;
  assign n12697 = n12688 & n12696 ;
  assign n12698 = ~n12695 & ~n12697 ;
  assign n12699 = n12693 & n12698 ;
  assign n12700 = n10521 & n10542 ;
  assign n12701 = ~n12699 & n12700 ;
  assign n12702 = n10521 & ~n10542 ;
  assign n12703 = n12699 & n12702 ;
  assign n12704 = ~n12701 & ~n12703 ;
  assign n12705 = \u1_u0_crc16_sum_reg[0]/P0001  & ~n4911 ;
  assign n12706 = ~n10519 & n12705 ;
  assign n12707 = \u1_u0_crc16_sum_reg[0]/P0001  & ~n7203 ;
  assign n12708 = ~n10553 & ~n12707 ;
  assign n12709 = ~n12706 & n12708 ;
  assign n12710 = n12704 & n12709 ;
  assign n12711 = \u1_u0_crc16_sum_reg[10]/P0001  & ~n7203 ;
  assign n12712 = \u1_u0_crc16_sum_reg[10]/P0001  & ~n4911 ;
  assign n12713 = ~n10519 & n12712 ;
  assign n12714 = ~n12711 & ~n12713 ;
  assign n12715 = \u1_u0_crc16_sum_reg[2]/P0001  & n7203 ;
  assign n12716 = ~n10520 & n12715 ;
  assign n12717 = ~n10553 & ~n12716 ;
  assign n12718 = n12714 & n12717 ;
  assign n12719 = \u1_u0_crc16_sum_reg[11]/P0001  & ~n7203 ;
  assign n12720 = \u1_u0_crc16_sum_reg[11]/P0001  & ~n4911 ;
  assign n12721 = ~n10519 & n12720 ;
  assign n12722 = ~n12719 & ~n12721 ;
  assign n12723 = \u1_u0_crc16_sum_reg[3]/P0001  & n7203 ;
  assign n12724 = ~n10520 & n12723 ;
  assign n12725 = ~n10553 & ~n12724 ;
  assign n12726 = n12722 & n12725 ;
  assign n12727 = \u1_u0_crc16_sum_reg[12]/P0001  & ~n7203 ;
  assign n12728 = \u1_u0_crc16_sum_reg[12]/P0001  & ~n4911 ;
  assign n12729 = ~n10519 & n12728 ;
  assign n12730 = ~n12727 & ~n12729 ;
  assign n12731 = \u1_u0_crc16_sum_reg[4]/P0001  & n7203 ;
  assign n12732 = ~n10520 & n12731 ;
  assign n12733 = ~n10553 & ~n12732 ;
  assign n12734 = n12730 & n12733 ;
  assign n12735 = \u1_u0_crc16_sum_reg[13]/P0001  & ~n7203 ;
  assign n12736 = \u1_u0_crc16_sum_reg[13]/P0001  & ~n4911 ;
  assign n12737 = ~n10519 & n12736 ;
  assign n12738 = ~n12735 & ~n12737 ;
  assign n12739 = \u1_u0_crc16_sum_reg[5]/P0001  & n7203 ;
  assign n12740 = ~n10520 & n12739 ;
  assign n12741 = ~n10553 & ~n12740 ;
  assign n12742 = n12738 & n12741 ;
  assign n12743 = \u1_u0_crc16_sum_reg[14]/P0001  & ~n7203 ;
  assign n12744 = \u1_u0_crc16_sum_reg[14]/P0001  & ~n4911 ;
  assign n12745 = ~n10519 & n12744 ;
  assign n12746 = ~n12743 & ~n12745 ;
  assign n12747 = \u1_u0_crc16_sum_reg[6]/P0001  & n7203 ;
  assign n12748 = ~n10520 & n12747 ;
  assign n12749 = ~n10553 & ~n12748 ;
  assign n12750 = n12746 & n12749 ;
  assign n12751 = n10521 & n12688 ;
  assign n12752 = \u1_u0_crc16_sum_reg[2]/P0001  & ~n4911 ;
  assign n12753 = ~n10519 & n12752 ;
  assign n12754 = \u1_u0_crc16_sum_reg[2]/P0001  & ~n7203 ;
  assign n12755 = ~n10553 & ~n12754 ;
  assign n12756 = ~n12753 & n12755 ;
  assign n12757 = ~n12751 & n12756 ;
  assign n12758 = \u1_u0_crc16_sum_reg[3]/P0001  & ~n7203 ;
  assign n12759 = \u1_u0_crc16_sum_reg[3]/P0001  & ~n4911 ;
  assign n12760 = ~n10519 & n12759 ;
  assign n12761 = ~n12758 & ~n12760 ;
  assign n12762 = \u0_rx_data_reg[5]/P0001  & ~\u0_rx_data_reg[6]/P0001  ;
  assign n12763 = ~\u0_rx_data_reg[5]/P0001  & \u0_rx_data_reg[6]/P0001  ;
  assign n12764 = ~n12762 & ~n12763 ;
  assign n12765 = ~n10527 & ~n12764 ;
  assign n12766 = n10527 & n12764 ;
  assign n12767 = ~n12765 & ~n12766 ;
  assign n12768 = n7203 & n12767 ;
  assign n12769 = ~n10520 & n12768 ;
  assign n12770 = ~n10553 & ~n12769 ;
  assign n12771 = n12761 & n12770 ;
  assign n12772 = n7203 & ~n10596 ;
  assign n12773 = ~n10520 & n12772 ;
  assign n12774 = \u1_u0_crc16_sum_reg[4]/P0001  & ~n4911 ;
  assign n12775 = ~n10519 & n12774 ;
  assign n12776 = \u1_u0_crc16_sum_reg[4]/P0001  & ~n7203 ;
  assign n12777 = ~n10553 & ~n12776 ;
  assign n12778 = ~n12775 & n12777 ;
  assign n12779 = ~n12773 & n12778 ;
  assign n12780 = \u0_rx_data_reg[3]/P0001  & ~\u0_rx_data_reg[4]/P0001  ;
  assign n12781 = ~n10524 & n12780 ;
  assign n12782 = ~\u0_rx_data_reg[3]/P0001  & ~\u0_rx_data_reg[4]/P0001  ;
  assign n12783 = n10524 & n12782 ;
  assign n12784 = ~n12781 & ~n12783 ;
  assign n12785 = ~\u0_rx_data_reg[3]/P0001  & \u0_rx_data_reg[4]/P0001  ;
  assign n12786 = ~n10524 & n12785 ;
  assign n12787 = \u0_rx_data_reg[3]/P0001  & \u0_rx_data_reg[4]/P0001  ;
  assign n12788 = n10524 & n12787 ;
  assign n12789 = ~n12786 & ~n12788 ;
  assign n12790 = n12784 & n12789 ;
  assign n12791 = n7203 & n12790 ;
  assign n12792 = ~n10520 & n12791 ;
  assign n12793 = \u1_u0_crc16_sum_reg[5]/P0001  & ~n7203 ;
  assign n12794 = \u1_u0_crc16_sum_reg[5]/P0001  & ~n4911 ;
  assign n12795 = ~n10519 & n12794 ;
  assign n12796 = ~n12793 & ~n12795 ;
  assign n12797 = ~n10553 & n12796 ;
  assign n12798 = ~n12792 & n12797 ;
  assign n12799 = \u1_u0_crc16_sum_reg[6]/P0001  & ~n7203 ;
  assign n12800 = \u1_u0_crc16_sum_reg[6]/P0001  & ~n4911 ;
  assign n12801 = ~n10519 & n12800 ;
  assign n12802 = ~n12799 & ~n12801 ;
  assign n12803 = ~n10491 & ~n10562 ;
  assign n12804 = n10491 & n10562 ;
  assign n12805 = ~n12803 & ~n12804 ;
  assign n12806 = n7203 & ~n12805 ;
  assign n12807 = ~n10520 & n12806 ;
  assign n12808 = ~n10553 & ~n12807 ;
  assign n12809 = n12802 & n12808 ;
  assign n12810 = \u1_u0_crc16_sum_reg[7]/P0001  & ~n7203 ;
  assign n12811 = \u1_u0_crc16_sum_reg[7]/P0001  & ~n4911 ;
  assign n12812 = ~n10519 & n12811 ;
  assign n12813 = ~n12810 & ~n12812 ;
  assign n12814 = \u0_rx_data_reg[1]/P0001  & ~\u0_rx_data_reg[2]/P0001  ;
  assign n12815 = ~\u0_rx_data_reg[1]/P0001  & \u0_rx_data_reg[2]/P0001  ;
  assign n12816 = ~n12814 & ~n12815 ;
  assign n12817 = ~n10530 & ~n12816 ;
  assign n12818 = n10530 & n12816 ;
  assign n12819 = ~n12817 & ~n12818 ;
  assign n12820 = n7203 & n12819 ;
  assign n12821 = ~n10520 & n12820 ;
  assign n12822 = ~n10553 & ~n12821 ;
  assign n12823 = n12813 & n12822 ;
  assign n12824 = ~\u1_u0_crc16_sum_reg[0]/P0001  & n10494 ;
  assign n12825 = \u1_u0_crc16_sum_reg[0]/P0001  & ~n10494 ;
  assign n12826 = ~n12824 & ~n12825 ;
  assign n12827 = ~n10564 & ~n12826 ;
  assign n12828 = n10564 & n12826 ;
  assign n12829 = ~n12827 & ~n12828 ;
  assign n12830 = n10521 & ~n12829 ;
  assign n12831 = \u1_u0_crc16_sum_reg[8]/P0001  & ~n4911 ;
  assign n12832 = ~n10519 & n12831 ;
  assign n12833 = \u1_u0_crc16_sum_reg[8]/P0001  & ~n7203 ;
  assign n12834 = ~n10553 & ~n12833 ;
  assign n12835 = ~n12832 & n12834 ;
  assign n12836 = ~n12830 & n12835 ;
  assign n12837 = \u1_u0_crc16_sum_reg[9]/P0001  & ~n7203 ;
  assign n12838 = \u1_u0_crc16_sum_reg[9]/P0001  & ~n4911 ;
  assign n12839 = ~n10519 & n12838 ;
  assign n12840 = ~n12837 & ~n12839 ;
  assign n12841 = ~\u0_rx_data_reg[0]/P0001  & ~\u1_u0_crc16_sum_reg[15]/P0001  ;
  assign n12842 = \u0_rx_data_reg[0]/P0001  & \u1_u0_crc16_sum_reg[15]/P0001  ;
  assign n12843 = ~n12841 & ~n12842 ;
  assign n12844 = ~\u1_u0_crc16_sum_reg[1]/P0001  & ~n12843 ;
  assign n12845 = \u1_u0_crc16_sum_reg[1]/P0001  & n12843 ;
  assign n12846 = ~n12844 & ~n12845 ;
  assign n12847 = n7203 & n12846 ;
  assign n12848 = ~n10520 & n12847 ;
  assign n12849 = ~n10553 & ~n12848 ;
  assign n12850 = n12840 & n12849 ;
  assign n12851 = ~\u4_buf0_reg[27]/P0001  & \u4_csr_reg[10]/P0001  ;
  assign n12852 = ~\u4_buf0_reg[26]/NET0131  & \u4_csr_reg[9]/NET0131  ;
  assign n12853 = ~n12851 & ~n12852 ;
  assign n12854 = ~\u4_buf0_reg[28]/P0001  & ~\u4_buf0_reg[29]/P0001  ;
  assign n12855 = \u4_buf0_reg[27]/P0001  & ~\u4_csr_reg[10]/P0001  ;
  assign n12856 = ~\u4_buf0_reg[30]/P0001  & ~n12855 ;
  assign n12857 = n12854 & n12856 ;
  assign n12858 = ~n12853 & n12857 ;
  assign n12859 = ~\u4_buf0_reg[25]/NET0131  & \u4_csr_reg[8]/P0001  ;
  assign n12860 = ~\u4_buf0_reg[24]/NET0131  & \u4_csr_reg[7]/P0001  ;
  assign n12861 = ~n12859 & ~n12860 ;
  assign n12862 = \u4_buf0_reg[23]/NET0131  & ~\u4_csr_reg[6]/NET0131  ;
  assign n12863 = \u4_buf0_reg[24]/NET0131  & ~\u4_csr_reg[7]/P0001  ;
  assign n12864 = ~n12862 & ~n12863 ;
  assign n12865 = n12861 & ~n12864 ;
  assign n12866 = \u4_buf0_reg[22]/NET0131  & ~\u4_csr_reg[5]/NET0131  ;
  assign n12867 = \u4_buf0_reg[21]/NET0131  & ~\u4_csr_reg[4]/NET0131  ;
  assign n12868 = ~n12866 & ~n12867 ;
  assign n12869 = ~\u4_buf0_reg[21]/NET0131  & \u4_csr_reg[4]/NET0131  ;
  assign n12870 = ~\u4_buf0_reg[20]/NET0131  & \u4_csr_reg[3]/P0001  ;
  assign n12871 = ~n12869 & ~n12870 ;
  assign n12872 = n12868 & ~n12871 ;
  assign n12873 = \u4_buf0_reg[18]/P0001  & ~\u4_csr_reg[1]/P0001  ;
  assign n12874 = ~\u4_buf0_reg[17]/NET0131  & \u4_csr_reg[0]/P0001  ;
  assign n12875 = ~n12873 & n12874 ;
  assign n12876 = ~\u4_buf0_reg[18]/P0001  & \u4_csr_reg[1]/P0001  ;
  assign n12877 = ~\u4_buf0_reg[19]/NET0131  & \u4_csr_reg[2]/NET0131  ;
  assign n12878 = ~n12876 & ~n12877 ;
  assign n12879 = ~n12875 & n12878 ;
  assign n12880 = \u4_buf0_reg[20]/NET0131  & ~\u4_csr_reg[3]/P0001  ;
  assign n12881 = \u4_buf0_reg[19]/NET0131  & ~\u4_csr_reg[2]/NET0131  ;
  assign n12882 = ~n12880 & ~n12881 ;
  assign n12883 = n12868 & n12882 ;
  assign n12884 = ~n12879 & n12883 ;
  assign n12885 = ~n12872 & ~n12884 ;
  assign n12886 = ~\u4_buf0_reg[23]/NET0131  & \u4_csr_reg[6]/NET0131  ;
  assign n12887 = ~\u4_buf0_reg[22]/NET0131  & \u4_csr_reg[5]/NET0131  ;
  assign n12888 = ~n12886 & ~n12887 ;
  assign n12889 = n12861 & n12888 ;
  assign n12890 = n12885 & n12889 ;
  assign n12891 = ~n12865 & ~n12890 ;
  assign n12892 = \u4_buf0_reg[25]/NET0131  & ~\u4_csr_reg[8]/P0001  ;
  assign n12893 = \u4_buf0_reg[26]/NET0131  & ~\u4_csr_reg[9]/NET0131  ;
  assign n12894 = ~n12892 & ~n12893 ;
  assign n12895 = n12857 & n12894 ;
  assign n12896 = n12891 & n12895 ;
  assign n12897 = ~n12858 & ~n12896 ;
  assign n12898 = \u4_u2_int_stat_reg[4]/P0001  & n5451 ;
  assign n12899 = ~\u1_u3_buf1_not_aloc_reg/P0001  & n12506 ;
  assign n12900 = ~n2793 & n12899 ;
  assign n12901 = ~n2794 & n12900 ;
  assign n12902 = n11311 & n12901 ;
  assign n12903 = ~n12898 & ~n12902 ;
  assign n12904 = ~\u4_u3_csr0_reg[5]/P0001  & ~\u4_u3_csr0_reg[6]/P0001  ;
  assign n12905 = ~\u4_u3_csr0_reg[3]/NET0131  & ~\u4_u3_csr0_reg[4]/P0001  ;
  assign n12906 = n12904 & n12905 ;
  assign n12907 = ~\u4_u3_csr0_reg[1]/P0001  & ~\u4_u3_csr0_reg[2]/P0001  ;
  assign n12908 = ~\u4_u3_csr0_reg[0]/P0001  & ~\u4_u3_csr0_reg[10]/P0001  ;
  assign n12909 = n12907 & n12908 ;
  assign n12910 = n12906 & n12909 ;
  assign n12911 = ~\u4_u3_csr0_reg[7]/P0001  & ~\u4_u3_csr0_reg[8]/P0001  ;
  assign n12912 = ~\u4_u3_csr0_reg[9]/P0001  & n12911 ;
  assign n12913 = n12910 & n12912 ;
  assign n12914 = n6268 & ~n6594 ;
  assign n12915 = ~n6593 & n12914 ;
  assign n12916 = ~\u4_u3_dma_in_cnt_reg[11]/P0001  & ~n6283 ;
  assign n12917 = n7222 & n12916 ;
  assign n12918 = ~n12915 & n12917 ;
  assign n12919 = ~n12913 & ~n12918 ;
  assign n12920 = \u4_u3_int_stat_reg[4]/P0001  & n5455 ;
  assign n12921 = n11568 & n12901 ;
  assign n12922 = ~n12920 & ~n12921 ;
  assign n12923 = ~\u4_u0_csr0_reg[5]/P0001  & ~\u4_u0_csr0_reg[6]/P0001  ;
  assign n12924 = ~\u4_u0_csr0_reg[3]/NET0131  & ~\u4_u0_csr0_reg[4]/P0001  ;
  assign n12925 = n12923 & n12924 ;
  assign n12926 = ~\u4_u0_csr0_reg[1]/P0001  & ~\u4_u0_csr0_reg[2]/P0001  ;
  assign n12927 = ~\u4_u0_csr0_reg[0]/P0001  & ~\u4_u0_csr0_reg[10]/P0001  ;
  assign n12928 = n12926 & n12927 ;
  assign n12929 = n12925 & n12928 ;
  assign n12930 = ~\u4_u0_csr0_reg[7]/P0001  & ~\u4_u0_csr0_reg[8]/P0001  ;
  assign n12931 = ~\u4_u0_csr0_reg[9]/P0001  & n12930 ;
  assign n12932 = n12929 & n12931 ;
  assign n12933 = n6326 & ~n6628 ;
  assign n12934 = ~n6627 & n12933 ;
  assign n12935 = ~\u4_u0_dma_in_cnt_reg[11]/P0001  & ~n6340 ;
  assign n12936 = n7243 & n12935 ;
  assign n12937 = ~n12934 & n12936 ;
  assign n12938 = ~n12932 & ~n12937 ;
  assign n12939 = \u4_u0_int_stat_reg[4]/P0001  & n5459 ;
  assign n12940 = n11816 & n12901 ;
  assign n12941 = ~n12939 & ~n12940 ;
  assign n12942 = ~\u4_u1_csr0_reg[5]/P0001  & ~\u4_u1_csr0_reg[6]/P0001  ;
  assign n12943 = ~\u4_u1_csr0_reg[3]/NET0131  & ~\u4_u1_csr0_reg[4]/P0001  ;
  assign n12944 = n12942 & n12943 ;
  assign n12945 = ~\u4_u1_csr0_reg[1]/P0001  & ~\u4_u1_csr0_reg[2]/P0001  ;
  assign n12946 = ~\u4_u1_csr0_reg[0]/P0001  & ~\u4_u1_csr0_reg[10]/P0001  ;
  assign n12947 = n12945 & n12946 ;
  assign n12948 = n12944 & n12947 ;
  assign n12949 = ~\u4_u1_csr0_reg[7]/P0001  & ~\u4_u1_csr0_reg[8]/P0001  ;
  assign n12950 = ~\u4_u1_csr0_reg[9]/P0001  & n12949 ;
  assign n12951 = n12948 & n12950 ;
  assign n12952 = n7275 & n7565 ;
  assign n12953 = ~n6404 & n12952 ;
  assign n12954 = n6656 & n12952 ;
  assign n12955 = ~n6655 & n12954 ;
  assign n12956 = ~n12953 & ~n12955 ;
  assign n12957 = ~n12951 & n12956 ;
  assign n12958 = \u4_u1_int_stat_reg[4]/P0001  & n5463 ;
  assign n12959 = n12050 & n12901 ;
  assign n12960 = ~n12958 & ~n12959 ;
  assign n12961 = \u0_u0_T1_gt_5_0_mS_reg/P0001  & \u0_u0_resume_req_s_reg/P0001  ;
  assign n12962 = \u0_u0_state_reg[9]/P0001  & ~n12961 ;
  assign n12963 = ~n5768 & n12962 ;
  assign n12964 = ~n6192 & ~n12963 ;
  assign n12965 = n12653 & ~n12964 ;
  assign n12966 = \u0_u0_state_reg[3]/P0001  & ~\u0_u0_state_reg[6]/NET0131  ;
  assign n12967 = n12965 & n12966 ;
  assign n12968 = ~\u0_u0_T1_gt_3_0_mS_reg/P0001  & \u0_u0_state_reg[9]/P0001  ;
  assign n12969 = ~n6150 & ~n12968 ;
  assign n12970 = n6133 & ~n12969 ;
  assign n12971 = n6132 & n12970 ;
  assign n12972 = ~\u0_u0_T2_gt_1_0_mS_reg/P0001  & n5746 ;
  assign n12973 = n5938 & n12972 ;
  assign n12974 = ~n12971 & ~n12973 ;
  assign n12975 = ~n12967 & n12974 ;
  assign n12976 = ~n6200 & n12975 ;
  assign n12977 = n5748 & ~n12976 ;
  assign n12978 = ~\u4_u2_dma_in_cnt_reg[11]/P0001  & ~n6419 ;
  assign n12979 = ~n6422 & n7284 ;
  assign n12980 = n12978 & n12979 ;
  assign n12981 = ~\u4_u2_csr0_reg[5]/P0001  & ~\u4_u2_csr0_reg[6]/P0001  ;
  assign n12982 = ~\u4_u2_csr0_reg[3]/NET0131  & ~\u4_u2_csr0_reg[4]/P0001  ;
  assign n12983 = n12981 & n12982 ;
  assign n12984 = ~\u4_u2_csr0_reg[1]/P0001  & ~\u4_u2_csr0_reg[2]/P0001  ;
  assign n12985 = ~\u4_u2_csr0_reg[0]/P0001  & ~\u4_u2_csr0_reg[10]/P0001  ;
  assign n12986 = n12984 & n12985 ;
  assign n12987 = n12983 & n12986 ;
  assign n12988 = ~\u4_u2_csr0_reg[7]/P0001  & ~\u4_u2_csr0_reg[8]/P0001  ;
  assign n12989 = ~\u4_u2_csr0_reg[9]/P0001  & n12988 ;
  assign n12990 = n12987 & n12989 ;
  assign n12991 = n6668 & n7284 ;
  assign n12992 = n12978 & n12991 ;
  assign n12993 = ~n12990 & ~n12992 ;
  assign n12994 = ~n12980 & n12993 ;
  assign n12995 = n6452 & n12993 ;
  assign n12996 = n6449 & n12995 ;
  assign n12997 = ~n12994 & ~n12996 ;
  assign n12998 = \u0_u0_state_reg[4]/NET0131  & n5765 ;
  assign n12999 = \OpMode_pad_o[1]_pad  & ~n12998 ;
  assign n13000 = \u0_u0_T2_wakeup_reg/P0001  & \u0_u0_state_reg[5]/P0001  ;
  assign n13001 = ~n12999 & ~n13000 ;
  assign n13002 = ~n12646 & ~n13000 ;
  assign n13003 = n12532 & n13002 ;
  assign n13004 = ~n13001 & ~n13003 ;
  assign n13005 = ~n5939 & ~n13004 ;
  assign n13006 = n12304 & n12596 ;
  assign n13007 = ~\u4_csr_reg[24]/P0001  & \u4_csr_reg[28]/P0001  ;
  assign n13008 = ~n13006 & ~n13007 ;
  assign n13009 = ~\u4_csr_reg[28]/P0001  & n12291 ;
  assign n13010 = n5555 & ~n12289 ;
  assign n13011 = n13009 & n13010 ;
  assign n13012 = \u4_csr_reg[26]/NET0131  & ~n13011 ;
  assign n13013 = n13008 & n13012 ;
  assign n13014 = ~\u4_csr_reg[26]/NET0131  & ~n12300 ;
  assign n13015 = \u1_u3_in_token_reg/NET0131  & ~\u4_csr_reg[26]/NET0131  ;
  assign n13016 = ~\u4_csr_reg[27]/NET0131  & n13015 ;
  assign n13017 = ~n13014 & ~n13016 ;
  assign n13018 = ~n12602 & ~n13017 ;
  assign n13019 = ~\u4_csr_reg[27]/NET0131  & ~n13018 ;
  assign n13020 = ~n13013 & n13019 ;
  assign n13021 = ~\u4_csr_reg[29]/P0001  & n12291 ;
  assign n13022 = n12289 & ~n13007 ;
  assign n13023 = ~n13021 & n13022 ;
  assign n13024 = ~n12289 & n12292 ;
  assign n13025 = ~n12291 & n13024 ;
  assign n13026 = ~n5555 & ~n13007 ;
  assign n13027 = n2363 & ~n13026 ;
  assign n13028 = ~n13025 & n13027 ;
  assign n13029 = ~n13023 & n13028 ;
  assign n13030 = ~\u1_u0_pid_reg[3]/NET0131  & n7806 ;
  assign n13031 = n13025 & ~n13030 ;
  assign n13032 = ~n13029 & ~n13031 ;
  assign n13033 = ~n13020 & n13032 ;
  assign n13034 = \u0_u0_idle_cnt1_reg[4]/P0001  & \u0_u0_idle_cnt1_reg[5]/P0001  ;
  assign n13035 = ~n12576 & n13034 ;
  assign n13036 = n11231 & ~n13035 ;
  assign n13037 = ~n8672 & ~n13036 ;
  assign n13038 = ~n8666 & n13037 ;
  assign n13039 = ~\u4_u3_buf0_orig_reg[25]/P0001  & n12412 ;
  assign n13040 = n12411 & n13039 ;
  assign n13041 = \u4_u3_buf0_orig_reg[26]/P0001  & ~n13040 ;
  assign n13042 = ~n12415 & ~n13041 ;
  assign n13043 = \sram_data_i[16]_pad  & \wb_addr_i[17]_pad  ;
  assign n13044 = \u4_dout_reg[16]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13045 = ~n13043 & ~n13044 ;
  assign n13046 = \sram_data_i[17]_pad  & \wb_addr_i[17]_pad  ;
  assign n13047 = \u4_dout_reg[17]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13048 = ~n13046 & ~n13047 ;
  assign n13049 = \sram_data_i[18]_pad  & \wb_addr_i[17]_pad  ;
  assign n13050 = \u4_dout_reg[18]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13051 = ~n13049 & ~n13050 ;
  assign n13052 = \sram_data_i[19]_pad  & \wb_addr_i[17]_pad  ;
  assign n13053 = \u4_dout_reg[19]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13054 = ~n13052 & ~n13053 ;
  assign n13055 = \sram_data_i[20]_pad  & \wb_addr_i[17]_pad  ;
  assign n13056 = \u4_dout_reg[20]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13057 = ~n13055 & ~n13056 ;
  assign n13058 = \sram_data_i[21]_pad  & \wb_addr_i[17]_pad  ;
  assign n13059 = \u4_dout_reg[21]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13060 = ~n13058 & ~n13059 ;
  assign n13061 = \sram_data_i[25]_pad  & \wb_addr_i[17]_pad  ;
  assign n13062 = \u4_dout_reg[25]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13063 = ~n13061 & ~n13062 ;
  assign n13064 = \sram_data_i[26]_pad  & \wb_addr_i[17]_pad  ;
  assign n13065 = \u4_dout_reg[26]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13066 = ~n13064 & ~n13065 ;
  assign n13067 = \sram_data_i[27]_pad  & \wb_addr_i[17]_pad  ;
  assign n13068 = \u4_dout_reg[27]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13069 = ~n13067 & ~n13068 ;
  assign n13070 = \sram_data_i[28]_pad  & \wb_addr_i[17]_pad  ;
  assign n13071 = \u4_dout_reg[28]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13072 = ~n13070 & ~n13071 ;
  assign n13073 = \sram_data_i[29]_pad  & \wb_addr_i[17]_pad  ;
  assign n13074 = \u4_dout_reg[29]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13075 = ~n13073 & ~n13074 ;
  assign n13076 = \sram_data_i[30]_pad  & \wb_addr_i[17]_pad  ;
  assign n13077 = \u4_dout_reg[30]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13078 = ~n13076 & ~n13077 ;
  assign n13079 = \sram_data_i[31]_pad  & \wb_addr_i[17]_pad  ;
  assign n13080 = \u4_dout_reg[31]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13081 = ~n13079 & ~n13080 ;
  assign n13082 = \sram_data_i[5]_pad  & \wb_addr_i[17]_pad  ;
  assign n13083 = \u4_dout_reg[5]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13084 = ~n13082 & ~n13083 ;
  assign n13085 = \sram_data_i[6]_pad  & \wb_addr_i[17]_pad  ;
  assign n13086 = \u4_dout_reg[6]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13087 = ~n13085 & ~n13086 ;
  assign n13088 = \sram_data_i[8]_pad  & \wb_addr_i[17]_pad  ;
  assign n13089 = \u4_dout_reg[8]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13090 = ~n13088 & ~n13089 ;
  assign n13091 = n12438 & n12441 ;
  assign n13092 = ~\u4_u0_buf0_orig_reg[23]/P0001  & ~\u4_u0_buf0_orig_reg[25]/P0001  ;
  assign n13093 = ~\u4_u0_buf0_orig_reg[24]/P0001  & n13092 ;
  assign n13094 = n12441 & n13093 ;
  assign n13095 = \u4_u0_buf0_orig_reg[26]/P0001  & ~n13094 ;
  assign n13096 = ~n13091 & ~n13095 ;
  assign n13097 = \sram_data_i[24]_pad  & \wb_addr_i[17]_pad  ;
  assign n13098 = \u4_dout_reg[24]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n13099 = ~n13097 & ~n13098 ;
  assign n13100 = ~\u4_u1_buf0_orig_reg[25]/P0001  & n12465 ;
  assign n13101 = n12464 & n13100 ;
  assign n13102 = \u4_u1_buf0_orig_reg[26]/P0001  & ~n13101 ;
  assign n13103 = ~n12468 & ~n13102 ;
  assign n13104 = ~\u4_u2_buf0_orig_reg[25]/P0001  & n12488 ;
  assign n13105 = n12487 & n13104 ;
  assign n13106 = \u4_u2_buf0_orig_reg[26]/P0001  & ~n13105 ;
  assign n13107 = ~n12491 & ~n13106 ;
  assign n13108 = ~\u4_u3_buf0_orig_reg[27]/P0001  & n12415 ;
  assign n13109 = \u4_u3_buf0_orig_reg[27]/P0001  & ~n12415 ;
  assign n13110 = ~n13108 & ~n13109 ;
  assign n13111 = ~\u4_u0_buf0_orig_reg[27]/P0001  & n13091 ;
  assign n13112 = \u4_u0_buf0_orig_reg[27]/P0001  & ~n13091 ;
  assign n13113 = ~n13111 & ~n13112 ;
  assign n13114 = ~\u4_u1_buf0_orig_reg[27]/P0001  & n12468 ;
  assign n13115 = \u4_u1_buf0_orig_reg[27]/P0001  & ~n12468 ;
  assign n13116 = ~n13114 & ~n13115 ;
  assign n13117 = ~n4438 & ~n4439 ;
  assign n13118 = \u1_u3_new_sizeb_reg[0]/P0001  & n3483 ;
  assign n13119 = ~n13117 & ~n13118 ;
  assign n13120 = n13117 & n13118 ;
  assign n13121 = ~n13119 & ~n13120 ;
  assign n13122 = ~\u4_u2_buf0_orig_reg[27]/P0001  & n12491 ;
  assign n13123 = \u4_u2_buf0_orig_reg[27]/P0001  & ~n12491 ;
  assign n13124 = ~n13122 & ~n13123 ;
  assign n13125 = ~\u1_u0_rxv1_reg/P0001  & ~n4911 ;
  assign n13126 = ~n10519 & n13125 ;
  assign n13127 = rst_i_pad & n7203 ;
  assign n13128 = rst_i_pad & \u1_u0_rxv1_reg/P0001  ;
  assign n13129 = ~n4936 & n13128 ;
  assign n13130 = ~n13127 & ~n13129 ;
  assign n13131 = ~n13126 & ~n13130 ;
  assign n13132 = n5764 & n5768 ;
  assign n13133 = ~n5762 & ~n13132 ;
  assign n13134 = n5758 & ~n13133 ;
  assign n13135 = ~\u0_u0_chirp_cnt_is_6_reg/P0001  & n13134 ;
  assign n13136 = ~\u0_u0_chirp_cnt_reg[0]/P0001  & ~n13135 ;
  assign n13137 = ~\u0_u0_chirp_cnt_is_6_reg/P0001  & \u0_u0_chirp_cnt_reg[0]/P0001  ;
  assign n13138 = n13134 & n13137 ;
  assign n13139 = ~\u0_u0_state_reg[10]/P0001  & ~n13138 ;
  assign n13140 = ~n13136 & n13139 ;
  assign n13141 = \u4_u2_csr1_reg[0]/P0001  & n5171 ;
  assign n13142 = n5156 & n13141 ;
  assign n13143 = \u4_u1_csr1_reg[0]/P0001  & n5175 ;
  assign n13144 = \u4_u0_csr1_reg[0]/P0001  & n5140 ;
  assign n13145 = ~n13143 & ~n13144 ;
  assign n13146 = ~n13142 & n13145 ;
  assign n13147 = \u4_u3_csr1_reg[0]/P0001  & n5195 ;
  assign n13148 = \u4_csr_reg[15]/NET0131  & n5198 ;
  assign n13149 = ~n13147 & ~n13148 ;
  assign n13150 = n13146 & n13149 ;
  assign n13151 = \u4_u2_csr1_reg[1]/P0001  & n5171 ;
  assign n13152 = n5156 & n13151 ;
  assign n13153 = \u4_u1_csr1_reg[1]/P0001  & n5175 ;
  assign n13154 = \u4_u0_csr1_reg[1]/P0001  & n5140 ;
  assign n13155 = ~n13153 & ~n13154 ;
  assign n13156 = ~n13152 & n13155 ;
  assign n13157 = \u4_u3_csr1_reg[1]/P0001  & n5195 ;
  assign n13158 = \u4_csr_reg[16]/P0001  & n5198 ;
  assign n13159 = ~n13157 & ~n13158 ;
  assign n13160 = n13156 & n13159 ;
  assign n13161 = \u4_u2_buf1_reg[5]/P0001  & n5171 ;
  assign n13162 = n5156 & n13161 ;
  assign n13163 = \u4_u1_buf1_reg[5]/P0001  & n5175 ;
  assign n13164 = \u4_u0_buf1_reg[5]/P0001  & n5140 ;
  assign n13165 = ~n13163 & ~n13164 ;
  assign n13166 = ~n13162 & n13165 ;
  assign n13167 = \u4_u3_buf1_reg[5]/P0001  & n5195 ;
  assign n13168 = \u4_buf1_reg[5]/P0001  & n5198 ;
  assign n13169 = ~n13167 & ~n13168 ;
  assign n13170 = n13166 & n13169 ;
  assign n13171 = \u4_u2_csr1_reg[2]/P0001  & n5171 ;
  assign n13172 = n5156 & n13171 ;
  assign n13173 = \u4_u1_csr1_reg[2]/P0001  & n5175 ;
  assign n13174 = \u4_u0_csr1_reg[2]/P0001  & n5140 ;
  assign n13175 = ~n13173 & ~n13174 ;
  assign n13176 = ~n13172 & n13175 ;
  assign n13177 = \u4_u3_csr1_reg[2]/P0001  & n5195 ;
  assign n13178 = \u4_csr_reg[17]/P0001  & n5198 ;
  assign n13179 = ~n13177 & ~n13178 ;
  assign n13180 = n13176 & n13179 ;
  assign n13181 = \u4_u2_csr0_reg[1]/P0001  & n5171 ;
  assign n13182 = n5156 & n13181 ;
  assign n13183 = \u4_u1_csr0_reg[1]/P0001  & n5175 ;
  assign n13184 = \u4_u0_csr0_reg[1]/P0001  & n5140 ;
  assign n13185 = ~n13183 & ~n13184 ;
  assign n13186 = ~n13182 & n13185 ;
  assign n13187 = \u4_u3_csr0_reg[1]/P0001  & n5195 ;
  assign n13188 = \u4_csr_reg[1]/P0001  & n5198 ;
  assign n13189 = ~n13187 & ~n13188 ;
  assign n13190 = n13186 & n13189 ;
  assign n13191 = \u4_u2_csr1_reg[7]/P0001  & n5171 ;
  assign n13192 = n5156 & n13191 ;
  assign n13193 = \u4_u1_csr1_reg[7]/P0001  & n5175 ;
  assign n13194 = \u4_u0_csr1_reg[7]/P0001  & n5140 ;
  assign n13195 = ~n13193 & ~n13194 ;
  assign n13196 = ~n13192 & n13195 ;
  assign n13197 = \u4_u3_csr1_reg[7]/P0001  & n5195 ;
  assign n13198 = \u4_csr_reg[22]/P0001  & n5198 ;
  assign n13199 = ~n13197 & ~n13198 ;
  assign n13200 = n13196 & n13199 ;
  assign n13201 = \u4_u2_csr1_reg[8]/P0001  & n5171 ;
  assign n13202 = n5156 & n13201 ;
  assign n13203 = \u4_u1_csr1_reg[8]/P0001  & n5175 ;
  assign n13204 = \u4_u0_csr1_reg[8]/P0001  & n5140 ;
  assign n13205 = ~n13203 & ~n13204 ;
  assign n13206 = ~n13202 & n13205 ;
  assign n13207 = \u4_u3_csr1_reg[8]/P0001  & n5195 ;
  assign n13208 = \u4_csr_reg[23]/P0001  & n5198 ;
  assign n13209 = ~n13207 & ~n13208 ;
  assign n13210 = n13206 & n13209 ;
  assign n13211 = \u4_u2_csr1_reg[9]/P0001  & n5171 ;
  assign n13212 = n5156 & n13211 ;
  assign n13213 = \u4_u1_csr1_reg[9]/P0001  & n5175 ;
  assign n13214 = \u4_u0_csr1_reg[9]/P0001  & n5140 ;
  assign n13215 = ~n13213 & ~n13214 ;
  assign n13216 = ~n13212 & n13215 ;
  assign n13217 = \u4_u3_csr1_reg[9]/P0001  & n5195 ;
  assign n13218 = \u4_csr_reg[24]/P0001  & n5198 ;
  assign n13219 = ~n13217 & ~n13218 ;
  assign n13220 = n13216 & n13219 ;
  assign n13221 = \u4_u2_csr1_reg[10]/P0001  & n5171 ;
  assign n13222 = n5156 & n13221 ;
  assign n13223 = \u4_u1_csr1_reg[10]/P0001  & n5175 ;
  assign n13224 = \u4_u0_csr1_reg[10]/P0001  & n5140 ;
  assign n13225 = ~n13223 & ~n13224 ;
  assign n13226 = ~n13222 & n13225 ;
  assign n13227 = \u4_u3_csr1_reg[10]/P0001  & n5195 ;
  assign n13228 = \u4_csr_reg[25]/P0001  & n5198 ;
  assign n13229 = ~n13227 & ~n13228 ;
  assign n13230 = n13226 & n13229 ;
  assign n13231 = \u4_u2_csr1_reg[11]/P0001  & n5171 ;
  assign n13232 = n5156 & n13231 ;
  assign n13233 = \u4_u1_csr1_reg[11]/P0001  & n5175 ;
  assign n13234 = \u4_u0_csr1_reg[11]/P0001  & n5140 ;
  assign n13235 = ~n13233 & ~n13234 ;
  assign n13236 = ~n13232 & n13235 ;
  assign n13237 = \u4_u3_csr1_reg[11]/P0001  & n5195 ;
  assign n13238 = \u4_csr_reg[26]/NET0131  & n5198 ;
  assign n13239 = ~n13237 & ~n13238 ;
  assign n13240 = n13236 & n13239 ;
  assign n13241 = \u4_u2_csr1_reg[12]/P0001  & n5171 ;
  assign n13242 = n5156 & n13241 ;
  assign n13243 = \u4_u1_csr1_reg[12]/P0001  & n5175 ;
  assign n13244 = \u4_u0_csr1_reg[12]/P0001  & n5140 ;
  assign n13245 = ~n13243 & ~n13244 ;
  assign n13246 = ~n13242 & n13245 ;
  assign n13247 = \u4_u3_csr1_reg[12]/P0001  & n5195 ;
  assign n13248 = \u4_csr_reg[27]/NET0131  & n5198 ;
  assign n13249 = ~n13247 & ~n13248 ;
  assign n13250 = n13246 & n13249 ;
  assign n13251 = \u4_u2_uc_dpd_reg[0]/P0001  & n5171 ;
  assign n13252 = n5156 & n13251 ;
  assign n13253 = \u4_u1_uc_dpd_reg[0]/P0001  & n5175 ;
  assign n13254 = \u4_u0_uc_dpd_reg[0]/P0001  & n5140 ;
  assign n13255 = ~n13253 & ~n13254 ;
  assign n13256 = ~n13252 & n13255 ;
  assign n13257 = \u4_u3_uc_dpd_reg[0]/P0001  & n5195 ;
  assign n13258 = \u4_csr_reg[28]/P0001  & n5198 ;
  assign n13259 = ~n13257 & ~n13258 ;
  assign n13260 = n13256 & n13259 ;
  assign n13261 = \u4_u2_uc_dpd_reg[1]/P0001  & n5171 ;
  assign n13262 = n5156 & n13261 ;
  assign n13263 = \u4_u1_uc_dpd_reg[1]/P0001  & n5175 ;
  assign n13264 = \u4_u0_uc_dpd_reg[1]/P0001  & n5140 ;
  assign n13265 = ~n13263 & ~n13264 ;
  assign n13266 = ~n13262 & n13265 ;
  assign n13267 = \u4_u3_uc_dpd_reg[1]/P0001  & n5195 ;
  assign n13268 = \u4_csr_reg[29]/P0001  & n5198 ;
  assign n13269 = ~n13267 & ~n13268 ;
  assign n13270 = n13266 & n13269 ;
  assign n13271 = \u4_u2_csr0_reg[2]/P0001  & n5171 ;
  assign n13272 = n5156 & n13271 ;
  assign n13273 = \u4_u1_csr0_reg[2]/P0001  & n5175 ;
  assign n13274 = \u4_u0_csr0_reg[2]/P0001  & n5140 ;
  assign n13275 = ~n13273 & ~n13274 ;
  assign n13276 = ~n13272 & n13275 ;
  assign n13277 = \u4_u3_csr0_reg[2]/P0001  & n5195 ;
  assign n13278 = \u4_csr_reg[2]/NET0131  & n5198 ;
  assign n13279 = ~n13277 & ~n13278 ;
  assign n13280 = n13276 & n13279 ;
  assign n13281 = \u4_u2_uc_bsel_reg[0]/P0001  & n5171 ;
  assign n13282 = n5156 & n13281 ;
  assign n13283 = \u4_u1_uc_bsel_reg[0]/P0001  & n5175 ;
  assign n13284 = \u4_u0_uc_bsel_reg[0]/P0001  & n5140 ;
  assign n13285 = ~n13283 & ~n13284 ;
  assign n13286 = ~n13282 & n13285 ;
  assign n13287 = \u4_u3_uc_bsel_reg[0]/P0001  & n5195 ;
  assign n13288 = \u4_csr_reg[30]/NET0131  & n5198 ;
  assign n13289 = ~n13287 & ~n13288 ;
  assign n13290 = n13286 & n13289 ;
  assign n13291 = \u4_u2_uc_bsel_reg[1]/P0001  & n5171 ;
  assign n13292 = n5156 & n13291 ;
  assign n13293 = \u4_u1_uc_bsel_reg[1]/P0001  & n5175 ;
  assign n13294 = \u4_u0_uc_bsel_reg[1]/P0001  & n5140 ;
  assign n13295 = ~n13293 & ~n13294 ;
  assign n13296 = ~n13292 & n13295 ;
  assign n13297 = \u4_u3_uc_bsel_reg[1]/P0001  & n5195 ;
  assign n13298 = \u4_csr_reg[31]/P0001  & n5198 ;
  assign n13299 = ~n13297 & ~n13298 ;
  assign n13300 = n13296 & n13299 ;
  assign n13301 = \u4_u2_csr0_reg[3]/NET0131  & n5171 ;
  assign n13302 = n5156 & n13301 ;
  assign n13303 = \u4_u1_csr0_reg[3]/NET0131  & n5175 ;
  assign n13304 = \u4_u0_csr0_reg[3]/NET0131  & n5140 ;
  assign n13305 = ~n13303 & ~n13304 ;
  assign n13306 = ~n13302 & n13305 ;
  assign n13307 = \u4_u3_csr0_reg[3]/NET0131  & n5195 ;
  assign n13308 = \u4_csr_reg[3]/P0001  & n5198 ;
  assign n13309 = ~n13307 & ~n13308 ;
  assign n13310 = n13306 & n13309 ;
  assign n13311 = \u4_u2_csr0_reg[4]/P0001  & n5171 ;
  assign n13312 = n5156 & n13311 ;
  assign n13313 = \u4_u1_csr0_reg[4]/P0001  & n5175 ;
  assign n13314 = \u4_u0_csr0_reg[4]/P0001  & n5140 ;
  assign n13315 = ~n13313 & ~n13314 ;
  assign n13316 = ~n13312 & n13315 ;
  assign n13317 = \u4_u3_csr0_reg[4]/P0001  & n5195 ;
  assign n13318 = \u4_csr_reg[4]/NET0131  & n5198 ;
  assign n13319 = ~n13317 & ~n13318 ;
  assign n13320 = n13316 & n13319 ;
  assign n13321 = \u4_u2_csr0_reg[5]/P0001  & n5171 ;
  assign n13322 = n5156 & n13321 ;
  assign n13323 = \u4_u1_csr0_reg[5]/P0001  & n5175 ;
  assign n13324 = \u4_u0_csr0_reg[5]/P0001  & n5140 ;
  assign n13325 = ~n13323 & ~n13324 ;
  assign n13326 = ~n13322 & n13325 ;
  assign n13327 = \u4_u3_csr0_reg[5]/P0001  & n5195 ;
  assign n13328 = \u4_csr_reg[5]/NET0131  & n5198 ;
  assign n13329 = ~n13327 & ~n13328 ;
  assign n13330 = n13326 & n13329 ;
  assign n13331 = \u4_u2_csr0_reg[6]/P0001  & n5171 ;
  assign n13332 = n5156 & n13331 ;
  assign n13333 = \u4_u1_csr0_reg[6]/P0001  & n5175 ;
  assign n13334 = \u4_u0_csr0_reg[6]/P0001  & n5140 ;
  assign n13335 = ~n13333 & ~n13334 ;
  assign n13336 = ~n13332 & n13335 ;
  assign n13337 = \u4_u3_csr0_reg[6]/P0001  & n5195 ;
  assign n13338 = \u4_csr_reg[6]/NET0131  & n5198 ;
  assign n13339 = ~n13337 & ~n13338 ;
  assign n13340 = n13336 & n13339 ;
  assign n13341 = \u4_u2_csr0_reg[7]/P0001  & n5171 ;
  assign n13342 = n5156 & n13341 ;
  assign n13343 = \u4_u1_csr0_reg[7]/P0001  & n5175 ;
  assign n13344 = \u4_u0_csr0_reg[7]/P0001  & n5140 ;
  assign n13345 = ~n13343 & ~n13344 ;
  assign n13346 = ~n13342 & n13345 ;
  assign n13347 = \u4_u3_csr0_reg[7]/P0001  & n5195 ;
  assign n13348 = \u4_csr_reg[7]/P0001  & n5198 ;
  assign n13349 = ~n13347 & ~n13348 ;
  assign n13350 = n13346 & n13349 ;
  assign n13351 = \u4_u2_csr0_reg[8]/P0001  & n5171 ;
  assign n13352 = n5156 & n13351 ;
  assign n13353 = \u4_u1_csr0_reg[8]/P0001  & n5175 ;
  assign n13354 = \u4_u0_csr0_reg[8]/P0001  & n5140 ;
  assign n13355 = ~n13353 & ~n13354 ;
  assign n13356 = ~n13352 & n13355 ;
  assign n13357 = \u4_u3_csr0_reg[8]/P0001  & n5195 ;
  assign n13358 = \u4_csr_reg[8]/P0001  & n5198 ;
  assign n13359 = ~n13357 & ~n13358 ;
  assign n13360 = n13356 & n13359 ;
  assign n13361 = \u4_u2_csr0_reg[9]/P0001  & n5171 ;
  assign n13362 = n5156 & n13361 ;
  assign n13363 = \u4_u1_csr0_reg[9]/P0001  & n5175 ;
  assign n13364 = \u4_u0_csr0_reg[9]/P0001  & n5140 ;
  assign n13365 = ~n13363 & ~n13364 ;
  assign n13366 = ~n13362 & n13365 ;
  assign n13367 = \u4_u3_csr0_reg[9]/P0001  & n5195 ;
  assign n13368 = \u4_csr_reg[9]/NET0131  & n5198 ;
  assign n13369 = ~n13367 & ~n13368 ;
  assign n13370 = n13366 & n13369 ;
  assign n13371 = \u4_u2_buf1_reg[24]/P0001  & n5171 ;
  assign n13372 = n5156 & n13371 ;
  assign n13373 = \u4_u1_buf1_reg[24]/P0001  & n5175 ;
  assign n13374 = \u4_u0_buf1_reg[24]/P0001  & n5140 ;
  assign n13375 = ~n13373 & ~n13374 ;
  assign n13376 = ~n13372 & n13375 ;
  assign n13377 = \u4_u3_buf1_reg[24]/P0001  & n5195 ;
  assign n13378 = \u4_buf1_reg[24]/NET0131  & n5198 ;
  assign n13379 = ~n13377 & ~n13378 ;
  assign n13380 = n13376 & n13379 ;
  assign n13381 = \u4_u2_buf0_reg[0]/P0001  & n5171 ;
  assign n13382 = n5156 & n13381 ;
  assign n13383 = \u4_u1_buf0_reg[0]/P0001  & n5175 ;
  assign n13384 = \u4_u0_buf0_reg[0]/P0001  & n5140 ;
  assign n13385 = ~n13383 & ~n13384 ;
  assign n13386 = ~n13382 & n13385 ;
  assign n13387 = \u4_u3_buf0_reg[0]/P0001  & n5195 ;
  assign n13388 = \u4_buf0_reg[0]/P0001  & n5198 ;
  assign n13389 = ~n13387 & ~n13388 ;
  assign n13390 = n13386 & n13389 ;
  assign n13391 = \u4_u2_buf0_reg[10]/P0001  & n5171 ;
  assign n13392 = n5156 & n13391 ;
  assign n13393 = \u4_u1_buf0_reg[10]/P0001  & n5175 ;
  assign n13394 = \u4_u0_buf0_reg[10]/P0001  & n5140 ;
  assign n13395 = ~n13393 & ~n13394 ;
  assign n13396 = ~n13392 & n13395 ;
  assign n13397 = \u4_u3_buf0_reg[10]/P0001  & n5195 ;
  assign n13398 = \u4_buf0_reg[10]/P0001  & n5198 ;
  assign n13399 = ~n13397 & ~n13398 ;
  assign n13400 = n13396 & n13399 ;
  assign n13401 = \u4_u2_buf0_reg[11]/P0001  & n5171 ;
  assign n13402 = n5156 & n13401 ;
  assign n13403 = \u4_u1_buf0_reg[11]/P0001  & n5175 ;
  assign n13404 = \u4_u0_buf0_reg[11]/P0001  & n5140 ;
  assign n13405 = ~n13403 & ~n13404 ;
  assign n13406 = ~n13402 & n13405 ;
  assign n13407 = \u4_u3_buf0_reg[11]/P0001  & n5195 ;
  assign n13408 = \u4_buf0_reg[11]/P0001  & n5198 ;
  assign n13409 = ~n13407 & ~n13408 ;
  assign n13410 = n13406 & n13409 ;
  assign n13411 = \u4_u2_buf0_reg[12]/P0001  & n5171 ;
  assign n13412 = n5156 & n13411 ;
  assign n13413 = \u4_u1_buf0_reg[12]/P0001  & n5175 ;
  assign n13414 = \u4_u0_buf0_reg[12]/P0001  & n5140 ;
  assign n13415 = ~n13413 & ~n13414 ;
  assign n13416 = ~n13412 & n13415 ;
  assign n13417 = \u4_u3_buf0_reg[12]/P0001  & n5195 ;
  assign n13418 = \u4_buf0_reg[12]/P0001  & n5198 ;
  assign n13419 = ~n13417 & ~n13418 ;
  assign n13420 = n13416 & n13419 ;
  assign n13421 = \u4_u2_buf0_reg[13]/P0001  & n5171 ;
  assign n13422 = n5156 & n13421 ;
  assign n13423 = \u4_u1_buf0_reg[13]/P0001  & n5175 ;
  assign n13424 = \u4_u0_buf0_reg[13]/P0001  & n5140 ;
  assign n13425 = ~n13423 & ~n13424 ;
  assign n13426 = ~n13422 & n13425 ;
  assign n13427 = \u4_u3_buf0_reg[13]/P0001  & n5195 ;
  assign n13428 = \u4_buf0_reg[13]/P0001  & n5198 ;
  assign n13429 = ~n13427 & ~n13428 ;
  assign n13430 = n13426 & n13429 ;
  assign n13431 = \u4_u2_buf0_reg[14]/P0001  & n5171 ;
  assign n13432 = n5156 & n13431 ;
  assign n13433 = \u4_u1_buf0_reg[14]/P0001  & n5175 ;
  assign n13434 = \u4_u0_buf0_reg[14]/P0001  & n5140 ;
  assign n13435 = ~n13433 & ~n13434 ;
  assign n13436 = ~n13432 & n13435 ;
  assign n13437 = \u4_u3_buf0_reg[14]/P0001  & n5195 ;
  assign n13438 = \u4_buf0_reg[14]/P0001  & n5198 ;
  assign n13439 = ~n13437 & ~n13438 ;
  assign n13440 = n13436 & n13439 ;
  assign n13441 = \u4_u2_buf0_reg[15]/P0001  & n5171 ;
  assign n13442 = n5156 & n13441 ;
  assign n13443 = \u4_u1_buf0_reg[15]/P0001  & n5175 ;
  assign n13444 = \u4_u0_buf0_reg[15]/P0001  & n5140 ;
  assign n13445 = ~n13443 & ~n13444 ;
  assign n13446 = ~n13442 & n13445 ;
  assign n13447 = \u4_u3_buf0_reg[15]/P0001  & n5195 ;
  assign n13448 = \u4_buf0_reg[15]/P0001  & n5198 ;
  assign n13449 = ~n13447 & ~n13448 ;
  assign n13450 = n13446 & n13449 ;
  assign n13451 = \u4_u2_buf0_reg[16]/P0001  & n5171 ;
  assign n13452 = n5156 & n13451 ;
  assign n13453 = \u4_u1_buf0_reg[16]/P0001  & n5175 ;
  assign n13454 = \u4_u0_buf0_reg[16]/P0001  & n5140 ;
  assign n13455 = ~n13453 & ~n13454 ;
  assign n13456 = ~n13452 & n13455 ;
  assign n13457 = \u4_u3_buf0_reg[16]/P0001  & n5195 ;
  assign n13458 = \u4_buf0_reg[16]/P0001  & n5198 ;
  assign n13459 = ~n13457 & ~n13458 ;
  assign n13460 = n13456 & n13459 ;
  assign n13461 = \u4_u2_buf0_reg[17]/P0001  & n5171 ;
  assign n13462 = n5156 & n13461 ;
  assign n13463 = \u4_u1_buf0_reg[17]/P0001  & n5175 ;
  assign n13464 = \u4_u0_buf0_reg[17]/P0001  & n5140 ;
  assign n13465 = ~n13463 & ~n13464 ;
  assign n13466 = ~n13462 & n13465 ;
  assign n13467 = \u4_u3_buf0_reg[17]/P0001  & n5195 ;
  assign n13468 = \u4_buf0_reg[17]/NET0131  & n5198 ;
  assign n13469 = ~n13467 & ~n13468 ;
  assign n13470 = n13466 & n13469 ;
  assign n13471 = \u4_u2_buf0_reg[18]/P0001  & n5171 ;
  assign n13472 = n5156 & n13471 ;
  assign n13473 = \u4_u1_buf0_reg[18]/P0001  & n5175 ;
  assign n13474 = \u4_u0_buf0_reg[18]/P0001  & n5140 ;
  assign n13475 = ~n13473 & ~n13474 ;
  assign n13476 = ~n13472 & n13475 ;
  assign n13477 = \u4_u3_buf0_reg[18]/P0001  & n5195 ;
  assign n13478 = \u4_buf0_reg[18]/P0001  & n5198 ;
  assign n13479 = ~n13477 & ~n13478 ;
  assign n13480 = n13476 & n13479 ;
  assign n13481 = \u4_u2_buf0_reg[19]/P0001  & n5171 ;
  assign n13482 = n5156 & n13481 ;
  assign n13483 = \u4_u1_buf0_reg[19]/P0001  & n5175 ;
  assign n13484 = \u4_u0_buf0_reg[19]/P0001  & n5140 ;
  assign n13485 = ~n13483 & ~n13484 ;
  assign n13486 = ~n13482 & n13485 ;
  assign n13487 = \u4_u3_buf0_reg[19]/P0001  & n5195 ;
  assign n13488 = \u4_buf0_reg[19]/NET0131  & n5198 ;
  assign n13489 = ~n13487 & ~n13488 ;
  assign n13490 = n13486 & n13489 ;
  assign n13491 = \u4_u2_buf1_reg[6]/P0001  & n5171 ;
  assign n13492 = n5156 & n13491 ;
  assign n13493 = \u4_u1_buf1_reg[6]/P0001  & n5175 ;
  assign n13494 = \u4_u0_buf1_reg[6]/P0001  & n5140 ;
  assign n13495 = ~n13493 & ~n13494 ;
  assign n13496 = ~n13492 & n13495 ;
  assign n13497 = \u4_u3_buf1_reg[6]/P0001  & n5195 ;
  assign n13498 = \u4_buf1_reg[6]/P0001  & n5198 ;
  assign n13499 = ~n13497 & ~n13498 ;
  assign n13500 = n13496 & n13499 ;
  assign n13501 = \u4_u2_buf0_reg[1]/P0001  & n5171 ;
  assign n13502 = n5156 & n13501 ;
  assign n13503 = \u4_u1_buf0_reg[1]/P0001  & n5175 ;
  assign n13504 = \u4_u0_buf0_reg[1]/P0001  & n5140 ;
  assign n13505 = ~n13503 & ~n13504 ;
  assign n13506 = ~n13502 & n13505 ;
  assign n13507 = \u4_u3_buf0_reg[1]/P0001  & n5195 ;
  assign n13508 = \u4_buf0_reg[1]/P0001  & n5198 ;
  assign n13509 = ~n13507 & ~n13508 ;
  assign n13510 = n13506 & n13509 ;
  assign n13511 = \u4_u2_buf0_reg[20]/P0001  & n5171 ;
  assign n13512 = n5156 & n13511 ;
  assign n13513 = \u4_u1_buf0_reg[20]/P0001  & n5175 ;
  assign n13514 = \u4_u0_buf0_reg[20]/P0001  & n5140 ;
  assign n13515 = ~n13513 & ~n13514 ;
  assign n13516 = ~n13512 & n13515 ;
  assign n13517 = \u4_u3_buf0_reg[20]/P0001  & n5195 ;
  assign n13518 = \u4_buf0_reg[20]/NET0131  & n5198 ;
  assign n13519 = ~n13517 & ~n13518 ;
  assign n13520 = n13516 & n13519 ;
  assign n13521 = \u4_u2_buf0_reg[21]/P0001  & n5171 ;
  assign n13522 = n5156 & n13521 ;
  assign n13523 = \u4_u1_buf0_reg[21]/P0001  & n5175 ;
  assign n13524 = \u4_u0_buf0_reg[21]/P0001  & n5140 ;
  assign n13525 = ~n13523 & ~n13524 ;
  assign n13526 = ~n13522 & n13525 ;
  assign n13527 = \u4_u3_buf0_reg[21]/P0001  & n5195 ;
  assign n13528 = \u4_buf0_reg[21]/NET0131  & n5198 ;
  assign n13529 = ~n13527 & ~n13528 ;
  assign n13530 = n13526 & n13529 ;
  assign n13531 = \u4_u2_buf0_reg[22]/P0001  & n5171 ;
  assign n13532 = n5156 & n13531 ;
  assign n13533 = \u4_u1_buf0_reg[22]/P0001  & n5175 ;
  assign n13534 = \u4_u0_buf0_reg[22]/P0001  & n5140 ;
  assign n13535 = ~n13533 & ~n13534 ;
  assign n13536 = ~n13532 & n13535 ;
  assign n13537 = \u4_u3_buf0_reg[22]/P0001  & n5195 ;
  assign n13538 = \u4_buf0_reg[22]/NET0131  & n5198 ;
  assign n13539 = ~n13537 & ~n13538 ;
  assign n13540 = n13536 & n13539 ;
  assign n13541 = \u4_u2_buf0_reg[23]/P0001  & n5171 ;
  assign n13542 = n5156 & n13541 ;
  assign n13543 = \u4_u1_buf0_reg[23]/P0001  & n5175 ;
  assign n13544 = \u4_u0_buf0_reg[23]/P0001  & n5140 ;
  assign n13545 = ~n13543 & ~n13544 ;
  assign n13546 = ~n13542 & n13545 ;
  assign n13547 = \u4_u3_buf0_reg[23]/P0001  & n5195 ;
  assign n13548 = \u4_buf0_reg[23]/NET0131  & n5198 ;
  assign n13549 = ~n13547 & ~n13548 ;
  assign n13550 = n13546 & n13549 ;
  assign n13551 = \u4_u2_buf0_reg[24]/P0001  & n5171 ;
  assign n13552 = n5156 & n13551 ;
  assign n13553 = \u4_u1_buf0_reg[24]/P0001  & n5175 ;
  assign n13554 = \u4_u0_buf0_reg[24]/P0001  & n5140 ;
  assign n13555 = ~n13553 & ~n13554 ;
  assign n13556 = ~n13552 & n13555 ;
  assign n13557 = \u4_u3_buf0_reg[24]/P0001  & n5195 ;
  assign n13558 = \u4_buf0_reg[24]/NET0131  & n5198 ;
  assign n13559 = ~n13557 & ~n13558 ;
  assign n13560 = n13556 & n13559 ;
  assign n13561 = \u4_u2_buf0_reg[25]/P0001  & n5171 ;
  assign n13562 = n5156 & n13561 ;
  assign n13563 = \u4_u1_buf0_reg[25]/P0001  & n5175 ;
  assign n13564 = \u4_u0_buf0_reg[25]/P0001  & n5140 ;
  assign n13565 = ~n13563 & ~n13564 ;
  assign n13566 = ~n13562 & n13565 ;
  assign n13567 = \u4_u3_buf0_reg[25]/P0001  & n5195 ;
  assign n13568 = \u4_buf0_reg[25]/NET0131  & n5198 ;
  assign n13569 = ~n13567 & ~n13568 ;
  assign n13570 = n13566 & n13569 ;
  assign n13571 = \u4_u2_buf0_reg[26]/P0001  & n5171 ;
  assign n13572 = n5156 & n13571 ;
  assign n13573 = \u4_u1_buf0_reg[26]/P0001  & n5175 ;
  assign n13574 = \u4_u0_buf0_reg[26]/P0001  & n5140 ;
  assign n13575 = ~n13573 & ~n13574 ;
  assign n13576 = ~n13572 & n13575 ;
  assign n13577 = \u4_u3_buf0_reg[26]/P0001  & n5195 ;
  assign n13578 = \u4_buf0_reg[26]/NET0131  & n5198 ;
  assign n13579 = ~n13577 & ~n13578 ;
  assign n13580 = n13576 & n13579 ;
  assign n13581 = \u4_u2_buf0_reg[27]/P0001  & n5171 ;
  assign n13582 = n5156 & n13581 ;
  assign n13583 = \u4_u1_buf0_reg[27]/P0001  & n5175 ;
  assign n13584 = \u4_u0_buf0_reg[27]/P0001  & n5140 ;
  assign n13585 = ~n13583 & ~n13584 ;
  assign n13586 = ~n13582 & n13585 ;
  assign n13587 = \u4_u3_buf0_reg[27]/P0001  & n5195 ;
  assign n13588 = \u4_buf0_reg[27]/P0001  & n5198 ;
  assign n13589 = ~n13587 & ~n13588 ;
  assign n13590 = n13586 & n13589 ;
  assign n13591 = \u4_u2_buf0_reg[28]/P0001  & n5171 ;
  assign n13592 = n5156 & n13591 ;
  assign n13593 = \u4_u1_buf0_reg[28]/P0001  & n5175 ;
  assign n13594 = \u4_u0_buf0_reg[28]/P0001  & n5140 ;
  assign n13595 = ~n13593 & ~n13594 ;
  assign n13596 = ~n13592 & n13595 ;
  assign n13597 = \u4_u3_buf0_reg[28]/P0001  & n5195 ;
  assign n13598 = \u4_buf0_reg[28]/P0001  & n5198 ;
  assign n13599 = ~n13597 & ~n13598 ;
  assign n13600 = n13596 & n13599 ;
  assign n13601 = \u4_u2_buf0_reg[29]/P0001  & n5171 ;
  assign n13602 = n5156 & n13601 ;
  assign n13603 = \u4_u1_buf0_reg[29]/P0001  & n5175 ;
  assign n13604 = \u4_u0_buf0_reg[29]/P0001  & n5140 ;
  assign n13605 = ~n13603 & ~n13604 ;
  assign n13606 = ~n13602 & n13605 ;
  assign n13607 = \u4_u3_buf0_reg[29]/P0001  & n5195 ;
  assign n13608 = \u4_buf0_reg[29]/P0001  & n5198 ;
  assign n13609 = ~n13607 & ~n13608 ;
  assign n13610 = n13606 & n13609 ;
  assign n13611 = \u4_u2_buf0_reg[2]/P0001  & n5171 ;
  assign n13612 = n5156 & n13611 ;
  assign n13613 = \u4_u1_buf0_reg[2]/P0001  & n5175 ;
  assign n13614 = \u4_u0_buf0_reg[2]/P0001  & n5140 ;
  assign n13615 = ~n13613 & ~n13614 ;
  assign n13616 = ~n13612 & n13615 ;
  assign n13617 = \u4_u3_buf0_reg[2]/P0001  & n5195 ;
  assign n13618 = \u4_buf0_reg[2]/P0001  & n5198 ;
  assign n13619 = ~n13617 & ~n13618 ;
  assign n13620 = n13616 & n13619 ;
  assign n13621 = \u4_u2_buf0_reg[30]/P0001  & n5171 ;
  assign n13622 = n5156 & n13621 ;
  assign n13623 = \u4_u1_buf0_reg[30]/P0001  & n5175 ;
  assign n13624 = \u4_u0_buf0_reg[30]/P0001  & n5140 ;
  assign n13625 = ~n13623 & ~n13624 ;
  assign n13626 = ~n13622 & n13625 ;
  assign n13627 = \u4_u3_buf0_reg[30]/P0001  & n5195 ;
  assign n13628 = \u4_buf0_reg[30]/P0001  & n5198 ;
  assign n13629 = ~n13627 & ~n13628 ;
  assign n13630 = n13626 & n13629 ;
  assign n13631 = \u4_u2_buf0_reg[31]/P0001  & n5171 ;
  assign n13632 = n5156 & n13631 ;
  assign n13633 = \u4_u1_buf0_reg[31]/P0001  & n5175 ;
  assign n13634 = \u4_u0_buf0_reg[31]/P0001  & n5140 ;
  assign n13635 = ~n13633 & ~n13634 ;
  assign n13636 = ~n13632 & n13635 ;
  assign n13637 = \u4_u3_buf0_reg[31]/P0001  & n5195 ;
  assign n13638 = \u4_buf0_reg[31]/P0001  & n5198 ;
  assign n13639 = ~n13637 & ~n13638 ;
  assign n13640 = n13636 & n13639 ;
  assign n13641 = \u4_u2_buf0_reg[3]/P0001  & n5171 ;
  assign n13642 = n5156 & n13641 ;
  assign n13643 = \u4_u1_buf0_reg[3]/P0001  & n5175 ;
  assign n13644 = \u4_u0_buf0_reg[3]/P0001  & n5140 ;
  assign n13645 = ~n13643 & ~n13644 ;
  assign n13646 = ~n13642 & n13645 ;
  assign n13647 = \u4_u3_buf0_reg[3]/P0001  & n5195 ;
  assign n13648 = \u4_buf0_reg[3]/P0001  & n5198 ;
  assign n13649 = ~n13647 & ~n13648 ;
  assign n13650 = n13646 & n13649 ;
  assign n13651 = \u4_u2_buf0_reg[4]/P0001  & n5171 ;
  assign n13652 = n5156 & n13651 ;
  assign n13653 = \u4_u1_buf0_reg[4]/P0001  & n5175 ;
  assign n13654 = \u4_u0_buf0_reg[4]/P0001  & n5140 ;
  assign n13655 = ~n13653 & ~n13654 ;
  assign n13656 = ~n13652 & n13655 ;
  assign n13657 = \u4_u3_buf0_reg[4]/P0001  & n5195 ;
  assign n13658 = \u4_buf0_reg[4]/P0001  & n5198 ;
  assign n13659 = ~n13657 & ~n13658 ;
  assign n13660 = n13656 & n13659 ;
  assign n13661 = \u4_u2_buf0_reg[5]/P0001  & n5171 ;
  assign n13662 = n5156 & n13661 ;
  assign n13663 = \u4_u1_buf0_reg[5]/P0001  & n5175 ;
  assign n13664 = \u4_u0_buf0_reg[5]/P0001  & n5140 ;
  assign n13665 = ~n13663 & ~n13664 ;
  assign n13666 = ~n13662 & n13665 ;
  assign n13667 = \u4_u3_buf0_reg[5]/P0001  & n5195 ;
  assign n13668 = \u4_buf0_reg[5]/P0001  & n5198 ;
  assign n13669 = ~n13667 & ~n13668 ;
  assign n13670 = n13666 & n13669 ;
  assign n13671 = \u4_u2_buf0_reg[6]/P0001  & n5171 ;
  assign n13672 = n5156 & n13671 ;
  assign n13673 = \u4_u1_buf0_reg[6]/P0001  & n5175 ;
  assign n13674 = \u4_u0_buf0_reg[6]/P0001  & n5140 ;
  assign n13675 = ~n13673 & ~n13674 ;
  assign n13676 = ~n13672 & n13675 ;
  assign n13677 = \u4_u3_buf0_reg[6]/P0001  & n5195 ;
  assign n13678 = \u4_buf0_reg[6]/P0001  & n5198 ;
  assign n13679 = ~n13677 & ~n13678 ;
  assign n13680 = n13676 & n13679 ;
  assign n13681 = \u4_u2_buf0_reg[7]/P0001  & n5171 ;
  assign n13682 = n5156 & n13681 ;
  assign n13683 = \u4_u1_buf0_reg[7]/P0001  & n5175 ;
  assign n13684 = \u4_u0_buf0_reg[7]/P0001  & n5140 ;
  assign n13685 = ~n13683 & ~n13684 ;
  assign n13686 = ~n13682 & n13685 ;
  assign n13687 = \u4_u3_buf0_reg[7]/P0001  & n5195 ;
  assign n13688 = \u4_buf0_reg[7]/P0001  & n5198 ;
  assign n13689 = ~n13687 & ~n13688 ;
  assign n13690 = n13686 & n13689 ;
  assign n13691 = \u4_u2_buf0_reg[8]/P0001  & n5171 ;
  assign n13692 = n5156 & n13691 ;
  assign n13693 = \u4_u1_buf0_reg[8]/P0001  & n5175 ;
  assign n13694 = \u4_u0_buf0_reg[8]/P0001  & n5140 ;
  assign n13695 = ~n13693 & ~n13694 ;
  assign n13696 = ~n13692 & n13695 ;
  assign n13697 = \u4_u3_buf0_reg[8]/P0001  & n5195 ;
  assign n13698 = \u4_buf0_reg[8]/P0001  & n5198 ;
  assign n13699 = ~n13697 & ~n13698 ;
  assign n13700 = n13696 & n13699 ;
  assign n13701 = \u4_u2_buf0_reg[9]/P0001  & n5171 ;
  assign n13702 = n5156 & n13701 ;
  assign n13703 = \u4_u1_buf0_reg[9]/P0001  & n5175 ;
  assign n13704 = \u4_u0_buf0_reg[9]/P0001  & n5140 ;
  assign n13705 = ~n13703 & ~n13704 ;
  assign n13706 = ~n13702 & n13705 ;
  assign n13707 = \u4_u3_buf0_reg[9]/P0001  & n5195 ;
  assign n13708 = \u4_buf0_reg[9]/P0001  & n5198 ;
  assign n13709 = ~n13707 & ~n13708 ;
  assign n13710 = n13706 & n13709 ;
  assign n13711 = \u4_u2_buf1_reg[0]/P0001  & n5171 ;
  assign n13712 = n5156 & n13711 ;
  assign n13713 = \u4_u1_buf1_reg[0]/P0001  & n5175 ;
  assign n13714 = \u4_u0_buf1_reg[0]/P0001  & n5140 ;
  assign n13715 = ~n13713 & ~n13714 ;
  assign n13716 = ~n13712 & n13715 ;
  assign n13717 = \u4_u3_buf1_reg[0]/P0001  & n5195 ;
  assign n13718 = \u4_buf1_reg[0]/P0001  & n5198 ;
  assign n13719 = ~n13717 & ~n13718 ;
  assign n13720 = n13716 & n13719 ;
  assign n13721 = \u4_u2_buf1_reg[10]/P0001  & n5171 ;
  assign n13722 = n5156 & n13721 ;
  assign n13723 = \u4_u1_buf1_reg[10]/P0001  & n5175 ;
  assign n13724 = \u4_u0_buf1_reg[10]/P0001  & n5140 ;
  assign n13725 = ~n13723 & ~n13724 ;
  assign n13726 = ~n13722 & n13725 ;
  assign n13727 = \u4_u3_buf1_reg[10]/P0001  & n5195 ;
  assign n13728 = \u4_buf1_reg[10]/P0001  & n5198 ;
  assign n13729 = ~n13727 & ~n13728 ;
  assign n13730 = n13726 & n13729 ;
  assign n13731 = \u4_u2_buf1_reg[11]/P0001  & n5171 ;
  assign n13732 = n5156 & n13731 ;
  assign n13733 = \u4_u1_buf1_reg[11]/P0001  & n5175 ;
  assign n13734 = \u4_u0_buf1_reg[11]/P0001  & n5140 ;
  assign n13735 = ~n13733 & ~n13734 ;
  assign n13736 = ~n13732 & n13735 ;
  assign n13737 = \u4_u3_buf1_reg[11]/P0001  & n5195 ;
  assign n13738 = \u4_buf1_reg[11]/P0001  & n5198 ;
  assign n13739 = ~n13737 & ~n13738 ;
  assign n13740 = n13736 & n13739 ;
  assign n13741 = \u4_u2_buf1_reg[12]/P0001  & n5171 ;
  assign n13742 = n5156 & n13741 ;
  assign n13743 = \u4_u1_buf1_reg[12]/P0001  & n5175 ;
  assign n13744 = \u4_u0_buf1_reg[12]/P0001  & n5140 ;
  assign n13745 = ~n13743 & ~n13744 ;
  assign n13746 = ~n13742 & n13745 ;
  assign n13747 = \u4_u3_buf1_reg[12]/P0001  & n5195 ;
  assign n13748 = \u4_buf1_reg[12]/P0001  & n5198 ;
  assign n13749 = ~n13747 & ~n13748 ;
  assign n13750 = n13746 & n13749 ;
  assign n13751 = \u4_u2_buf1_reg[13]/P0001  & n5171 ;
  assign n13752 = n5156 & n13751 ;
  assign n13753 = \u4_u1_buf1_reg[13]/P0001  & n5175 ;
  assign n13754 = \u4_u0_buf1_reg[13]/P0001  & n5140 ;
  assign n13755 = ~n13753 & ~n13754 ;
  assign n13756 = ~n13752 & n13755 ;
  assign n13757 = \u4_u3_buf1_reg[13]/P0001  & n5195 ;
  assign n13758 = \u4_buf1_reg[13]/P0001  & n5198 ;
  assign n13759 = ~n13757 & ~n13758 ;
  assign n13760 = n13756 & n13759 ;
  assign n13761 = \u4_u2_buf1_reg[14]/P0001  & n5171 ;
  assign n13762 = n5156 & n13761 ;
  assign n13763 = \u4_u1_buf1_reg[14]/P0001  & n5175 ;
  assign n13764 = \u4_u0_buf1_reg[14]/P0001  & n5140 ;
  assign n13765 = ~n13763 & ~n13764 ;
  assign n13766 = ~n13762 & n13765 ;
  assign n13767 = \u4_u3_buf1_reg[14]/P0001  & n5195 ;
  assign n13768 = \u4_buf1_reg[14]/P0001  & n5198 ;
  assign n13769 = ~n13767 & ~n13768 ;
  assign n13770 = n13766 & n13769 ;
  assign n13771 = \u4_u2_buf1_reg[15]/P0001  & n5171 ;
  assign n13772 = n5156 & n13771 ;
  assign n13773 = \u4_u1_buf1_reg[15]/P0001  & n5175 ;
  assign n13774 = \u4_u0_buf1_reg[15]/P0001  & n5140 ;
  assign n13775 = ~n13773 & ~n13774 ;
  assign n13776 = ~n13772 & n13775 ;
  assign n13777 = \u4_u3_buf1_reg[15]/P0001  & n5195 ;
  assign n13778 = \u4_buf1_reg[15]/P0001  & n5198 ;
  assign n13779 = ~n13777 & ~n13778 ;
  assign n13780 = n13776 & n13779 ;
  assign n13781 = \u4_u2_buf1_reg[16]/P0001  & n5171 ;
  assign n13782 = n5156 & n13781 ;
  assign n13783 = \u4_u1_buf1_reg[16]/P0001  & n5175 ;
  assign n13784 = \u4_u0_buf1_reg[16]/P0001  & n5140 ;
  assign n13785 = ~n13783 & ~n13784 ;
  assign n13786 = ~n13782 & n13785 ;
  assign n13787 = \u4_u3_buf1_reg[16]/P0001  & n5195 ;
  assign n13788 = \u4_buf1_reg[16]/P0001  & n5198 ;
  assign n13789 = ~n13787 & ~n13788 ;
  assign n13790 = n13786 & n13789 ;
  assign n13791 = \u4_u2_buf1_reg[17]/P0001  & n5171 ;
  assign n13792 = n5156 & n13791 ;
  assign n13793 = \u4_u1_buf1_reg[17]/P0001  & n5175 ;
  assign n13794 = \u4_u0_buf1_reg[17]/P0001  & n5140 ;
  assign n13795 = ~n13793 & ~n13794 ;
  assign n13796 = ~n13792 & n13795 ;
  assign n13797 = \u4_u3_buf1_reg[17]/P0001  & n5195 ;
  assign n13798 = \u4_buf1_reg[17]/NET0131  & n5198 ;
  assign n13799 = ~n13797 & ~n13798 ;
  assign n13800 = n13796 & n13799 ;
  assign n13801 = \u4_u2_buf1_reg[18]/P0001  & n5171 ;
  assign n13802 = n5156 & n13801 ;
  assign n13803 = \u4_u1_buf1_reg[18]/P0001  & n5175 ;
  assign n13804 = \u4_u0_buf1_reg[18]/P0001  & n5140 ;
  assign n13805 = ~n13803 & ~n13804 ;
  assign n13806 = ~n13802 & n13805 ;
  assign n13807 = \u4_u3_buf1_reg[18]/P0001  & n5195 ;
  assign n13808 = \u4_buf1_reg[18]/P0001  & n5198 ;
  assign n13809 = ~n13807 & ~n13808 ;
  assign n13810 = n13806 & n13809 ;
  assign n13811 = \u4_u2_buf1_reg[19]/P0001  & n5171 ;
  assign n13812 = n5156 & n13811 ;
  assign n13813 = \u4_u1_buf1_reg[19]/P0001  & n5175 ;
  assign n13814 = \u4_u0_buf1_reg[19]/P0001  & n5140 ;
  assign n13815 = ~n13813 & ~n13814 ;
  assign n13816 = ~n13812 & n13815 ;
  assign n13817 = \u4_u3_buf1_reg[19]/P0001  & n5195 ;
  assign n13818 = \u4_buf1_reg[19]/NET0131  & n5198 ;
  assign n13819 = ~n13817 & ~n13818 ;
  assign n13820 = n13816 & n13819 ;
  assign n13821 = \u4_u2_buf1_reg[1]/P0001  & n5171 ;
  assign n13822 = n5156 & n13821 ;
  assign n13823 = \u4_u1_buf1_reg[1]/P0001  & n5175 ;
  assign n13824 = \u4_u0_buf1_reg[1]/P0001  & n5140 ;
  assign n13825 = ~n13823 & ~n13824 ;
  assign n13826 = ~n13822 & n13825 ;
  assign n13827 = \u4_u3_buf1_reg[1]/P0001  & n5195 ;
  assign n13828 = \u4_buf1_reg[1]/P0001  & n5198 ;
  assign n13829 = ~n13827 & ~n13828 ;
  assign n13830 = n13826 & n13829 ;
  assign n13831 = \u4_u2_buf1_reg[20]/P0001  & n5171 ;
  assign n13832 = n5156 & n13831 ;
  assign n13833 = \u4_u1_buf1_reg[20]/P0001  & n5175 ;
  assign n13834 = \u4_u0_buf1_reg[20]/P0001  & n5140 ;
  assign n13835 = ~n13833 & ~n13834 ;
  assign n13836 = ~n13832 & n13835 ;
  assign n13837 = \u4_u3_buf1_reg[20]/P0001  & n5195 ;
  assign n13838 = \u4_buf1_reg[20]/NET0131  & n5198 ;
  assign n13839 = ~n13837 & ~n13838 ;
  assign n13840 = n13836 & n13839 ;
  assign n13841 = \u4_u2_buf1_reg[21]/P0001  & n5171 ;
  assign n13842 = n5156 & n13841 ;
  assign n13843 = \u4_u1_buf1_reg[21]/P0001  & n5175 ;
  assign n13844 = \u4_u0_buf1_reg[21]/P0001  & n5140 ;
  assign n13845 = ~n13843 & ~n13844 ;
  assign n13846 = ~n13842 & n13845 ;
  assign n13847 = \u4_u3_buf1_reg[21]/P0001  & n5195 ;
  assign n13848 = \u4_buf1_reg[21]/NET0131  & n5198 ;
  assign n13849 = ~n13847 & ~n13848 ;
  assign n13850 = n13846 & n13849 ;
  assign n13851 = \u4_u2_buf1_reg[22]/P0001  & n5171 ;
  assign n13852 = n5156 & n13851 ;
  assign n13853 = \u4_u1_buf1_reg[22]/P0001  & n5175 ;
  assign n13854 = \u4_u0_buf1_reg[22]/P0001  & n5140 ;
  assign n13855 = ~n13853 & ~n13854 ;
  assign n13856 = ~n13852 & n13855 ;
  assign n13857 = \u4_u3_buf1_reg[22]/P0001  & n5195 ;
  assign n13858 = \u4_buf1_reg[22]/NET0131  & n5198 ;
  assign n13859 = ~n13857 & ~n13858 ;
  assign n13860 = n13856 & n13859 ;
  assign n13861 = \u4_u2_buf1_reg[23]/P0001  & n5171 ;
  assign n13862 = n5156 & n13861 ;
  assign n13863 = \u4_u1_buf1_reg[23]/P0001  & n5175 ;
  assign n13864 = \u4_u0_buf1_reg[23]/P0001  & n5140 ;
  assign n13865 = ~n13863 & ~n13864 ;
  assign n13866 = ~n13862 & n13865 ;
  assign n13867 = \u4_u3_buf1_reg[23]/P0001  & n5195 ;
  assign n13868 = \u4_buf1_reg[23]/NET0131  & n5198 ;
  assign n13869 = ~n13867 & ~n13868 ;
  assign n13870 = n13866 & n13869 ;
  assign n13871 = \u4_u2_buf1_reg[25]/P0001  & n5171 ;
  assign n13872 = n5156 & n13871 ;
  assign n13873 = \u4_u1_buf1_reg[25]/P0001  & n5175 ;
  assign n13874 = \u4_u0_buf1_reg[25]/P0001  & n5140 ;
  assign n13875 = ~n13873 & ~n13874 ;
  assign n13876 = ~n13872 & n13875 ;
  assign n13877 = \u4_u3_buf1_reg[25]/P0001  & n5195 ;
  assign n13878 = \u4_buf1_reg[25]/NET0131  & n5198 ;
  assign n13879 = ~n13877 & ~n13878 ;
  assign n13880 = n13876 & n13879 ;
  assign n13881 = \u4_u2_buf1_reg[3]/P0001  & n5171 ;
  assign n13882 = n5156 & n13881 ;
  assign n13883 = \u4_u1_buf1_reg[3]/P0001  & n5175 ;
  assign n13884 = \u4_u0_buf1_reg[3]/P0001  & n5140 ;
  assign n13885 = ~n13883 & ~n13884 ;
  assign n13886 = ~n13882 & n13885 ;
  assign n13887 = \u4_u3_buf1_reg[3]/P0001  & n5195 ;
  assign n13888 = \u4_buf1_reg[3]/P0001  & n5198 ;
  assign n13889 = ~n13887 & ~n13888 ;
  assign n13890 = n13886 & n13889 ;
  assign n13891 = \u4_u2_buf1_reg[26]/P0001  & n5171 ;
  assign n13892 = n5156 & n13891 ;
  assign n13893 = \u4_u1_buf1_reg[26]/P0001  & n5175 ;
  assign n13894 = \u4_u0_buf1_reg[26]/P0001  & n5140 ;
  assign n13895 = ~n13893 & ~n13894 ;
  assign n13896 = ~n13892 & n13895 ;
  assign n13897 = \u4_u3_buf1_reg[26]/P0001  & n5195 ;
  assign n13898 = \u4_buf1_reg[26]/NET0131  & n5198 ;
  assign n13899 = ~n13897 & ~n13898 ;
  assign n13900 = n13896 & n13899 ;
  assign n13901 = \u4_u2_buf1_reg[27]/P0001  & n5171 ;
  assign n13902 = n5156 & n13901 ;
  assign n13903 = \u4_u1_buf1_reg[27]/P0001  & n5175 ;
  assign n13904 = \u4_u0_buf1_reg[27]/P0001  & n5140 ;
  assign n13905 = ~n13903 & ~n13904 ;
  assign n13906 = ~n13902 & n13905 ;
  assign n13907 = \u4_u3_buf1_reg[27]/P0001  & n5195 ;
  assign n13908 = \u4_buf1_reg[27]/P0001  & n5198 ;
  assign n13909 = ~n13907 & ~n13908 ;
  assign n13910 = n13906 & n13909 ;
  assign n13911 = \u4_u2_buf1_reg[28]/P0001  & n5171 ;
  assign n13912 = n5156 & n13911 ;
  assign n13913 = \u4_u1_buf1_reg[28]/P0001  & n5175 ;
  assign n13914 = \u4_u0_buf1_reg[28]/P0001  & n5140 ;
  assign n13915 = ~n13913 & ~n13914 ;
  assign n13916 = ~n13912 & n13915 ;
  assign n13917 = \u4_u3_buf1_reg[28]/P0001  & n5195 ;
  assign n13918 = \u4_buf1_reg[28]/P0001  & n5198 ;
  assign n13919 = ~n13917 & ~n13918 ;
  assign n13920 = n13916 & n13919 ;
  assign n13921 = \u4_u2_buf1_reg[29]/P0001  & n5171 ;
  assign n13922 = n5156 & n13921 ;
  assign n13923 = \u4_u1_buf1_reg[29]/P0001  & n5175 ;
  assign n13924 = \u4_u0_buf1_reg[29]/P0001  & n5140 ;
  assign n13925 = ~n13923 & ~n13924 ;
  assign n13926 = ~n13922 & n13925 ;
  assign n13927 = \u4_u3_buf1_reg[29]/P0001  & n5195 ;
  assign n13928 = \u4_buf1_reg[29]/P0001  & n5198 ;
  assign n13929 = ~n13927 & ~n13928 ;
  assign n13930 = n13926 & n13929 ;
  assign n13931 = \u4_u2_buf1_reg[2]/P0001  & n5171 ;
  assign n13932 = n5156 & n13931 ;
  assign n13933 = \u4_u1_buf1_reg[2]/P0001  & n5175 ;
  assign n13934 = \u4_u0_buf1_reg[2]/P0001  & n5140 ;
  assign n13935 = ~n13933 & ~n13934 ;
  assign n13936 = ~n13932 & n13935 ;
  assign n13937 = \u4_u3_buf1_reg[2]/P0001  & n5195 ;
  assign n13938 = \u4_buf1_reg[2]/P0001  & n5198 ;
  assign n13939 = ~n13937 & ~n13938 ;
  assign n13940 = n13936 & n13939 ;
  assign n13941 = \u4_u2_buf1_reg[30]/P0001  & n5171 ;
  assign n13942 = n5156 & n13941 ;
  assign n13943 = \u4_u1_buf1_reg[30]/P0001  & n5175 ;
  assign n13944 = \u4_u0_buf1_reg[30]/P0001  & n5140 ;
  assign n13945 = ~n13943 & ~n13944 ;
  assign n13946 = ~n13942 & n13945 ;
  assign n13947 = \u4_u3_buf1_reg[30]/P0001  & n5195 ;
  assign n13948 = \u4_buf1_reg[30]/P0001  & n5198 ;
  assign n13949 = ~n13947 & ~n13948 ;
  assign n13950 = n13946 & n13949 ;
  assign n13951 = \u4_u2_buf1_reg[31]/P0001  & n5171 ;
  assign n13952 = n5156 & n13951 ;
  assign n13953 = \u4_u1_buf1_reg[31]/P0001  & n5175 ;
  assign n13954 = \u4_u0_buf1_reg[31]/P0001  & n5140 ;
  assign n13955 = ~n13953 & ~n13954 ;
  assign n13956 = ~n13952 & n13955 ;
  assign n13957 = \u4_u3_buf1_reg[31]/P0001  & n5195 ;
  assign n13958 = \u4_buf1_reg[31]/P0001  & n5198 ;
  assign n13959 = ~n13957 & ~n13958 ;
  assign n13960 = n13956 & n13959 ;
  assign n13961 = \u4_u2_buf1_reg[4]/P0001  & n5171 ;
  assign n13962 = n5156 & n13961 ;
  assign n13963 = \u4_u1_buf1_reg[4]/P0001  & n5175 ;
  assign n13964 = \u4_u0_buf1_reg[4]/P0001  & n5140 ;
  assign n13965 = ~n13963 & ~n13964 ;
  assign n13966 = ~n13962 & n13965 ;
  assign n13967 = \u4_u3_buf1_reg[4]/P0001  & n5195 ;
  assign n13968 = \u4_buf1_reg[4]/P0001  & n5198 ;
  assign n13969 = ~n13967 & ~n13968 ;
  assign n13970 = n13966 & n13969 ;
  assign n13971 = \u4_u2_buf1_reg[7]/P0001  & n5171 ;
  assign n13972 = n5156 & n13971 ;
  assign n13973 = \u4_u1_buf1_reg[7]/P0001  & n5175 ;
  assign n13974 = \u4_u0_buf1_reg[7]/P0001  & n5140 ;
  assign n13975 = ~n13973 & ~n13974 ;
  assign n13976 = ~n13972 & n13975 ;
  assign n13977 = \u4_u3_buf1_reg[7]/P0001  & n5195 ;
  assign n13978 = \u4_buf1_reg[7]/P0001  & n5198 ;
  assign n13979 = ~n13977 & ~n13978 ;
  assign n13980 = n13976 & n13979 ;
  assign n13981 = \u4_u2_buf1_reg[8]/P0001  & n5171 ;
  assign n13982 = n5156 & n13981 ;
  assign n13983 = \u4_u1_buf1_reg[8]/P0001  & n5175 ;
  assign n13984 = \u4_u0_buf1_reg[8]/P0001  & n5140 ;
  assign n13985 = ~n13983 & ~n13984 ;
  assign n13986 = ~n13982 & n13985 ;
  assign n13987 = \u4_u3_buf1_reg[8]/P0001  & n5195 ;
  assign n13988 = \u4_buf1_reg[8]/P0001  & n5198 ;
  assign n13989 = ~n13987 & ~n13988 ;
  assign n13990 = n13986 & n13989 ;
  assign n13991 = \u4_u2_buf1_reg[9]/P0001  & n5171 ;
  assign n13992 = n5156 & n13991 ;
  assign n13993 = \u4_u1_buf1_reg[9]/P0001  & n5175 ;
  assign n13994 = \u4_u0_buf1_reg[9]/P0001  & n5140 ;
  assign n13995 = ~n13993 & ~n13994 ;
  assign n13996 = ~n13992 & n13995 ;
  assign n13997 = \u4_u3_buf1_reg[9]/P0001  & n5195 ;
  assign n13998 = \u4_buf1_reg[9]/P0001  & n5198 ;
  assign n13999 = ~n13997 & ~n13998 ;
  assign n14000 = n13996 & n13999 ;
  assign n14001 = \u4_u2_csr0_reg[0]/P0001  & n5171 ;
  assign n14002 = n5156 & n14001 ;
  assign n14003 = \u4_u1_csr0_reg[0]/P0001  & n5175 ;
  assign n14004 = \u4_u0_csr0_reg[0]/P0001  & n5140 ;
  assign n14005 = ~n14003 & ~n14004 ;
  assign n14006 = ~n14002 & n14005 ;
  assign n14007 = \u4_u3_csr0_reg[0]/P0001  & n5195 ;
  assign n14008 = \u4_csr_reg[0]/P0001  & n5198 ;
  assign n14009 = ~n14007 & ~n14008 ;
  assign n14010 = n14006 & n14009 ;
  assign n14011 = \u4_u2_csr0_reg[10]/P0001  & n5171 ;
  assign n14012 = n5156 & n14011 ;
  assign n14013 = \u4_u1_csr0_reg[10]/P0001  & n5175 ;
  assign n14014 = \u4_u0_csr0_reg[10]/P0001  & n5140 ;
  assign n14015 = ~n14013 & ~n14014 ;
  assign n14016 = ~n14012 & n14015 ;
  assign n14017 = \u4_u3_csr0_reg[10]/P0001  & n5195 ;
  assign n14018 = \u4_csr_reg[10]/P0001  & n5198 ;
  assign n14019 = ~n14017 & ~n14018 ;
  assign n14020 = n14016 & n14019 ;
  assign n14021 = \u4_u2_csr0_reg[11]/P0001  & n5171 ;
  assign n14022 = n5156 & n14021 ;
  assign n14023 = \u4_u1_csr0_reg[11]/P0001  & n5175 ;
  assign n14024 = \u4_u0_csr0_reg[11]/P0001  & n5140 ;
  assign n14025 = ~n14023 & ~n14024 ;
  assign n14026 = ~n14022 & n14025 ;
  assign n14027 = \u4_u3_csr0_reg[11]/P0001  & n5195 ;
  assign n14028 = \u4_csr_reg[11]/P0001  & n5198 ;
  assign n14029 = ~n14027 & ~n14028 ;
  assign n14030 = n14026 & n14029 ;
  assign n14031 = \u4_u2_csr0_reg[12]/P0001  & n5171 ;
  assign n14032 = n5156 & n14031 ;
  assign n14033 = \u4_u1_csr0_reg[12]/P0001  & n5175 ;
  assign n14034 = \u4_u0_csr0_reg[12]/P0001  & n5140 ;
  assign n14035 = ~n14033 & ~n14034 ;
  assign n14036 = ~n14032 & n14035 ;
  assign n14037 = \u4_u3_csr0_reg[12]/P0001  & n5195 ;
  assign n14038 = \u4_csr_reg[12]/P0001  & n5198 ;
  assign n14039 = ~n14037 & ~n14038 ;
  assign n14040 = n14036 & n14039 ;
  assign n14041 = ~\u1_u2_mack_r_reg/P0001  & ~\u1_u2_state_reg[2]/NET0131  ;
  assign n14042 = ~\u1_u3_abort_reg/P0001  & ~n14041 ;
  assign n14043 = n4106 & n14042 ;
  assign n14044 = ~\u1_u2_rx_data_done_r2_reg/P0001  & \u1_u2_state_reg[2]/NET0131  ;
  assign n14045 = ~\u1_u3_abort_reg/P0001  & n14044 ;
  assign n14046 = n11572 & n14045 ;
  assign n14047 = ~n14043 & ~n14046 ;
  assign n14048 = rst_i_pad & ~n14047 ;
  assign n14049 = n11231 & ~n13034 ;
  assign n14050 = ~n8672 & n14049 ;
  assign n14051 = ~n8666 & n14050 ;
  assign n14052 = ~\u0_u0_chirp_cnt_reg[1]/P0001  & ~n13138 ;
  assign n14053 = ~\u0_u0_chirp_cnt_is_6_reg/P0001  & \u0_u0_chirp_cnt_reg[1]/P0001  ;
  assign n14054 = \u0_u0_chirp_cnt_reg[0]/P0001  & n14053 ;
  assign n14055 = n13134 & n14054 ;
  assign n14056 = ~\u0_u0_state_reg[10]/P0001  & ~n14055 ;
  assign n14057 = ~n14052 & n14056 ;
  assign n14058 = \u0_u0_chirp_cnt_reg[2]/P0001  & ~\u0_u0_state_reg[10]/P0001  ;
  assign n14059 = ~n14055 & n14058 ;
  assign n14060 = ~\u0_u0_chirp_cnt_reg[2]/P0001  & ~\u0_u0_state_reg[10]/P0001  ;
  assign n14061 = n14054 & n14060 ;
  assign n14062 = n13134 & n14061 ;
  assign n14063 = ~n14059 & ~n14062 ;
  assign n14064 = n2564 & n8864 ;
  assign n14065 = n2560 & n14064 ;
  assign n14066 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[0]_pad  ;
  assign n14067 = n8820 & n14066 ;
  assign n14068 = n14065 & n14067 ;
  assign n14069 = rst_i_pad & \u4_funct_adr_reg[0]/P0001  ;
  assign n14070 = ~\wb_addr_i[4]_pad  & n8820 ;
  assign n14071 = rst_i_pad & n2564 ;
  assign n14072 = n8864 & n14071 ;
  assign n14073 = n2560 & n14072 ;
  assign n14074 = n14070 & n14073 ;
  assign n14075 = ~n14069 & ~n14074 ;
  assign n14076 = ~n14068 & ~n14075 ;
  assign n14077 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[1]_pad  ;
  assign n14078 = n8820 & n14077 ;
  assign n14079 = n14065 & n14078 ;
  assign n14080 = rst_i_pad & \u4_funct_adr_reg[1]/P0001  ;
  assign n14081 = ~n14074 & ~n14080 ;
  assign n14082 = ~n14079 & ~n14081 ;
  assign n14083 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[2]_pad  ;
  assign n14084 = n8820 & n14083 ;
  assign n14085 = n14065 & n14084 ;
  assign n14086 = rst_i_pad & \u4_funct_adr_reg[2]/P0001  ;
  assign n14087 = ~n14074 & ~n14086 ;
  assign n14088 = ~n14085 & ~n14087 ;
  assign n14089 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[3]_pad  ;
  assign n14090 = n8820 & n14089 ;
  assign n14091 = n14065 & n14090 ;
  assign n14092 = rst_i_pad & \u4_funct_adr_reg[3]/P0001  ;
  assign n14093 = ~n14074 & ~n14092 ;
  assign n14094 = ~n14091 & ~n14093 ;
  assign n14095 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[4]_pad  ;
  assign n14096 = n8820 & n14095 ;
  assign n14097 = n14065 & n14096 ;
  assign n14098 = rst_i_pad & \u4_funct_adr_reg[4]/P0001  ;
  assign n14099 = ~n14074 & ~n14098 ;
  assign n14100 = ~n14097 & ~n14099 ;
  assign n14101 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[5]_pad  ;
  assign n14102 = n8820 & n14101 ;
  assign n14103 = n14065 & n14102 ;
  assign n14104 = rst_i_pad & \u4_funct_adr_reg[5]/P0001  ;
  assign n14105 = ~n14074 & ~n14104 ;
  assign n14106 = ~n14103 & ~n14105 ;
  assign n14107 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[6]_pad  ;
  assign n14108 = n8820 & n14107 ;
  assign n14109 = n14065 & n14108 ;
  assign n14110 = rst_i_pad & \u4_funct_adr_reg[6]/P0001  ;
  assign n14111 = ~n14074 & ~n14110 ;
  assign n14112 = ~n14109 & ~n14111 ;
  assign n14113 = n2568 & n14066 ;
  assign n14114 = n14065 & n14113 ;
  assign n14115 = rst_i_pad & \u4_inta_msk_reg[0]/P0001  ;
  assign n14116 = ~\wb_addr_i[4]_pad  & n2568 ;
  assign n14117 = n14073 & n14116 ;
  assign n14118 = ~n14115 & ~n14117 ;
  assign n14119 = ~n14114 & ~n14118 ;
  assign n14120 = n2568 & n14077 ;
  assign n14121 = n14065 & n14120 ;
  assign n14122 = rst_i_pad & \u4_inta_msk_reg[1]/P0001  ;
  assign n14123 = ~n14117 & ~n14122 ;
  assign n14124 = ~n14121 & ~n14123 ;
  assign n14125 = n2568 & n14083 ;
  assign n14126 = n14065 & n14125 ;
  assign n14127 = rst_i_pad & \u4_inta_msk_reg[2]/P0001  ;
  assign n14128 = ~n14117 & ~n14127 ;
  assign n14129 = ~n14126 & ~n14128 ;
  assign n14130 = n2568 & n14089 ;
  assign n14131 = n14065 & n14130 ;
  assign n14132 = rst_i_pad & \u4_inta_msk_reg[3]/P0001  ;
  assign n14133 = ~n14117 & ~n14132 ;
  assign n14134 = ~n14131 & ~n14133 ;
  assign n14135 = n2568 & n14095 ;
  assign n14136 = n14065 & n14135 ;
  assign n14137 = rst_i_pad & \u4_inta_msk_reg[4]/P0001  ;
  assign n14138 = ~n14117 & ~n14137 ;
  assign n14139 = ~n14136 & ~n14138 ;
  assign n14140 = n2568 & n14101 ;
  assign n14141 = n14065 & n14140 ;
  assign n14142 = rst_i_pad & \u4_inta_msk_reg[5]/P0001  ;
  assign n14143 = ~n14117 & ~n14142 ;
  assign n14144 = ~n14141 & ~n14143 ;
  assign n14145 = n2568 & n14107 ;
  assign n14146 = n14065 & n14145 ;
  assign n14147 = rst_i_pad & \u4_inta_msk_reg[6]/P0001  ;
  assign n14148 = ~n14117 & ~n14147 ;
  assign n14149 = ~n14146 & ~n14148 ;
  assign n14150 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[7]_pad  ;
  assign n14151 = n2568 & n14150 ;
  assign n14152 = n14065 & n14151 ;
  assign n14153 = rst_i_pad & \u4_inta_msk_reg[7]/P0001  ;
  assign n14154 = ~n14117 & ~n14153 ;
  assign n14155 = ~n14152 & ~n14154 ;
  assign n14156 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[8]_pad  ;
  assign n14157 = n2568 & n14156 ;
  assign n14158 = n14065 & n14157 ;
  assign n14159 = rst_i_pad & \u4_inta_msk_reg[8]/P0001  ;
  assign n14160 = ~n14117 & ~n14159 ;
  assign n14161 = ~n14158 & ~n14160 ;
  assign n14162 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[16]_pad  ;
  assign n14163 = n2568 & n14162 ;
  assign n14164 = n14065 & n14163 ;
  assign n14165 = rst_i_pad & \u4_intb_msk_reg[0]/P0001  ;
  assign n14166 = ~n14117 & ~n14165 ;
  assign n14167 = ~n14164 & ~n14166 ;
  assign n14168 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[17]_pad  ;
  assign n14169 = n2568 & n14168 ;
  assign n14170 = n14065 & n14169 ;
  assign n14171 = rst_i_pad & \u4_intb_msk_reg[1]/P0001  ;
  assign n14172 = ~n14117 & ~n14171 ;
  assign n14173 = ~n14170 & ~n14172 ;
  assign n14174 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[18]_pad  ;
  assign n14175 = n2568 & n14174 ;
  assign n14176 = n14065 & n14175 ;
  assign n14177 = rst_i_pad & \u4_intb_msk_reg[2]/P0001  ;
  assign n14178 = ~n14117 & ~n14177 ;
  assign n14179 = ~n14176 & ~n14178 ;
  assign n14180 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[19]_pad  ;
  assign n14181 = n2568 & n14180 ;
  assign n14182 = n14065 & n14181 ;
  assign n14183 = rst_i_pad & \u4_intb_msk_reg[3]/P0001  ;
  assign n14184 = ~n14117 & ~n14183 ;
  assign n14185 = ~n14182 & ~n14184 ;
  assign n14186 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[20]_pad  ;
  assign n14187 = n2568 & n14186 ;
  assign n14188 = n14065 & n14187 ;
  assign n14189 = rst_i_pad & \u4_intb_msk_reg[4]/P0001  ;
  assign n14190 = ~n14117 & ~n14189 ;
  assign n14191 = ~n14188 & ~n14190 ;
  assign n14192 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[21]_pad  ;
  assign n14193 = n2568 & n14192 ;
  assign n14194 = n14065 & n14193 ;
  assign n14195 = rst_i_pad & \u4_intb_msk_reg[5]/P0001  ;
  assign n14196 = ~n14117 & ~n14195 ;
  assign n14197 = ~n14194 & ~n14196 ;
  assign n14198 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[22]_pad  ;
  assign n14199 = n2568 & n14198 ;
  assign n14200 = n14065 & n14199 ;
  assign n14201 = rst_i_pad & \u4_intb_msk_reg[6]/P0001  ;
  assign n14202 = ~n14117 & ~n14201 ;
  assign n14203 = ~n14200 & ~n14202 ;
  assign n14204 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[23]_pad  ;
  assign n14205 = n2568 & n14204 ;
  assign n14206 = n14065 & n14205 ;
  assign n14207 = rst_i_pad & \u4_intb_msk_reg[7]/P0001  ;
  assign n14208 = ~n14117 & ~n14207 ;
  assign n14209 = ~n14206 & ~n14208 ;
  assign n14210 = ~\wb_addr_i[4]_pad  & ~\wb_data_i[24]_pad  ;
  assign n14211 = n2568 & n14210 ;
  assign n14212 = n14065 & n14211 ;
  assign n14213 = rst_i_pad & \u4_intb_msk_reg[8]/P0001  ;
  assign n14214 = ~n14117 & ~n14213 ;
  assign n14215 = ~n14212 & ~n14214 ;
  assign n14216 = \u1_u3_rx_ack_to_cnt_reg[4]/P0001  & \u1_u3_rx_ack_to_cnt_reg[6]/P0001  ;
  assign n14217 = \u1_u3_rx_ack_to_cnt_reg[5]/P0001  & n14216 ;
  assign n14218 = n12632 & n14217 ;
  assign n14219 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & \u1_u3_rx_ack_to_cnt_reg[7]/P0001  ;
  assign n14220 = ~n14218 & n14219 ;
  assign n14221 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & \u1_u3_rx_ack_to_cnt_reg[5]/P0001  ;
  assign n14222 = n14216 & n14221 ;
  assign n14223 = n12632 & n14222 ;
  assign n14224 = ~\u1_u3_rx_ack_to_cnt_reg[7]/P0001  & n14223 ;
  assign n14225 = ~n14220 & ~n14224 ;
  assign n14226 = \u1_u3_tx_data_to_cnt_reg[4]/P0001  & \u1_u3_tx_data_to_cnt_reg[6]/P0001  ;
  assign n14227 = \u1_u3_tx_data_to_cnt_reg[5]/P0001  & n14226 ;
  assign n14228 = n12665 & n14227 ;
  assign n14229 = ~\u0_rx_active_reg/P0001  & \u1_u3_tx_data_to_cnt_reg[7]/P0001  ;
  assign n14230 = ~n14228 & n14229 ;
  assign n14231 = ~\u0_rx_active_reg/P0001  & \u1_u3_tx_data_to_cnt_reg[5]/P0001  ;
  assign n14232 = n14226 & n14231 ;
  assign n14233 = n12665 & n14232 ;
  assign n14234 = ~\u1_u3_tx_data_to_cnt_reg[7]/P0001  & n14233 ;
  assign n14235 = ~n14230 & ~n14234 ;
  assign n14236 = ~\u4_int_srcb_reg[1]/P0001  & ~\u4_pid_cs_err_r_reg/P0001  ;
  assign n14237 = n5667 & ~n14236 ;
  assign n14238 = ~\u4_int_srcb_reg[7]/P0001  & ~\u4_rx_err_r_reg/P0001  ;
  assign n14239 = n5667 & ~n14238 ;
  assign n14240 = ~\u4_int_srcb_reg[8]/P0001  & ~\u4_usb_reset_r_reg/P0001  ;
  assign n14241 = n5667 & ~n14240 ;
  assign n14242 = n5743 & n5761 ;
  assign n14243 = n5742 & n14242 ;
  assign n14244 = n5757 & n14243 ;
  assign n14245 = \u0_u0_state_reg[13]/NET0131  & ~n5766 ;
  assign n14246 = ~n5760 & n14245 ;
  assign n14247 = ~\u0_u0_chirp_cnt_is_6_reg/P0001  & ~n14246 ;
  assign n14248 = n14244 & ~n14247 ;
  assign n14249 = \u0_u0_state_reg[13]/NET0131  & n12368 ;
  assign n14250 = n12643 & n14249 ;
  assign n14251 = n5746 & n14250 ;
  assign n14252 = ~n5766 & n14251 ;
  assign n14253 = n5743 & n5764 ;
  assign n14254 = n5742 & n14253 ;
  assign n14255 = n5757 & n14254 ;
  assign n14256 = ~n5768 & n14245 ;
  assign n14257 = ~\u0_u0_chirp_cnt_is_6_reg/P0001  & ~n14256 ;
  assign n14258 = n14255 & ~n14257 ;
  assign n14259 = ~n14252 & ~n14258 ;
  assign n14260 = ~n14248 & n14259 ;
  assign n14261 = n5748 & ~n14260 ;
  assign n14262 = ~n5768 & ~n12961 ;
  assign n14263 = n5748 & n6173 ;
  assign n14264 = ~n6192 & n14263 ;
  assign n14265 = n14262 & n14264 ;
  assign n14266 = n12653 & n14265 ;
  assign n14267 = \u0_u0_state_reg[3]/P0001  & n6178 ;
  assign n14268 = ~n6198 & n14267 ;
  assign n14269 = ~n8667 & ~n14268 ;
  assign n14270 = ~n8670 & n14269 ;
  assign n14271 = n5748 & n6132 ;
  assign n14272 = ~n14270 & n14271 ;
  assign n14273 = ~n14266 & ~n14272 ;
  assign n14274 = ~resume_req_i_pad & ~\resume_req_r_reg/P0001  ;
  assign n14275 = rst_i_pad & ~\suspend_clr_wr_reg/P0001  ;
  assign n14276 = ~n14274 & n14275 ;
  assign n14277 = ~n9110 & ~n9149 ;
  assign n14278 = \u4_u0_buf0_orig_reg[30]/NET0131  & ~\u4_u0_dma_out_cnt_reg[11]/P0001  ;
  assign n14279 = ~\u4_u0_buf0_orig_reg[30]/NET0131  & \u4_u0_dma_out_cnt_reg[11]/P0001  ;
  assign n14280 = ~n14278 & ~n14279 ;
  assign n14281 = ~n9148 & n14280 ;
  assign n14282 = ~n14277 & n14281 ;
  assign n14283 = ~n9151 & n14281 ;
  assign n14284 = n9146 & n14283 ;
  assign n14285 = ~n14282 & ~n14284 ;
  assign n14286 = ~n9148 & ~n14277 ;
  assign n14287 = ~n9148 & ~n9151 ;
  assign n14288 = n9146 & n14287 ;
  assign n14289 = ~n14286 & ~n14288 ;
  assign n14290 = ~n14280 & n14289 ;
  assign n14291 = n14285 & ~n14290 ;
  assign n14292 = ~n9061 & ~n9100 ;
  assign n14293 = ~n9097 & n14292 ;
  assign n14294 = ~n9100 & n9102 ;
  assign n14295 = \u4_u3_buf0_orig_reg[30]/NET0131  & ~\u4_u3_dma_out_cnt_reg[11]/P0001  ;
  assign n14296 = ~\u4_u3_buf0_orig_reg[30]/NET0131  & \u4_u3_dma_out_cnt_reg[11]/P0001  ;
  assign n14297 = ~n14295 & ~n14296 ;
  assign n14298 = ~n9099 & n14297 ;
  assign n14299 = ~n14294 & n14298 ;
  assign n14300 = ~n14293 & n14299 ;
  assign n14301 = ~n9099 & ~n14294 ;
  assign n14302 = ~n14293 & n14301 ;
  assign n14303 = ~n14297 & ~n14302 ;
  assign n14304 = ~n14300 & ~n14303 ;
  assign n14305 = \sram_data_i[10]_pad  & \wb_addr_i[17]_pad  ;
  assign n14306 = \u4_dout_reg[10]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n14307 = ~n14305 & ~n14306 ;
  assign n14308 = \sram_data_i[11]_pad  & \wb_addr_i[17]_pad  ;
  assign n14309 = \u4_dout_reg[11]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n14310 = ~n14308 & ~n14309 ;
  assign n14311 = \sram_data_i[9]_pad  & \wb_addr_i[17]_pad  ;
  assign n14312 = \u4_dout_reg[9]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n14313 = ~n14311 & ~n14312 ;
  assign n14314 = \u0_u0_idle_cnt1_reg[2]/P0001  & \u0_u0_idle_cnt1_reg[3]/P0001  ;
  assign n14315 = n11227 & n14314 ;
  assign n14316 = ~\u0_u0_idle_cnt1_reg[4]/P0001  & n14315 ;
  assign n14317 = \u0_u0_idle_cnt1_reg[4]/P0001  & ~n14315 ;
  assign n14318 = ~n14316 & ~n14317 ;
  assign n14319 = ~n9159 & ~n9198 ;
  assign n14320 = ~n9195 & n14319 ;
  assign n14321 = ~n9198 & n9200 ;
  assign n14322 = \u4_u1_buf0_orig_reg[30]/NET0131  & ~\u4_u1_dma_out_cnt_reg[11]/P0001  ;
  assign n14323 = ~\u4_u1_buf0_orig_reg[30]/NET0131  & \u4_u1_dma_out_cnt_reg[11]/P0001  ;
  assign n14324 = ~n14322 & ~n14323 ;
  assign n14325 = ~n9197 & n14324 ;
  assign n14326 = ~n14321 & n14325 ;
  assign n14327 = ~n14320 & n14326 ;
  assign n14328 = ~n9197 & ~n14321 ;
  assign n14329 = ~n14320 & n14328 ;
  assign n14330 = ~n14324 & ~n14329 ;
  assign n14331 = ~n14327 & ~n14330 ;
  assign n14332 = ~n9208 & ~n9247 ;
  assign n14333 = \u4_u2_buf0_orig_reg[30]/NET0131  & ~\u4_u2_dma_out_cnt_reg[11]/P0001  ;
  assign n14334 = ~\u4_u2_buf0_orig_reg[30]/NET0131  & \u4_u2_dma_out_cnt_reg[11]/P0001  ;
  assign n14335 = ~n14333 & ~n14334 ;
  assign n14336 = ~n9246 & n14335 ;
  assign n14337 = ~n14332 & n14336 ;
  assign n14338 = ~n9249 & n14336 ;
  assign n14339 = n9244 & n14338 ;
  assign n14340 = ~n14337 & ~n14339 ;
  assign n14341 = ~n9246 & ~n14332 ;
  assign n14342 = ~n9246 & ~n9249 ;
  assign n14343 = n9244 & n14342 ;
  assign n14344 = ~n14341 & ~n14343 ;
  assign n14345 = ~n14335 & n14344 ;
  assign n14346 = n14340 & ~n14345 ;
  assign n14347 = ~n9214 & ~n9240 ;
  assign n14348 = n9215 & ~n14347 ;
  assign n14349 = n9235 & ~n14347 ;
  assign n14350 = n9232 & n14349 ;
  assign n14351 = ~n14348 & ~n14350 ;
  assign n14352 = n9232 & n9235 ;
  assign n14353 = ~n9215 & n14347 ;
  assign n14354 = ~n14352 & n14353 ;
  assign n14355 = n14351 & ~n14354 ;
  assign n14356 = ~n9067 & ~n9093 ;
  assign n14357 = n9068 & ~n14356 ;
  assign n14358 = n9088 & ~n14356 ;
  assign n14359 = n9085 & n14358 ;
  assign n14360 = ~n14357 & ~n14359 ;
  assign n14361 = n9085 & n9088 ;
  assign n14362 = ~n9068 & n14356 ;
  assign n14363 = ~n14361 & n14362 ;
  assign n14364 = n14360 & ~n14363 ;
  assign n14365 = ~n9116 & ~n9142 ;
  assign n14366 = n9117 & ~n14365 ;
  assign n14367 = n9137 & ~n14365 ;
  assign n14368 = n9134 & n14367 ;
  assign n14369 = ~n14366 & ~n14368 ;
  assign n14370 = n9134 & n9137 ;
  assign n14371 = ~n9117 & n14365 ;
  assign n14372 = ~n14370 & n14371 ;
  assign n14373 = n14369 & ~n14372 ;
  assign n14374 = ~n9165 & ~n9191 ;
  assign n14375 = n9166 & ~n14374 ;
  assign n14376 = n9186 & ~n14374 ;
  assign n14377 = n9183 & n14376 ;
  assign n14378 = ~n14375 & ~n14377 ;
  assign n14379 = n9183 & n9186 ;
  assign n14380 = ~n9166 & n14374 ;
  assign n14381 = ~n14379 & n14380 ;
  assign n14382 = n14378 & ~n14381 ;
  assign n14383 = ~\u1_u3_adr_reg[0]/P0001  & n3483 ;
  assign n14384 = ~n5705 & ~n14383 ;
  assign n14385 = ~\u4_u3_buf0_orig_reg[23]/P0001  & n12411 ;
  assign n14386 = \u4_u3_buf0_orig_reg[23]/P0001  & ~n12411 ;
  assign n14387 = ~n14385 & ~n14386 ;
  assign n14388 = ~\u4_u0_buf0_orig_reg[23]/P0001  & n12441 ;
  assign n14389 = \u4_u0_buf0_orig_reg[23]/P0001  & ~n12441 ;
  assign n14390 = ~n14388 & ~n14389 ;
  assign n14391 = ~\u4_u1_buf0_orig_reg[23]/P0001  & n12464 ;
  assign n14392 = \u4_u1_buf0_orig_reg[23]/P0001  & ~n12464 ;
  assign n14393 = ~n14391 & ~n14392 ;
  assign n14394 = ~\u4_u2_buf0_orig_reg[23]/P0001  & n12487 ;
  assign n14395 = \u4_u2_buf0_orig_reg[23]/P0001  & ~n12487 ;
  assign n14396 = ~n14394 & ~n14395 ;
  assign n14397 = ~\wb_data_i[24]_pad  & n8820 ;
  assign n14398 = n2635 & n14397 ;
  assign n14399 = rst_i_pad & \u4_u2_iena_reg[0]/P0001  ;
  assign n14400 = rst_i_pad & n8820 ;
  assign n14401 = n2635 & n14400 ;
  assign n14402 = ~n14399 & ~n14401 ;
  assign n14403 = ~n14398 & ~n14402 ;
  assign n14404 = ~\wb_data_i[25]_pad  & n8820 ;
  assign n14405 = n2635 & n14404 ;
  assign n14406 = rst_i_pad & \u4_u2_iena_reg[1]/P0001  ;
  assign n14407 = ~n14401 & ~n14406 ;
  assign n14408 = ~n14405 & ~n14407 ;
  assign n14409 = ~\wb_data_i[26]_pad  & n8820 ;
  assign n14410 = n2635 & n14409 ;
  assign n14411 = rst_i_pad & \u4_u2_iena_reg[2]/P0001  ;
  assign n14412 = ~n14401 & ~n14411 ;
  assign n14413 = ~n14410 & ~n14412 ;
  assign n14414 = ~\wb_data_i[27]_pad  & n8820 ;
  assign n14415 = n2635 & n14414 ;
  assign n14416 = rst_i_pad & \u4_u2_iena_reg[3]/P0001  ;
  assign n14417 = ~n14401 & ~n14416 ;
  assign n14418 = ~n14415 & ~n14417 ;
  assign n14419 = ~\wb_data_i[28]_pad  & n8820 ;
  assign n14420 = n2635 & n14419 ;
  assign n14421 = rst_i_pad & \u4_u2_iena_reg[4]/P0001  ;
  assign n14422 = ~n14401 & ~n14421 ;
  assign n14423 = ~n14420 & ~n14422 ;
  assign n14424 = ~\wb_data_i[29]_pad  & n8820 ;
  assign n14425 = n2635 & n14424 ;
  assign n14426 = rst_i_pad & \u4_u2_iena_reg[5]/P0001  ;
  assign n14427 = ~n14401 & ~n14426 ;
  assign n14428 = ~n14425 & ~n14427 ;
  assign n14429 = ~\wb_data_i[16]_pad  & n8820 ;
  assign n14430 = n2635 & n14429 ;
  assign n14431 = rst_i_pad & \u4_u2_ienb_reg[0]/P0001  ;
  assign n14432 = ~n14401 & ~n14431 ;
  assign n14433 = ~n14430 & ~n14432 ;
  assign n14434 = ~\wb_data_i[17]_pad  & n8820 ;
  assign n14435 = n2635 & n14434 ;
  assign n14436 = rst_i_pad & \u4_u2_ienb_reg[1]/P0001  ;
  assign n14437 = ~n14401 & ~n14436 ;
  assign n14438 = ~n14435 & ~n14437 ;
  assign n14439 = ~\wb_data_i[18]_pad  & n8820 ;
  assign n14440 = n2635 & n14439 ;
  assign n14441 = rst_i_pad & \u4_u2_ienb_reg[2]/P0001  ;
  assign n14442 = ~n14401 & ~n14441 ;
  assign n14443 = ~n14440 & ~n14442 ;
  assign n14444 = ~\wb_data_i[19]_pad  & n8820 ;
  assign n14445 = n2635 & n14444 ;
  assign n14446 = rst_i_pad & \u4_u2_ienb_reg[3]/P0001  ;
  assign n14447 = ~n14401 & ~n14446 ;
  assign n14448 = ~n14445 & ~n14447 ;
  assign n14449 = ~\wb_data_i[20]_pad  & n8820 ;
  assign n14450 = n2635 & n14449 ;
  assign n14451 = rst_i_pad & \u4_u2_ienb_reg[4]/P0001  ;
  assign n14452 = ~n14401 & ~n14451 ;
  assign n14453 = ~n14450 & ~n14452 ;
  assign n14454 = ~\wb_data_i[21]_pad  & n8820 ;
  assign n14455 = n2635 & n14454 ;
  assign n14456 = rst_i_pad & \u4_u2_ienb_reg[5]/P0001  ;
  assign n14457 = ~n14401 & ~n14456 ;
  assign n14458 = ~n14455 & ~n14457 ;
  assign n14459 = \u4_u2_int_stat_reg[1]/P0001  & n5451 ;
  assign n14460 = \u4_u2_ep_match_r_reg/P0001  & ~n4912 ;
  assign n14461 = n4911 & n14460 ;
  assign n14462 = n5451 & n14461 ;
  assign n14463 = ~n4935 & n14462 ;
  assign n14464 = ~n14459 & ~n14463 ;
  assign n14465 = ~\wb_data_i[13]_pad  & n8816 ;
  assign n14466 = n2635 & n14465 ;
  assign n14467 = rst_i_pad & \u4_u2_ots_stop_reg/P0001  ;
  assign n14468 = rst_i_pad & n8816 ;
  assign n14469 = n2635 & n14468 ;
  assign n14470 = ~n14467 & ~n14469 ;
  assign n14471 = ~n14466 & ~n14470 ;
  assign n14472 = \u4_u3_buf0_orig_reg[9]/P0001  & ~n2572 ;
  assign n14473 = n11558 & ~n14472 ;
  assign n14474 = \u4_u3_buf0_orig_reg[7]/P0001  & ~n2572 ;
  assign n14475 = n3063 & ~n14474 ;
  assign n14476 = \u4_u3_buf0_orig_reg[0]/P0001  & ~n2572 ;
  assign n14477 = n11316 & ~n14476 ;
  assign n14478 = \u4_u3_buf0_orig_reg[10]/P0001  & ~n2572 ;
  assign n14479 = n2651 & ~n14478 ;
  assign n14480 = \u4_u3_buf0_orig_reg[11]/P0001  & ~n2572 ;
  assign n14481 = n2846 & ~n14480 ;
  assign n14482 = \u4_u3_buf0_orig_reg[12]/P0001  & ~n2572 ;
  assign n14483 = n11327 & ~n14482 ;
  assign n14484 = \u4_u3_buf0_orig_reg[14]/P0001  & ~n2572 ;
  assign n14485 = n2571 & ~n14484 ;
  assign n14486 = \u4_u3_buf0_orig_reg[15]/P0001  & ~n2572 ;
  assign n14487 = n2857 & ~n14486 ;
  assign n14488 = \u4_u3_buf0_orig_reg[16]/P0001  & ~n2572 ;
  assign n14489 = n11338 & ~n14488 ;
  assign n14490 = \u4_u3_buf0_orig_reg[17]/P0001  & ~n2572 ;
  assign n14491 = n11349 & ~n14490 ;
  assign n14492 = \u4_u3_buf0_orig_reg[18]/P0001  & ~n2572 ;
  assign n14493 = n11360 & ~n14492 ;
  assign n14494 = \u4_u3_buf0_orig_reg[19]/P0001  & ~n2572 ;
  assign n14495 = n11371 & ~n14494 ;
  assign n14496 = \u4_u3_buf0_orig_reg[1]/P0001  & ~n2572 ;
  assign n14497 = n11382 & ~n14496 ;
  assign n14498 = \u4_u3_buf0_orig_reg[20]/P0001  & ~n2572 ;
  assign n14499 = n11393 & ~n14498 ;
  assign n14500 = \u4_u3_buf0_orig_reg[22]/P0001  & ~n2572 ;
  assign n14501 = n11415 & ~n14500 ;
  assign n14502 = \u4_u3_buf0_orig_reg[23]/P0001  & ~n2572 ;
  assign n14503 = n11426 & ~n14502 ;
  assign n14504 = \u4_u3_buf0_orig_reg[24]/P0001  & ~n2572 ;
  assign n14505 = n11437 & ~n14504 ;
  assign n14506 = \u4_u3_buf0_orig_reg[25]/P0001  & ~n2572 ;
  assign n14507 = n11448 & ~n14506 ;
  assign n14508 = \u4_u3_buf0_orig_reg[26]/P0001  & ~n2572 ;
  assign n14509 = n11459 & ~n14508 ;
  assign n14510 = \u4_u3_buf0_orig_reg[27]/P0001  & ~n2572 ;
  assign n14511 = n11470 & ~n14510 ;
  assign n14512 = \u4_u3_buf0_orig_reg[28]/P0001  & ~n2572 ;
  assign n14513 = n11481 & ~n14512 ;
  assign n14514 = \u4_u3_buf0_orig_reg[29]/NET0131  & ~n2572 ;
  assign n14515 = n11492 & ~n14514 ;
  assign n14516 = \u4_u3_buf0_orig_reg[2]/P0001  & ~n2572 ;
  assign n14517 = n11503 & ~n14516 ;
  assign n14518 = \u4_u3_buf0_orig_reg[30]/NET0131  & ~n2572 ;
  assign n14519 = n11514 & ~n14518 ;
  assign n14520 = \u4_u3_buf0_orig_reg[31]/P0001  & ~n2572 ;
  assign n14521 = n11525 & ~n14520 ;
  assign n14522 = \u4_u3_buf0_orig_reg[3]/P0001  & ~n2572 ;
  assign n14523 = n11536 & ~n14522 ;
  assign n14524 = \u4_u3_buf0_orig_reg[4]/P0001  & ~n2572 ;
  assign n14525 = n3041 & ~n14524 ;
  assign n14526 = \u4_u3_buf0_orig_reg[5]/P0001  & ~n2572 ;
  assign n14527 = n3052 & ~n14526 ;
  assign n14528 = \u4_u3_buf0_orig_reg[6]/P0001  & ~n2572 ;
  assign n14529 = n2877 & ~n14528 ;
  assign n14530 = ~\wb_data_i[15]_pad  & n8816 ;
  assign n14531 = n2635 & n14530 ;
  assign n14532 = rst_i_pad & \u4_u2_csr1_reg[0]/P0001  ;
  assign n14533 = ~n14469 & ~n14532 ;
  assign n14534 = ~n14531 & ~n14533 ;
  assign n14535 = ~\wb_data_i[0]_pad  & n8816 ;
  assign n14536 = n2567 & n14535 ;
  assign n14537 = rst_i_pad & \u4_u3_csr0_reg[0]/P0001  ;
  assign n14538 = n2567 & n14468 ;
  assign n14539 = ~n14537 & ~n14538 ;
  assign n14540 = ~n14536 & ~n14539 ;
  assign n14541 = ~\wb_data_i[10]_pad  & n8816 ;
  assign n14542 = n2567 & n14541 ;
  assign n14543 = rst_i_pad & \u4_u3_csr0_reg[10]/P0001  ;
  assign n14544 = ~n14538 & ~n14543 ;
  assign n14545 = ~n14542 & ~n14544 ;
  assign n14546 = ~\wb_data_i[11]_pad  & n8816 ;
  assign n14547 = n2567 & n14546 ;
  assign n14548 = rst_i_pad & \u4_u3_csr0_reg[11]/P0001  ;
  assign n14549 = ~n14538 & ~n14548 ;
  assign n14550 = ~n14547 & ~n14549 ;
  assign n14551 = ~\wb_data_i[12]_pad  & n8816 ;
  assign n14552 = n2567 & n14551 ;
  assign n14553 = rst_i_pad & \u4_u3_csr0_reg[12]/P0001  ;
  assign n14554 = ~n14538 & ~n14553 ;
  assign n14555 = ~n14552 & ~n14554 ;
  assign n14556 = ~\wb_data_i[1]_pad  & n8816 ;
  assign n14557 = n2567 & n14556 ;
  assign n14558 = rst_i_pad & \u4_u3_csr0_reg[1]/P0001  ;
  assign n14559 = ~n14538 & ~n14558 ;
  assign n14560 = ~n14557 & ~n14559 ;
  assign n14561 = ~\wb_data_i[2]_pad  & n8816 ;
  assign n14562 = n2567 & n14561 ;
  assign n14563 = rst_i_pad & \u4_u3_csr0_reg[2]/P0001  ;
  assign n14564 = ~n14538 & ~n14563 ;
  assign n14565 = ~n14562 & ~n14564 ;
  assign n14566 = ~\wb_data_i[3]_pad  & n8816 ;
  assign n14567 = n2567 & n14566 ;
  assign n14568 = rst_i_pad & \u4_u3_csr0_reg[3]/NET0131  ;
  assign n14569 = ~n14538 & ~n14568 ;
  assign n14570 = ~n14567 & ~n14569 ;
  assign n14571 = ~\wb_data_i[4]_pad  & n8816 ;
  assign n14572 = n2567 & n14571 ;
  assign n14573 = rst_i_pad & \u4_u3_csr0_reg[4]/P0001  ;
  assign n14574 = ~n14538 & ~n14573 ;
  assign n14575 = ~n14572 & ~n14574 ;
  assign n14576 = ~\wb_data_i[5]_pad  & n8816 ;
  assign n14577 = n2567 & n14576 ;
  assign n14578 = rst_i_pad & \u4_u3_csr0_reg[5]/P0001  ;
  assign n14579 = ~n14538 & ~n14578 ;
  assign n14580 = ~n14577 & ~n14579 ;
  assign n14581 = ~\wb_data_i[6]_pad  & n8816 ;
  assign n14582 = n2567 & n14581 ;
  assign n14583 = rst_i_pad & \u4_u3_csr0_reg[6]/P0001  ;
  assign n14584 = ~n14538 & ~n14583 ;
  assign n14585 = ~n14582 & ~n14584 ;
  assign n14586 = ~\wb_data_i[7]_pad  & n8816 ;
  assign n14587 = n2567 & n14586 ;
  assign n14588 = rst_i_pad & \u4_u3_csr0_reg[7]/P0001  ;
  assign n14589 = ~n14538 & ~n14588 ;
  assign n14590 = ~n14587 & ~n14589 ;
  assign n14591 = ~\wb_data_i[8]_pad  & n8816 ;
  assign n14592 = n2567 & n14591 ;
  assign n14593 = rst_i_pad & \u4_u3_csr0_reg[8]/P0001  ;
  assign n14594 = ~n14538 & ~n14593 ;
  assign n14595 = ~n14592 & ~n14594 ;
  assign n14596 = ~\wb_data_i[9]_pad  & n8816 ;
  assign n14597 = n2567 & n14596 ;
  assign n14598 = rst_i_pad & \u4_u3_csr0_reg[9]/P0001  ;
  assign n14599 = ~n14538 & ~n14598 ;
  assign n14600 = ~n14597 & ~n14599 ;
  assign n14601 = n2567 & n14530 ;
  assign n14602 = rst_i_pad & \u4_u3_csr1_reg[0]/P0001  ;
  assign n14603 = ~n14538 & ~n14602 ;
  assign n14604 = ~n14601 & ~n14603 ;
  assign n14605 = ~\wb_data_i[25]_pad  & n8816 ;
  assign n14606 = n2567 & n14605 ;
  assign n14607 = rst_i_pad & \u4_u3_csr1_reg[10]/P0001  ;
  assign n14608 = ~n14538 & ~n14607 ;
  assign n14609 = ~n14606 & ~n14608 ;
  assign n14610 = ~\wb_data_i[26]_pad  & n8816 ;
  assign n14611 = n2567 & n14610 ;
  assign n14612 = rst_i_pad & \u4_u3_csr1_reg[11]/P0001  ;
  assign n14613 = ~n14538 & ~n14612 ;
  assign n14614 = ~n14611 & ~n14613 ;
  assign n14615 = ~\wb_data_i[27]_pad  & n8816 ;
  assign n14616 = n2567 & n14615 ;
  assign n14617 = rst_i_pad & \u4_u3_csr1_reg[12]/P0001  ;
  assign n14618 = ~n14538 & ~n14617 ;
  assign n14619 = ~n14616 & ~n14618 ;
  assign n14620 = ~\wb_data_i[16]_pad  & n8816 ;
  assign n14621 = n2567 & n14620 ;
  assign n14622 = rst_i_pad & \u4_u3_csr1_reg[1]/P0001  ;
  assign n14623 = ~n14538 & ~n14622 ;
  assign n14624 = ~n14621 & ~n14623 ;
  assign n14625 = ~\wb_data_i[17]_pad  & n8816 ;
  assign n14626 = n2567 & n14625 ;
  assign n14627 = rst_i_pad & \u4_u3_csr1_reg[2]/P0001  ;
  assign n14628 = ~n14538 & ~n14627 ;
  assign n14629 = ~n14626 & ~n14628 ;
  assign n14630 = ~\wb_data_i[18]_pad  & n8816 ;
  assign n14631 = n2567 & n14630 ;
  assign n14632 = rst_i_pad & \u4_u3_csr1_reg[3]/P0001  ;
  assign n14633 = ~n14538 & ~n14632 ;
  assign n14634 = ~n14631 & ~n14633 ;
  assign n14635 = ~\wb_data_i[19]_pad  & n8816 ;
  assign n14636 = n2567 & n14635 ;
  assign n14637 = rst_i_pad & \u4_u3_csr1_reg[4]/P0001  ;
  assign n14638 = ~n14538 & ~n14637 ;
  assign n14639 = ~n14636 & ~n14638 ;
  assign n14640 = ~\wb_data_i[20]_pad  & n8816 ;
  assign n14641 = n2567 & n14640 ;
  assign n14642 = rst_i_pad & \u4_u3_csr1_reg[5]/P0001  ;
  assign n14643 = ~n14538 & ~n14642 ;
  assign n14644 = ~n14641 & ~n14643 ;
  assign n14645 = ~\wb_data_i[21]_pad  & n8816 ;
  assign n14646 = n2567 & n14645 ;
  assign n14647 = rst_i_pad & \u4_u3_csr1_reg[6]/P0001  ;
  assign n14648 = ~n14538 & ~n14647 ;
  assign n14649 = ~n14646 & ~n14648 ;
  assign n14650 = ~\wb_data_i[24]_pad  & n8816 ;
  assign n14651 = n2567 & n14650 ;
  assign n14652 = rst_i_pad & \u4_u3_csr1_reg[9]/P0001  ;
  assign n14653 = ~n14538 & ~n14652 ;
  assign n14654 = ~n14651 & ~n14653 ;
  assign n14655 = \u4_u3_buf0_orig_reg[13]/P0001  & ~n2572 ;
  assign n14656 = n2722 & ~n14655 ;
  assign n14657 = \u4_u1_csr1_reg[7]/P0001  & n8816 ;
  assign n14658 = \u4_u1_buf1_reg[22]/P0001  & n2731 ;
  assign n14659 = \u4_u1_buf0_reg[22]/P0001  & n2568 ;
  assign n14660 = ~n14658 & ~n14659 ;
  assign n14661 = ~n14657 & n14660 ;
  assign n14662 = n8866 & ~n14661 ;
  assign n14663 = \u4_u3_csr1_reg[7]/P0001  & n8816 ;
  assign n14664 = \u4_u3_buf1_reg[22]/P0001  & n2731 ;
  assign n14665 = \u4_u3_buf0_reg[22]/P0001  & n2568 ;
  assign n14666 = ~n14664 & ~n14665 ;
  assign n14667 = ~n14663 & n14666 ;
  assign n14668 = n8836 & ~n14667 ;
  assign n14669 = ~n14662 & ~n14668 ;
  assign n14670 = \u4_u2_csr1_reg[7]/P0001  & n8816 ;
  assign n14671 = \u4_u2_buf1_reg[22]/P0001  & n2731 ;
  assign n14672 = \u4_u2_buf0_reg[22]/P0001  & n2568 ;
  assign n14673 = ~n14671 & ~n14672 ;
  assign n14674 = ~n14670 & n14673 ;
  assign n14675 = n8826 & ~n14674 ;
  assign n14676 = n14669 & ~n14675 ;
  assign n14677 = \u1_frame_no_r_reg[6]/P0001  & \wb_addr_i[4]_pad  ;
  assign n14678 = n8816 & n14677 ;
  assign n14679 = \u4_intb_msk_reg[6]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n14680 = n2568 & n14679 ;
  assign n14681 = \u4_int_srcb_reg[2]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n14682 = n2731 & n14681 ;
  assign n14683 = ~n14680 & ~n14682 ;
  assign n14684 = ~n14678 & n14683 ;
  assign n14685 = n8864 & ~n14684 ;
  assign n14686 = \u4_u0_csr1_reg[7]/P0001  & n8816 ;
  assign n14687 = \u4_u0_buf1_reg[22]/P0001  & n2731 ;
  assign n14688 = \u4_u0_buf0_reg[22]/P0001  & n2568 ;
  assign n14689 = ~n14687 & ~n14688 ;
  assign n14690 = ~n14686 & n14689 ;
  assign n14691 = n8815 & ~n14690 ;
  assign n14692 = ~n14685 & ~n14691 ;
  assign n14693 = n14676 & n14692 ;
  assign n14694 = \u4_u3_buf0_orig_reg[8]/P0001  & ~n2572 ;
  assign n14695 = n11547 & ~n14694 ;
  assign n14696 = n2567 & n14397 ;
  assign n14697 = rst_i_pad & \u4_u3_iena_reg[0]/P0001  ;
  assign n14698 = n2567 & n14400 ;
  assign n14699 = ~n14697 & ~n14698 ;
  assign n14700 = ~n14696 & ~n14699 ;
  assign n14701 = n2567 & n14404 ;
  assign n14702 = rst_i_pad & \u4_u3_iena_reg[1]/P0001  ;
  assign n14703 = ~n14698 & ~n14702 ;
  assign n14704 = ~n14701 & ~n14703 ;
  assign n14705 = n2567 & n14409 ;
  assign n14706 = rst_i_pad & \u4_u3_iena_reg[2]/P0001  ;
  assign n14707 = ~n14698 & ~n14706 ;
  assign n14708 = ~n14705 & ~n14707 ;
  assign n14709 = n2567 & n14414 ;
  assign n14710 = rst_i_pad & \u4_u3_iena_reg[3]/P0001  ;
  assign n14711 = ~n14698 & ~n14710 ;
  assign n14712 = ~n14709 & ~n14711 ;
  assign n14713 = n2567 & n14419 ;
  assign n14714 = rst_i_pad & \u4_u3_iena_reg[4]/P0001  ;
  assign n14715 = ~n14698 & ~n14714 ;
  assign n14716 = ~n14713 & ~n14715 ;
  assign n14717 = n2567 & n14424 ;
  assign n14718 = rst_i_pad & \u4_u3_iena_reg[5]/P0001  ;
  assign n14719 = ~n14698 & ~n14718 ;
  assign n14720 = ~n14717 & ~n14719 ;
  assign n14721 = n2567 & n14429 ;
  assign n14722 = rst_i_pad & \u4_u3_ienb_reg[0]/P0001  ;
  assign n14723 = ~n14698 & ~n14722 ;
  assign n14724 = ~n14721 & ~n14723 ;
  assign n14725 = n2567 & n14439 ;
  assign n14726 = rst_i_pad & \u4_u3_ienb_reg[2]/P0001  ;
  assign n14727 = ~n14698 & ~n14726 ;
  assign n14728 = ~n14725 & ~n14727 ;
  assign n14729 = n2567 & n14444 ;
  assign n14730 = rst_i_pad & \u4_u3_ienb_reg[3]/P0001  ;
  assign n14731 = ~n14698 & ~n14730 ;
  assign n14732 = ~n14729 & ~n14731 ;
  assign n14733 = n2567 & n14434 ;
  assign n14734 = rst_i_pad & \u4_u3_ienb_reg[1]/P0001  ;
  assign n14735 = ~n14698 & ~n14734 ;
  assign n14736 = ~n14733 & ~n14735 ;
  assign n14737 = n2567 & n14449 ;
  assign n14738 = rst_i_pad & \u4_u3_ienb_reg[4]/P0001  ;
  assign n14739 = ~n14698 & ~n14738 ;
  assign n14740 = ~n14737 & ~n14739 ;
  assign n14741 = n2567 & n14454 ;
  assign n14742 = rst_i_pad & \u4_u3_ienb_reg[5]/P0001  ;
  assign n14743 = ~n14698 & ~n14742 ;
  assign n14744 = ~n14741 & ~n14743 ;
  assign n14745 = \u4_u3_int_stat_reg[1]/P0001  & n5455 ;
  assign n14746 = \u4_u3_ep_match_r_reg/P0001  & ~n4912 ;
  assign n14747 = n4911 & n14746 ;
  assign n14748 = n5455 & n14747 ;
  assign n14749 = ~n4935 & n14748 ;
  assign n14750 = ~n14745 & ~n14749 ;
  assign n14751 = n2567 & n14465 ;
  assign n14752 = rst_i_pad & \u4_u3_ots_stop_reg/P0001  ;
  assign n14753 = ~n14538 & ~n14752 ;
  assign n14754 = ~n14751 & ~n14753 ;
  assign n14755 = \u4_u1_csr0_reg[7]/P0001  & n8816 ;
  assign n14756 = \u4_u1_buf1_reg[7]/P0001  & n2731 ;
  assign n14757 = \u4_u1_buf0_reg[7]/P0001  & n2568 ;
  assign n14758 = ~n14756 & ~n14757 ;
  assign n14759 = ~n14755 & n14758 ;
  assign n14760 = n8866 & ~n14759 ;
  assign n14761 = \u4_u3_csr0_reg[7]/P0001  & n8816 ;
  assign n14762 = \u4_u3_buf1_reg[7]/P0001  & n2731 ;
  assign n14763 = \u4_u3_buf0_reg[7]/P0001  & n2568 ;
  assign n14764 = ~n14762 & ~n14763 ;
  assign n14765 = ~n14761 & n14764 ;
  assign n14766 = n8836 & ~n14765 ;
  assign n14767 = ~n14760 & ~n14766 ;
  assign n14768 = \u4_u2_csr0_reg[7]/P0001  & n8816 ;
  assign n14769 = \u4_u2_buf1_reg[7]/P0001  & n2731 ;
  assign n14770 = \u4_u2_buf0_reg[7]/P0001  & n2568 ;
  assign n14771 = ~n14769 & ~n14770 ;
  assign n14772 = ~n14768 & n14771 ;
  assign n14773 = n8826 & ~n14772 ;
  assign n14774 = n14767 & ~n14773 ;
  assign n14775 = \u4_utmi_vend_stat_r_reg[7]/P0001  & \wb_addr_i[4]_pad  ;
  assign n14776 = n8820 & n14775 ;
  assign n14777 = \u4_inta_msk_reg[7]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n14778 = n2568 & n14777 ;
  assign n14779 = \u1_sof_time_reg[7]/P0001  & \wb_addr_i[4]_pad  ;
  assign n14780 = n8816 & n14779 ;
  assign n14781 = ~n14778 & ~n14780 ;
  assign n14782 = ~n14776 & n14781 ;
  assign n14783 = n8864 & ~n14782 ;
  assign n14784 = \u4_u0_csr0_reg[7]/P0001  & n8816 ;
  assign n14785 = \u4_u0_buf1_reg[7]/P0001  & n2731 ;
  assign n14786 = \u4_u0_buf0_reg[7]/P0001  & n2568 ;
  assign n14787 = ~n14785 & ~n14786 ;
  assign n14788 = ~n14784 & n14787 ;
  assign n14789 = n8815 & ~n14788 ;
  assign n14790 = ~n14783 & ~n14789 ;
  assign n14791 = n14774 & n14790 ;
  assign n14792 = \u4_u0_buf0_orig_reg[0]/P0001  & ~n2590 ;
  assign n14793 = n11580 & ~n14792 ;
  assign n14794 = \u4_u0_buf0_orig_reg[10]/P0001  & ~n2590 ;
  assign n14795 = n2661 & ~n14794 ;
  assign n14796 = \u4_u0_buf0_orig_reg[11]/P0001  & ~n2590 ;
  assign n14797 = n2887 & ~n14796 ;
  assign n14798 = \u4_u0_buf0_orig_reg[12]/P0001  & ~n2590 ;
  assign n14799 = n11590 & ~n14798 ;
  assign n14800 = \u4_u0_buf0_orig_reg[13]/P0001  & ~n2590 ;
  assign n14801 = n2745 & ~n14800 ;
  assign n14802 = \u4_u0_buf0_orig_reg[14]/P0001  & ~n2590 ;
  assign n14803 = n2589 & ~n14802 ;
  assign n14804 = \u4_u0_buf0_orig_reg[15]/P0001  & ~n2590 ;
  assign n14805 = n2897 & ~n14804 ;
  assign n14806 = \u4_u0_buf0_orig_reg[16]/P0001  & ~n2590 ;
  assign n14807 = n11600 & ~n14806 ;
  assign n14808 = \u4_u0_buf0_orig_reg[17]/P0001  & ~n2590 ;
  assign n14809 = n11610 & ~n14808 ;
  assign n14810 = \u4_u0_buf0_orig_reg[18]/P0001  & ~n2590 ;
  assign n14811 = n11620 & ~n14810 ;
  assign n14812 = \u4_u0_buf0_orig_reg[19]/P0001  & ~n2590 ;
  assign n14813 = n11630 & ~n14812 ;
  assign n14814 = \u4_u0_buf0_orig_reg[1]/P0001  & ~n2590 ;
  assign n14815 = n11640 & ~n14814 ;
  assign n14816 = \u4_u0_buf0_orig_reg[20]/P0001  & ~n2590 ;
  assign n14817 = n11650 & ~n14816 ;
  assign n14818 = \u4_u0_buf0_orig_reg[21]/P0001  & ~n2590 ;
  assign n14819 = n11660 & ~n14818 ;
  assign n14820 = \u4_u0_buf0_orig_reg[22]/P0001  & ~n2590 ;
  assign n14821 = n11670 & ~n14820 ;
  assign n14822 = \u4_u0_buf0_orig_reg[23]/P0001  & ~n2590 ;
  assign n14823 = n11680 & ~n14822 ;
  assign n14824 = \u4_u0_buf0_orig_reg[24]/P0001  & ~n2590 ;
  assign n14825 = n11690 & ~n14824 ;
  assign n14826 = \u4_u0_buf0_orig_reg[25]/P0001  & ~n2590 ;
  assign n14827 = n11700 & ~n14826 ;
  assign n14828 = \u4_u0_buf0_orig_reg[26]/P0001  & ~n2590 ;
  assign n14829 = n11710 & ~n14828 ;
  assign n14830 = \u4_u0_buf0_orig_reg[27]/P0001  & ~n2590 ;
  assign n14831 = n11720 & ~n14830 ;
  assign n14832 = \u4_u0_buf0_orig_reg[28]/P0001  & ~n2590 ;
  assign n14833 = n11730 & ~n14832 ;
  assign n14834 = \u4_u0_buf0_orig_reg[29]/NET0131  & ~n2590 ;
  assign n14835 = n11740 & ~n14834 ;
  assign n14836 = \u4_u0_buf0_orig_reg[2]/P0001  & ~n2590 ;
  assign n14837 = n11750 & ~n14836 ;
  assign n14838 = \u4_u0_buf0_orig_reg[30]/NET0131  & ~n2590 ;
  assign n14839 = n11760 & ~n14838 ;
  assign n14840 = \u4_u0_buf0_orig_reg[31]/P0001  & ~n2590 ;
  assign n14841 = n11770 & ~n14840 ;
  assign n14842 = \u4_u0_buf0_orig_reg[3]/P0001  & ~n2590 ;
  assign n14843 = n11780 & ~n14842 ;
  assign n14844 = \u4_u0_buf0_orig_reg[4]/P0001  & ~n2590 ;
  assign n14845 = n3100 & ~n14844 ;
  assign n14846 = \u4_u0_buf0_orig_reg[5]/P0001  & ~n2590 ;
  assign n14847 = n3110 & ~n14846 ;
  assign n14848 = \u4_u0_buf0_orig_reg[6]/P0001  & ~n2590 ;
  assign n14849 = n2907 & ~n14848 ;
  assign n14850 = \u4_u0_buf0_orig_reg[7]/P0001  & ~n2590 ;
  assign n14851 = n3120 & ~n14850 ;
  assign n14852 = \u4_u0_buf0_orig_reg[8]/P0001  & ~n2590 ;
  assign n14853 = n11790 & ~n14852 ;
  assign n14854 = \u4_u0_buf0_orig_reg[9]/P0001  & ~n2590 ;
  assign n14855 = n11800 & ~n14854 ;
  assign n14856 = \u4_u1_csr1_reg[8]/P0001  & n8816 ;
  assign n14857 = \u4_u1_buf1_reg[23]/P0001  & n2731 ;
  assign n14858 = \u4_u1_buf0_reg[23]/P0001  & n2568 ;
  assign n14859 = ~n14857 & ~n14858 ;
  assign n14860 = ~n14856 & n14859 ;
  assign n14861 = n8866 & ~n14860 ;
  assign n14862 = \u4_u2_csr1_reg[8]/P0001  & n8816 ;
  assign n14863 = \u4_u2_buf1_reg[23]/P0001  & n2731 ;
  assign n14864 = \u4_u2_buf0_reg[23]/P0001  & n2568 ;
  assign n14865 = ~n14863 & ~n14864 ;
  assign n14866 = ~n14862 & n14865 ;
  assign n14867 = n8826 & ~n14866 ;
  assign n14868 = ~n14861 & ~n14867 ;
  assign n14869 = \u4_u3_csr1_reg[8]/P0001  & n8816 ;
  assign n14870 = \u4_u3_buf1_reg[23]/P0001  & n2731 ;
  assign n14871 = \u4_u3_buf0_reg[23]/P0001  & n2568 ;
  assign n14872 = ~n14870 & ~n14871 ;
  assign n14873 = ~n14869 & n14872 ;
  assign n14874 = n8836 & ~n14873 ;
  assign n14875 = n14868 & ~n14874 ;
  assign n14876 = \u1_frame_no_r_reg[7]/P0001  & \wb_addr_i[4]_pad  ;
  assign n14877 = n8816 & n14876 ;
  assign n14878 = \u4_intb_msk_reg[7]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n14879 = n2568 & n14878 ;
  assign n14880 = \u4_int_srcb_reg[3]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n14881 = n2731 & n14880 ;
  assign n14882 = ~n14879 & ~n14881 ;
  assign n14883 = ~n14877 & n14882 ;
  assign n14884 = n8864 & ~n14883 ;
  assign n14885 = \u4_u0_csr1_reg[8]/P0001  & n8816 ;
  assign n14886 = \u4_u0_buf1_reg[23]/P0001  & n2731 ;
  assign n14887 = \u4_u0_buf0_reg[23]/P0001  & n2568 ;
  assign n14888 = ~n14886 & ~n14887 ;
  assign n14889 = ~n14885 & n14888 ;
  assign n14890 = n8815 & ~n14889 ;
  assign n14891 = ~n14884 & ~n14890 ;
  assign n14892 = n14875 & n14891 ;
  assign n14893 = ~\u0_rx_err_reg/P0001  & \u1_u0_rxv2_reg/P0001  ;
  assign n14894 = n7202 & n14893 ;
  assign n14895 = ~n10520 & n14894 ;
  assign n14896 = n2587 & n14535 ;
  assign n14897 = rst_i_pad & \u4_u0_csr0_reg[0]/P0001  ;
  assign n14898 = n2587 & n14468 ;
  assign n14899 = ~n14897 & ~n14898 ;
  assign n14900 = ~n14896 & ~n14899 ;
  assign n14901 = n2587 & n14541 ;
  assign n14902 = rst_i_pad & \u4_u0_csr0_reg[10]/P0001  ;
  assign n14903 = ~n14898 & ~n14902 ;
  assign n14904 = ~n14901 & ~n14903 ;
  assign n14905 = n2587 & n14546 ;
  assign n14906 = rst_i_pad & \u4_u0_csr0_reg[11]/P0001  ;
  assign n14907 = ~n14898 & ~n14906 ;
  assign n14908 = ~n14905 & ~n14907 ;
  assign n14909 = n2587 & n14551 ;
  assign n14910 = rst_i_pad & \u4_u0_csr0_reg[12]/P0001  ;
  assign n14911 = ~n14898 & ~n14910 ;
  assign n14912 = ~n14909 & ~n14911 ;
  assign n14913 = n2587 & n14556 ;
  assign n14914 = rst_i_pad & \u4_u0_csr0_reg[1]/P0001  ;
  assign n14915 = ~n14898 & ~n14914 ;
  assign n14916 = ~n14913 & ~n14915 ;
  assign n14917 = n2587 & n14561 ;
  assign n14918 = rst_i_pad & \u4_u0_csr0_reg[2]/P0001  ;
  assign n14919 = ~n14898 & ~n14918 ;
  assign n14920 = ~n14917 & ~n14919 ;
  assign n14921 = n2587 & n14566 ;
  assign n14922 = rst_i_pad & \u4_u0_csr0_reg[3]/NET0131  ;
  assign n14923 = ~n14898 & ~n14922 ;
  assign n14924 = ~n14921 & ~n14923 ;
  assign n14925 = n2587 & n14571 ;
  assign n14926 = rst_i_pad & \u4_u0_csr0_reg[4]/P0001  ;
  assign n14927 = ~n14898 & ~n14926 ;
  assign n14928 = ~n14925 & ~n14927 ;
  assign n14929 = n2587 & n14576 ;
  assign n14930 = rst_i_pad & \u4_u0_csr0_reg[5]/P0001  ;
  assign n14931 = ~n14898 & ~n14930 ;
  assign n14932 = ~n14929 & ~n14931 ;
  assign n14933 = n2587 & n14581 ;
  assign n14934 = rst_i_pad & \u4_u0_csr0_reg[6]/P0001  ;
  assign n14935 = ~n14898 & ~n14934 ;
  assign n14936 = ~n14933 & ~n14935 ;
  assign n14937 = n2587 & n14586 ;
  assign n14938 = rst_i_pad & \u4_u0_csr0_reg[7]/P0001  ;
  assign n14939 = ~n14898 & ~n14938 ;
  assign n14940 = ~n14937 & ~n14939 ;
  assign n14941 = n2587 & n14591 ;
  assign n14942 = rst_i_pad & \u4_u0_csr0_reg[8]/P0001  ;
  assign n14943 = ~n14898 & ~n14942 ;
  assign n14944 = ~n14941 & ~n14943 ;
  assign n14945 = n2587 & n14596 ;
  assign n14946 = rst_i_pad & \u4_u0_csr0_reg[9]/P0001  ;
  assign n14947 = ~n14898 & ~n14946 ;
  assign n14948 = ~n14945 & ~n14947 ;
  assign n14949 = n2587 & n14530 ;
  assign n14950 = rst_i_pad & \u4_u0_csr1_reg[0]/P0001  ;
  assign n14951 = ~n14898 & ~n14950 ;
  assign n14952 = ~n14949 & ~n14951 ;
  assign n14953 = n2587 & n14605 ;
  assign n14954 = rst_i_pad & \u4_u0_csr1_reg[10]/P0001  ;
  assign n14955 = ~n14898 & ~n14954 ;
  assign n14956 = ~n14953 & ~n14955 ;
  assign n14957 = n2587 & n14610 ;
  assign n14958 = rst_i_pad & \u4_u0_csr1_reg[11]/P0001  ;
  assign n14959 = ~n14898 & ~n14958 ;
  assign n14960 = ~n14957 & ~n14959 ;
  assign n14961 = n2587 & n14615 ;
  assign n14962 = rst_i_pad & \u4_u0_csr1_reg[12]/P0001  ;
  assign n14963 = ~n14898 & ~n14962 ;
  assign n14964 = ~n14961 & ~n14963 ;
  assign n14965 = n2587 & n14620 ;
  assign n14966 = rst_i_pad & \u4_u0_csr1_reg[1]/P0001  ;
  assign n14967 = ~n14898 & ~n14966 ;
  assign n14968 = ~n14965 & ~n14967 ;
  assign n14969 = n2587 & n14625 ;
  assign n14970 = rst_i_pad & \u4_u0_csr1_reg[2]/P0001  ;
  assign n14971 = ~n14898 & ~n14970 ;
  assign n14972 = ~n14969 & ~n14971 ;
  assign n14973 = n2587 & n14630 ;
  assign n14974 = rst_i_pad & \u4_u0_csr1_reg[3]/P0001  ;
  assign n14975 = ~n14898 & ~n14974 ;
  assign n14976 = ~n14973 & ~n14975 ;
  assign n14977 = n2587 & n14635 ;
  assign n14978 = rst_i_pad & \u4_u0_csr1_reg[4]/P0001  ;
  assign n14979 = ~n14898 & ~n14978 ;
  assign n14980 = ~n14977 & ~n14979 ;
  assign n14981 = n2587 & n14640 ;
  assign n14982 = rst_i_pad & \u4_u0_csr1_reg[5]/P0001  ;
  assign n14983 = ~n14898 & ~n14982 ;
  assign n14984 = ~n14981 & ~n14983 ;
  assign n14985 = n2587 & n14645 ;
  assign n14986 = rst_i_pad & \u4_u0_csr1_reg[6]/P0001  ;
  assign n14987 = ~n14898 & ~n14986 ;
  assign n14988 = ~n14985 & ~n14987 ;
  assign n14989 = n2587 & n14650 ;
  assign n14990 = rst_i_pad & \u4_u0_csr1_reg[9]/P0001  ;
  assign n14991 = ~n14898 & ~n14990 ;
  assign n14992 = ~n14989 & ~n14991 ;
  assign n14993 = \u4_u3_buf0_orig_reg[21]/P0001  & ~n2572 ;
  assign n14994 = n11404 & ~n14993 ;
  assign n14995 = n2587 & n14397 ;
  assign n14996 = rst_i_pad & \u4_u0_iena_reg[0]/P0001  ;
  assign n14997 = n2587 & n14400 ;
  assign n14998 = ~n14996 & ~n14997 ;
  assign n14999 = ~n14995 & ~n14998 ;
  assign n15000 = n2587 & n14404 ;
  assign n15001 = rst_i_pad & \u4_u0_iena_reg[1]/P0001  ;
  assign n15002 = ~n14997 & ~n15001 ;
  assign n15003 = ~n15000 & ~n15002 ;
  assign n15004 = n2587 & n14409 ;
  assign n15005 = rst_i_pad & \u4_u0_iena_reg[2]/P0001  ;
  assign n15006 = ~n14997 & ~n15005 ;
  assign n15007 = ~n15004 & ~n15006 ;
  assign n15008 = n2587 & n14414 ;
  assign n15009 = rst_i_pad & \u4_u0_iena_reg[3]/P0001  ;
  assign n15010 = ~n14997 & ~n15009 ;
  assign n15011 = ~n15008 & ~n15010 ;
  assign n15012 = n2587 & n14419 ;
  assign n15013 = rst_i_pad & \u4_u0_iena_reg[4]/P0001  ;
  assign n15014 = ~n14997 & ~n15013 ;
  assign n15015 = ~n15012 & ~n15014 ;
  assign n15016 = n2587 & n14424 ;
  assign n15017 = rst_i_pad & \u4_u0_iena_reg[5]/P0001  ;
  assign n15018 = ~n14997 & ~n15017 ;
  assign n15019 = ~n15016 & ~n15018 ;
  assign n15020 = n2587 & n14429 ;
  assign n15021 = rst_i_pad & \u4_u0_ienb_reg[0]/P0001  ;
  assign n15022 = ~n14997 & ~n15021 ;
  assign n15023 = ~n15020 & ~n15022 ;
  assign n15024 = n2587 & n14434 ;
  assign n15025 = rst_i_pad & \u4_u0_ienb_reg[1]/P0001  ;
  assign n15026 = ~n14997 & ~n15025 ;
  assign n15027 = ~n15024 & ~n15026 ;
  assign n15028 = n2587 & n14439 ;
  assign n15029 = rst_i_pad & \u4_u0_ienb_reg[2]/P0001  ;
  assign n15030 = ~n14997 & ~n15029 ;
  assign n15031 = ~n15028 & ~n15030 ;
  assign n15032 = n2587 & n14444 ;
  assign n15033 = rst_i_pad & \u4_u0_ienb_reg[3]/P0001  ;
  assign n15034 = ~n14997 & ~n15033 ;
  assign n15035 = ~n15032 & ~n15034 ;
  assign n15036 = n2587 & n14449 ;
  assign n15037 = rst_i_pad & \u4_u0_ienb_reg[4]/P0001  ;
  assign n15038 = ~n14997 & ~n15037 ;
  assign n15039 = ~n15036 & ~n15038 ;
  assign n15040 = n2587 & n14454 ;
  assign n15041 = rst_i_pad & \u4_u0_ienb_reg[5]/P0001  ;
  assign n15042 = ~n14997 & ~n15041 ;
  assign n15043 = ~n15040 & ~n15042 ;
  assign n15044 = \u4_u0_int_stat_reg[1]/P0001  & n5459 ;
  assign n15045 = \u4_u0_ep_match_r_reg/P0001  & ~n4912 ;
  assign n15046 = n4911 & n15045 ;
  assign n15047 = n5459 & n15046 ;
  assign n15048 = ~n4935 & n15047 ;
  assign n15049 = ~n15044 & ~n15048 ;
  assign n15050 = n2587 & n14465 ;
  assign n15051 = rst_i_pad & \u4_u0_ots_stop_reg/P0001  ;
  assign n15052 = ~n14898 & ~n15051 ;
  assign n15053 = ~n15050 & ~n15052 ;
  assign n15054 = \u4_u1_buf0_orig_reg[0]/P0001  & ~n2623 ;
  assign n15055 = n11820 & ~n15054 ;
  assign n15056 = \u4_u1_buf0_orig_reg[10]/P0001  & ~n2623 ;
  assign n15057 = n2671 & ~n15056 ;
  assign n15058 = \u4_u1_buf0_orig_reg[11]/P0001  & ~n2623 ;
  assign n15059 = n2925 & ~n15058 ;
  assign n15060 = \u4_u1_buf0_orig_reg[12]/P0001  & ~n2623 ;
  assign n15061 = n11830 & ~n15060 ;
  assign n15062 = \u4_u1_buf0_orig_reg[13]/P0001  & ~n2623 ;
  assign n15063 = n2765 & ~n15062 ;
  assign n15064 = \u4_u1_buf0_orig_reg[14]/P0001  & ~n2623 ;
  assign n15065 = n2622 & ~n15064 ;
  assign n15066 = \u4_u1_buf0_orig_reg[15]/P0001  & ~n2623 ;
  assign n15067 = n2935 & ~n15066 ;
  assign n15068 = \u4_u1_buf0_orig_reg[16]/P0001  & ~n2623 ;
  assign n15069 = n11840 & ~n15068 ;
  assign n15070 = \u4_u1_buf0_orig_reg[17]/P0001  & ~n2623 ;
  assign n15071 = n11850 & ~n15070 ;
  assign n15072 = \u4_u1_buf0_orig_reg[18]/P0001  & ~n2623 ;
  assign n15073 = n11860 & ~n15072 ;
  assign n15074 = \u4_u1_buf0_orig_reg[19]/P0001  & ~n2623 ;
  assign n15075 = n11870 & ~n15074 ;
  assign n15076 = \u4_u1_buf0_orig_reg[1]/P0001  & ~n2623 ;
  assign n15077 = n11880 & ~n15076 ;
  assign n15078 = \u4_u1_buf0_orig_reg[20]/P0001  & ~n2623 ;
  assign n15079 = n11890 & ~n15078 ;
  assign n15080 = \u4_u1_buf0_orig_reg[21]/P0001  & ~n2623 ;
  assign n15081 = n11900 & ~n15080 ;
  assign n15082 = \u4_u1_buf0_orig_reg[22]/P0001  & ~n2623 ;
  assign n15083 = n11910 & ~n15082 ;
  assign n15084 = \u4_u1_buf0_orig_reg[23]/P0001  & ~n2623 ;
  assign n15085 = n11920 & ~n15084 ;
  assign n15086 = \u4_u1_buf0_orig_reg[24]/P0001  & ~n2623 ;
  assign n15087 = n11930 & ~n15086 ;
  assign n15088 = \u4_u1_buf0_orig_reg[25]/P0001  & ~n2623 ;
  assign n15089 = n11940 & ~n15088 ;
  assign n15090 = \u4_u1_buf0_orig_reg[26]/P0001  & ~n2623 ;
  assign n15091 = n11950 & ~n15090 ;
  assign n15092 = \u4_u1_buf0_orig_reg[27]/P0001  & ~n2623 ;
  assign n15093 = n11960 & ~n15092 ;
  assign n15094 = \u4_u1_buf0_orig_reg[28]/P0001  & ~n2623 ;
  assign n15095 = n11970 & ~n15094 ;
  assign n15096 = \u4_u1_buf0_orig_reg[29]/NET0131  & ~n2623 ;
  assign n15097 = n11980 & ~n15096 ;
  assign n15098 = \u4_u1_buf0_orig_reg[2]/P0001  & ~n2623 ;
  assign n15099 = n11990 & ~n15098 ;
  assign n15100 = \u4_u1_buf0_orig_reg[30]/NET0131  & ~n2623 ;
  assign n15101 = n12000 & ~n15100 ;
  assign n15102 = \u4_u1_buf0_orig_reg[31]/P0001  & ~n2623 ;
  assign n15103 = n12010 & ~n15102 ;
  assign n15104 = \u4_u1_buf0_orig_reg[3]/P0001  & ~n2623 ;
  assign n15105 = n12020 & ~n15104 ;
  assign n15106 = \u4_u1_buf0_orig_reg[4]/P0001  & ~n2623 ;
  assign n15107 = n3154 & ~n15106 ;
  assign n15108 = \u4_u1_buf0_orig_reg[5]/P0001  & ~n2623 ;
  assign n15109 = n3164 & ~n15108 ;
  assign n15110 = \u4_u1_buf0_orig_reg[6]/P0001  & ~n2623 ;
  assign n15111 = n2953 & ~n15110 ;
  assign n15112 = \u4_u1_buf0_orig_reg[7]/P0001  & ~n2623 ;
  assign n15113 = n3174 & ~n15112 ;
  assign n15114 = \u4_u1_buf0_orig_reg[8]/P0001  & ~n2623 ;
  assign n15115 = n12030 & ~n15114 ;
  assign n15116 = \u4_u1_buf0_orig_reg[9]/P0001  & ~n2623 ;
  assign n15117 = n12040 & ~n15116 ;
  assign n15118 = ~\u1_u2_word_done_r_reg/P0001  & ~n8180 ;
  assign n15119 = n2620 & n14535 ;
  assign n15120 = rst_i_pad & \u4_u1_csr0_reg[0]/P0001  ;
  assign n15121 = n2620 & n14468 ;
  assign n15122 = ~n15120 & ~n15121 ;
  assign n15123 = ~n15119 & ~n15122 ;
  assign n15124 = n2620 & n14541 ;
  assign n15125 = rst_i_pad & \u4_u1_csr0_reg[10]/P0001  ;
  assign n15126 = ~n15121 & ~n15125 ;
  assign n15127 = ~n15124 & ~n15126 ;
  assign n15128 = n2620 & n14546 ;
  assign n15129 = rst_i_pad & \u4_u1_csr0_reg[11]/P0001  ;
  assign n15130 = ~n15121 & ~n15129 ;
  assign n15131 = ~n15128 & ~n15130 ;
  assign n15132 = n2620 & n14551 ;
  assign n15133 = rst_i_pad & \u4_u1_csr0_reg[12]/P0001  ;
  assign n15134 = ~n15121 & ~n15133 ;
  assign n15135 = ~n15132 & ~n15134 ;
  assign n15136 = n2620 & n14556 ;
  assign n15137 = rst_i_pad & \u4_u1_csr0_reg[1]/P0001  ;
  assign n15138 = ~n15121 & ~n15137 ;
  assign n15139 = ~n15136 & ~n15138 ;
  assign n15140 = n2620 & n14561 ;
  assign n15141 = rst_i_pad & \u4_u1_csr0_reg[2]/P0001  ;
  assign n15142 = ~n15121 & ~n15141 ;
  assign n15143 = ~n15140 & ~n15142 ;
  assign n15144 = n2620 & n14566 ;
  assign n15145 = rst_i_pad & \u4_u1_csr0_reg[3]/NET0131  ;
  assign n15146 = ~n15121 & ~n15145 ;
  assign n15147 = ~n15144 & ~n15146 ;
  assign n15148 = \u1_u3_rx_ack_to_cnt_reg[2]/P0001  & n12630 ;
  assign n15149 = ~\u1_u3_rx_ack_to_cnt_reg[3]/P0001  & ~n15148 ;
  assign n15150 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & ~n12632 ;
  assign n15151 = ~n15149 & n15150 ;
  assign n15152 = n2620 & n14571 ;
  assign n15153 = rst_i_pad & \u4_u1_csr0_reg[4]/P0001  ;
  assign n15154 = ~n15121 & ~n15153 ;
  assign n15155 = ~n15152 & ~n15154 ;
  assign n15156 = n2620 & n14576 ;
  assign n15157 = rst_i_pad & \u4_u1_csr0_reg[5]/P0001  ;
  assign n15158 = ~n15121 & ~n15157 ;
  assign n15159 = ~n15156 & ~n15158 ;
  assign n15160 = n2620 & n14581 ;
  assign n15161 = rst_i_pad & \u4_u1_csr0_reg[6]/P0001  ;
  assign n15162 = ~n15121 & ~n15161 ;
  assign n15163 = ~n15160 & ~n15162 ;
  assign n15164 = n2620 & n14586 ;
  assign n15165 = rst_i_pad & \u4_u1_csr0_reg[7]/P0001  ;
  assign n15166 = ~n15121 & ~n15165 ;
  assign n15167 = ~n15164 & ~n15166 ;
  assign n15168 = n2620 & n14591 ;
  assign n15169 = rst_i_pad & \u4_u1_csr0_reg[8]/P0001  ;
  assign n15170 = ~n15121 & ~n15169 ;
  assign n15171 = ~n15168 & ~n15170 ;
  assign n15172 = n2620 & n14596 ;
  assign n15173 = rst_i_pad & \u4_u1_csr0_reg[9]/P0001  ;
  assign n15174 = ~n15121 & ~n15173 ;
  assign n15175 = ~n15172 & ~n15174 ;
  assign n15176 = n2620 & n14530 ;
  assign n15177 = rst_i_pad & \u4_u1_csr1_reg[0]/P0001  ;
  assign n15178 = ~n15121 & ~n15177 ;
  assign n15179 = ~n15176 & ~n15178 ;
  assign n15180 = n2620 & n14605 ;
  assign n15181 = rst_i_pad & \u4_u1_csr1_reg[10]/P0001  ;
  assign n15182 = ~n15121 & ~n15181 ;
  assign n15183 = ~n15180 & ~n15182 ;
  assign n15184 = n2620 & n14610 ;
  assign n15185 = rst_i_pad & \u4_u1_csr1_reg[11]/P0001  ;
  assign n15186 = ~n15121 & ~n15185 ;
  assign n15187 = ~n15184 & ~n15186 ;
  assign n15188 = n2620 & n14615 ;
  assign n15189 = rst_i_pad & \u4_u1_csr1_reg[12]/P0001  ;
  assign n15190 = ~n15121 & ~n15189 ;
  assign n15191 = ~n15188 & ~n15190 ;
  assign n15192 = n2620 & n14620 ;
  assign n15193 = rst_i_pad & \u4_u1_csr1_reg[1]/P0001  ;
  assign n15194 = ~n15121 & ~n15193 ;
  assign n15195 = ~n15192 & ~n15194 ;
  assign n15196 = n2620 & n14625 ;
  assign n15197 = rst_i_pad & \u4_u1_csr1_reg[2]/P0001  ;
  assign n15198 = ~n15121 & ~n15197 ;
  assign n15199 = ~n15196 & ~n15198 ;
  assign n15200 = n2620 & n14630 ;
  assign n15201 = rst_i_pad & \u4_u1_csr1_reg[3]/P0001  ;
  assign n15202 = ~n15121 & ~n15201 ;
  assign n15203 = ~n15200 & ~n15202 ;
  assign n15204 = n2620 & n14635 ;
  assign n15205 = rst_i_pad & \u4_u1_csr1_reg[4]/P0001  ;
  assign n15206 = ~n15121 & ~n15205 ;
  assign n15207 = ~n15204 & ~n15206 ;
  assign n15208 = n2620 & n14640 ;
  assign n15209 = rst_i_pad & \u4_u1_csr1_reg[5]/P0001  ;
  assign n15210 = ~n15121 & ~n15209 ;
  assign n15211 = ~n15208 & ~n15210 ;
  assign n15212 = n2620 & n14645 ;
  assign n15213 = rst_i_pad & \u4_u1_csr1_reg[6]/P0001  ;
  assign n15214 = ~n15121 & ~n15213 ;
  assign n15215 = ~n15212 & ~n15214 ;
  assign n15216 = n2620 & n14650 ;
  assign n15217 = rst_i_pad & \u4_u1_csr1_reg[9]/P0001  ;
  assign n15218 = ~n15121 & ~n15217 ;
  assign n15219 = ~n15216 & ~n15218 ;
  assign n15220 = ~n5760 & ~n5766 ;
  assign n15221 = n5761 & n15220 ;
  assign n15222 = ~n13132 & ~n15221 ;
  assign n15223 = n5758 & n5773 ;
  assign n15224 = ~n15222 & n15223 ;
  assign n15225 = \u1_u3_tx_data_to_cnt_reg[2]/P0001  & n12663 ;
  assign n15226 = ~\u1_u3_tx_data_to_cnt_reg[3]/P0001  & ~n15225 ;
  assign n15227 = ~\u0_rx_active_reg/P0001  & ~n12665 ;
  assign n15228 = ~n15226 & n15227 ;
  assign n15229 = n6173 & ~n6192 ;
  assign n15230 = \u0_u0_state_reg[4]/NET0131  & ~n12961 ;
  assign n15231 = ~n5768 & ~n15230 ;
  assign n15232 = n15229 & ~n15231 ;
  assign n15233 = n12653 & n15232 ;
  assign n15234 = ~n5765 & n6144 ;
  assign n15235 = n6143 & n15234 ;
  assign n15236 = ~\u0_u0_T2_gt_1_0_mS_reg/P0001  & ~\u0_u0_state_reg[4]/NET0131  ;
  assign n15237 = ~\u0_u0_state_reg[10]/P0001  & \u0_u0_state_reg[7]/NET0131  ;
  assign n15238 = n5736 & n15237 ;
  assign n15239 = n5735 & n15238 ;
  assign n15240 = n5746 & n15239 ;
  assign n15241 = ~n15236 & n15240 ;
  assign n15242 = ~n15235 & ~n15241 ;
  assign n15243 = ~n15233 & n15242 ;
  assign n15244 = n5748 & ~n15243 ;
  assign n15245 = n2620 & n14397 ;
  assign n15246 = rst_i_pad & \u4_u1_iena_reg[0]/P0001  ;
  assign n15247 = n2620 & n14400 ;
  assign n15248 = ~n15246 & ~n15247 ;
  assign n15249 = ~n15245 & ~n15248 ;
  assign n15250 = n2620 & n14404 ;
  assign n15251 = rst_i_pad & \u4_u1_iena_reg[1]/P0001  ;
  assign n15252 = ~n15247 & ~n15251 ;
  assign n15253 = ~n15250 & ~n15252 ;
  assign n15254 = n2620 & n14409 ;
  assign n15255 = rst_i_pad & \u4_u1_iena_reg[2]/P0001  ;
  assign n15256 = ~n15247 & ~n15255 ;
  assign n15257 = ~n15254 & ~n15256 ;
  assign n15258 = n2620 & n14414 ;
  assign n15259 = rst_i_pad & \u4_u1_iena_reg[3]/P0001  ;
  assign n15260 = ~n15247 & ~n15259 ;
  assign n15261 = ~n15258 & ~n15260 ;
  assign n15262 = n2620 & n14419 ;
  assign n15263 = rst_i_pad & \u4_u1_iena_reg[4]/P0001  ;
  assign n15264 = ~n15247 & ~n15263 ;
  assign n15265 = ~n15262 & ~n15264 ;
  assign n15266 = n2620 & n14424 ;
  assign n15267 = rst_i_pad & \u4_u1_iena_reg[5]/P0001  ;
  assign n15268 = ~n15247 & ~n15267 ;
  assign n15269 = ~n15266 & ~n15268 ;
  assign n15270 = n2620 & n14429 ;
  assign n15271 = rst_i_pad & \u4_u1_ienb_reg[0]/P0001  ;
  assign n15272 = ~n15247 & ~n15271 ;
  assign n15273 = ~n15270 & ~n15272 ;
  assign n15274 = n2620 & n14434 ;
  assign n15275 = rst_i_pad & \u4_u1_ienb_reg[1]/P0001  ;
  assign n15276 = ~n15247 & ~n15275 ;
  assign n15277 = ~n15274 & ~n15276 ;
  assign n15278 = n2620 & n14439 ;
  assign n15279 = rst_i_pad & \u4_u1_ienb_reg[2]/P0001  ;
  assign n15280 = ~n15247 & ~n15279 ;
  assign n15281 = ~n15278 & ~n15280 ;
  assign n15282 = n2620 & n14444 ;
  assign n15283 = rst_i_pad & \u4_u1_ienb_reg[3]/P0001  ;
  assign n15284 = ~n15247 & ~n15283 ;
  assign n15285 = ~n15282 & ~n15284 ;
  assign n15286 = n2620 & n14449 ;
  assign n15287 = rst_i_pad & \u4_u1_ienb_reg[4]/P0001  ;
  assign n15288 = ~n15247 & ~n15287 ;
  assign n15289 = ~n15286 & ~n15288 ;
  assign n15290 = n2620 & n14454 ;
  assign n15291 = rst_i_pad & \u4_u1_ienb_reg[5]/P0001  ;
  assign n15292 = ~n15247 & ~n15291 ;
  assign n15293 = ~n15290 & ~n15292 ;
  assign n15294 = \u4_u1_int_stat_reg[1]/P0001  & n5463 ;
  assign n15295 = \u4_u1_ep_match_r_reg/P0001  & ~n4912 ;
  assign n15296 = n4911 & n15295 ;
  assign n15297 = n5463 & n15296 ;
  assign n15298 = ~n4935 & n15297 ;
  assign n15299 = ~n15294 & ~n15298 ;
  assign n15300 = n2620 & n14465 ;
  assign n15301 = rst_i_pad & \u4_u1_ots_stop_reg/P0001  ;
  assign n15302 = ~n15121 & ~n15301 ;
  assign n15303 = ~n15300 & ~n15302 ;
  assign n15304 = \u4_u2_buf0_orig_reg[0]/P0001  & ~n2638 ;
  assign n15305 = n12054 & ~n15304 ;
  assign n15306 = \u4_u2_buf0_orig_reg[10]/P0001  & ~n2638 ;
  assign n15307 = n2681 & ~n15306 ;
  assign n15308 = \u4_u2_buf0_orig_reg[11]/P0001  & ~n2638 ;
  assign n15309 = n2963 & ~n15308 ;
  assign n15310 = \u4_u2_buf0_orig_reg[12]/P0001  & ~n2638 ;
  assign n15311 = n12064 & ~n15310 ;
  assign n15312 = \u4_u2_buf0_orig_reg[13]/P0001  & ~n2638 ;
  assign n15313 = n2801 & ~n15312 ;
  assign n15314 = \u4_u2_buf0_orig_reg[14]/P0001  & ~n2638 ;
  assign n15315 = n2637 & ~n15314 ;
  assign n15316 = \u4_u2_buf0_orig_reg[15]/P0001  & ~n2638 ;
  assign n15317 = n2973 & ~n15316 ;
  assign n15318 = \u4_u2_buf0_orig_reg[16]/P0001  & ~n2638 ;
  assign n15319 = n12074 & ~n15318 ;
  assign n15320 = \u4_u2_buf0_orig_reg[17]/P0001  & ~n2638 ;
  assign n15321 = n12084 & ~n15320 ;
  assign n15322 = \u4_u2_buf0_orig_reg[18]/P0001  & ~n2638 ;
  assign n15323 = n12094 & ~n15322 ;
  assign n15324 = \u4_u2_buf0_orig_reg[19]/P0001  & ~n2638 ;
  assign n15325 = n12104 & ~n15324 ;
  assign n15326 = \u4_u2_buf0_orig_reg[1]/P0001  & ~n2638 ;
  assign n15327 = n12114 & ~n15326 ;
  assign n15328 = \u4_u2_buf0_orig_reg[20]/P0001  & ~n2638 ;
  assign n15329 = n12124 & ~n15328 ;
  assign n15330 = \u4_u2_buf0_orig_reg[21]/P0001  & ~n2638 ;
  assign n15331 = n12134 & ~n15330 ;
  assign n15332 = \u4_u2_buf0_orig_reg[22]/P0001  & ~n2638 ;
  assign n15333 = n12144 & ~n15332 ;
  assign n15334 = \u4_u2_buf0_orig_reg[23]/P0001  & ~n2638 ;
  assign n15335 = n12154 & ~n15334 ;
  assign n15336 = \u4_u2_buf0_orig_reg[24]/P0001  & ~n2638 ;
  assign n15337 = n12164 & ~n15336 ;
  assign n15338 = \u4_u2_buf0_orig_reg[25]/P0001  & ~n2638 ;
  assign n15339 = n12174 & ~n15338 ;
  assign n15340 = \u4_u2_buf0_orig_reg[26]/P0001  & ~n2638 ;
  assign n15341 = n12184 & ~n15340 ;
  assign n15342 = \u4_u2_buf0_orig_reg[27]/P0001  & ~n2638 ;
  assign n15343 = n12194 & ~n15342 ;
  assign n15344 = \u4_u2_buf0_orig_reg[28]/P0001  & ~n2638 ;
  assign n15345 = n12204 & ~n15344 ;
  assign n15346 = \u4_u2_buf0_orig_reg[29]/NET0131  & ~n2638 ;
  assign n15347 = n12214 & ~n15346 ;
  assign n15348 = \u4_u2_buf0_orig_reg[2]/P0001  & ~n2638 ;
  assign n15349 = n12224 & ~n15348 ;
  assign n15350 = \u4_u2_buf0_orig_reg[30]/NET0131  & ~n2638 ;
  assign n15351 = n12234 & ~n15350 ;
  assign n15352 = \u4_u2_buf0_orig_reg[31]/P0001  & ~n2638 ;
  assign n15353 = n12244 & ~n15352 ;
  assign n15354 = \u4_u2_buf0_orig_reg[3]/P0001  & ~n2638 ;
  assign n15355 = n12254 & ~n15354 ;
  assign n15356 = \u4_u2_buf0_orig_reg[4]/P0001  & ~n2638 ;
  assign n15357 = n3208 & ~n15356 ;
  assign n15358 = \u4_u2_buf0_orig_reg[5]/P0001  & ~n2638 ;
  assign n15359 = n3218 & ~n15358 ;
  assign n15360 = \u4_u2_buf0_orig_reg[6]/P0001  & ~n2638 ;
  assign n15361 = n2991 & ~n15360 ;
  assign n15362 = \u4_u2_buf0_orig_reg[7]/P0001  & ~n2638 ;
  assign n15363 = n3228 & ~n15362 ;
  assign n15364 = \u4_u2_buf0_orig_reg[8]/P0001  & ~n2638 ;
  assign n15365 = n12264 & ~n15364 ;
  assign n15366 = \u4_u2_buf0_orig_reg[9]/P0001  & ~n2638 ;
  assign n15367 = n12274 & ~n15366 ;
  assign n15368 = n2635 & n14535 ;
  assign n15369 = rst_i_pad & \u4_u2_csr0_reg[0]/P0001  ;
  assign n15370 = ~n14469 & ~n15369 ;
  assign n15371 = ~n15368 & ~n15370 ;
  assign n15372 = n2635 & n14541 ;
  assign n15373 = rst_i_pad & \u4_u2_csr0_reg[10]/P0001  ;
  assign n15374 = ~n14469 & ~n15373 ;
  assign n15375 = ~n15372 & ~n15374 ;
  assign n15376 = n2635 & n14546 ;
  assign n15377 = rst_i_pad & \u4_u2_csr0_reg[11]/P0001  ;
  assign n15378 = ~n14469 & ~n15377 ;
  assign n15379 = ~n15376 & ~n15378 ;
  assign n15380 = n2635 & n14551 ;
  assign n15381 = rst_i_pad & \u4_u2_csr0_reg[12]/P0001  ;
  assign n15382 = ~n14469 & ~n15381 ;
  assign n15383 = ~n15380 & ~n15382 ;
  assign n15384 = n2635 & n14556 ;
  assign n15385 = rst_i_pad & \u4_u2_csr0_reg[1]/P0001  ;
  assign n15386 = ~n14469 & ~n15385 ;
  assign n15387 = ~n15384 & ~n15386 ;
  assign n15388 = n2635 & n14561 ;
  assign n15389 = rst_i_pad & \u4_u2_csr0_reg[2]/P0001  ;
  assign n15390 = ~n14469 & ~n15389 ;
  assign n15391 = ~n15388 & ~n15390 ;
  assign n15392 = n2635 & n14566 ;
  assign n15393 = rst_i_pad & \u4_u2_csr0_reg[3]/NET0131  ;
  assign n15394 = ~n14469 & ~n15393 ;
  assign n15395 = ~n15392 & ~n15394 ;
  assign n15396 = n2635 & n14571 ;
  assign n15397 = rst_i_pad & \u4_u2_csr0_reg[4]/P0001  ;
  assign n15398 = ~n14469 & ~n15397 ;
  assign n15399 = ~n15396 & ~n15398 ;
  assign n15400 = n2635 & n14576 ;
  assign n15401 = rst_i_pad & \u4_u2_csr0_reg[5]/P0001  ;
  assign n15402 = ~n14469 & ~n15401 ;
  assign n15403 = ~n15400 & ~n15402 ;
  assign n15404 = n2635 & n14581 ;
  assign n15405 = rst_i_pad & \u4_u2_csr0_reg[6]/P0001  ;
  assign n15406 = ~n14469 & ~n15405 ;
  assign n15407 = ~n15404 & ~n15406 ;
  assign n15408 = n2635 & n14586 ;
  assign n15409 = rst_i_pad & \u4_u2_csr0_reg[7]/P0001  ;
  assign n15410 = ~n14469 & ~n15409 ;
  assign n15411 = ~n15408 & ~n15410 ;
  assign n15412 = n2635 & n14591 ;
  assign n15413 = rst_i_pad & \u4_u2_csr0_reg[8]/P0001  ;
  assign n15414 = ~n14469 & ~n15413 ;
  assign n15415 = ~n15412 & ~n15414 ;
  assign n15416 = n2635 & n14596 ;
  assign n15417 = rst_i_pad & \u4_u2_csr0_reg[9]/P0001  ;
  assign n15418 = ~n14469 & ~n15417 ;
  assign n15419 = ~n15416 & ~n15418 ;
  assign n15420 = n2635 & n14605 ;
  assign n15421 = rst_i_pad & \u4_u2_csr1_reg[10]/P0001  ;
  assign n15422 = ~n14469 & ~n15421 ;
  assign n15423 = ~n15420 & ~n15422 ;
  assign n15424 = n2635 & n14610 ;
  assign n15425 = rst_i_pad & \u4_u2_csr1_reg[11]/P0001  ;
  assign n15426 = ~n14469 & ~n15425 ;
  assign n15427 = ~n15424 & ~n15426 ;
  assign n15428 = n2635 & n14615 ;
  assign n15429 = rst_i_pad & \u4_u2_csr1_reg[12]/P0001  ;
  assign n15430 = ~n14469 & ~n15429 ;
  assign n15431 = ~n15428 & ~n15430 ;
  assign n15432 = n2635 & n14620 ;
  assign n15433 = rst_i_pad & \u4_u2_csr1_reg[1]/P0001  ;
  assign n15434 = ~n14469 & ~n15433 ;
  assign n15435 = ~n15432 & ~n15434 ;
  assign n15436 = n2635 & n14625 ;
  assign n15437 = rst_i_pad & \u4_u2_csr1_reg[2]/P0001  ;
  assign n15438 = ~n14469 & ~n15437 ;
  assign n15439 = ~n15436 & ~n15438 ;
  assign n15440 = n2635 & n14630 ;
  assign n15441 = rst_i_pad & \u4_u2_csr1_reg[3]/P0001  ;
  assign n15442 = ~n14469 & ~n15441 ;
  assign n15443 = ~n15440 & ~n15442 ;
  assign n15444 = n2635 & n14635 ;
  assign n15445 = rst_i_pad & \u4_u2_csr1_reg[4]/P0001  ;
  assign n15446 = ~n14469 & ~n15445 ;
  assign n15447 = ~n15444 & ~n15446 ;
  assign n15448 = n2635 & n14640 ;
  assign n15449 = rst_i_pad & \u4_u2_csr1_reg[5]/P0001  ;
  assign n15450 = ~n14469 & ~n15449 ;
  assign n15451 = ~n15448 & ~n15450 ;
  assign n15452 = n2635 & n14645 ;
  assign n15453 = rst_i_pad & \u4_u2_csr1_reg[6]/P0001  ;
  assign n15454 = ~n14469 & ~n15453 ;
  assign n15455 = ~n15452 & ~n15454 ;
  assign n15456 = n2635 & n14650 ;
  assign n15457 = rst_i_pad & \u4_u2_csr1_reg[9]/P0001  ;
  assign n15458 = ~n14469 & ~n15457 ;
  assign n15459 = ~n15456 & ~n15458 ;
  assign n15460 = n7742 & ~n7749 ;
  assign n15461 = n7726 & n7729 ;
  assign n15462 = n15460 & n15461 ;
  assign n15463 = n7799 & n15462 ;
  assign n15464 = n7733 & n7752 ;
  assign n15465 = n7718 & n15464 ;
  assign n15466 = n7795 & n15465 ;
  assign n15467 = n15463 & n15466 ;
  assign n15468 = ~\u4_csr_reg[26]/NET0131  & \u4_csr_reg[27]/NET0131  ;
  assign n15469 = \u1_u3_state_reg[9]/P0001  & \u4_csr_reg[15]/NET0131  ;
  assign n15470 = n15468 & n15469 ;
  assign n15471 = ~n15467 & n15470 ;
  assign n15472 = \u0_u0_state_reg[14]/P0001  & ~n5760 ;
  assign n15473 = ~n5766 & ~n15472 ;
  assign n15474 = n14244 & ~n15473 ;
  assign n15475 = \u0_u0_state_reg[14]/P0001  & ~n5768 ;
  assign n15476 = ~n5766 & ~n15475 ;
  assign n15477 = n14255 & ~n15476 ;
  assign n15478 = ~n15474 & ~n15477 ;
  assign n15479 = n5773 & ~n15478 ;
  assign n15480 = \u1_u3_out_to_small_reg/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n15481 = ~\u4_u2_int_stat_reg[6]/P0001  & ~n15480 ;
  assign n15482 = n5451 & ~n15481 ;
  assign n15483 = \u1_u3_out_to_small_reg/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n15484 = ~\u4_u0_int_stat_reg[6]/P0001  & ~n15483 ;
  assign n15485 = n5459 & ~n15484 ;
  assign n15486 = \u1_u3_out_to_small_reg/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n15487 = ~\u4_u1_int_stat_reg[6]/P0001  & ~n15486 ;
  assign n15488 = n5463 & ~n15487 ;
  assign n15489 = n2587 & n8816 ;
  assign n15490 = \u1_u3_out_to_small_reg/P0001  & \u4_u0_ots_stop_reg/P0001  ;
  assign n15491 = rst_i_pad & ~n15490 ;
  assign n15492 = \u4_u0_csr1_reg[8]/P0001  & n15491 ;
  assign n15493 = ~n15489 & n15492 ;
  assign n15494 = rst_i_pad & \wb_data_i[23]_pad  ;
  assign n15495 = n8816 & n15494 ;
  assign n15496 = n2587 & n15495 ;
  assign n15497 = ~n15493 & ~n15496 ;
  assign n15498 = ~\u0_u0_usb_suspend_reg/P0001  & n8671 ;
  assign n15499 = \u0_u0_state_reg[3]/P0001  & ~n6192 ;
  assign n15500 = ~n15498 & n15499 ;
  assign n15501 = n12335 & n12341 ;
  assign n15502 = ~\u0_u0_state_reg[0]/NET0131  & ~\u0_u0_state_reg[9]/P0001  ;
  assign n15503 = n5743 & n15502 ;
  assign n15504 = ~n6145 & n15503 ;
  assign n15505 = n15501 & n15504 ;
  assign n15506 = n5734 & n15505 ;
  assign n15507 = ~\u0_u0_state_reg[3]/P0001  & ~n15506 ;
  assign n15508 = ~n6157 & ~n15498 ;
  assign n15509 = n15507 & n15508 ;
  assign n15510 = ~n15500 & ~n15509 ;
  assign n15511 = n2635 & n8816 ;
  assign n15512 = \u1_u3_out_to_small_reg/P0001  & \u4_u2_ots_stop_reg/P0001  ;
  assign n15513 = rst_i_pad & ~n15512 ;
  assign n15514 = \u4_u2_csr1_reg[8]/P0001  & n15513 ;
  assign n15515 = ~n15511 & n15514 ;
  assign n15516 = n2635 & n15495 ;
  assign n15517 = ~n15515 & ~n15516 ;
  assign n15518 = \u4_u0_csr0_reg[4]/P0001  & n8816 ;
  assign n15519 = \u4_u0_buf1_reg[4]/P0001  & n2731 ;
  assign n15520 = ~n15518 & ~n15519 ;
  assign n15521 = \u4_u0_int_stat_reg[4]/P0001  & n8820 ;
  assign n15522 = \u4_u0_buf0_reg[4]/P0001  & n2568 ;
  assign n15523 = ~n15521 & ~n15522 ;
  assign n15524 = n15520 & n15523 ;
  assign n15525 = n8815 & ~n15524 ;
  assign n15526 = \u4_u2_buf0_reg[4]/P0001  & n2568 ;
  assign n15527 = \u4_u2_csr0_reg[4]/P0001  & n8816 ;
  assign n15528 = ~n15526 & ~n15527 ;
  assign n15529 = \u4_u2_buf1_reg[4]/P0001  & n2731 ;
  assign n15530 = \u4_u2_int_stat_reg[4]/P0001  & n8820 ;
  assign n15531 = ~n15529 & ~n15530 ;
  assign n15532 = n15528 & n15531 ;
  assign n15533 = n8826 & ~n15532 ;
  assign n15534 = ~n15525 & ~n15533 ;
  assign n15535 = \u4_u3_csr0_reg[4]/P0001  & n8816 ;
  assign n15536 = \u4_u3_buf1_reg[4]/P0001  & n2731 ;
  assign n15537 = ~n15535 & ~n15536 ;
  assign n15538 = \u4_u3_int_stat_reg[4]/P0001  & n8820 ;
  assign n15539 = \u4_u3_buf0_reg[4]/P0001  & n2568 ;
  assign n15540 = ~n15538 & ~n15539 ;
  assign n15541 = n15537 & n15540 ;
  assign n15542 = n8836 & ~n15541 ;
  assign n15543 = n15534 & ~n15542 ;
  assign n15544 = \u4_funct_adr_reg[4]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n15545 = n8820 & n15544 ;
  assign n15546 = \u4_inta_msk_reg[4]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n15547 = n2568 & n15546 ;
  assign n15548 = ~n15545 & ~n15547 ;
  assign n15549 = \LineState_r_reg[1]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n15550 = n8816 & n15549 ;
  assign n15551 = \u4_utmi_vend_stat_r_reg[4]/P0001  & \wb_addr_i[4]_pad  ;
  assign n15552 = n8820 & n15551 ;
  assign n15553 = \u1_sof_time_reg[4]/P0001  & \wb_addr_i[4]_pad  ;
  assign n15554 = n8816 & n15553 ;
  assign n15555 = ~n15552 & ~n15554 ;
  assign n15556 = ~n15550 & n15555 ;
  assign n15557 = n15548 & n15556 ;
  assign n15558 = n8864 & ~n15557 ;
  assign n15559 = \u4_u1_csr0_reg[4]/P0001  & n8816 ;
  assign n15560 = \u4_u1_buf1_reg[4]/P0001  & n2731 ;
  assign n15561 = ~n15559 & ~n15560 ;
  assign n15562 = \u4_u1_int_stat_reg[4]/P0001  & n8820 ;
  assign n15563 = \u4_u1_buf0_reg[4]/P0001  & n2568 ;
  assign n15564 = ~n15562 & ~n15563 ;
  assign n15565 = n15561 & n15564 ;
  assign n15566 = n8866 & ~n15565 ;
  assign n15567 = ~n15558 & ~n15566 ;
  assign n15568 = n15543 & n15567 ;
  assign n15569 = n2567 & n15495 ;
  assign n15570 = n2567 & n8816 ;
  assign n15571 = \u1_u3_out_to_small_reg/P0001  & \u4_u3_ots_stop_reg/P0001  ;
  assign n15572 = rst_i_pad & ~n15571 ;
  assign n15573 = \u4_u3_csr1_reg[8]/P0001  & n15572 ;
  assign n15574 = ~n15570 & n15573 ;
  assign n15575 = ~n15569 & ~n15574 ;
  assign n15576 = \u0_u0_idle_cnt1_reg[6]/P0001  & \u0_u0_idle_cnt1_reg[7]/P0001  ;
  assign n15577 = n13034 & n15576 ;
  assign n15578 = n14315 & n15577 ;
  assign n15579 = ~n11231 & ~n15578 ;
  assign n15580 = n13034 & n14315 ;
  assign n15581 = ~n11231 & ~n15576 ;
  assign n15582 = \u0_u0_idle_cnt1_reg[6]/P0001  & n15581 ;
  assign n15583 = ~n15580 & n15582 ;
  assign n15584 = n15579 & ~n15583 ;
  assign n15585 = n2620 & n8816 ;
  assign n15586 = \u1_u3_out_to_small_reg/P0001  & \u4_u1_ots_stop_reg/P0001  ;
  assign n15587 = rst_i_pad & ~n15586 ;
  assign n15588 = \u4_u1_csr1_reg[8]/P0001  & n15587 ;
  assign n15589 = ~n15585 & n15588 ;
  assign n15590 = n2620 & n15495 ;
  assign n15591 = ~n15589 & ~n15590 ;
  assign n15592 = rst_i_pad & \wb_data_i[22]_pad  ;
  assign n15593 = n8816 & n15592 ;
  assign n15594 = n2567 & n15593 ;
  assign n15595 = ~\u4_u3_csr1_reg[7]/P0001  & ~n15571 ;
  assign n15596 = rst_i_pad & ~n15595 ;
  assign n15597 = ~n15570 & n15596 ;
  assign n15598 = ~n15594 & ~n15597 ;
  assign n15599 = n2587 & n15593 ;
  assign n15600 = ~\u4_u0_csr1_reg[7]/P0001  & ~n15490 ;
  assign n15601 = rst_i_pad & ~n15600 ;
  assign n15602 = ~n15489 & n15601 ;
  assign n15603 = ~n15599 & ~n15602 ;
  assign n15604 = n2620 & n15593 ;
  assign n15605 = ~\u4_u1_csr1_reg[7]/P0001  & ~n15586 ;
  assign n15606 = rst_i_pad & ~n15605 ;
  assign n15607 = ~n15585 & n15606 ;
  assign n15608 = ~n15604 & ~n15607 ;
  assign n15609 = n2635 & n15593 ;
  assign n15610 = ~\u4_u2_csr1_reg[7]/P0001  & ~n15512 ;
  assign n15611 = rst_i_pad & ~n15610 ;
  assign n15612 = ~n15511 & n15611 ;
  assign n15613 = ~n15609 & ~n15612 ;
  assign n15614 = \sram_data_i[12]_pad  & \wb_addr_i[17]_pad  ;
  assign n15615 = \u4_dout_reg[12]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n15616 = ~n15614 & ~n15615 ;
  assign n15617 = \sram_data_i[13]_pad  & \wb_addr_i[17]_pad  ;
  assign n15618 = \u4_dout_reg[13]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n15619 = ~n15617 & ~n15618 ;
  assign n15620 = \sram_data_i[15]_pad  & \wb_addr_i[17]_pad  ;
  assign n15621 = \u4_dout_reg[15]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n15622 = ~n15620 & ~n15621 ;
  assign n15623 = ~VControl_Load_pad_o_pad & \u4_utmi_vend_wr_r_reg/P0001  ;
  assign n15624 = rst_i_pad & n15623 ;
  assign n15625 = rst_i_pad & \wb_addr_i[4]_pad  ;
  assign n15626 = n8820 & n15625 ;
  assign n15627 = n14065 & n15626 ;
  assign n15628 = ~n15624 & ~n15627 ;
  assign n15629 = \u0_u0_mode_hs_reg/P0001  & n5765 ;
  assign n15630 = ~\u0_u0_mode_hs_reg/P0001  & n5759 ;
  assign n15631 = ~n15629 & ~n15630 ;
  assign n15632 = \u0_u0_idle_long_reg/P0001  & \u0_u0_ls_idle_r_reg/P0001  ;
  assign n15633 = n15631 & ~n15632 ;
  assign n15634 = ~\u0_u0_idle_long_reg/P0001  & ~\u0_u0_ls_idle_r_reg/P0001  ;
  assign n15635 = rst_i_pad & ~n15634 ;
  assign n15636 = ~n15633 & n15635 ;
  assign n15637 = \u4_u0_uc_bsel_reg[1]/P0001  & n8816 ;
  assign n15638 = \u4_u0_buf1_reg[31]/P0001  & n2731 ;
  assign n15639 = \u4_u0_buf0_reg[31]/P0001  & n2568 ;
  assign n15640 = ~n15638 & ~n15639 ;
  assign n15641 = ~n15637 & n15640 ;
  assign n15642 = n8815 & ~n15641 ;
  assign n15643 = \u4_u1_uc_bsel_reg[1]/P0001  & n8816 ;
  assign n15644 = \u4_u1_buf1_reg[31]/P0001  & n2731 ;
  assign n15645 = \u4_u1_buf0_reg[31]/P0001  & n2568 ;
  assign n15646 = ~n15644 & ~n15645 ;
  assign n15647 = ~n15643 & n15646 ;
  assign n15648 = n8866 & ~n15647 ;
  assign n15649 = ~n15642 & ~n15648 ;
  assign n15650 = \u1_mfm_cnt_reg[3]/P0001  & \wb_addr_i[4]_pad  ;
  assign n15651 = n8816 & n15650 ;
  assign n15652 = n8864 & n15651 ;
  assign n15653 = \u4_u3_uc_bsel_reg[1]/P0001  & n8816 ;
  assign n15654 = \u4_u3_buf1_reg[31]/P0001  & n2731 ;
  assign n15655 = \u4_u3_buf0_reg[31]/P0001  & n2568 ;
  assign n15656 = ~n15654 & ~n15655 ;
  assign n15657 = ~n15653 & n15656 ;
  assign n15658 = n8836 & ~n15657 ;
  assign n15659 = ~n15652 & ~n15658 ;
  assign n15660 = \u4_u2_uc_bsel_reg[1]/P0001  & n8816 ;
  assign n15661 = \u4_u2_buf1_reg[31]/P0001  & n2731 ;
  assign n15662 = \u4_u2_buf0_reg[31]/P0001  & n2568 ;
  assign n15663 = ~n15661 & ~n15662 ;
  assign n15664 = ~n15660 & n15663 ;
  assign n15665 = n8826 & ~n15664 ;
  assign n15666 = n15659 & ~n15665 ;
  assign n15667 = n15649 & n15666 ;
  assign n15668 = \u4_u0_uc_bsel_reg[0]/P0001  & n8816 ;
  assign n15669 = \u4_u0_buf1_reg[30]/P0001  & n2731 ;
  assign n15670 = \u4_u0_buf0_reg[30]/P0001  & n2568 ;
  assign n15671 = ~n15669 & ~n15670 ;
  assign n15672 = ~n15668 & n15671 ;
  assign n15673 = n8815 & ~n15672 ;
  assign n15674 = \u4_u1_uc_bsel_reg[0]/P0001  & n8816 ;
  assign n15675 = \u4_u1_buf1_reg[30]/P0001  & n2731 ;
  assign n15676 = \u4_u1_buf0_reg[30]/P0001  & n2568 ;
  assign n15677 = ~n15675 & ~n15676 ;
  assign n15678 = ~n15674 & n15677 ;
  assign n15679 = n8866 & ~n15678 ;
  assign n15680 = ~n15673 & ~n15679 ;
  assign n15681 = \u1_mfm_cnt_reg[2]/P0001  & \wb_addr_i[4]_pad  ;
  assign n15682 = n8816 & n15681 ;
  assign n15683 = n8864 & n15682 ;
  assign n15684 = \u4_u3_uc_bsel_reg[0]/P0001  & n8816 ;
  assign n15685 = \u4_u3_buf1_reg[30]/P0001  & n2731 ;
  assign n15686 = \u4_u3_buf0_reg[30]/P0001  & n2568 ;
  assign n15687 = ~n15685 & ~n15686 ;
  assign n15688 = ~n15684 & n15687 ;
  assign n15689 = n8836 & ~n15688 ;
  assign n15690 = ~n15683 & ~n15689 ;
  assign n15691 = \u4_u2_uc_bsel_reg[0]/P0001  & n8816 ;
  assign n15692 = \u4_u2_buf1_reg[30]/P0001  & n2731 ;
  assign n15693 = \u4_u2_buf0_reg[30]/P0001  & n2568 ;
  assign n15694 = ~n15692 & ~n15693 ;
  assign n15695 = ~n15691 & n15694 ;
  assign n15696 = n8826 & ~n15695 ;
  assign n15697 = n15690 & ~n15696 ;
  assign n15698 = n15680 & n15697 ;
  assign n15699 = \u4_u2_iena_reg[5]/P0001  & n8820 ;
  assign n15700 = \u4_u2_buf0_reg[29]/P0001  & n2568 ;
  assign n15701 = ~n15699 & ~n15700 ;
  assign n15702 = \u4_u2_buf1_reg[29]/P0001  & n2731 ;
  assign n15703 = \u4_u2_uc_dpd_reg[1]/P0001  & n8816 ;
  assign n15704 = ~n15702 & ~n15703 ;
  assign n15705 = n15701 & n15704 ;
  assign n15706 = n8826 & ~n15705 ;
  assign n15707 = \u4_u0_buf1_reg[29]/P0001  & n2731 ;
  assign n15708 = \u4_u0_iena_reg[5]/P0001  & n8820 ;
  assign n15709 = ~n15707 & ~n15708 ;
  assign n15710 = \u4_u0_buf0_reg[29]/P0001  & n2568 ;
  assign n15711 = \u4_u0_uc_dpd_reg[1]/P0001  & n8816 ;
  assign n15712 = ~n15710 & ~n15711 ;
  assign n15713 = n15709 & n15712 ;
  assign n15714 = n8815 & ~n15713 ;
  assign n15715 = ~n15706 & ~n15714 ;
  assign n15716 = \u1_mfm_cnt_reg[1]/P0001  & \wb_addr_i[4]_pad  ;
  assign n15717 = n8816 & n15716 ;
  assign n15718 = n8864 & n15717 ;
  assign n15719 = \u4_u3_buf0_reg[29]/P0001  & n2568 ;
  assign n15720 = \u4_u3_uc_dpd_reg[1]/P0001  & n8816 ;
  assign n15721 = ~n15719 & ~n15720 ;
  assign n15722 = \u4_u3_iena_reg[5]/P0001  & n8820 ;
  assign n15723 = \u4_u3_buf1_reg[29]/P0001  & n2731 ;
  assign n15724 = ~n15722 & ~n15723 ;
  assign n15725 = n15721 & n15724 ;
  assign n15726 = n8836 & ~n15725 ;
  assign n15727 = ~n15718 & ~n15726 ;
  assign n15728 = \u4_u1_buf0_reg[29]/P0001  & n2568 ;
  assign n15729 = \u4_u1_buf1_reg[29]/P0001  & n2731 ;
  assign n15730 = ~n15728 & ~n15729 ;
  assign n15731 = \u4_u1_uc_dpd_reg[1]/P0001  & n8816 ;
  assign n15732 = \u4_u1_iena_reg[5]/P0001  & n8820 ;
  assign n15733 = ~n15731 & ~n15732 ;
  assign n15734 = n15730 & n15733 ;
  assign n15735 = n8866 & ~n15734 ;
  assign n15736 = n15727 & ~n15735 ;
  assign n15737 = n15715 & n15736 ;
  assign n15738 = \u1_u3_uc_bsel_set_reg/P0001  & \u4_u2_ep_match_r_reg/P0001  ;
  assign n15739 = rst_i_pad & \u4_u2_uc_bsel_reg[0]/P0001  ;
  assign n15740 = ~n15738 & n15739 ;
  assign n15741 = rst_i_pad & \u1_u3_idin_reg[0]/P0001  ;
  assign n15742 = n15738 & n15741 ;
  assign n15743 = ~n15740 & ~n15742 ;
  assign n15744 = rst_i_pad & \u4_u2_uc_bsel_reg[1]/P0001  ;
  assign n15745 = ~n15738 & n15744 ;
  assign n15746 = rst_i_pad & \u1_u3_idin_reg[1]/P0001  ;
  assign n15747 = n15738 & n15746 ;
  assign n15748 = ~n15745 & ~n15747 ;
  assign n15749 = rst_i_pad & \u4_u2_uc_dpd_reg[1]/P0001  ;
  assign n15750 = ~n15738 & n15749 ;
  assign n15751 = rst_i_pad & \u1_u3_idin_reg[3]/P0001  ;
  assign n15752 = n15738 & n15751 ;
  assign n15753 = ~n15750 & ~n15752 ;
  assign n15754 = \u4_u3_csr1_reg[12]/P0001  & n8816 ;
  assign n15755 = \u4_u3_buf1_reg[27]/P0001  & n2731 ;
  assign n15756 = ~n15754 & ~n15755 ;
  assign n15757 = \u4_u3_iena_reg[3]/P0001  & n8820 ;
  assign n15758 = \u4_u3_buf0_reg[27]/P0001  & n2568 ;
  assign n15759 = ~n15757 & ~n15758 ;
  assign n15760 = n15756 & n15759 ;
  assign n15761 = n8836 & ~n15760 ;
  assign n15762 = \u4_u2_iena_reg[3]/P0001  & n8820 ;
  assign n15763 = \u4_u2_buf1_reg[27]/P0001  & n2731 ;
  assign n15764 = ~n15762 & ~n15763 ;
  assign n15765 = \u4_u2_buf0_reg[27]/P0001  & n2568 ;
  assign n15766 = \u4_u2_csr1_reg[12]/P0001  & n8816 ;
  assign n15767 = ~n15765 & ~n15766 ;
  assign n15768 = n15764 & n15767 ;
  assign n15769 = n8826 & ~n15768 ;
  assign n15770 = ~n15761 & ~n15769 ;
  assign n15771 = \u4_int_srcb_reg[7]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n15772 = n2731 & n15771 ;
  assign n15773 = n8864 & n15772 ;
  assign n15774 = \u4_u1_buf0_reg[27]/P0001  & n2568 ;
  assign n15775 = \u4_u1_csr1_reg[12]/P0001  & n8816 ;
  assign n15776 = ~n15774 & ~n15775 ;
  assign n15777 = \u4_u1_buf1_reg[27]/P0001  & n2731 ;
  assign n15778 = \u4_u1_iena_reg[3]/P0001  & n8820 ;
  assign n15779 = ~n15777 & ~n15778 ;
  assign n15780 = n15776 & n15779 ;
  assign n15781 = n8866 & ~n15780 ;
  assign n15782 = ~n15773 & ~n15781 ;
  assign n15783 = \u4_u0_iena_reg[3]/P0001  & n8820 ;
  assign n15784 = \u4_u0_buf1_reg[27]/P0001  & n2731 ;
  assign n15785 = ~n15783 & ~n15784 ;
  assign n15786 = \u4_u0_csr1_reg[12]/P0001  & n8816 ;
  assign n15787 = \u4_u0_buf0_reg[27]/P0001  & n2568 ;
  assign n15788 = ~n15786 & ~n15787 ;
  assign n15789 = n15785 & n15788 ;
  assign n15790 = n8815 & ~n15789 ;
  assign n15791 = n15782 & ~n15790 ;
  assign n15792 = n15770 & n15791 ;
  assign n15793 = \u1_u3_uc_bsel_set_reg/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n15794 = rst_i_pad & \u4_u3_uc_bsel_reg[0]/P0001  ;
  assign n15795 = ~n15793 & n15794 ;
  assign n15796 = n15741 & n15793 ;
  assign n15797 = ~n15795 & ~n15796 ;
  assign n15798 = rst_i_pad & \u4_u3_uc_bsel_reg[1]/P0001  ;
  assign n15799 = ~n15793 & n15798 ;
  assign n15800 = n15746 & n15793 ;
  assign n15801 = ~n15799 & ~n15800 ;
  assign n15802 = rst_i_pad & \u4_u3_uc_dpd_reg[0]/P0001  ;
  assign n15803 = ~n15793 & n15802 ;
  assign n15804 = rst_i_pad & \u1_u3_idin_reg[2]/P0001  ;
  assign n15805 = n15793 & n15804 ;
  assign n15806 = ~n15803 & ~n15805 ;
  assign n15807 = \u4_u1_buf1_reg[8]/P0001  & n2731 ;
  assign n15808 = \u4_u1_csr0_reg[8]/P0001  & n8816 ;
  assign n15809 = \u4_u1_buf0_reg[8]/P0001  & n2568 ;
  assign n15810 = ~n15808 & ~n15809 ;
  assign n15811 = ~n15807 & n15810 ;
  assign n15812 = n8866 & ~n15811 ;
  assign n15813 = \u4_u2_buf1_reg[8]/P0001  & n2731 ;
  assign n15814 = \u4_u2_buf0_reg[8]/P0001  & n2568 ;
  assign n15815 = \u4_u2_csr0_reg[8]/P0001  & n8816 ;
  assign n15816 = ~n15814 & ~n15815 ;
  assign n15817 = ~n15813 & n15816 ;
  assign n15818 = n8826 & ~n15817 ;
  assign n15819 = ~n15812 & ~n15818 ;
  assign n15820 = \u4_u0_buf1_reg[8]/P0001  & n2731 ;
  assign n15821 = \u4_u0_buf0_reg[8]/P0001  & n2568 ;
  assign n15822 = \u4_u0_csr0_reg[8]/P0001  & n8816 ;
  assign n15823 = ~n15821 & ~n15822 ;
  assign n15824 = ~n15820 & n15823 ;
  assign n15825 = n8815 & ~n15824 ;
  assign n15826 = \u4_u3_buf1_reg[8]/P0001  & n2731 ;
  assign n15827 = \u4_u3_csr0_reg[8]/P0001  & n8816 ;
  assign n15828 = \u4_u3_buf0_reg[8]/P0001  & n2568 ;
  assign n15829 = ~n15827 & ~n15828 ;
  assign n15830 = ~n15826 & n15829 ;
  assign n15831 = n8836 & ~n15830 ;
  assign n15832 = ~n15825 & ~n15831 ;
  assign n15833 = \u1_sof_time_reg[8]/P0001  & \wb_addr_i[4]_pad  ;
  assign n15834 = n8816 & n15833 ;
  assign n15835 = \u4_inta_msk_reg[8]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n15836 = n2568 & n15835 ;
  assign n15837 = ~n15834 & ~n15836 ;
  assign n15838 = n8864 & ~n15837 ;
  assign n15839 = n15832 & ~n15838 ;
  assign n15840 = n15819 & n15839 ;
  assign n15841 = rst_i_pad & \u4_u2_uc_dpd_reg[0]/P0001  ;
  assign n15842 = ~n15738 & n15841 ;
  assign n15843 = n15738 & n15804 ;
  assign n15844 = ~n15842 & ~n15843 ;
  assign n15845 = rst_i_pad & \u4_u3_uc_dpd_reg[1]/P0001  ;
  assign n15846 = ~n15793 & n15845 ;
  assign n15847 = n15751 & n15793 ;
  assign n15848 = ~n15846 & ~n15847 ;
  assign n15849 = \u1_u3_uc_bsel_set_reg/P0001  & \u4_u0_ep_match_r_reg/P0001  ;
  assign n15850 = rst_i_pad & \u4_u0_uc_bsel_reg[0]/P0001  ;
  assign n15851 = ~n15849 & n15850 ;
  assign n15852 = n15741 & n15849 ;
  assign n15853 = ~n15851 & ~n15852 ;
  assign n15854 = rst_i_pad & \u4_u0_uc_bsel_reg[1]/P0001  ;
  assign n15855 = ~n15849 & n15854 ;
  assign n15856 = n15746 & n15849 ;
  assign n15857 = ~n15855 & ~n15856 ;
  assign n15858 = rst_i_pad & \u4_u0_uc_dpd_reg[0]/P0001  ;
  assign n15859 = ~n15849 & n15858 ;
  assign n15860 = n15804 & n15849 ;
  assign n15861 = ~n15859 & ~n15860 ;
  assign n15862 = rst_i_pad & \u4_u0_uc_dpd_reg[1]/P0001  ;
  assign n15863 = ~n15849 & n15862 ;
  assign n15864 = n15751 & n15849 ;
  assign n15865 = ~n15863 & ~n15864 ;
  assign n15866 = ~\u1_u0_pid_reg[2]/NET0131  & n7806 ;
  assign n15867 = n13025 & ~n15866 ;
  assign n15868 = ~n12304 & ~n13009 ;
  assign n15869 = n2363 & ~n15868 ;
  assign n15870 = ~\u4_csr_reg[28]/P0001  & n2361 ;
  assign n15871 = n12304 & n15870 ;
  assign n15872 = ~n15869 & ~n15871 ;
  assign n15873 = n5555 & ~n13025 ;
  assign n15874 = ~n15872 & n15873 ;
  assign n15875 = ~n15867 & ~n15874 ;
  assign n15876 = n5748 & n6157 ;
  assign n15877 = ~\u0_u0_me_cnt_100_ms_reg/P0001  & n5748 ;
  assign n15878 = n8663 & n15877 ;
  assign n15879 = ~n15876 & ~n15878 ;
  assign n15880 = \u1_u3_uc_bsel_set_reg/P0001  & \u4_u1_ep_match_r_reg/P0001  ;
  assign n15881 = rst_i_pad & \u4_u1_uc_bsel_reg[0]/P0001  ;
  assign n15882 = ~n15880 & n15881 ;
  assign n15883 = n15741 & n15880 ;
  assign n15884 = ~n15882 & ~n15883 ;
  assign n15885 = rst_i_pad & \u4_u1_uc_bsel_reg[1]/P0001  ;
  assign n15886 = ~n15880 & n15885 ;
  assign n15887 = n15746 & n15880 ;
  assign n15888 = ~n15886 & ~n15887 ;
  assign n15889 = rst_i_pad & \u4_u1_uc_dpd_reg[0]/P0001  ;
  assign n15890 = ~n15880 & n15889 ;
  assign n15891 = n15804 & n15880 ;
  assign n15892 = ~n15890 & ~n15891 ;
  assign n15893 = rst_i_pad & \u4_u1_uc_dpd_reg[1]/P0001  ;
  assign n15894 = ~n15880 & n15893 ;
  assign n15895 = n15751 & n15880 ;
  assign n15896 = ~n15894 & ~n15895 ;
  assign n15897 = ~\u1_u3_new_sizeb_reg[0]/P0001  & ~n3483 ;
  assign n15898 = ~n4440 & ~n15897 ;
  assign n15899 = ~\u0_u0_T2_wakeup_reg/P0001  & n6137 ;
  assign n15900 = n6143 & n15899 ;
  assign n15901 = ~\u0_u0_state_reg[5]/P0001  & ~n12961 ;
  assign n15902 = ~n5768 & ~n15901 ;
  assign n15903 = n15229 & n15902 ;
  assign n15904 = n12653 & n15903 ;
  assign n15905 = ~n15900 & ~n15904 ;
  assign n15906 = n5748 & ~n15905 ;
  assign n15907 = ~\u0_u0_T2_gt_1_0_mS_reg/P0001  & n15240 ;
  assign n15908 = ~n6167 & ~n15907 ;
  assign n15909 = n5748 & ~n15908 ;
  assign n15910 = \u4_intb_msk_reg[0]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n15911 = n2568 & n15910 ;
  assign n15912 = \u1_frame_no_r_reg[0]/P0001  & \wb_addr_i[4]_pad  ;
  assign n15913 = n8816 & n15912 ;
  assign n15914 = ~n15911 & ~n15913 ;
  assign n15915 = n8864 & ~n15914 ;
  assign n15916 = \u4_u1_csr1_reg[1]/P0001  & n8816 ;
  assign n15917 = \u4_u1_buf1_reg[16]/P0001  & n2731 ;
  assign n15918 = ~n15916 & ~n15917 ;
  assign n15919 = \u4_u1_ienb_reg[0]/P0001  & n8820 ;
  assign n15920 = \u4_u1_buf0_reg[16]/P0001  & n2568 ;
  assign n15921 = ~n15919 & ~n15920 ;
  assign n15922 = n15918 & n15921 ;
  assign n15923 = n8866 & ~n15922 ;
  assign n15924 = ~n15915 & ~n15923 ;
  assign n15925 = \u4_u3_buf0_reg[16]/P0001  & n2568 ;
  assign n15926 = \u4_u3_csr1_reg[1]/P0001  & n8816 ;
  assign n15927 = ~n15925 & ~n15926 ;
  assign n15928 = \u4_u3_buf1_reg[16]/P0001  & n2731 ;
  assign n15929 = \u4_u3_ienb_reg[0]/P0001  & n8820 ;
  assign n15930 = ~n15928 & ~n15929 ;
  assign n15931 = n15927 & n15930 ;
  assign n15932 = n8836 & ~n15931 ;
  assign n15933 = \u4_u0_csr1_reg[1]/P0001  & n8816 ;
  assign n15934 = \u4_u0_buf1_reg[16]/P0001  & n2731 ;
  assign n15935 = ~n15933 & ~n15934 ;
  assign n15936 = \u4_u0_ienb_reg[0]/P0001  & n8820 ;
  assign n15937 = \u4_u0_buf0_reg[16]/P0001  & n2568 ;
  assign n15938 = ~n15936 & ~n15937 ;
  assign n15939 = n15935 & n15938 ;
  assign n15940 = n8815 & ~n15939 ;
  assign n15941 = ~n15932 & ~n15940 ;
  assign n15942 = \u4_u2_csr1_reg[1]/P0001  & n8816 ;
  assign n15943 = \u4_u2_buf1_reg[16]/P0001  & n2731 ;
  assign n15944 = ~n15942 & ~n15943 ;
  assign n15945 = \u4_u2_ienb_reg[0]/P0001  & n8820 ;
  assign n15946 = \u4_u2_buf0_reg[16]/P0001  & n2568 ;
  assign n15947 = ~n15945 & ~n15946 ;
  assign n15948 = n15944 & n15947 ;
  assign n15949 = n8826 & ~n15948 ;
  assign n15950 = n15941 & ~n15949 ;
  assign n15951 = n15924 & n15950 ;
  assign n15952 = \u4_intb_msk_reg[1]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n15953 = n2568 & n15952 ;
  assign n15954 = \u1_frame_no_r_reg[1]/P0001  & \wb_addr_i[4]_pad  ;
  assign n15955 = n8816 & n15954 ;
  assign n15956 = ~n15953 & ~n15955 ;
  assign n15957 = n8864 & ~n15956 ;
  assign n15958 = \u4_u1_csr1_reg[2]/P0001  & n8816 ;
  assign n15959 = \u4_u1_buf1_reg[17]/P0001  & n2731 ;
  assign n15960 = ~n15958 & ~n15959 ;
  assign n15961 = \u4_u1_ienb_reg[1]/P0001  & n8820 ;
  assign n15962 = \u4_u1_buf0_reg[17]/P0001  & n2568 ;
  assign n15963 = ~n15961 & ~n15962 ;
  assign n15964 = n15960 & n15963 ;
  assign n15965 = n8866 & ~n15964 ;
  assign n15966 = ~n15957 & ~n15965 ;
  assign n15967 = \u4_u3_csr1_reg[2]/P0001  & n8816 ;
  assign n15968 = \u4_u3_buf0_reg[17]/P0001  & n2568 ;
  assign n15969 = ~n15967 & ~n15968 ;
  assign n15970 = \u4_u3_ienb_reg[1]/P0001  & n8820 ;
  assign n15971 = \u4_u3_buf1_reg[17]/P0001  & n2731 ;
  assign n15972 = ~n15970 & ~n15971 ;
  assign n15973 = n15969 & n15972 ;
  assign n15974 = n8836 & ~n15973 ;
  assign n15975 = \u4_u0_csr1_reg[2]/P0001  & n8816 ;
  assign n15976 = \u4_u0_buf1_reg[17]/P0001  & n2731 ;
  assign n15977 = ~n15975 & ~n15976 ;
  assign n15978 = \u4_u0_ienb_reg[1]/P0001  & n8820 ;
  assign n15979 = \u4_u0_buf0_reg[17]/P0001  & n2568 ;
  assign n15980 = ~n15978 & ~n15979 ;
  assign n15981 = n15977 & n15980 ;
  assign n15982 = n8815 & ~n15981 ;
  assign n15983 = ~n15974 & ~n15982 ;
  assign n15984 = \u4_u2_csr1_reg[2]/P0001  & n8816 ;
  assign n15985 = \u4_u2_buf1_reg[17]/P0001  & n2731 ;
  assign n15986 = ~n15984 & ~n15985 ;
  assign n15987 = \u4_u2_ienb_reg[1]/P0001  & n8820 ;
  assign n15988 = \u4_u2_buf0_reg[17]/P0001  & n2568 ;
  assign n15989 = ~n15987 & ~n15988 ;
  assign n15990 = n15986 & n15989 ;
  assign n15991 = n8826 & ~n15990 ;
  assign n15992 = n15983 & ~n15991 ;
  assign n15993 = n15966 & n15992 ;
  assign n15994 = \u4_intb_msk_reg[2]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n15995 = n2568 & n15994 ;
  assign n15996 = \u1_frame_no_r_reg[2]/P0001  & \wb_addr_i[4]_pad  ;
  assign n15997 = n8816 & n15996 ;
  assign n15998 = ~n15995 & ~n15997 ;
  assign n15999 = n8864 & ~n15998 ;
  assign n16000 = \u4_u1_csr1_reg[3]/P0001  & n8816 ;
  assign n16001 = \u4_u1_buf1_reg[18]/P0001  & n2731 ;
  assign n16002 = ~n16000 & ~n16001 ;
  assign n16003 = \u4_u1_ienb_reg[2]/P0001  & n8820 ;
  assign n16004 = \u4_u1_buf0_reg[18]/P0001  & n2568 ;
  assign n16005 = ~n16003 & ~n16004 ;
  assign n16006 = n16002 & n16005 ;
  assign n16007 = n8866 & ~n16006 ;
  assign n16008 = ~n15999 & ~n16007 ;
  assign n16009 = \u4_u2_buf0_reg[18]/P0001  & n2568 ;
  assign n16010 = \u4_u2_csr1_reg[3]/P0001  & n8816 ;
  assign n16011 = ~n16009 & ~n16010 ;
  assign n16012 = \u4_u2_buf1_reg[18]/P0001  & n2731 ;
  assign n16013 = \u4_u2_ienb_reg[2]/P0001  & n8820 ;
  assign n16014 = ~n16012 & ~n16013 ;
  assign n16015 = n16011 & n16014 ;
  assign n16016 = n8826 & ~n16015 ;
  assign n16017 = \u4_u0_csr1_reg[3]/P0001  & n8816 ;
  assign n16018 = \u4_u0_buf1_reg[18]/P0001  & n2731 ;
  assign n16019 = ~n16017 & ~n16018 ;
  assign n16020 = \u4_u0_ienb_reg[2]/P0001  & n8820 ;
  assign n16021 = \u4_u0_buf0_reg[18]/P0001  & n2568 ;
  assign n16022 = ~n16020 & ~n16021 ;
  assign n16023 = n16019 & n16022 ;
  assign n16024 = n8815 & ~n16023 ;
  assign n16025 = ~n16016 & ~n16024 ;
  assign n16026 = \u4_u3_csr1_reg[3]/P0001  & n8816 ;
  assign n16027 = \u4_u3_buf1_reg[18]/P0001  & n2731 ;
  assign n16028 = ~n16026 & ~n16027 ;
  assign n16029 = \u4_u3_ienb_reg[2]/P0001  & n8820 ;
  assign n16030 = \u4_u3_buf0_reg[18]/P0001  & n2568 ;
  assign n16031 = ~n16029 & ~n16030 ;
  assign n16032 = n16028 & n16031 ;
  assign n16033 = n8836 & ~n16032 ;
  assign n16034 = n16025 & ~n16033 ;
  assign n16035 = n16008 & n16034 ;
  assign n16036 = \u4_intb_msk_reg[3]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16037 = n2568 & n16036 ;
  assign n16038 = \u1_frame_no_r_reg[3]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16039 = n8816 & n16038 ;
  assign n16040 = ~n16037 & ~n16039 ;
  assign n16041 = n8864 & ~n16040 ;
  assign n16042 = \u4_u1_csr1_reg[4]/P0001  & n8816 ;
  assign n16043 = \u4_u1_buf1_reg[19]/P0001  & n2731 ;
  assign n16044 = ~n16042 & ~n16043 ;
  assign n16045 = \u4_u1_ienb_reg[3]/P0001  & n8820 ;
  assign n16046 = \u4_u1_buf0_reg[19]/P0001  & n2568 ;
  assign n16047 = ~n16045 & ~n16046 ;
  assign n16048 = n16044 & n16047 ;
  assign n16049 = n8866 & ~n16048 ;
  assign n16050 = ~n16041 & ~n16049 ;
  assign n16051 = \u4_u2_buf0_reg[19]/P0001  & n2568 ;
  assign n16052 = \u4_u2_csr1_reg[4]/P0001  & n8816 ;
  assign n16053 = ~n16051 & ~n16052 ;
  assign n16054 = \u4_u2_buf1_reg[19]/P0001  & n2731 ;
  assign n16055 = \u4_u2_ienb_reg[3]/P0001  & n8820 ;
  assign n16056 = ~n16054 & ~n16055 ;
  assign n16057 = n16053 & n16056 ;
  assign n16058 = n8826 & ~n16057 ;
  assign n16059 = \u4_u0_csr1_reg[4]/P0001  & n8816 ;
  assign n16060 = \u4_u0_buf1_reg[19]/P0001  & n2731 ;
  assign n16061 = ~n16059 & ~n16060 ;
  assign n16062 = \u4_u0_ienb_reg[3]/P0001  & n8820 ;
  assign n16063 = \u4_u0_buf0_reg[19]/P0001  & n2568 ;
  assign n16064 = ~n16062 & ~n16063 ;
  assign n16065 = n16061 & n16064 ;
  assign n16066 = n8815 & ~n16065 ;
  assign n16067 = ~n16058 & ~n16066 ;
  assign n16068 = \u4_u3_csr1_reg[4]/P0001  & n8816 ;
  assign n16069 = \u4_u3_buf1_reg[19]/P0001  & n2731 ;
  assign n16070 = ~n16068 & ~n16069 ;
  assign n16071 = \u4_u3_ienb_reg[3]/P0001  & n8820 ;
  assign n16072 = \u4_u3_buf0_reg[19]/P0001  & n2568 ;
  assign n16073 = ~n16071 & ~n16072 ;
  assign n16074 = n16070 & n16073 ;
  assign n16075 = n8836 & ~n16074 ;
  assign n16076 = n16067 & ~n16075 ;
  assign n16077 = n16050 & n16076 ;
  assign n16078 = \u4_int_srcb_reg[5]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16079 = n2731 & n16078 ;
  assign n16080 = \u1_frame_no_r_reg[9]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16081 = n8816 & n16080 ;
  assign n16082 = ~n16079 & ~n16081 ;
  assign n16083 = n8864 & ~n16082 ;
  assign n16084 = \u4_u1_csr1_reg[10]/P0001  & n8816 ;
  assign n16085 = \u4_u1_buf1_reg[25]/P0001  & n2731 ;
  assign n16086 = ~n16084 & ~n16085 ;
  assign n16087 = \u4_u1_iena_reg[1]/P0001  & n8820 ;
  assign n16088 = \u4_u1_buf0_reg[25]/P0001  & n2568 ;
  assign n16089 = ~n16087 & ~n16088 ;
  assign n16090 = n16086 & n16089 ;
  assign n16091 = n8866 & ~n16090 ;
  assign n16092 = ~n16083 & ~n16091 ;
  assign n16093 = \u4_u3_buf0_reg[25]/P0001  & n2568 ;
  assign n16094 = \u4_u3_csr1_reg[10]/P0001  & n8816 ;
  assign n16095 = ~n16093 & ~n16094 ;
  assign n16096 = \u4_u3_buf1_reg[25]/P0001  & n2731 ;
  assign n16097 = \u4_u3_iena_reg[1]/P0001  & n8820 ;
  assign n16098 = ~n16096 & ~n16097 ;
  assign n16099 = n16095 & n16098 ;
  assign n16100 = n8836 & ~n16099 ;
  assign n16101 = \u4_u0_csr1_reg[10]/P0001  & n8816 ;
  assign n16102 = \u4_u0_buf1_reg[25]/P0001  & n2731 ;
  assign n16103 = ~n16101 & ~n16102 ;
  assign n16104 = \u4_u0_iena_reg[1]/P0001  & n8820 ;
  assign n16105 = \u4_u0_buf0_reg[25]/P0001  & n2568 ;
  assign n16106 = ~n16104 & ~n16105 ;
  assign n16107 = n16103 & n16106 ;
  assign n16108 = n8815 & ~n16107 ;
  assign n16109 = ~n16100 & ~n16108 ;
  assign n16110 = \u4_u2_csr1_reg[10]/P0001  & n8816 ;
  assign n16111 = \u4_u2_buf1_reg[25]/P0001  & n2731 ;
  assign n16112 = ~n16110 & ~n16111 ;
  assign n16113 = \u4_u2_iena_reg[1]/P0001  & n8820 ;
  assign n16114 = \u4_u2_buf0_reg[25]/P0001  & n2568 ;
  assign n16115 = ~n16113 & ~n16114 ;
  assign n16116 = n16112 & n16115 ;
  assign n16117 = n8826 & ~n16116 ;
  assign n16118 = n16109 & ~n16117 ;
  assign n16119 = n16092 & n16118 ;
  assign n16120 = \u4_int_srcb_reg[6]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16121 = n2731 & n16120 ;
  assign n16122 = \u1_frame_no_r_reg[10]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16123 = n8816 & n16122 ;
  assign n16124 = ~n16121 & ~n16123 ;
  assign n16125 = n8864 & ~n16124 ;
  assign n16126 = \u4_u1_iena_reg[2]/P0001  & n8820 ;
  assign n16127 = \u4_u1_buf1_reg[26]/P0001  & n2731 ;
  assign n16128 = ~n16126 & ~n16127 ;
  assign n16129 = \u4_u1_csr1_reg[11]/P0001  & n8816 ;
  assign n16130 = \u4_u1_buf0_reg[26]/P0001  & n2568 ;
  assign n16131 = ~n16129 & ~n16130 ;
  assign n16132 = n16128 & n16131 ;
  assign n16133 = n8866 & ~n16132 ;
  assign n16134 = ~n16125 & ~n16133 ;
  assign n16135 = \u4_u3_buf0_reg[26]/P0001  & n2568 ;
  assign n16136 = \u4_u3_csr1_reg[11]/P0001  & n8816 ;
  assign n16137 = ~n16135 & ~n16136 ;
  assign n16138 = \u4_u3_buf1_reg[26]/P0001  & n2731 ;
  assign n16139 = \u4_u3_iena_reg[2]/P0001  & n8820 ;
  assign n16140 = ~n16138 & ~n16139 ;
  assign n16141 = n16137 & n16140 ;
  assign n16142 = n8836 & ~n16141 ;
  assign n16143 = \u4_u0_iena_reg[2]/P0001  & n8820 ;
  assign n16144 = \u4_u0_buf1_reg[26]/P0001  & n2731 ;
  assign n16145 = ~n16143 & ~n16144 ;
  assign n16146 = \u4_u0_csr1_reg[11]/P0001  & n8816 ;
  assign n16147 = \u4_u0_buf0_reg[26]/P0001  & n2568 ;
  assign n16148 = ~n16146 & ~n16147 ;
  assign n16149 = n16145 & n16148 ;
  assign n16150 = n8815 & ~n16149 ;
  assign n16151 = ~n16142 & ~n16150 ;
  assign n16152 = \u4_u2_iena_reg[2]/P0001  & n8820 ;
  assign n16153 = \u4_u2_buf1_reg[26]/P0001  & n2731 ;
  assign n16154 = ~n16152 & ~n16153 ;
  assign n16155 = \u4_u2_csr1_reg[11]/P0001  & n8816 ;
  assign n16156 = \u4_u2_buf0_reg[26]/P0001  & n2568 ;
  assign n16157 = ~n16155 & ~n16156 ;
  assign n16158 = n16154 & n16157 ;
  assign n16159 = n8826 & ~n16158 ;
  assign n16160 = n16151 & ~n16159 ;
  assign n16161 = n16134 & n16160 ;
  assign n16162 = \u4_int_srcb_reg[8]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16163 = n2731 & n16162 ;
  assign n16164 = \u1_mfm_cnt_reg[0]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16165 = n8816 & n16164 ;
  assign n16166 = ~n16163 & ~n16165 ;
  assign n16167 = n8864 & ~n16166 ;
  assign n16168 = \u4_u1_iena_reg[4]/P0001  & n8820 ;
  assign n16169 = \u4_u1_buf1_reg[28]/P0001  & n2731 ;
  assign n16170 = ~n16168 & ~n16169 ;
  assign n16171 = \u4_u1_uc_dpd_reg[0]/P0001  & n8816 ;
  assign n16172 = \u4_u1_buf0_reg[28]/P0001  & n2568 ;
  assign n16173 = ~n16171 & ~n16172 ;
  assign n16174 = n16170 & n16173 ;
  assign n16175 = n8866 & ~n16174 ;
  assign n16176 = ~n16167 & ~n16175 ;
  assign n16177 = \u4_u2_iena_reg[4]/P0001  & n8820 ;
  assign n16178 = \u4_u2_buf0_reg[28]/P0001  & n2568 ;
  assign n16179 = ~n16177 & ~n16178 ;
  assign n16180 = \u4_u2_uc_dpd_reg[0]/P0001  & n8816 ;
  assign n16181 = \u4_u2_buf1_reg[28]/P0001  & n2731 ;
  assign n16182 = ~n16180 & ~n16181 ;
  assign n16183 = n16179 & n16182 ;
  assign n16184 = n8826 & ~n16183 ;
  assign n16185 = \u4_u0_iena_reg[4]/P0001  & n8820 ;
  assign n16186 = \u4_u0_buf1_reg[28]/P0001  & n2731 ;
  assign n16187 = ~n16185 & ~n16186 ;
  assign n16188 = \u4_u0_uc_dpd_reg[0]/P0001  & n8816 ;
  assign n16189 = \u4_u0_buf0_reg[28]/P0001  & n2568 ;
  assign n16190 = ~n16188 & ~n16189 ;
  assign n16191 = n16187 & n16190 ;
  assign n16192 = n8815 & ~n16191 ;
  assign n16193 = ~n16184 & ~n16192 ;
  assign n16194 = \u4_u3_iena_reg[4]/P0001  & n8820 ;
  assign n16195 = \u4_u3_buf1_reg[28]/P0001  & n2731 ;
  assign n16196 = ~n16194 & ~n16195 ;
  assign n16197 = \u4_u3_uc_dpd_reg[0]/P0001  & n8816 ;
  assign n16198 = \u4_u3_buf0_reg[28]/P0001  & n2568 ;
  assign n16199 = ~n16197 & ~n16198 ;
  assign n16200 = n16196 & n16199 ;
  assign n16201 = n8836 & ~n16200 ;
  assign n16202 = n16193 & ~n16201 ;
  assign n16203 = n16176 & n16202 ;
  assign n16204 = \u4_u2_buf0_reg[21]/P0001  & n2568 ;
  assign n16205 = \u4_u2_csr1_reg[6]/P0001  & n8816 ;
  assign n16206 = ~n16204 & ~n16205 ;
  assign n16207 = \u4_u2_buf1_reg[21]/P0001  & n2731 ;
  assign n16208 = \u4_u2_ienb_reg[5]/P0001  & n8820 ;
  assign n16209 = ~n16207 & ~n16208 ;
  assign n16210 = n16206 & n16209 ;
  assign n16211 = n8826 & ~n16210 ;
  assign n16212 = \u4_u3_csr1_reg[6]/P0001  & n8816 ;
  assign n16213 = \u4_u3_buf1_reg[21]/P0001  & n2731 ;
  assign n16214 = ~n16212 & ~n16213 ;
  assign n16215 = \u4_u3_ienb_reg[5]/P0001  & n8820 ;
  assign n16216 = \u4_u3_buf0_reg[21]/P0001  & n2568 ;
  assign n16217 = ~n16215 & ~n16216 ;
  assign n16218 = n16214 & n16217 ;
  assign n16219 = n8836 & ~n16218 ;
  assign n16220 = ~n16211 & ~n16219 ;
  assign n16221 = \u4_u0_csr1_reg[6]/P0001  & n8816 ;
  assign n16222 = \u4_u0_buf1_reg[21]/P0001  & n2731 ;
  assign n16223 = ~n16221 & ~n16222 ;
  assign n16224 = \u4_u0_ienb_reg[5]/P0001  & n8820 ;
  assign n16225 = \u4_u0_buf0_reg[21]/P0001  & n2568 ;
  assign n16226 = ~n16224 & ~n16225 ;
  assign n16227 = n16223 & n16226 ;
  assign n16228 = n8815 & ~n16227 ;
  assign n16229 = n16220 & ~n16228 ;
  assign n16230 = \u1_frame_no_r_reg[5]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16231 = n8816 & n16230 ;
  assign n16232 = \u4_intb_msk_reg[5]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16233 = n2568 & n16232 ;
  assign n16234 = \u4_int_srcb_reg[1]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16235 = n2731 & n16234 ;
  assign n16236 = ~n16233 & ~n16235 ;
  assign n16237 = ~n16231 & n16236 ;
  assign n16238 = n8864 & ~n16237 ;
  assign n16239 = \u4_u1_csr1_reg[6]/P0001  & n8816 ;
  assign n16240 = \u4_u1_buf1_reg[21]/P0001  & n2731 ;
  assign n16241 = ~n16239 & ~n16240 ;
  assign n16242 = \u4_u1_ienb_reg[5]/P0001  & n8820 ;
  assign n16243 = \u4_u1_buf0_reg[21]/P0001  & n2568 ;
  assign n16244 = ~n16242 & ~n16243 ;
  assign n16245 = n16241 & n16244 ;
  assign n16246 = n8866 & ~n16245 ;
  assign n16247 = ~n16238 & ~n16246 ;
  assign n16248 = n16229 & n16247 ;
  assign n16249 = \u4_u3_buf0_reg[24]/P0001  & n2568 ;
  assign n16250 = \u4_u3_csr1_reg[9]/P0001  & n8816 ;
  assign n16251 = ~n16249 & ~n16250 ;
  assign n16252 = \u4_u3_buf1_reg[24]/P0001  & n2731 ;
  assign n16253 = \u4_u3_iena_reg[0]/P0001  & n8820 ;
  assign n16254 = ~n16252 & ~n16253 ;
  assign n16255 = n16251 & n16254 ;
  assign n16256 = n8836 & ~n16255 ;
  assign n16257 = \u4_u2_csr1_reg[9]/P0001  & n8816 ;
  assign n16258 = \u4_u2_buf1_reg[24]/P0001  & n2731 ;
  assign n16259 = ~n16257 & ~n16258 ;
  assign n16260 = \u4_u2_iena_reg[0]/P0001  & n8820 ;
  assign n16261 = \u4_u2_buf0_reg[24]/P0001  & n2568 ;
  assign n16262 = ~n16260 & ~n16261 ;
  assign n16263 = n16259 & n16262 ;
  assign n16264 = n8826 & ~n16263 ;
  assign n16265 = ~n16256 & ~n16264 ;
  assign n16266 = \u4_u0_csr1_reg[9]/P0001  & n8816 ;
  assign n16267 = \u4_u0_buf1_reg[24]/P0001  & n2731 ;
  assign n16268 = ~n16266 & ~n16267 ;
  assign n16269 = \u4_u0_iena_reg[0]/P0001  & n8820 ;
  assign n16270 = \u4_u0_buf0_reg[24]/P0001  & n2568 ;
  assign n16271 = ~n16269 & ~n16270 ;
  assign n16272 = n16268 & n16271 ;
  assign n16273 = n8815 & ~n16272 ;
  assign n16274 = n16265 & ~n16273 ;
  assign n16275 = \u1_frame_no_r_reg[8]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16276 = n8816 & n16275 ;
  assign n16277 = \u4_intb_msk_reg[8]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16278 = n2568 & n16277 ;
  assign n16279 = \u4_int_srcb_reg[4]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16280 = n2731 & n16279 ;
  assign n16281 = ~n16278 & ~n16280 ;
  assign n16282 = ~n16276 & n16281 ;
  assign n16283 = n8864 & ~n16282 ;
  assign n16284 = \u4_u1_csr1_reg[9]/P0001  & n8816 ;
  assign n16285 = \u4_u1_buf1_reg[24]/P0001  & n2731 ;
  assign n16286 = ~n16284 & ~n16285 ;
  assign n16287 = \u4_u1_iena_reg[0]/P0001  & n8820 ;
  assign n16288 = \u4_u1_buf0_reg[24]/P0001  & n2568 ;
  assign n16289 = ~n16287 & ~n16288 ;
  assign n16290 = n16286 & n16289 ;
  assign n16291 = n8866 & ~n16290 ;
  assign n16292 = ~n16283 & ~n16291 ;
  assign n16293 = n16274 & n16292 ;
  assign n16294 = \u4_u3_buf0_reg[20]/P0001  & n2568 ;
  assign n16295 = \u4_u3_csr1_reg[5]/P0001  & n8816 ;
  assign n16296 = ~n16294 & ~n16295 ;
  assign n16297 = \u4_u3_buf1_reg[20]/P0001  & n2731 ;
  assign n16298 = \u4_u3_ienb_reg[4]/P0001  & n8820 ;
  assign n16299 = ~n16297 & ~n16298 ;
  assign n16300 = n16296 & n16299 ;
  assign n16301 = n8836 & ~n16300 ;
  assign n16302 = \u4_u2_csr1_reg[5]/P0001  & n8816 ;
  assign n16303 = \u4_u2_buf1_reg[20]/P0001  & n2731 ;
  assign n16304 = ~n16302 & ~n16303 ;
  assign n16305 = \u4_u2_ienb_reg[4]/P0001  & n8820 ;
  assign n16306 = \u4_u2_buf0_reg[20]/P0001  & n2568 ;
  assign n16307 = ~n16305 & ~n16306 ;
  assign n16308 = n16304 & n16307 ;
  assign n16309 = n8826 & ~n16308 ;
  assign n16310 = ~n16301 & ~n16309 ;
  assign n16311 = \u4_u0_csr1_reg[5]/P0001  & n8816 ;
  assign n16312 = \u4_u0_buf1_reg[20]/P0001  & n2731 ;
  assign n16313 = ~n16311 & ~n16312 ;
  assign n16314 = \u4_u0_ienb_reg[4]/P0001  & n8820 ;
  assign n16315 = \u4_u0_buf0_reg[20]/P0001  & n2568 ;
  assign n16316 = ~n16314 & ~n16315 ;
  assign n16317 = n16313 & n16316 ;
  assign n16318 = n8815 & ~n16317 ;
  assign n16319 = n16310 & ~n16318 ;
  assign n16320 = \u1_frame_no_r_reg[4]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16321 = n8816 & n16320 ;
  assign n16322 = \u4_intb_msk_reg[4]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16323 = n2568 & n16322 ;
  assign n16324 = \u4_int_srcb_reg[0]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16325 = n2731 & n16324 ;
  assign n16326 = ~n16323 & ~n16325 ;
  assign n16327 = ~n16321 & n16326 ;
  assign n16328 = n8864 & ~n16327 ;
  assign n16329 = \u4_u1_csr1_reg[5]/P0001  & n8816 ;
  assign n16330 = \u4_u1_buf1_reg[20]/P0001  & n2731 ;
  assign n16331 = ~n16329 & ~n16330 ;
  assign n16332 = \u4_u1_ienb_reg[4]/P0001  & n8820 ;
  assign n16333 = \u4_u1_buf0_reg[20]/P0001  & n2568 ;
  assign n16334 = ~n16332 & ~n16333 ;
  assign n16335 = n16331 & n16334 ;
  assign n16336 = n8866 & ~n16335 ;
  assign n16337 = ~n16328 & ~n16336 ;
  assign n16338 = n16319 & n16337 ;
  assign n16339 = \u1_u3_out_to_small_reg/P0001  & \u4_u3_ep_match_r_reg/P0001  ;
  assign n16340 = ~\u4_u3_int_stat_reg[6]/P0001  & ~n16339 ;
  assign n16341 = n5455 & ~n16340 ;
  assign n16342 = ~n6195 & ~n6198 ;
  assign n16343 = n5748 & n6178 ;
  assign n16344 = n16342 & n16343 ;
  assign n16345 = n6132 & n16344 ;
  assign n16346 = \u0_u0_state_reg[2]/NET0131  & ~n8668 ;
  assign n16347 = ~n6150 & n16346 ;
  assign n16348 = ~n6147 & ~n16347 ;
  assign n16349 = n5748 & ~n16348 ;
  assign n16350 = n6134 & n16349 ;
  assign n16351 = ~n16345 & ~n16350 ;
  assign n16352 = \u4_u3_buf0_reg[5]/P0001  & n2568 ;
  assign n16353 = \u4_u3_csr0_reg[5]/P0001  & n8816 ;
  assign n16354 = ~n16352 & ~n16353 ;
  assign n16355 = \u4_u3_buf1_reg[5]/P0001  & n2731 ;
  assign n16356 = \u4_u3_int_stat_reg[5]/P0001  & n8820 ;
  assign n16357 = ~n16355 & ~n16356 ;
  assign n16358 = n16354 & n16357 ;
  assign n16359 = n8836 & ~n16358 ;
  assign n16360 = \u4_u2_csr0_reg[5]/P0001  & n8816 ;
  assign n16361 = \u4_u2_buf1_reg[5]/P0001  & n2731 ;
  assign n16362 = ~n16360 & ~n16361 ;
  assign n16363 = \u4_u2_int_stat_reg[5]/P0001  & n8820 ;
  assign n16364 = \u4_u2_buf0_reg[5]/P0001  & n2568 ;
  assign n16365 = ~n16363 & ~n16364 ;
  assign n16366 = n16362 & n16365 ;
  assign n16367 = n8826 & ~n16366 ;
  assign n16368 = ~n16359 & ~n16367 ;
  assign n16369 = \u4_u0_csr0_reg[5]/P0001  & n8816 ;
  assign n16370 = \u4_u0_buf1_reg[5]/P0001  & n2731 ;
  assign n16371 = ~n16369 & ~n16370 ;
  assign n16372 = \u4_u0_int_stat_reg[5]/P0001  & n8820 ;
  assign n16373 = \u4_u0_buf0_reg[5]/P0001  & n2568 ;
  assign n16374 = ~n16372 & ~n16373 ;
  assign n16375 = n16371 & n16374 ;
  assign n16376 = n8815 & ~n16375 ;
  assign n16377 = n16368 & ~n16376 ;
  assign n16378 = \u1_sof_time_reg[5]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16379 = n8816 & n16378 ;
  assign n16380 = \u4_funct_adr_reg[5]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16381 = n8820 & n16380 ;
  assign n16382 = ~n16379 & ~n16381 ;
  assign n16383 = \u4_utmi_vend_stat_r_reg[5]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16384 = n8820 & n16383 ;
  assign n16385 = \u4_inta_msk_reg[5]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16386 = n2568 & n16385 ;
  assign n16387 = ~n16384 & ~n16386 ;
  assign n16388 = n16382 & n16387 ;
  assign n16389 = n8864 & ~n16388 ;
  assign n16390 = \u4_u1_csr0_reg[5]/P0001  & n8816 ;
  assign n16391 = \u4_u1_buf1_reg[5]/P0001  & n2731 ;
  assign n16392 = ~n16390 & ~n16391 ;
  assign n16393 = \u4_u1_int_stat_reg[5]/P0001  & n8820 ;
  assign n16394 = \u4_u1_buf0_reg[5]/P0001  & n2568 ;
  assign n16395 = ~n16393 & ~n16394 ;
  assign n16396 = n16392 & n16395 ;
  assign n16397 = n8866 & ~n16396 ;
  assign n16398 = ~n16389 & ~n16397 ;
  assign n16399 = n16377 & n16398 ;
  assign n16400 = \u4_u3_buf0_reg[6]/P0001  & n2568 ;
  assign n16401 = \u4_u3_csr0_reg[6]/P0001  & n8816 ;
  assign n16402 = ~n16400 & ~n16401 ;
  assign n16403 = \u4_u3_buf1_reg[6]/P0001  & n2731 ;
  assign n16404 = \u4_u3_int_stat_reg[6]/P0001  & n8820 ;
  assign n16405 = ~n16403 & ~n16404 ;
  assign n16406 = n16402 & n16405 ;
  assign n16407 = n8836 & ~n16406 ;
  assign n16408 = \u4_u2_csr0_reg[6]/P0001  & n8816 ;
  assign n16409 = \u4_u2_buf1_reg[6]/P0001  & n2731 ;
  assign n16410 = ~n16408 & ~n16409 ;
  assign n16411 = \u4_u2_int_stat_reg[6]/P0001  & n8820 ;
  assign n16412 = \u4_u2_buf0_reg[6]/P0001  & n2568 ;
  assign n16413 = ~n16411 & ~n16412 ;
  assign n16414 = n16410 & n16413 ;
  assign n16415 = n8826 & ~n16414 ;
  assign n16416 = ~n16407 & ~n16415 ;
  assign n16417 = \u4_u0_csr0_reg[6]/P0001  & n8816 ;
  assign n16418 = \u4_u0_buf1_reg[6]/P0001  & n2731 ;
  assign n16419 = ~n16417 & ~n16418 ;
  assign n16420 = \u4_u0_int_stat_reg[6]/P0001  & n8820 ;
  assign n16421 = \u4_u0_buf0_reg[6]/P0001  & n2568 ;
  assign n16422 = ~n16420 & ~n16421 ;
  assign n16423 = n16419 & n16422 ;
  assign n16424 = n8815 & ~n16423 ;
  assign n16425 = n16416 & ~n16424 ;
  assign n16426 = \u4_funct_adr_reg[6]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16427 = n8820 & n16426 ;
  assign n16428 = \u1_sof_time_reg[6]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16429 = n8816 & n16428 ;
  assign n16430 = ~n16427 & ~n16429 ;
  assign n16431 = \u4_utmi_vend_stat_r_reg[6]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16432 = n8820 & n16431 ;
  assign n16433 = \u4_inta_msk_reg[6]/P0001  & ~\wb_addr_i[4]_pad  ;
  assign n16434 = n2568 & n16433 ;
  assign n16435 = ~n16432 & ~n16434 ;
  assign n16436 = n16430 & n16435 ;
  assign n16437 = n8864 & ~n16436 ;
  assign n16438 = \u4_u1_csr0_reg[6]/P0001  & n8816 ;
  assign n16439 = \u4_u1_buf1_reg[6]/P0001  & n2731 ;
  assign n16440 = ~n16438 & ~n16439 ;
  assign n16441 = \u4_u1_int_stat_reg[6]/P0001  & n8820 ;
  assign n16442 = \u4_u1_buf0_reg[6]/P0001  & n2568 ;
  assign n16443 = ~n16441 & ~n16442 ;
  assign n16444 = n16440 & n16443 ;
  assign n16445 = n8866 & ~n16444 ;
  assign n16446 = ~n16437 & ~n16445 ;
  assign n16447 = n16425 & n16446 ;
  assign n16448 = ~\u5_state_reg[3]/P0001  & ~\u5_wb_req_s1_reg/P0001  ;
  assign n16449 = rst_i_pad & ~n8183 ;
  assign n16450 = ~n16448 & n16449 ;
  assign n16451 = n8182 & n16450 ;
  assign n16452 = \sram_data_i[14]_pad  & \wb_addr_i[17]_pad  ;
  assign n16453 = \u4_dout_reg[14]/P0001  & ~\wb_addr_i[17]_pad  ;
  assign n16454 = ~n16452 & ~n16453 ;
  assign n16455 = ~n9218 & ~n9229 ;
  assign n16456 = ~n9228 & n16455 ;
  assign n16457 = ~n9217 & ~n9234 ;
  assign n16458 = ~n9220 & ~n16457 ;
  assign n16459 = ~n16456 & n16458 ;
  assign n16460 = n9220 & n16457 ;
  assign n16461 = n16455 & n16457 ;
  assign n16462 = ~n9228 & n16461 ;
  assign n16463 = ~n16460 & ~n16462 ;
  assign n16464 = ~n16459 & n16463 ;
  assign n16465 = ~n9215 & ~n9240 ;
  assign n16466 = ~n14352 & n16465 ;
  assign n16467 = ~n9211 & ~n9239 ;
  assign n16468 = ~n9214 & ~n16467 ;
  assign n16469 = ~n16466 & n16468 ;
  assign n16470 = n9214 & n16467 ;
  assign n16471 = n16465 & n16467 ;
  assign n16472 = ~n14352 & n16471 ;
  assign n16473 = ~n16470 & ~n16472 ;
  assign n16474 = ~n16469 & n16473 ;
  assign n16475 = ~n9071 & ~n9082 ;
  assign n16476 = ~n9081 & n16475 ;
  assign n16477 = ~n9070 & ~n9087 ;
  assign n16478 = ~n9073 & ~n16477 ;
  assign n16479 = ~n16476 & n16478 ;
  assign n16480 = n9073 & n16477 ;
  assign n16481 = n16475 & n16477 ;
  assign n16482 = ~n9081 & n16481 ;
  assign n16483 = ~n16480 & ~n16482 ;
  assign n16484 = ~n16479 & n16483 ;
  assign n16485 = ~n9068 & ~n9093 ;
  assign n16486 = ~n14361 & n16485 ;
  assign n16487 = ~n9064 & ~n9092 ;
  assign n16488 = ~n9067 & ~n16487 ;
  assign n16489 = ~n16486 & n16488 ;
  assign n16490 = n9067 & n16487 ;
  assign n16491 = n16485 & n16487 ;
  assign n16492 = ~n14361 & n16491 ;
  assign n16493 = ~n16490 & ~n16492 ;
  assign n16494 = ~n16489 & n16493 ;
  assign n16495 = ~n9120 & ~n9131 ;
  assign n16496 = ~n9130 & n16495 ;
  assign n16497 = ~n9119 & ~n9136 ;
  assign n16498 = ~n9122 & ~n16497 ;
  assign n16499 = ~n16496 & n16498 ;
  assign n16500 = n9122 & n16497 ;
  assign n16501 = n16495 & n16497 ;
  assign n16502 = ~n9130 & n16501 ;
  assign n16503 = ~n16500 & ~n16502 ;
  assign n16504 = ~n16499 & n16503 ;
  assign n16505 = ~n9117 & ~n9142 ;
  assign n16506 = ~n14370 & n16505 ;
  assign n16507 = ~n9113 & ~n9141 ;
  assign n16508 = ~n9116 & ~n16507 ;
  assign n16509 = ~n16506 & n16508 ;
  assign n16510 = n9116 & n16507 ;
  assign n16511 = n16505 & n16507 ;
  assign n16512 = ~n14370 & n16511 ;
  assign n16513 = ~n16510 & ~n16512 ;
  assign n16514 = ~n16509 & n16513 ;
  assign n16515 = ~n9169 & ~n9180 ;
  assign n16516 = ~n9179 & n16515 ;
  assign n16517 = ~n9168 & ~n9185 ;
  assign n16518 = ~n9171 & ~n16517 ;
  assign n16519 = ~n16516 & n16518 ;
  assign n16520 = n9171 & n16517 ;
  assign n16521 = n16515 & n16517 ;
  assign n16522 = ~n9179 & n16521 ;
  assign n16523 = ~n16520 & ~n16522 ;
  assign n16524 = ~n16519 & n16523 ;
  assign n16525 = ~n9166 & ~n9191 ;
  assign n16526 = ~n14379 & n16525 ;
  assign n16527 = ~n9162 & ~n9190 ;
  assign n16528 = ~n9165 & ~n16527 ;
  assign n16529 = ~n16526 & n16528 ;
  assign n16530 = n9165 & n16527 ;
  assign n16531 = n16525 & n16527 ;
  assign n16532 = ~n14379 & n16531 ;
  assign n16533 = ~n16530 & ~n16532 ;
  assign n16534 = ~n16529 & n16533 ;
  assign n16535 = rst_i_pad & \u0_tx_ready_reg/NET0131  ;
  assign n16536 = n1850 & n16535 ;
  assign n16537 = n1835 & n16536 ;
  assign n16538 = rst_i_pad & ~\u0_tx_ready_reg/NET0131  ;
  assign n16539 = n1834 & n16538 ;
  assign n16540 = n1838 & n16539 ;
  assign n16541 = ~n16537 & ~n16540 ;
  assign n16542 = ~\u0_u0_state_reg[3]/P0001  & ~n6157 ;
  assign n16543 = ~n15506 & n16542 ;
  assign n16544 = ~n15499 & ~n16543 ;
  assign n16545 = \u4_u1_csr0_reg[10]/P0001  & n8816 ;
  assign n16546 = \u4_u1_buf1_reg[10]/P0001  & n2731 ;
  assign n16547 = \u4_u1_buf0_reg[10]/P0001  & n2568 ;
  assign n16548 = ~n16546 & ~n16547 ;
  assign n16549 = ~n16545 & n16548 ;
  assign n16550 = n8866 & ~n16549 ;
  assign n16551 = \u4_u3_csr0_reg[10]/P0001  & n8816 ;
  assign n16552 = \u4_u3_buf1_reg[10]/P0001  & n2731 ;
  assign n16553 = \u4_u3_buf0_reg[10]/P0001  & n2568 ;
  assign n16554 = ~n16552 & ~n16553 ;
  assign n16555 = ~n16551 & n16554 ;
  assign n16556 = n8836 & ~n16555 ;
  assign n16557 = ~n16550 & ~n16556 ;
  assign n16558 = \u1_sof_time_reg[10]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16559 = n8816 & n16558 ;
  assign n16560 = n8864 & n16559 ;
  assign n16561 = \u4_u0_csr0_reg[10]/P0001  & n8816 ;
  assign n16562 = \u4_u0_buf1_reg[10]/P0001  & n2731 ;
  assign n16563 = \u4_u0_buf0_reg[10]/P0001  & n2568 ;
  assign n16564 = ~n16562 & ~n16563 ;
  assign n16565 = ~n16561 & n16564 ;
  assign n16566 = n8815 & ~n16565 ;
  assign n16567 = ~n16560 & ~n16566 ;
  assign n16568 = \u4_u2_csr0_reg[10]/P0001  & n8816 ;
  assign n16569 = \u4_u2_buf1_reg[10]/P0001  & n2731 ;
  assign n16570 = \u4_u2_buf0_reg[10]/P0001  & n2568 ;
  assign n16571 = ~n16569 & ~n16570 ;
  assign n16572 = ~n16568 & n16571 ;
  assign n16573 = n8826 & ~n16572 ;
  assign n16574 = n16567 & ~n16573 ;
  assign n16575 = n16557 & n16574 ;
  assign n16576 = \u4_u1_csr0_reg[11]/P0001  & n8816 ;
  assign n16577 = \u4_u1_buf1_reg[11]/P0001  & n2731 ;
  assign n16578 = \u4_u1_buf0_reg[11]/P0001  & n2568 ;
  assign n16579 = ~n16577 & ~n16578 ;
  assign n16580 = ~n16576 & n16579 ;
  assign n16581 = n8866 & ~n16580 ;
  assign n16582 = \u4_u3_csr0_reg[11]/P0001  & n8816 ;
  assign n16583 = \u4_u3_buf1_reg[11]/P0001  & n2731 ;
  assign n16584 = \u4_u3_buf0_reg[11]/P0001  & n2568 ;
  assign n16585 = ~n16583 & ~n16584 ;
  assign n16586 = ~n16582 & n16585 ;
  assign n16587 = n8836 & ~n16586 ;
  assign n16588 = ~n16581 & ~n16587 ;
  assign n16589 = \u1_sof_time_reg[11]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16590 = n8816 & n16589 ;
  assign n16591 = n8864 & n16590 ;
  assign n16592 = \u4_u0_csr0_reg[11]/P0001  & n8816 ;
  assign n16593 = \u4_u0_buf1_reg[11]/P0001  & n2731 ;
  assign n16594 = \u4_u0_buf0_reg[11]/P0001  & n2568 ;
  assign n16595 = ~n16593 & ~n16594 ;
  assign n16596 = ~n16592 & n16595 ;
  assign n16597 = n8815 & ~n16596 ;
  assign n16598 = ~n16591 & ~n16597 ;
  assign n16599 = \u4_u2_csr0_reg[11]/P0001  & n8816 ;
  assign n16600 = \u4_u2_buf1_reg[11]/P0001  & n2731 ;
  assign n16601 = \u4_u2_buf0_reg[11]/P0001  & n2568 ;
  assign n16602 = ~n16600 & ~n16601 ;
  assign n16603 = ~n16599 & n16602 ;
  assign n16604 = n8826 & ~n16603 ;
  assign n16605 = n16598 & ~n16604 ;
  assign n16606 = n16588 & n16605 ;
  assign n16607 = \u4_u1_csr0_reg[9]/P0001  & n8816 ;
  assign n16608 = \u4_u1_buf1_reg[9]/P0001  & n2731 ;
  assign n16609 = \u4_u1_buf0_reg[9]/P0001  & n2568 ;
  assign n16610 = ~n16608 & ~n16609 ;
  assign n16611 = ~n16607 & n16610 ;
  assign n16612 = n8866 & ~n16611 ;
  assign n16613 = \u4_u3_csr0_reg[9]/P0001  & n8816 ;
  assign n16614 = \u4_u3_buf1_reg[9]/P0001  & n2731 ;
  assign n16615 = \u4_u3_buf0_reg[9]/P0001  & n2568 ;
  assign n16616 = ~n16614 & ~n16615 ;
  assign n16617 = ~n16613 & n16616 ;
  assign n16618 = n8836 & ~n16617 ;
  assign n16619 = ~n16612 & ~n16618 ;
  assign n16620 = \u1_sof_time_reg[9]/P0001  & \wb_addr_i[4]_pad  ;
  assign n16621 = n8816 & n16620 ;
  assign n16622 = n8864 & n16621 ;
  assign n16623 = \u4_u0_csr0_reg[9]/P0001  & n8816 ;
  assign n16624 = \u4_u0_buf1_reg[9]/P0001  & n2731 ;
  assign n16625 = \u4_u0_buf0_reg[9]/P0001  & n2568 ;
  assign n16626 = ~n16624 & ~n16625 ;
  assign n16627 = ~n16623 & n16626 ;
  assign n16628 = n8815 & ~n16627 ;
  assign n16629 = ~n16622 & ~n16628 ;
  assign n16630 = \u4_u2_csr0_reg[9]/P0001  & n8816 ;
  assign n16631 = \u4_u2_buf1_reg[9]/P0001  & n2731 ;
  assign n16632 = \u4_u2_buf0_reg[9]/P0001  & n2568 ;
  assign n16633 = ~n16631 & ~n16632 ;
  assign n16634 = ~n16630 & n16633 ;
  assign n16635 = n8826 & ~n16634 ;
  assign n16636 = n16629 & ~n16635 ;
  assign n16637 = n16619 & n16636 ;
  assign n16638 = \u1_u3_rx_ack_to_cnt_reg[4]/P0001  & \u1_u3_rx_ack_to_cnt_reg[5]/P0001  ;
  assign n16639 = n12632 & n16638 ;
  assign n16640 = ~\u1_u3_rx_ack_to_cnt_reg[6]/P0001  & ~n16639 ;
  assign n16641 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & ~n14218 ;
  assign n16642 = ~n16640 & n16641 ;
  assign n16643 = \u1_u3_tx_data_to_cnt_reg[4]/P0001  & \u1_u3_tx_data_to_cnt_reg[5]/P0001  ;
  assign n16644 = n12665 & n16643 ;
  assign n16645 = ~\u1_u3_tx_data_to_cnt_reg[6]/P0001  & ~n16644 ;
  assign n16646 = ~\u0_rx_active_reg/P0001  & ~n14228 ;
  assign n16647 = ~n16645 & n16646 ;
  assign n16648 = ~\u0_u0_state_reg[6]/NET0131  & ~n5765 ;
  assign n16649 = n6144 & ~n16648 ;
  assign n16650 = n6143 & n16649 ;
  assign n16651 = ~\u0_u0_T2_gt_100_uS_reg/P0001  & n12655 ;
  assign n16652 = n12653 & n16651 ;
  assign n16653 = ~n16650 & ~n16652 ;
  assign n16654 = n5748 & ~n16653 ;
  assign n16655 = ~\u4_u3_buf0_orig_reg[21]/P0001  & ~n12409 ;
  assign n16656 = \u4_u3_buf0_orig_reg[22]/P0001  & ~n16655 ;
  assign n16657 = ~n12411 & ~n16656 ;
  assign n16658 = \u5_wb_req_s1_reg/P0001  & ~wb_we_i_pad ;
  assign n16659 = ~\wb_addr_i[4]_pad  & n2731 ;
  assign n16660 = n8864 & n16659 ;
  assign n16661 = n2560 & n16660 ;
  assign n16662 = n16658 & n16661 ;
  assign n16663 = ~\u4_u0_buf0_orig_reg[21]/P0001  & ~n12439 ;
  assign n16664 = \u4_u0_buf0_orig_reg[22]/P0001  & ~n16663 ;
  assign n16665 = ~n12441 & ~n16664 ;
  assign n16666 = ~\u4_u1_buf0_orig_reg[21]/P0001  & ~n12462 ;
  assign n16667 = \u4_u1_buf0_orig_reg[22]/P0001  & ~n16666 ;
  assign n16668 = ~n12464 & ~n16667 ;
  assign n16669 = ~\u4_u2_buf0_orig_reg[21]/P0001  & ~n12485 ;
  assign n16670 = \u4_u2_buf0_orig_reg[22]/P0001  & ~n16669 ;
  assign n16671 = ~n12487 & ~n16670 ;
  assign n16672 = \u0_u0_idle_cnt1_reg[2]/P0001  & n11227 ;
  assign n16673 = ~\u0_u0_idle_cnt1_reg[3]/P0001  & ~n16672 ;
  assign n16674 = ~n14315 & ~n16673 ;
  assign n16675 = ~n9166 & ~n9184 ;
  assign n16676 = ~n9185 & ~n16675 ;
  assign n16677 = n9183 & n16676 ;
  assign n16678 = n9183 & ~n9185 ;
  assign n16679 = n16675 & ~n16678 ;
  assign n16680 = ~n16677 & ~n16679 ;
  assign n16681 = ~n9068 & ~n9086 ;
  assign n16682 = ~n9087 & ~n16681 ;
  assign n16683 = n9085 & n16682 ;
  assign n16684 = n9085 & ~n9087 ;
  assign n16685 = n16681 & ~n16684 ;
  assign n16686 = ~n16683 & ~n16685 ;
  assign n16687 = ~n9117 & ~n9135 ;
  assign n16688 = ~n9136 & ~n16687 ;
  assign n16689 = n9134 & n16688 ;
  assign n16690 = n9134 & ~n9136 ;
  assign n16691 = n16687 & ~n16690 ;
  assign n16692 = ~n16689 & ~n16691 ;
  assign n16693 = ~n9215 & ~n9233 ;
  assign n16694 = ~n9234 & ~n16693 ;
  assign n16695 = n9232 & n16694 ;
  assign n16696 = n9232 & ~n9234 ;
  assign n16697 = n16693 & ~n16696 ;
  assign n16698 = ~n16695 & ~n16697 ;
  assign n16699 = \u4_buf0_reg[13]/P0001  & \u4_buf0_reg[14]/P0001  ;
  assign n16700 = \u4_buf0_reg[11]/P0001  & n16699 ;
  assign n16701 = \u4_buf0_reg[0]/P0001  & \u4_buf0_reg[10]/P0001  ;
  assign n16702 = \u4_buf0_reg[12]/P0001  & n16701 ;
  assign n16703 = n16700 & n16702 ;
  assign n16704 = \u4_buf0_reg[5]/P0001  & \u4_buf0_reg[6]/P0001  ;
  assign n16705 = \u4_buf0_reg[3]/P0001  & \u4_buf0_reg[4]/P0001  ;
  assign n16706 = n16704 & n16705 ;
  assign n16707 = \u4_buf0_reg[1]/P0001  & \u4_buf0_reg[2]/P0001  ;
  assign n16708 = \u4_buf0_reg[15]/P0001  & \u4_buf0_reg[16]/P0001  ;
  assign n16709 = n16707 & n16708 ;
  assign n16710 = n16706 & n16709 ;
  assign n16711 = \u4_buf0_reg[7]/P0001  & \u4_buf0_reg[8]/P0001  ;
  assign n16712 = \u4_buf0_reg[9]/P0001  & n16711 ;
  assign n16713 = n16710 & n16712 ;
  assign n16714 = n16703 & n16713 ;
  assign n16715 = ~\u4_buf0_reg[31]/P0001  & ~n16714 ;
  assign n16716 = \u4_buf1_reg[13]/P0001  & \u4_buf1_reg[14]/P0001  ;
  assign n16717 = \u4_buf1_reg[11]/P0001  & n16716 ;
  assign n16718 = \u4_buf1_reg[0]/P0001  & \u4_buf1_reg[10]/P0001  ;
  assign n16719 = \u4_buf1_reg[12]/P0001  & n16718 ;
  assign n16720 = n16717 & n16719 ;
  assign n16721 = \u4_buf1_reg[5]/P0001  & \u4_buf1_reg[6]/P0001  ;
  assign n16722 = \u4_buf1_reg[3]/P0001  & \u4_buf1_reg[4]/P0001  ;
  assign n16723 = n16721 & n16722 ;
  assign n16724 = \u4_buf1_reg[1]/P0001  & \u4_buf1_reg[2]/P0001  ;
  assign n16725 = \u4_buf1_reg[15]/P0001  & \u4_buf1_reg[16]/P0001  ;
  assign n16726 = n16724 & n16725 ;
  assign n16727 = n16723 & n16726 ;
  assign n16728 = \u4_buf1_reg[7]/P0001  & \u4_buf1_reg[8]/P0001  ;
  assign n16729 = \u4_buf1_reg[9]/P0001  & n16728 ;
  assign n16730 = n16727 & n16729 ;
  assign n16731 = n16720 & n16730 ;
  assign n16732 = ~\u4_buf1_reg[31]/P0001  & ~n16731 ;
  assign n16733 = ~\u1_u0_state_reg[2]/P0001  & n7207 ;
  assign n16734 = ~\u0_rx_data_reg[0]/P0001  & n7202 ;
  assign n16735 = n16733 & n16734 ;
  assign n16736 = rst_i_pad & \u1_u0_pid_reg[0]/NET0131  ;
  assign n16737 = rst_i_pad & n7202 ;
  assign n16738 = n16733 & n16737 ;
  assign n16739 = ~n16736 & ~n16738 ;
  assign n16740 = ~n16735 & ~n16739 ;
  assign n16741 = ~\u0_rx_data_reg[1]/P0001  & n7202 ;
  assign n16742 = n16733 & n16741 ;
  assign n16743 = rst_i_pad & \u1_u0_pid_reg[1]/NET0131  ;
  assign n16744 = ~n16738 & ~n16743 ;
  assign n16745 = ~n16742 & ~n16744 ;
  assign n16746 = ~\u0_rx_data_reg[2]/P0001  & n7202 ;
  assign n16747 = n16733 & n16746 ;
  assign n16748 = rst_i_pad & \u1_u0_pid_reg[2]/NET0131  ;
  assign n16749 = ~n16738 & ~n16748 ;
  assign n16750 = ~n16747 & ~n16749 ;
  assign n16751 = ~\u0_rx_data_reg[3]/P0001  & n7202 ;
  assign n16752 = n16733 & n16751 ;
  assign n16753 = rst_i_pad & \u1_u0_pid_reg[3]/NET0131  ;
  assign n16754 = ~n16738 & ~n16753 ;
  assign n16755 = ~n16752 & ~n16754 ;
  assign n16756 = \u4_u0_csr0_reg[12]/P0001  & n8816 ;
  assign n16757 = \u4_u0_buf1_reg[12]/P0001  & n2731 ;
  assign n16758 = \u4_u0_buf0_reg[12]/P0001  & n2568 ;
  assign n16759 = ~n16757 & ~n16758 ;
  assign n16760 = ~n16756 & n16759 ;
  assign n16761 = n8815 & ~n16760 ;
  assign n16762 = \u4_u3_csr0_reg[12]/P0001  & n8816 ;
  assign n16763 = \u4_u3_buf1_reg[12]/P0001  & n2731 ;
  assign n16764 = \u4_u3_buf0_reg[12]/P0001  & n2568 ;
  assign n16765 = ~n16763 & ~n16764 ;
  assign n16766 = ~n16762 & n16765 ;
  assign n16767 = n8836 & ~n16766 ;
  assign n16768 = ~n16761 & ~n16767 ;
  assign n16769 = \u4_u2_csr0_reg[12]/P0001  & n8816 ;
  assign n16770 = \u4_u2_buf1_reg[12]/P0001  & n2731 ;
  assign n16771 = \u4_u2_buf0_reg[12]/P0001  & n2568 ;
  assign n16772 = ~n16770 & ~n16771 ;
  assign n16773 = ~n16769 & n16772 ;
  assign n16774 = n8826 & ~n16773 ;
  assign n16775 = \u4_u1_csr0_reg[12]/P0001  & n8816 ;
  assign n16776 = \u4_u1_buf1_reg[12]/P0001  & n2731 ;
  assign n16777 = \u4_u1_buf0_reg[12]/P0001  & n2568 ;
  assign n16778 = ~n16776 & ~n16777 ;
  assign n16779 = ~n16775 & n16778 ;
  assign n16780 = n8866 & ~n16779 ;
  assign n16781 = ~n16774 & ~n16780 ;
  assign n16782 = n16768 & n16781 ;
  assign n16783 = \u4_u2_ots_stop_reg/P0001  & n8816 ;
  assign n16784 = \u4_u2_buf1_reg[13]/P0001  & n2731 ;
  assign n16785 = \u4_u2_buf0_reg[13]/P0001  & n2568 ;
  assign n16786 = ~n16784 & ~n16785 ;
  assign n16787 = ~n16783 & n16786 ;
  assign n16788 = n8826 & ~n16787 ;
  assign n16789 = \u4_u0_ots_stop_reg/P0001  & n8816 ;
  assign n16790 = \u4_u0_buf1_reg[13]/P0001  & n2731 ;
  assign n16791 = \u4_u0_buf0_reg[13]/P0001  & n2568 ;
  assign n16792 = ~n16790 & ~n16791 ;
  assign n16793 = ~n16789 & n16792 ;
  assign n16794 = n8815 & ~n16793 ;
  assign n16795 = ~n16788 & ~n16794 ;
  assign n16796 = \u4_u3_ots_stop_reg/P0001  & n8816 ;
  assign n16797 = \u4_u3_buf1_reg[13]/P0001  & n2731 ;
  assign n16798 = \u4_u3_buf0_reg[13]/P0001  & n2568 ;
  assign n16799 = ~n16797 & ~n16798 ;
  assign n16800 = ~n16796 & n16799 ;
  assign n16801 = n8836 & ~n16800 ;
  assign n16802 = \u4_u1_ots_stop_reg/P0001  & n8816 ;
  assign n16803 = \u4_u1_buf1_reg[13]/P0001  & n2731 ;
  assign n16804 = \u4_u1_buf0_reg[13]/P0001  & n2568 ;
  assign n16805 = ~n16803 & ~n16804 ;
  assign n16806 = ~n16802 & n16805 ;
  assign n16807 = n8866 & ~n16806 ;
  assign n16808 = ~n16801 & ~n16807 ;
  assign n16809 = n16795 & n16808 ;
  assign n16810 = \u4_u2_csr1_reg[0]/P0001  & n8816 ;
  assign n16811 = \u4_u2_buf1_reg[15]/P0001  & n2731 ;
  assign n16812 = \u4_u2_buf0_reg[15]/P0001  & n2568 ;
  assign n16813 = ~n16811 & ~n16812 ;
  assign n16814 = ~n16810 & n16813 ;
  assign n16815 = n8826 & ~n16814 ;
  assign n16816 = \u4_u0_csr1_reg[0]/P0001  & n8816 ;
  assign n16817 = \u4_u0_buf1_reg[15]/P0001  & n2731 ;
  assign n16818 = \u4_u0_buf0_reg[15]/P0001  & n2568 ;
  assign n16819 = ~n16817 & ~n16818 ;
  assign n16820 = ~n16816 & n16819 ;
  assign n16821 = n8815 & ~n16820 ;
  assign n16822 = ~n16815 & ~n16821 ;
  assign n16823 = \u4_u3_csr1_reg[0]/P0001  & n8816 ;
  assign n16824 = \u4_u3_buf1_reg[15]/P0001  & n2731 ;
  assign n16825 = \u4_u3_buf0_reg[15]/P0001  & n2568 ;
  assign n16826 = ~n16824 & ~n16825 ;
  assign n16827 = ~n16823 & n16826 ;
  assign n16828 = n8836 & ~n16827 ;
  assign n16829 = \u4_u1_csr1_reg[0]/P0001  & n8816 ;
  assign n16830 = \u4_u1_buf1_reg[15]/P0001  & n2731 ;
  assign n16831 = \u4_u1_buf0_reg[15]/P0001  & n2568 ;
  assign n16832 = ~n16830 & ~n16831 ;
  assign n16833 = ~n16829 & n16832 ;
  assign n16834 = n8866 & ~n16833 ;
  assign n16835 = ~n16828 & ~n16834 ;
  assign n16836 = n16822 & n16835 ;
  assign n16837 = \u1_u3_rx_ack_to_cnt_reg[4]/P0001  & n12632 ;
  assign n16838 = ~\u1_u3_rx_ack_to_cnt_reg[5]/P0001  & ~n16837 ;
  assign n16839 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & ~n16639 ;
  assign n16840 = ~n16838 & n16839 ;
  assign n16841 = n7202 & n16733 ;
  assign n16842 = \u1_u0_pid_reg[4]/P0001  & ~n16841 ;
  assign n16843 = \u0_rx_data_reg[4]/P0001  & n7202 ;
  assign n16844 = n16733 & n16843 ;
  assign n16845 = rst_i_pad & ~n16844 ;
  assign n16846 = ~n16842 & n16845 ;
  assign n16847 = \u1_u0_pid_reg[5]/P0001  & ~n16841 ;
  assign n16848 = \u0_rx_data_reg[5]/P0001  & n7202 ;
  assign n16849 = n16733 & n16848 ;
  assign n16850 = rst_i_pad & ~n16849 ;
  assign n16851 = ~n16847 & n16850 ;
  assign n16852 = \u1_u0_pid_reg[6]/P0001  & ~n16841 ;
  assign n16853 = \u0_rx_data_reg[6]/P0001  & n7202 ;
  assign n16854 = n16733 & n16853 ;
  assign n16855 = rst_i_pad & ~n16854 ;
  assign n16856 = ~n16852 & n16855 ;
  assign n16857 = \u1_u0_pid_reg[7]/P0001  & ~n16841 ;
  assign n16858 = \u0_rx_data_reg[7]/P0001  & n7202 ;
  assign n16859 = n16733 & n16858 ;
  assign n16860 = rst_i_pad & ~n16859 ;
  assign n16861 = ~n16857 & n16860 ;
  assign n16862 = n7198 & n7200 ;
  assign n16863 = ~\u1_u0_token_valid_r1_reg/P0001  & ~n16862 ;
  assign n16864 = n8820 & n16658 ;
  assign n16865 = n2560 & n16864 ;
  assign n16866 = n8815 & n16865 ;
  assign n16867 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & \u1_u3_rx_ack_to_cnt_reg[2]/P0001  ;
  assign n16868 = ~n12630 & n16867 ;
  assign n16869 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & ~\u1_u3_rx_ack_to_cnt_reg[2]/P0001  ;
  assign n16870 = \u1_u3_rx_ack_to_cnt_reg[0]/P0001  & \u1_u3_rx_ack_to_cnt_reg[1]/P0001  ;
  assign n16871 = n16869 & n16870 ;
  assign n16872 = ~n16868 & ~n16871 ;
  assign n16873 = ~\u0_rx_active_reg/P0001  & \u1_u3_tx_data_to_cnt_reg[2]/P0001  ;
  assign n16874 = ~n12663 & n16873 ;
  assign n16875 = ~\u0_rx_active_reg/P0001  & ~\u1_u3_tx_data_to_cnt_reg[2]/P0001  ;
  assign n16876 = \u1_u3_tx_data_to_cnt_reg[0]/P0001  & \u1_u3_tx_data_to_cnt_reg[1]/P0001  ;
  assign n16877 = n16875 & n16876 ;
  assign n16878 = ~n16874 & ~n16877 ;
  assign n16879 = \u1_u3_tx_data_to_cnt_reg[4]/P0001  & n12665 ;
  assign n16880 = ~\u1_u3_tx_data_to_cnt_reg[5]/P0001  & ~n16879 ;
  assign n16881 = ~\u0_rx_active_reg/P0001  & ~n16644 ;
  assign n16882 = ~n16880 & n16881 ;
  assign n16883 = n8866 & n16865 ;
  assign n16884 = ~\u4_u0_inta_reg/P0001  & ~\u4_u0_intb_reg/P0001  ;
  assign n16885 = ~\u4_u1_inta_reg/P0001  & ~\u4_u1_intb_reg/P0001  ;
  assign n16886 = ~\u4_u2_inta_reg/P0001  & ~\u4_u2_intb_reg/P0001  ;
  assign n16887 = ~\u4_u3_inta_reg/P0001  & ~\u4_u3_intb_reg/P0001  ;
  assign n16888 = n8826 & n16865 ;
  assign n16889 = ~\u0_u0_me_ps2_reg[4]/P0001  & n7078 ;
  assign n16890 = ~\u0_u0_me_ps2_0_5_ms_reg/P0001  & \u0_u0_me_ps2_reg[3]/P0001  ;
  assign n16891 = ~\u0_u0_me_ps2_reg[2]/P0001  & ~\u0_u0_me_ps2_reg[5]/P0001  ;
  assign n16892 = n16890 & n16891 ;
  assign n16893 = n16889 & n16892 ;
  assign n16894 = n6696 & n16893 ;
  assign n16895 = n12415 & n12416 ;
  assign n16896 = \u4_u3_buf0_orig_reg[28]/P0001  & ~n13108 ;
  assign n16897 = ~n16895 & ~n16896 ;
  assign n16898 = n12468 & n12469 ;
  assign n16899 = \u4_u1_buf0_orig_reg[28]/P0001  & ~n13114 ;
  assign n16900 = ~n16898 & ~n16899 ;
  assign n16901 = n12447 & n13091 ;
  assign n16902 = \u4_u0_buf0_orig_reg[28]/P0001  & ~n13111 ;
  assign n16903 = ~n16901 & ~n16902 ;
  assign n16904 = \u0_u0_idle_cnt1_reg[6]/P0001  & ~n15580 ;
  assign n16905 = ~\u0_u0_idle_cnt1_reg[6]/P0001  & n13034 ;
  assign n16906 = n14315 & n16905 ;
  assign n16907 = ~n16904 & ~n16906 ;
  assign n16908 = n12491 & n12492 ;
  assign n16909 = \u4_u2_buf0_orig_reg[28]/P0001  & ~n13122 ;
  assign n16910 = ~n16908 & ~n16909 ;
  assign n16911 = ~n9077 & ~n9079 ;
  assign n16912 = ~n9078 & ~n9082 ;
  assign n16913 = ~n16911 & ~n16912 ;
  assign n16914 = n16911 & n16912 ;
  assign n16915 = ~n16913 & ~n16914 ;
  assign n16916 = ~n9081 & ~n9082 ;
  assign n16917 = ~n9071 & ~n9073 ;
  assign n16918 = ~n16916 & ~n16917 ;
  assign n16919 = ~n9082 & n16917 ;
  assign n16920 = ~n9081 & n16919 ;
  assign n16921 = ~n16918 & ~n16920 ;
  assign n16922 = \u4_u2_buf0_orig_reg[29]/NET0131  & ~n16908 ;
  assign n16923 = ~n12496 & ~n16922 ;
  assign n16924 = \u4_u0_buf0_orig_reg[29]/NET0131  & ~n16901 ;
  assign n16925 = ~n12445 & ~n16924 ;
  assign n16926 = \u4_u3_buf0_orig_reg[29]/NET0131  & ~n16895 ;
  assign n16927 = ~n12420 & ~n16926 ;
  assign n16928 = ~n9126 & ~n9128 ;
  assign n16929 = ~n9127 & ~n9131 ;
  assign n16930 = ~n16928 & ~n16929 ;
  assign n16931 = n16928 & n16929 ;
  assign n16932 = ~n16930 & ~n16931 ;
  assign n16933 = ~n9130 & ~n9131 ;
  assign n16934 = ~n9120 & ~n9122 ;
  assign n16935 = ~n16933 & ~n16934 ;
  assign n16936 = ~n9131 & n16934 ;
  assign n16937 = ~n9130 & n16936 ;
  assign n16938 = ~n16935 & ~n16937 ;
  assign n16939 = \u4_u1_buf0_orig_reg[29]/NET0131  & ~n16898 ;
  assign n16940 = ~n12473 & ~n16939 ;
  assign n16941 = ~n9175 & ~n9177 ;
  assign n16942 = ~n9176 & ~n9180 ;
  assign n16943 = ~n16941 & ~n16942 ;
  assign n16944 = n16941 & n16942 ;
  assign n16945 = ~n16943 & ~n16944 ;
  assign n16946 = ~n9179 & ~n9180 ;
  assign n16947 = ~n9169 & ~n9171 ;
  assign n16948 = ~n16946 & ~n16947 ;
  assign n16949 = ~n9180 & n16947 ;
  assign n16950 = ~n9179 & n16949 ;
  assign n16951 = ~n16948 & ~n16950 ;
  assign n16952 = ~n9224 & ~n9226 ;
  assign n16953 = ~n9225 & ~n9229 ;
  assign n16954 = ~n16952 & ~n16953 ;
  assign n16955 = n16952 & n16953 ;
  assign n16956 = ~n16954 & ~n16955 ;
  assign n16957 = ~n9228 & ~n9229 ;
  assign n16958 = ~n9218 & ~n9220 ;
  assign n16959 = ~n16957 & ~n16958 ;
  assign n16960 = ~n9229 & n16958 ;
  assign n16961 = ~n9228 & n16960 ;
  assign n16962 = ~n16959 & ~n16961 ;
  assign n16963 = \u4_buf1_reg[0]/P0001  & n2793 ;
  assign n16964 = \u4_buf1_reg[0]/P0001  & ~n2789 ;
  assign n16965 = n2788 & n16964 ;
  assign n16966 = ~n16963 & ~n16965 ;
  assign n16967 = n2788 & ~n2789 ;
  assign n16968 = \u4_buf0_reg[0]/P0001  & ~n2793 ;
  assign n16969 = ~n16967 & n16968 ;
  assign n16970 = n16966 & ~n16969 ;
  assign n16971 = \u4_buf1_reg[10]/P0001  & n2793 ;
  assign n16972 = \u4_buf1_reg[10]/P0001  & ~n2789 ;
  assign n16973 = n2788 & n16972 ;
  assign n16974 = ~n16971 & ~n16973 ;
  assign n16975 = \u4_buf0_reg[10]/P0001  & ~n2793 ;
  assign n16976 = ~n16967 & n16975 ;
  assign n16977 = n16974 & ~n16976 ;
  assign n16978 = \u4_buf1_reg[11]/P0001  & n2793 ;
  assign n16979 = \u4_buf1_reg[11]/P0001  & ~n2789 ;
  assign n16980 = n2788 & n16979 ;
  assign n16981 = ~n16978 & ~n16980 ;
  assign n16982 = \u4_buf0_reg[11]/P0001  & ~n2793 ;
  assign n16983 = ~n16967 & n16982 ;
  assign n16984 = n16981 & ~n16983 ;
  assign n16985 = \u4_buf1_reg[12]/P0001  & n2793 ;
  assign n16986 = \u4_buf1_reg[12]/P0001  & ~n2789 ;
  assign n16987 = n2788 & n16986 ;
  assign n16988 = ~n16985 & ~n16987 ;
  assign n16989 = \u4_buf0_reg[12]/P0001  & ~n2793 ;
  assign n16990 = ~n16967 & n16989 ;
  assign n16991 = n16988 & ~n16990 ;
  assign n16992 = \u4_buf1_reg[13]/P0001  & n2793 ;
  assign n16993 = \u4_buf1_reg[13]/P0001  & ~n2789 ;
  assign n16994 = n2788 & n16993 ;
  assign n16995 = ~n16992 & ~n16994 ;
  assign n16996 = \u4_buf0_reg[13]/P0001  & ~n2793 ;
  assign n16997 = ~n16967 & n16996 ;
  assign n16998 = n16995 & ~n16997 ;
  assign n16999 = \u4_buf1_reg[14]/P0001  & n2793 ;
  assign n17000 = \u4_buf1_reg[14]/P0001  & ~n2789 ;
  assign n17001 = n2788 & n17000 ;
  assign n17002 = ~n16999 & ~n17001 ;
  assign n17003 = \u4_buf0_reg[14]/P0001  & ~n2793 ;
  assign n17004 = ~n16967 & n17003 ;
  assign n17005 = n17002 & ~n17004 ;
  assign n17006 = \u4_buf1_reg[16]/P0001  & n2793 ;
  assign n17007 = \u4_buf1_reg[16]/P0001  & ~n2789 ;
  assign n17008 = n2788 & n17007 ;
  assign n17009 = ~n17006 & ~n17008 ;
  assign n17010 = \u4_buf0_reg[16]/P0001  & ~n2793 ;
  assign n17011 = ~n16967 & n17010 ;
  assign n17012 = n17009 & ~n17011 ;
  assign n17013 = \u4_buf1_reg[1]/P0001  & n2793 ;
  assign n17014 = \u4_buf1_reg[1]/P0001  & ~n2789 ;
  assign n17015 = n2788 & n17014 ;
  assign n17016 = ~n17013 & ~n17015 ;
  assign n17017 = \u4_buf0_reg[1]/P0001  & ~n2793 ;
  assign n17018 = ~n16967 & n17017 ;
  assign n17019 = n17016 & ~n17018 ;
  assign n17020 = \u4_buf1_reg[2]/P0001  & n2793 ;
  assign n17021 = \u4_buf1_reg[2]/P0001  & ~n2789 ;
  assign n17022 = n2788 & n17021 ;
  assign n17023 = ~n17020 & ~n17022 ;
  assign n17024 = \u4_buf0_reg[2]/P0001  & ~n2793 ;
  assign n17025 = ~n16967 & n17024 ;
  assign n17026 = n17023 & ~n17025 ;
  assign n17027 = \u4_buf1_reg[3]/P0001  & n2793 ;
  assign n17028 = \u4_buf1_reg[3]/P0001  & ~n2789 ;
  assign n17029 = n2788 & n17028 ;
  assign n17030 = ~n17027 & ~n17029 ;
  assign n17031 = \u4_buf0_reg[3]/P0001  & ~n2793 ;
  assign n17032 = ~n16967 & n17031 ;
  assign n17033 = n17030 & ~n17032 ;
  assign n17034 = \u4_buf1_reg[4]/P0001  & n2793 ;
  assign n17035 = \u4_buf1_reg[4]/P0001  & ~n2789 ;
  assign n17036 = n2788 & n17035 ;
  assign n17037 = ~n17034 & ~n17036 ;
  assign n17038 = \u4_buf0_reg[4]/P0001  & ~n2793 ;
  assign n17039 = ~n16967 & n17038 ;
  assign n17040 = n17037 & ~n17039 ;
  assign n17041 = \u4_buf1_reg[5]/P0001  & n2793 ;
  assign n17042 = \u4_buf1_reg[5]/P0001  & ~n2789 ;
  assign n17043 = n2788 & n17042 ;
  assign n17044 = ~n17041 & ~n17043 ;
  assign n17045 = \u4_buf0_reg[5]/P0001  & ~n2793 ;
  assign n17046 = ~n16967 & n17045 ;
  assign n17047 = n17044 & ~n17046 ;
  assign n17048 = \u4_buf1_reg[6]/P0001  & n2793 ;
  assign n17049 = \u4_buf1_reg[6]/P0001  & ~n2789 ;
  assign n17050 = n2788 & n17049 ;
  assign n17051 = ~n17048 & ~n17050 ;
  assign n17052 = \u4_buf0_reg[6]/P0001  & ~n2793 ;
  assign n17053 = ~n16967 & n17052 ;
  assign n17054 = n17051 & ~n17053 ;
  assign n17055 = \u4_buf1_reg[7]/P0001  & n2793 ;
  assign n17056 = \u4_buf1_reg[7]/P0001  & ~n2789 ;
  assign n17057 = n2788 & n17056 ;
  assign n17058 = ~n17055 & ~n17057 ;
  assign n17059 = \u4_buf0_reg[7]/P0001  & ~n2793 ;
  assign n17060 = ~n16967 & n17059 ;
  assign n17061 = n17058 & ~n17060 ;
  assign n17062 = \u4_buf1_reg[8]/P0001  & n2793 ;
  assign n17063 = \u4_buf1_reg[8]/P0001  & ~n2789 ;
  assign n17064 = n2788 & n17063 ;
  assign n17065 = ~n17062 & ~n17064 ;
  assign n17066 = \u4_buf0_reg[8]/P0001  & ~n2793 ;
  assign n17067 = ~n16967 & n17066 ;
  assign n17068 = n17065 & ~n17067 ;
  assign n17069 = \u4_buf1_reg[9]/P0001  & n2793 ;
  assign n17070 = \u4_buf1_reg[9]/P0001  & ~n2789 ;
  assign n17071 = n2788 & n17070 ;
  assign n17072 = ~n17069 & ~n17071 ;
  assign n17073 = \u4_buf0_reg[9]/P0001  & ~n2793 ;
  assign n17074 = ~n16967 & n17073 ;
  assign n17075 = n17072 & ~n17074 ;
  assign n17076 = \u4_buf1_reg[15]/P0001  & n2793 ;
  assign n17077 = \u4_buf1_reg[15]/P0001  & ~n2789 ;
  assign n17078 = n2788 & n17077 ;
  assign n17079 = ~n17076 & ~n17078 ;
  assign n17080 = \u4_buf0_reg[15]/P0001  & ~n2793 ;
  assign n17081 = ~n16967 & n17080 ;
  assign n17082 = n17079 & ~n17081 ;
  assign n17083 = ~\u1_u3_in_token_reg/NET0131  & ~n2350 ;
  assign n17084 = ~n2355 & ~n17083 ;
  assign n17085 = \u1_u0_pid_reg[2]/NET0131  & ~\u1_u3_in_token_reg/NET0131  ;
  assign n17086 = rst_i_pad & ~n17085 ;
  assign n17087 = ~n5016 & n17086 ;
  assign n17088 = n17084 & n17087 ;
  assign n17089 = n5734 & n6154 ;
  assign n17090 = n5746 & n17089 ;
  assign n17091 = \u0_u0_me_cnt_100_ms_reg/P0001  & \u0_u0_state_reg[8]/NET0131  ;
  assign n17092 = ~\u0_u0_usb_attached_reg/P0001  & ~n17091 ;
  assign n17093 = ~n17090 & ~n17092 ;
  assign n17094 = ~\u1_u3_rx_ack_to_cnt_reg[4]/P0001  & \u1_u3_rx_ack_to_cnt_reg[5]/P0001  ;
  assign n17095 = ~\u0_u0_mode_hs_reg/P0001  & ~\u1_u3_rx_ack_to_cnt_reg[1]/P0001  ;
  assign n17096 = n17094 & n17095 ;
  assign n17097 = \u1_u3_rx_ack_to_cnt_reg[4]/P0001  & ~\u1_u3_rx_ack_to_cnt_reg[5]/P0001  ;
  assign n17098 = \u0_u0_mode_hs_reg/P0001  & \u1_u3_rx_ack_to_cnt_reg[1]/P0001  ;
  assign n17099 = n17097 & n17098 ;
  assign n17100 = ~n17096 & ~n17099 ;
  assign n17101 = ~\u1_u3_rx_ack_to_cnt_reg[0]/P0001  & \u1_u3_rx_ack_to_cnt_reg[2]/P0001  ;
  assign n17102 = ~\u1_u3_rx_ack_to_cnt_reg[3]/P0001  & ~\u1_u3_rx_ack_to_cnt_reg[6]/P0001  ;
  assign n17103 = n17101 & n17102 ;
  assign n17104 = ~\u1_u3_rx_ack_to_cnt_reg[7]/P0001  & n17103 ;
  assign n17105 = ~n17100 & n17104 ;
  assign n17106 = ~\u1_u3_tx_data_to_cnt_reg[4]/P0001  & \u1_u3_tx_data_to_cnt_reg[5]/P0001  ;
  assign n17107 = ~\u0_u0_mode_hs_reg/P0001  & ~\u1_u3_tx_data_to_cnt_reg[1]/P0001  ;
  assign n17108 = n17106 & n17107 ;
  assign n17109 = \u1_u3_tx_data_to_cnt_reg[4]/P0001  & ~\u1_u3_tx_data_to_cnt_reg[5]/P0001  ;
  assign n17110 = \u0_u0_mode_hs_reg/P0001  & \u1_u3_tx_data_to_cnt_reg[1]/P0001  ;
  assign n17111 = n17109 & n17110 ;
  assign n17112 = ~n17108 & ~n17111 ;
  assign n17113 = ~\u1_u3_tx_data_to_cnt_reg[0]/P0001  & \u1_u3_tx_data_to_cnt_reg[2]/P0001  ;
  assign n17114 = ~\u1_u3_tx_data_to_cnt_reg[3]/P0001  & ~\u1_u3_tx_data_to_cnt_reg[6]/P0001  ;
  assign n17115 = n17113 & n17114 ;
  assign n17116 = ~\u1_u3_tx_data_to_cnt_reg[7]/P0001  & n17115 ;
  assign n17117 = ~n17112 & n17116 ;
  assign n17118 = ~\u0_u0_me_ps_reg[6]/P0001  & \u0_u0_me_ps_reg[7]/P0001  ;
  assign n17119 = \u0_u0_me_ps_reg[4]/P0001  & ~\u0_u0_me_ps_reg[5]/P0001  ;
  assign n17120 = n17118 & n17119 ;
  assign n17121 = \u0_u0_me_ps_reg[2]/P0001  & ~\u0_u0_me_ps_reg[3]/P0001  ;
  assign n17122 = n7086 & n17121 ;
  assign n17123 = n17120 & n17122 ;
  assign n17124 = n2795 & n4401 ;
  assign n17125 = ~n2795 & n4401 ;
  assign n17126 = rst_i_pad & n5016 ;
  assign n17127 = ~\u1_u0_pid_reg[2]/NET0131  & n2350 ;
  assign n17128 = rst_i_pad & \u1_u3_setup_token_reg/P0001  ;
  assign n17129 = ~n17127 & n17128 ;
  assign n17130 = ~n17126 & ~n17129 ;
  assign n17131 = \u4_u2_buf1_reg[14]/P0001  & n2731 ;
  assign n17132 = \u4_u2_buf0_reg[14]/P0001  & n2568 ;
  assign n17133 = ~n17131 & ~n17132 ;
  assign n17134 = n8826 & ~n17133 ;
  assign n17135 = \u4_u3_buf1_reg[14]/P0001  & n2731 ;
  assign n17136 = \u4_u3_buf0_reg[14]/P0001  & n2568 ;
  assign n17137 = ~n17135 & ~n17136 ;
  assign n17138 = n8836 & ~n17137 ;
  assign n17139 = ~n17134 & ~n17138 ;
  assign n17140 = \u4_u1_buf1_reg[14]/P0001  & n2731 ;
  assign n17141 = \u4_u1_buf0_reg[14]/P0001  & n2568 ;
  assign n17142 = ~n17140 & ~n17141 ;
  assign n17143 = n8866 & ~n17142 ;
  assign n17144 = \u4_u0_buf1_reg[14]/P0001  & n2731 ;
  assign n17145 = \u4_u0_buf0_reg[14]/P0001  & n2568 ;
  assign n17146 = ~n17144 & ~n17145 ;
  assign n17147 = n8815 & ~n17146 ;
  assign n17148 = ~n17143 & ~n17147 ;
  assign n17149 = n17139 & n17148 ;
  assign n17150 = ~\u1_u2_sizd_c_reg[0]/P0001  & n3433 ;
  assign n17151 = n3435 & n17150 ;
  assign n17152 = n3432 & n17151 ;
  assign n17153 = ~\u1_u2_rx_data_done_r_reg/P0001  & ~n17152 ;
  assign n17154 = n8836 & n16865 ;
  assign n17155 = n12411 & n12412 ;
  assign n17156 = \u4_u3_buf0_orig_reg[24]/P0001  & ~n14385 ;
  assign n17157 = ~n17155 & ~n17156 ;
  assign n17158 = n12464 & n12465 ;
  assign n17159 = \u4_u1_buf0_orig_reg[25]/P0001  & ~n17158 ;
  assign n17160 = ~n13101 & ~n17159 ;
  assign n17161 = n12436 & n12441 ;
  assign n17162 = \u4_u0_buf0_orig_reg[24]/P0001  & ~n14388 ;
  assign n17163 = ~n17161 & ~n17162 ;
  assign n17164 = \u4_u0_buf0_orig_reg[25]/P0001  & ~n17161 ;
  assign n17165 = ~n13094 & ~n17164 ;
  assign n17166 = \u4_u3_buf0_orig_reg[25]/P0001  & ~n17155 ;
  assign n17167 = ~n13040 & ~n17166 ;
  assign n17168 = \u4_u1_buf0_orig_reg[24]/P0001  & ~n14391 ;
  assign n17169 = ~n17158 & ~n17168 ;
  assign n17170 = n12487 & n12488 ;
  assign n17171 = \u4_u2_buf0_orig_reg[24]/P0001  & ~n14394 ;
  assign n17172 = ~n17170 & ~n17171 ;
  assign n17173 = \u4_u2_buf0_orig_reg[25]/P0001  & ~n17170 ;
  assign n17174 = ~n13105 & ~n17173 ;
  assign n17175 = \u4_u0_buf0_orig_reg[21]/P0001  & n12439 ;
  assign n17176 = ~n16663 & ~n17175 ;
  assign n17177 = \u4_u1_buf0_orig_reg[21]/P0001  & n12462 ;
  assign n17178 = ~n16666 & ~n17177 ;
  assign n17179 = \u4_u2_buf0_orig_reg[21]/P0001  & n12485 ;
  assign n17180 = ~n16669 & ~n17179 ;
  assign n17181 = \u4_u3_buf0_orig_reg[21]/P0001  & n12409 ;
  assign n17182 = ~n16655 & ~n17181 ;
  assign n17183 = \u1_u3_out_token_reg/NET0131  & ~n2352 ;
  assign n17184 = n5017 & ~n17183 ;
  assign n17185 = rst_i_pad & ~n17184 ;
  assign n17186 = ~\u0_u0_mode_hs_reg/P0001  & ~\u0_u0_state_reg[13]/NET0131  ;
  assign n17187 = ~\u0_u0_state_reg[13]/NET0131  & n5754 ;
  assign n17188 = n5746 & n17187 ;
  assign n17189 = ~n17186 & ~n17188 ;
  assign n17190 = ~\u0_u0_idle_cnt1_reg[2]/P0001  & \u0_u0_idle_cnt1_reg[3]/P0001  ;
  assign n17191 = ~\u0_u0_idle_cnt1_reg[0]/P0001  & \u0_u0_idle_cnt1_reg[1]/P0001  ;
  assign n17192 = n17190 & n17191 ;
  assign n17193 = n15577 & n17192 ;
  assign n17194 = \u4_u3_iena_reg[5]/P0001  & \u4_u3_int_stat_reg[6]/P0001  ;
  assign n17195 = \u4_u3_iena_reg[2]/P0001  & \u4_u3_int_stat_reg[2]/P0001  ;
  assign n17196 = \u4_u3_iena_reg[1]/P0001  & \u4_u3_int_stat_reg[1]/P0001  ;
  assign n17197 = ~n17195 & ~n17196 ;
  assign n17198 = ~n17194 & n17197 ;
  assign n17199 = \u4_u3_iena_reg[0]/P0001  & \u4_u3_int_stat_reg[0]/P0001  ;
  assign n17200 = \u4_u3_iena_reg[4]/P0001  & \u4_u3_int_stat_reg[5]/P0001  ;
  assign n17201 = ~n17199 & ~n17200 ;
  assign n17202 = ~\u4_u3_int_stat_reg[3]/P0001  & ~\u4_u3_int_stat_reg[4]/P0001  ;
  assign n17203 = \u4_u3_iena_reg[3]/P0001  & ~n17202 ;
  assign n17204 = n17201 & ~n17203 ;
  assign n17205 = n17198 & n17204 ;
  assign n17206 = \u4_u3_ienb_reg[1]/P0001  & \u4_u3_int_stat_reg[1]/P0001  ;
  assign n17207 = \u4_u3_ienb_reg[2]/P0001  & \u4_u3_int_stat_reg[2]/P0001  ;
  assign n17208 = \u4_u3_ienb_reg[0]/P0001  & \u4_u3_int_stat_reg[0]/P0001  ;
  assign n17209 = ~n17207 & ~n17208 ;
  assign n17210 = ~n17206 & n17209 ;
  assign n17211 = \u4_u3_ienb_reg[3]/P0001  & ~n17202 ;
  assign n17212 = \u4_u3_ienb_reg[4]/P0001  & \u4_u3_int_stat_reg[5]/P0001  ;
  assign n17213 = \u4_u3_ienb_reg[5]/P0001  & \u4_u3_int_stat_reg[6]/P0001  ;
  assign n17214 = ~n17212 & ~n17213 ;
  assign n17215 = ~n17211 & n17214 ;
  assign n17216 = n17210 & n17215 ;
  assign n17217 = \u4_u0_ienb_reg[5]/P0001  & \u4_u0_int_stat_reg[6]/P0001  ;
  assign n17218 = \u4_u0_ienb_reg[4]/P0001  & \u4_u0_int_stat_reg[5]/P0001  ;
  assign n17219 = \u4_u0_ienb_reg[1]/P0001  & \u4_u0_int_stat_reg[1]/P0001  ;
  assign n17220 = ~n17218 & ~n17219 ;
  assign n17221 = ~n17217 & n17220 ;
  assign n17222 = \u4_u0_ienb_reg[0]/P0001  & \u4_u0_int_stat_reg[0]/P0001  ;
  assign n17223 = \u4_u0_ienb_reg[2]/P0001  & \u4_u0_int_stat_reg[2]/P0001  ;
  assign n17224 = ~n17222 & ~n17223 ;
  assign n17225 = ~\u4_u0_int_stat_reg[3]/P0001  & ~\u4_u0_int_stat_reg[4]/P0001  ;
  assign n17226 = \u4_u0_ienb_reg[3]/P0001  & ~n17225 ;
  assign n17227 = n17224 & ~n17226 ;
  assign n17228 = n17221 & n17227 ;
  assign n17229 = \u4_u0_iena_reg[5]/P0001  & \u4_u0_int_stat_reg[6]/P0001  ;
  assign n17230 = \u4_u0_iena_reg[1]/P0001  & \u4_u0_int_stat_reg[1]/P0001  ;
  assign n17231 = \u4_u0_iena_reg[0]/P0001  & \u4_u0_int_stat_reg[0]/P0001  ;
  assign n17232 = ~n17230 & ~n17231 ;
  assign n17233 = ~n17229 & n17232 ;
  assign n17234 = \u4_u0_iena_reg[3]/P0001  & ~n17225 ;
  assign n17235 = \u4_u0_iena_reg[2]/P0001  & \u4_u0_int_stat_reg[2]/P0001  ;
  assign n17236 = \u4_u0_iena_reg[4]/P0001  & \u4_u0_int_stat_reg[5]/P0001  ;
  assign n17237 = ~n17235 & ~n17236 ;
  assign n17238 = ~n17234 & n17237 ;
  assign n17239 = n17233 & n17238 ;
  assign n17240 = \u4_u1_iena_reg[5]/P0001  & \u4_u1_int_stat_reg[6]/P0001  ;
  assign n17241 = \u4_u1_iena_reg[2]/P0001  & \u4_u1_int_stat_reg[2]/P0001  ;
  assign n17242 = \u4_u1_iena_reg[1]/P0001  & \u4_u1_int_stat_reg[1]/P0001  ;
  assign n17243 = ~n17241 & ~n17242 ;
  assign n17244 = ~n17240 & n17243 ;
  assign n17245 = \u4_u1_iena_reg[0]/P0001  & \u4_u1_int_stat_reg[0]/P0001  ;
  assign n17246 = \u4_u1_iena_reg[4]/P0001  & \u4_u1_int_stat_reg[5]/P0001  ;
  assign n17247 = ~n17245 & ~n17246 ;
  assign n17248 = ~\u4_u1_int_stat_reg[3]/P0001  & ~\u4_u1_int_stat_reg[4]/P0001  ;
  assign n17249 = \u4_u1_iena_reg[3]/P0001  & ~n17248 ;
  assign n17250 = n17247 & ~n17249 ;
  assign n17251 = n17244 & n17250 ;
  assign n17252 = \u4_u1_ienb_reg[5]/P0001  & \u4_u1_int_stat_reg[6]/P0001  ;
  assign n17253 = \u4_u1_ienb_reg[1]/P0001  & \u4_u1_int_stat_reg[1]/P0001  ;
  assign n17254 = \u4_u1_ienb_reg[0]/P0001  & \u4_u1_int_stat_reg[0]/P0001  ;
  assign n17255 = ~n17253 & ~n17254 ;
  assign n17256 = ~n17252 & n17255 ;
  assign n17257 = \u4_u1_ienb_reg[3]/P0001  & ~n17248 ;
  assign n17258 = \u4_u1_ienb_reg[2]/P0001  & \u4_u1_int_stat_reg[2]/P0001  ;
  assign n17259 = \u4_u1_ienb_reg[4]/P0001  & \u4_u1_int_stat_reg[5]/P0001  ;
  assign n17260 = ~n17258 & ~n17259 ;
  assign n17261 = ~n17257 & n17260 ;
  assign n17262 = n17256 & n17261 ;
  assign n17263 = \u4_u2_ienb_reg[1]/P0001  & \u4_u2_int_stat_reg[1]/P0001  ;
  assign n17264 = \u4_u2_ienb_reg[2]/P0001  & \u4_u2_int_stat_reg[2]/P0001  ;
  assign n17265 = \u4_u2_ienb_reg[0]/P0001  & \u4_u2_int_stat_reg[0]/P0001  ;
  assign n17266 = ~n17264 & ~n17265 ;
  assign n17267 = ~n17263 & n17266 ;
  assign n17268 = \u4_u2_ienb_reg[4]/P0001  & \u4_u2_int_stat_reg[5]/P0001  ;
  assign n17269 = \u4_u2_ienb_reg[5]/P0001  & \u4_u2_int_stat_reg[6]/P0001  ;
  assign n17270 = ~n17268 & ~n17269 ;
  assign n17271 = ~\u4_u2_int_stat_reg[3]/P0001  & ~\u4_u2_int_stat_reg[4]/P0001  ;
  assign n17272 = \u4_u2_ienb_reg[3]/P0001  & ~n17271 ;
  assign n17273 = n17270 & ~n17272 ;
  assign n17274 = n17267 & n17273 ;
  assign n17275 = \u4_u2_iena_reg[5]/P0001  & \u4_u2_int_stat_reg[6]/P0001  ;
  assign n17276 = \u4_u2_iena_reg[2]/P0001  & \u4_u2_int_stat_reg[2]/P0001  ;
  assign n17277 = \u4_u2_iena_reg[1]/P0001  & \u4_u2_int_stat_reg[1]/P0001  ;
  assign n17278 = ~n17276 & ~n17277 ;
  assign n17279 = ~n17275 & n17278 ;
  assign n17280 = \u4_u2_iena_reg[3]/P0001  & ~n17271 ;
  assign n17281 = \u4_u2_iena_reg[0]/P0001  & \u4_u2_int_stat_reg[0]/P0001  ;
  assign n17282 = \u4_u2_iena_reg[4]/P0001  & \u4_u2_int_stat_reg[5]/P0001  ;
  assign n17283 = ~n17281 & ~n17282 ;
  assign n17284 = ~n17280 & n17283 ;
  assign n17285 = n17279 & n17284 ;
  assign n17286 = n12488 & n12492 ;
  assign n17287 = ~\u4_u2_buf0_orig_reg[29]/NET0131  & ~\u4_u2_buf0_orig_reg[30]/NET0131  ;
  assign n17288 = n12486 & n12489 ;
  assign n17289 = n17287 & n17288 ;
  assign n17290 = n17286 & n17289 ;
  assign n17291 = n7848 & ~n17290 ;
  assign n17292 = ~\u4_u1_buf0_orig_reg[30]/NET0131  & n12465 ;
  assign n17293 = n12470 & n17292 ;
  assign n17294 = n12463 & n12466 ;
  assign n17295 = n17293 & n17294 ;
  assign n17296 = n8778 & ~n17295 ;
  assign n17297 = n12412 & n12416 ;
  assign n17298 = ~\u4_u3_buf0_orig_reg[29]/NET0131  & ~\u4_u3_buf0_orig_reg[30]/NET0131  ;
  assign n17299 = n12410 & n12413 ;
  assign n17300 = n17298 & n17299 ;
  assign n17301 = n17297 & n17300 ;
  assign n17302 = n7917 & ~n17301 ;
  assign n17303 = n12438 & n12440 ;
  assign n17304 = n12449 & n17303 ;
  assign n17305 = n8716 & ~n17304 ;
  assign n17306 = n7462 & n7868 ;
  assign n17307 = n4355 & ~n17306 ;
  assign n17308 = n7362 & n8734 ;
  assign n17309 = n4377 & ~n17308 ;
  assign n17310 = n7312 & n7933 ;
  assign n17311 = n4366 & ~n17310 ;
  assign n17312 = n7412 & n8798 ;
  assign n17313 = n4388 & ~n17312 ;
  assign n17314 = ~n11230 & ~n13034 ;
  assign n17315 = ~n14317 & ~n17314 ;
  assign n17316 = \u0_u0_idle_cnt1_reg[4]/P0001  & ~\u0_u0_idle_cnt1_reg[5]/P0001  ;
  assign n17317 = ~n14315 & n17316 ;
  assign n17318 = ~n17315 & ~n17317 ;
  assign n17319 = ~n11228 & ~n16672 ;
  assign n17320 = ~n9222 & ~n9226 ;
  assign n17321 = ~n9223 & ~n17320 ;
  assign n17322 = n9223 & n17320 ;
  assign n17323 = ~n17321 & ~n17322 ;
  assign n17324 = ~n9075 & ~n9079 ;
  assign n17325 = ~n9076 & ~n17324 ;
  assign n17326 = n9076 & n17324 ;
  assign n17327 = ~n17325 & ~n17326 ;
  assign n17328 = ~n9124 & ~n9128 ;
  assign n17329 = ~n9125 & ~n17328 ;
  assign n17330 = n9125 & n17328 ;
  assign n17331 = ~n17329 & ~n17330 ;
  assign n17332 = ~n9173 & ~n9177 ;
  assign n17333 = ~n9174 & ~n17332 ;
  assign n17334 = n9174 & n17332 ;
  assign n17335 = ~n17333 & ~n17334 ;
  assign n17336 = ~\u4_u3_dma_ack_clr1_reg/P0001  & \u4_u3_dma_ack_wr1_reg/P0001  ;
  assign n17337 = ~\dma_ack_i[3]_pad  & ~n17336 ;
  assign n17338 = rst_i_pad & ~n17337 ;
  assign n17339 = ~\u4_u0_dma_ack_clr1_reg/P0001  & \u4_u0_dma_ack_wr1_reg/P0001  ;
  assign n17340 = ~\dma_ack_i[0]_pad  & ~n17339 ;
  assign n17341 = rst_i_pad & ~n17340 ;
  assign n17342 = ~\u4_u1_dma_ack_clr1_reg/P0001  & \u4_u1_dma_ack_wr1_reg/P0001  ;
  assign n17343 = ~\dma_ack_i[1]_pad  & ~n17342 ;
  assign n17344 = rst_i_pad & ~n17343 ;
  assign n17345 = ~\u4_u2_dma_ack_clr1_reg/P0001  & \u4_u2_dma_ack_wr1_reg/P0001  ;
  assign n17346 = ~\dma_ack_i[2]_pad  & ~n17345 ;
  assign n17347 = rst_i_pad & ~n17346 ;
  assign n17348 = ~\u1_u3_tx_data_to_cnt_reg[0]/P0001  & ~\u1_u3_tx_data_to_cnt_reg[1]/P0001  ;
  assign n17349 = ~\u0_rx_active_reg/P0001  & ~n12663 ;
  assign n17350 = ~n17348 & n17349 ;
  assign n17351 = ~\u1_u3_rx_ack_to_cnt_reg[0]/P0001  & ~\u1_u3_rx_ack_to_cnt_reg[1]/P0001  ;
  assign n17352 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & ~n12630 ;
  assign n17353 = ~n17351 & n17352 ;
  assign n17354 = ~\u1_u3_rx_ack_to_clr_reg/P0001  & ~\u1_u3_rx_ack_to_cnt_reg[0]/P0001  ;
  assign n17355 = \u1_hms_cnt_reg[4]/P0001  & n6488 ;
  assign n17356 = n6480 & n17355 ;
  assign n17357 = n12610 & n12624 ;
  assign n17358 = \u1_u0_pid_reg[2]/NET0131  & \u1_u0_pid_reg[6]/P0001  ;
  assign n17359 = \u1_u0_pid_reg[3]/NET0131  & \u1_u0_pid_reg[7]/P0001  ;
  assign n17360 = ~n17358 & ~n17359 ;
  assign n17361 = ~\u1_u0_pid_reg[2]/NET0131  & ~\u1_u0_pid_reg[6]/P0001  ;
  assign n17362 = ~\u1_u0_pid_reg[3]/NET0131  & ~\u1_u0_pid_reg[7]/P0001  ;
  assign n17363 = ~n17361 & ~n17362 ;
  assign n17364 = n17360 & n17363 ;
  assign n17365 = \u1_u0_pid_reg[0]/NET0131  & ~\u1_u0_pid_reg[4]/P0001  ;
  assign n17366 = ~\u1_u0_pid_reg[0]/NET0131  & \u1_u0_pid_reg[4]/P0001  ;
  assign n17367 = ~n17365 & ~n17366 ;
  assign n17368 = \u1_u0_pid_reg[1]/NET0131  & ~\u1_u0_pid_reg[5]/P0001  ;
  assign n17369 = ~\u1_u0_pid_reg[1]/NET0131  & \u1_u0_pid_reg[5]/P0001  ;
  assign n17370 = ~n17368 & ~n17369 ;
  assign n17371 = ~n17367 & ~n17370 ;
  assign n17372 = n17364 & n17371 ;
  assign n17373 = ~\u0_u0_resume_req_s_reg/P0001  & \u0_u0_usb_suspend_reg/P0001  ;
  assign n17374 = ~\LineState_pad_i[0]_pad  & \LineState_pad_i[1]_pad  ;
  assign n17375 = ~n17373 & ~n17374 ;
  assign n17376 = \u4_u2_r2_reg/P0001  & ~\u4_u2_r4_reg/P0001  ;
  assign n17377 = ~\u4_u2_r1_reg/P0001  & ~n17376 ;
  assign n17378 = rst_i_pad & ~n17377 ;
  assign n17379 = \u4_u3_r2_reg/P0001  & ~\u4_u3_r4_reg/P0001  ;
  assign n17380 = ~\u4_u3_r1_reg/P0001  & ~n17379 ;
  assign n17381 = rst_i_pad & ~n17380 ;
  assign n17382 = \u4_u0_r2_reg/P0001  & ~\u4_u0_r4_reg/P0001  ;
  assign n17383 = ~\u4_u0_r1_reg/P0001  & ~n17382 ;
  assign n17384 = rst_i_pad & ~n17383 ;
  assign n17385 = \u4_u1_r2_reg/P0001  & ~\u4_u1_r4_reg/P0001  ;
  assign n17386 = ~\u4_u1_r1_reg/P0001  & ~n17385 ;
  assign n17387 = rst_i_pad & ~n17386 ;
  assign n17388 = n2366 & n12506 ;
  assign n17389 = ~\u0_rx_active_reg/P0001  & ~\u1_u3_tx_data_to_cnt_reg[0]/P0001  ;
  assign n17390 = ~\u4_u1_buf0_orig_reg[19]/P0001  & ~\u4_u1_buf0_orig_reg[20]/P0001  ;
  assign n17391 = ~n12462 & ~n17390 ;
  assign n17392 = ~n11227 & ~n12574 ;
  assign n17393 = ~\u1_u2_state_reg[4]/NET0131  & n4060 ;
  assign n17394 = \u4_u3_r5_reg/NET0131  & ~n6281 ;
  assign n17395 = \u4_u0_r5_reg/NET0131  & ~n6281 ;
  assign n17396 = \u4_u2_r5_reg/NET0131  & ~n6281 ;
  assign n17397 = \u1_u2_state_reg[1]/NET0131  & n4189 ;
  assign n17398 = ~TxValid_pad_o_pad & ~n2373 ;
  assign n17399 = ~\u0_u0_chirp_cnt_reg[0]/P0001  & \u0_u0_chirp_cnt_reg[1]/P0001  ;
  assign n17400 = \u0_u0_chirp_cnt_reg[2]/P0001  & n17399 ;
  assign n17401 = \u4_u1_r5_reg/NET0131  & ~n6281 ;
  assign n17402 = ~n8697 & ~n9125 ;
  assign n17403 = ~n7894 & ~n9076 ;
  assign n17404 = ~n7828 & ~n9223 ;
  assign n17405 = ~n8758 & ~n9174 ;
  assign n17406 = ~\u4_u3_buf0_orig_reg[19]/P0001  & ~\u4_u3_buf0_orig_reg[20]/P0001  ;
  assign n17407 = ~n12409 & ~n17406 ;
  assign n17408 = ~\u4_u0_buf0_orig_reg[19]/P0001  & ~\u4_u0_buf0_orig_reg[20]/P0001  ;
  assign n17409 = ~n12439 & ~n17408 ;
  assign n17410 = ~\u4_u2_buf0_orig_reg[19]/P0001  & ~\u4_u2_buf0_orig_reg[20]/P0001  ;
  assign n17411 = ~n12485 & ~n17410 ;
  assign n17412 = \u1_u3_new_size_reg[11]/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n17413 = \u1_u3_buffer_done_reg/P0001  & ~\u1_u3_out_to_small_r_reg/P0001  ;
  assign n17414 = ~\u1_u2_adr_cw_reg[0]/NET0131  & \u1_u2_mack_r_reg/P0001  ;
  assign n17415 = wb_cyc_i_pad & wb_stb_i_pad ;
  assign n17416 = RxError_pad_i_pad & rst_i_pad ;
  assign n17417 = RxActive_pad_i_pad & rst_i_pad ;
  assign n17418 = RxValid_pad_i_pad & rst_i_pad ;
  assign n17419 = \u1_u2_adr_cw_reg[0]/NET0131  & \u1_u2_mack_r_reg/P0001  ;
  assign n17420 = ~n3437 & n3439 ;
  assign n17421 = \u1_u2_sizd_c_reg[1]/P0001  & ~n3423 ;
  assign n17422 = ~n17420 & n17421 ;
  assign n17423 = n3679 & ~n17422 ;
  assign n17424 = ~\u1_u2_tx_dma_en_r_reg/P0001  & ~n3460 ;
  assign n17425 = ~n17423 & n17424 ;
  assign n17426 = rst_i_pad & ~n17425 ;
  assign n17427 = ~n5497 & ~n17424 ;
  assign n17428 = n17426 & ~n17427 ;
  assign n17429 = \u4_csr_reg[2]/NET0131  & ~n3617 ;
  assign n17430 = ~n3671 & ~n17429 ;
  assign n17431 = ~\u2_wack_r_reg/P0001  & ~n8189 ;
  assign n17432 = ~n8184 & n17431 ;
  assign n17433 = ~\u1_u2_word_done_r_reg/P0001  & ~n17432 ;
  assign n17434 = ~n8180 & n17433 ;
  assign n17435 = \u1_u2_adr_cw_reg[0]/NET0131  & ~n17434 ;
  assign n17436 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[2]_pad  ;
  assign n17437 = ~n17432 & n17436 ;
  assign n17438 = ~n8180 & n17437 ;
  assign n17439 = ~n17435 & ~n17438 ;
  assign n17440 = \u1_u2_adr_cw_reg[10]/P0001  & ~n17434 ;
  assign n17441 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[12]_pad  ;
  assign n17442 = ~n17432 & n17441 ;
  assign n17443 = ~n8180 & n17442 ;
  assign n17444 = ~n17440 & ~n17443 ;
  assign n17445 = \u1_u2_adr_cw_reg[11]/P0001  & ~n17434 ;
  assign n17446 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[13]_pad  ;
  assign n17447 = ~n17432 & n17446 ;
  assign n17448 = ~n8180 & n17447 ;
  assign n17449 = ~n17445 & ~n17448 ;
  assign n17450 = \u1_u2_adr_cw_reg[12]/P0001  & ~n17434 ;
  assign n17451 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[14]_pad  ;
  assign n17452 = ~n17432 & n17451 ;
  assign n17453 = ~n8180 & n17452 ;
  assign n17454 = ~n17450 & ~n17453 ;
  assign n17455 = \u1_u2_adr_cw_reg[13]/P0001  & ~n17434 ;
  assign n17456 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[15]_pad  ;
  assign n17457 = ~n17432 & n17456 ;
  assign n17458 = ~n8180 & n17457 ;
  assign n17459 = ~n17455 & ~n17458 ;
  assign n17460 = \u1_u2_adr_cw_reg[14]/P0001  & ~n17434 ;
  assign n17461 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[16]_pad  ;
  assign n17462 = ~n17432 & n17461 ;
  assign n17463 = ~n8180 & n17462 ;
  assign n17464 = ~n17460 & ~n17463 ;
  assign n17465 = \u1_u2_adr_cw_reg[1]/P0001  & ~n17434 ;
  assign n17466 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[3]_pad  ;
  assign n17467 = ~n17432 & n17466 ;
  assign n17468 = ~n8180 & n17467 ;
  assign n17469 = ~n17465 & ~n17468 ;
  assign n17470 = \u1_u2_adr_cw_reg[2]/P0001  & ~n17434 ;
  assign n17471 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[4]_pad  ;
  assign n17472 = ~n17432 & n17471 ;
  assign n17473 = ~n8180 & n17472 ;
  assign n17474 = ~n17470 & ~n17473 ;
  assign n17475 = \u1_u2_adr_cw_reg[3]/NET0131  & ~n17434 ;
  assign n17476 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[5]_pad  ;
  assign n17477 = ~n17432 & n17476 ;
  assign n17478 = ~n8180 & n17477 ;
  assign n17479 = ~n17475 & ~n17478 ;
  assign n17480 = \u1_u2_adr_cw_reg[4]/P0001  & ~n17434 ;
  assign n17481 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[6]_pad  ;
  assign n17482 = ~n17432 & n17481 ;
  assign n17483 = ~n8180 & n17482 ;
  assign n17484 = ~n17480 & ~n17483 ;
  assign n17485 = \u1_u2_adr_cw_reg[5]/NET0131  & ~n17434 ;
  assign n17486 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[7]_pad  ;
  assign n17487 = ~n17432 & n17486 ;
  assign n17488 = ~n8180 & n17487 ;
  assign n17489 = ~n17485 & ~n17488 ;
  assign n17490 = \u1_u2_adr_cw_reg[6]/NET0131  & ~n17434 ;
  assign n17491 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[8]_pad  ;
  assign n17492 = ~n17432 & n17491 ;
  assign n17493 = ~n8180 & n17492 ;
  assign n17494 = ~n17490 & ~n17493 ;
  assign n17495 = \u1_u2_adr_cw_reg[7]/NET0131  & ~n17434 ;
  assign n17496 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[9]_pad  ;
  assign n17497 = ~n17432 & n17496 ;
  assign n17498 = ~n8180 & n17497 ;
  assign n17499 = ~n17495 & ~n17498 ;
  assign n17500 = \u1_u2_adr_cw_reg[8]/P0001  & ~n17434 ;
  assign n17501 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[10]_pad  ;
  assign n17502 = ~n17432 & n17501 ;
  assign n17503 = ~n8180 & n17502 ;
  assign n17504 = ~n17500 & ~n17503 ;
  assign n17505 = \u1_u2_adr_cw_reg[9]/NET0131  & ~n17434 ;
  assign n17506 = ~\u1_u2_word_done_r_reg/P0001  & \wb_addr_i[11]_pad  ;
  assign n17507 = ~n17432 & n17506 ;
  assign n17508 = ~n8180 & n17507 ;
  assign n17509 = ~n17505 & ~n17508 ;
  assign n17510 = \u1_u2_dout_r_reg[0]/P0001  & ~n17434 ;
  assign n17511 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[0]_pad  ;
  assign n17512 = ~n17432 & n17511 ;
  assign n17513 = ~n8180 & n17512 ;
  assign n17514 = ~n17510 & ~n17513 ;
  assign n17515 = \u1_u2_dout_r_reg[10]/P0001  & ~n17434 ;
  assign n17516 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[10]_pad  ;
  assign n17517 = ~n17432 & n17516 ;
  assign n17518 = ~n8180 & n17517 ;
  assign n17519 = ~n17515 & ~n17518 ;
  assign n17520 = \u1_u2_dout_r_reg[11]/P0001  & ~n17434 ;
  assign n17521 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[11]_pad  ;
  assign n17522 = ~n17432 & n17521 ;
  assign n17523 = ~n8180 & n17522 ;
  assign n17524 = ~n17520 & ~n17523 ;
  assign n17525 = \u1_u2_dout_r_reg[12]/P0001  & ~n17434 ;
  assign n17526 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[12]_pad  ;
  assign n17527 = ~n17432 & n17526 ;
  assign n17528 = ~n8180 & n17527 ;
  assign n17529 = ~n17525 & ~n17528 ;
  assign n17530 = \u1_u2_dout_r_reg[13]/P0001  & ~n17434 ;
  assign n17531 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[13]_pad  ;
  assign n17532 = ~n17432 & n17531 ;
  assign n17533 = ~n8180 & n17532 ;
  assign n17534 = ~n17530 & ~n17533 ;
  assign n17535 = \u1_u2_dout_r_reg[14]/P0001  & ~n17434 ;
  assign n17536 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[14]_pad  ;
  assign n17537 = ~n17432 & n17536 ;
  assign n17538 = ~n8180 & n17537 ;
  assign n17539 = ~n17535 & ~n17538 ;
  assign n17540 = \u1_u2_dout_r_reg[15]/P0001  & ~n17434 ;
  assign n17541 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[15]_pad  ;
  assign n17542 = ~n17432 & n17541 ;
  assign n17543 = ~n8180 & n17542 ;
  assign n17544 = ~n17540 & ~n17543 ;
  assign n17545 = \u1_u2_dout_r_reg[16]/P0001  & ~n17434 ;
  assign n17546 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[16]_pad  ;
  assign n17547 = ~n17432 & n17546 ;
  assign n17548 = ~n8180 & n17547 ;
  assign n17549 = ~n17545 & ~n17548 ;
  assign n17550 = \u1_u2_dout_r_reg[17]/P0001  & ~n17434 ;
  assign n17551 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[17]_pad  ;
  assign n17552 = ~n17432 & n17551 ;
  assign n17553 = ~n8180 & n17552 ;
  assign n17554 = ~n17550 & ~n17553 ;
  assign n17555 = \u1_u2_dout_r_reg[18]/P0001  & ~n17434 ;
  assign n17556 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[18]_pad  ;
  assign n17557 = ~n17432 & n17556 ;
  assign n17558 = ~n8180 & n17557 ;
  assign n17559 = ~n17555 & ~n17558 ;
  assign n17560 = \u1_u2_dout_r_reg[19]/P0001  & ~n17434 ;
  assign n17561 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[19]_pad  ;
  assign n17562 = ~n17432 & n17561 ;
  assign n17563 = ~n8180 & n17562 ;
  assign n17564 = ~n17560 & ~n17563 ;
  assign n17565 = \u1_u2_dout_r_reg[1]/P0001  & ~n17434 ;
  assign n17566 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[1]_pad  ;
  assign n17567 = ~n17432 & n17566 ;
  assign n17568 = ~n8180 & n17567 ;
  assign n17569 = ~n17565 & ~n17568 ;
  assign n17570 = \u1_u2_dout_r_reg[20]/P0001  & ~n17434 ;
  assign n17571 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[20]_pad  ;
  assign n17572 = ~n17432 & n17571 ;
  assign n17573 = ~n8180 & n17572 ;
  assign n17574 = ~n17570 & ~n17573 ;
  assign n17575 = \u1_u2_dout_r_reg[21]/P0001  & ~n17434 ;
  assign n17576 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[21]_pad  ;
  assign n17577 = ~n17432 & n17576 ;
  assign n17578 = ~n8180 & n17577 ;
  assign n17579 = ~n17575 & ~n17578 ;
  assign n17580 = \u1_u2_dout_r_reg[22]/P0001  & ~n17434 ;
  assign n17581 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[22]_pad  ;
  assign n17582 = ~n17432 & n17581 ;
  assign n17583 = ~n8180 & n17582 ;
  assign n17584 = ~n17580 & ~n17583 ;
  assign n17585 = \u1_u2_dout_r_reg[23]/P0001  & ~n17434 ;
  assign n17586 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[23]_pad  ;
  assign n17587 = ~n17432 & n17586 ;
  assign n17588 = ~n8180 & n17587 ;
  assign n17589 = ~n17585 & ~n17588 ;
  assign n17590 = \u1_u2_dout_r_reg[24]/P0001  & ~n17434 ;
  assign n17591 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[24]_pad  ;
  assign n17592 = ~n17432 & n17591 ;
  assign n17593 = ~n8180 & n17592 ;
  assign n17594 = ~n17590 & ~n17593 ;
  assign n17595 = \u1_u2_dout_r_reg[25]/P0001  & ~n17434 ;
  assign n17596 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[25]_pad  ;
  assign n17597 = ~n17432 & n17596 ;
  assign n17598 = ~n8180 & n17597 ;
  assign n17599 = ~n17595 & ~n17598 ;
  assign n17600 = \u1_u2_dout_r_reg[26]/P0001  & ~n17434 ;
  assign n17601 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[26]_pad  ;
  assign n17602 = ~n17432 & n17601 ;
  assign n17603 = ~n8180 & n17602 ;
  assign n17604 = ~n17600 & ~n17603 ;
  assign n17605 = \u1_u2_dout_r_reg[27]/P0001  & ~n17434 ;
  assign n17606 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[27]_pad  ;
  assign n17607 = ~n17432 & n17606 ;
  assign n17608 = ~n8180 & n17607 ;
  assign n17609 = ~n17605 & ~n17608 ;
  assign n17610 = \u1_u2_dout_r_reg[28]/P0001  & ~n17434 ;
  assign n17611 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[28]_pad  ;
  assign n17612 = ~n17432 & n17611 ;
  assign n17613 = ~n8180 & n17612 ;
  assign n17614 = ~n17610 & ~n17613 ;
  assign n17615 = \u1_u2_dout_r_reg[29]/P0001  & ~n17434 ;
  assign n17616 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[29]_pad  ;
  assign n17617 = ~n17432 & n17616 ;
  assign n17618 = ~n8180 & n17617 ;
  assign n17619 = ~n17615 & ~n17618 ;
  assign n17620 = \u1_u2_dout_r_reg[2]/P0001  & ~n17434 ;
  assign n17621 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[2]_pad  ;
  assign n17622 = ~n17432 & n17621 ;
  assign n17623 = ~n8180 & n17622 ;
  assign n17624 = ~n17620 & ~n17623 ;
  assign n17625 = \u1_u2_dout_r_reg[30]/P0001  & ~n17434 ;
  assign n17626 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[30]_pad  ;
  assign n17627 = ~n17432 & n17626 ;
  assign n17628 = ~n8180 & n17627 ;
  assign n17629 = ~n17625 & ~n17628 ;
  assign n17630 = \u1_u2_dout_r_reg[31]/P0001  & ~n17434 ;
  assign n17631 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[31]_pad  ;
  assign n17632 = ~n17432 & n17631 ;
  assign n17633 = ~n8180 & n17632 ;
  assign n17634 = ~n17630 & ~n17633 ;
  assign n17635 = \u1_u2_dout_r_reg[3]/P0001  & ~n17434 ;
  assign n17636 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[3]_pad  ;
  assign n17637 = ~n17432 & n17636 ;
  assign n17638 = ~n8180 & n17637 ;
  assign n17639 = ~n17635 & ~n17638 ;
  assign n17640 = \u1_u2_dout_r_reg[4]/P0001  & ~n17434 ;
  assign n17641 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[4]_pad  ;
  assign n17642 = ~n17432 & n17641 ;
  assign n17643 = ~n8180 & n17642 ;
  assign n17644 = ~n17640 & ~n17643 ;
  assign n17645 = \u1_u2_dout_r_reg[5]/P0001  & ~n17434 ;
  assign n17646 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[5]_pad  ;
  assign n17647 = ~n17432 & n17646 ;
  assign n17648 = ~n8180 & n17647 ;
  assign n17649 = ~n17645 & ~n17648 ;
  assign n17650 = \u1_u2_dout_r_reg[6]/P0001  & ~n17434 ;
  assign n17651 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[6]_pad  ;
  assign n17652 = ~n17432 & n17651 ;
  assign n17653 = ~n8180 & n17652 ;
  assign n17654 = ~n17650 & ~n17653 ;
  assign n17655 = \u1_u2_dout_r_reg[7]/P0001  & ~n17434 ;
  assign n17656 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[7]_pad  ;
  assign n17657 = ~n17432 & n17656 ;
  assign n17658 = ~n8180 & n17657 ;
  assign n17659 = ~n17655 & ~n17658 ;
  assign n17660 = \u1_u2_dout_r_reg[8]/P0001  & ~n17434 ;
  assign n17661 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[8]_pad  ;
  assign n17662 = ~n17432 & n17661 ;
  assign n17663 = ~n8180 & n17662 ;
  assign n17664 = ~n17660 & ~n17663 ;
  assign n17665 = \u1_u2_dout_r_reg[9]/P0001  & ~n17434 ;
  assign n17666 = ~\u1_u2_word_done_r_reg/P0001  & \wb_data_i[9]_pad  ;
  assign n17667 = ~n17432 & n17666 ;
  assign n17668 = ~n8180 & n17667 ;
  assign n17669 = ~n17665 & ~n17668 ;
  assign n17670 = \u1_u2_mwe_reg/P0001  & \u1_u2_word_done_r_reg/P0001  ;
  assign n17671 = ~\u1_u2_mack_r_reg/P0001  & \u1_u2_mwe_reg/P0001  ;
  assign n17672 = ~n8179 & n17671 ;
  assign n17673 = ~n17670 & ~n17672 ;
  assign n17674 = n2557 & n2558 ;
  assign n17675 = n9843 & n17674 ;
  assign n17676 = n9850 & ~n17675 ;
  assign n17677 = n8193 & ~n17676 ;
  assign n17678 = n17673 & ~n17677 ;
  assign n17679 = \wb_addr_i[4]_pad  & n8820 ;
  assign n17680 = n14065 & n17679 ;
  assign n17681 = \u4_utmi_vend_ctrl_r_reg[0]/P0001  & ~n17680 ;
  assign n17682 = \wb_data_i[0]_pad  & n17679 ;
  assign n17683 = n14065 & n17682 ;
  assign n17684 = ~n17681 & ~n17683 ;
  assign n17685 = \u4_utmi_vend_ctrl_r_reg[1]/P0001  & ~n17680 ;
  assign n17686 = \wb_data_i[1]_pad  & n17679 ;
  assign n17687 = n14065 & n17686 ;
  assign n17688 = ~n17685 & ~n17687 ;
  assign n17689 = \u4_utmi_vend_ctrl_r_reg[2]/P0001  & ~n17680 ;
  assign n17690 = \wb_data_i[2]_pad  & n17679 ;
  assign n17691 = n14065 & n17690 ;
  assign n17692 = ~n17689 & ~n17691 ;
  assign n17693 = \u4_utmi_vend_ctrl_r_reg[3]/P0001  & ~n17680 ;
  assign n17694 = \wb_addr_i[4]_pad  & \wb_data_i[3]_pad  ;
  assign n17695 = n8820 & n17694 ;
  assign n17696 = n14065 & n17695 ;
  assign n17697 = ~n17693 & ~n17696 ;
  assign \dma_req_o[6]_pad  = 1'b0 ;
  assign \g37425/_0_  = ~n1878 ;
  assign \g37426/_0_  = ~n1936 ;
  assign \g37432/_0_  = ~n1998 ;
  assign \g37433/_0_  = ~n2056 ;
  assign \g37439/_0_  = ~n2298 ;
  assign \g37440/_0_  = ~n2349 ;
  assign \g37444/_00_  = ~n2395 ;
  assign \g37448/_0_  = ~n2420 ;
  assign \g37450/_0_  = ~n2426 ;
  assign \g37454/_0_  = ~n2458 ;
  assign \g37473/_0_  = ~n2472 ;
  assign \g37474/_0_  = ~n2487 ;
  assign \g37475/_0_  = ~n2499 ;
  assign \g37476/_0_  = ~n2517 ;
  assign \g37477/_0_  = ~n2529 ;
  assign \g37478/_0_  = ~n2543 ;
  assign \g37479/_0_  = ~n2555 ;
  assign \g37488/_0_  = ~n2582 ;
  assign \g37489/_0_  = ~n2601 ;
  assign \g37490/_0_  = ~n2618 ;
  assign \g37491/_0_  = ~n2633 ;
  assign \g37492/_0_  = ~n2648 ;
  assign \g37517/_0_  = ~n2659 ;
  assign \g37518/_0_  = ~n2669 ;
  assign \g37519/_0_  = ~n2679 ;
  assign \g37520/_0_  = ~n2689 ;
  assign \g37521/_0_  = ~n2702 ;
  assign \g37522/_0_  = n2719 ;
  assign \g37540/_0_  = ~n2730 ;
  assign \g37542/_0_  = ~n2743 ;
  assign \g37543/_0_  = ~n2753 ;
  assign \g37545/_0_  = ~n2763 ;
  assign \g37546/_0_  = ~n2773 ;
  assign \g37548/_0_  = ~n2783 ;
  assign \g37549/_0_  = ~n2799 ;
  assign \g37550/_0_  = ~n2809 ;
  assign \g37551/_0_  = ~n2819 ;
  assign \g37556/_0_  = n2835 ;
  assign \g37589/_0_  = ~n2843 ;
  assign \g37591/_0_  = ~n2854 ;
  assign \g37592/_0_  = ~n2865 ;
  assign \g37593/_0_  = ~n2874 ;
  assign \g37594/_0_  = ~n2885 ;
  assign \g37596/_0_  = ~n2895 ;
  assign \g37597/_0_  = ~n2905 ;
  assign \g37598/_0_  = ~n2915 ;
  assign \g37599/_0_  = ~n2923 ;
  assign \g37601/_0_  = ~n2933 ;
  assign \g37603/_0_  = ~n2943 ;
  assign \g37604/_0_  = ~n2951 ;
  assign \g37605/_0_  = ~n2961 ;
  assign \g37607/_0_  = ~n2971 ;
  assign \g37608/_0_  = ~n2981 ;
  assign \g37609/_0_  = ~n2989 ;
  assign \g37610/_0_  = ~n2999 ;
  assign \g37645/_0_  = ~n3008 ;
  assign \g37648/_0_  = ~n3016 ;
  assign \g37650/_0_  = ~n3024 ;
  assign \g37653/_0_  = ~n3032 ;
  assign \g37664/_3_  = ~n3038 ;
  assign \g37703/_0_  = ~n3049 ;
  assign \g37704/_0_  = ~n3060 ;
  assign \g37706/_0_  = ~n3071 ;
  assign \g37708/_0_  = ~n3080 ;
  assign \g37709/_0_  = ~n3089 ;
  assign \g37711/_0_  = ~n3098 ;
  assign \g37714/_0_  = ~n3108 ;
  assign \g37715/_0_  = ~n3118 ;
  assign \g37717/_0_  = ~n3128 ;
  assign \g37718/_0_  = ~n3136 ;
  assign \g37719/_0_  = ~n3144 ;
  assign \g37720/_0_  = ~n3152 ;
  assign \g37723/_0_  = ~n3162 ;
  assign \g37724/_0_  = ~n3172 ;
  assign \g37726/_0_  = ~n3182 ;
  assign \g37728/_0_  = ~n3190 ;
  assign \g37729/_0_  = ~n3198 ;
  assign \g37730/_0_  = ~n3206 ;
  assign \g37731/_0_  = ~n3216 ;
  assign \g37732/_0_  = ~n3226 ;
  assign \g37733/_0_  = ~n3236 ;
  assign \g37735/_0_  = ~n3244 ;
  assign \g37736/_0_  = ~n3252 ;
  assign \g37737/_0_  = ~n3260 ;
  assign \g37856/_0_  = ~n3269 ;
  assign \g37857/_0_  = ~n3278 ;
  assign \g37859/_0_  = ~n3287 ;
  assign \g37868/_0_  = ~n3295 ;
  assign \g37869/_0_  = ~n3303 ;
  assign \g37870/_0_  = ~n3311 ;
  assign \g37872/_0_  = n3360 ;
  assign \g37886/_0_  = ~n3368 ;
  assign \g37887/_0_  = ~n3376 ;
  assign \g37889/_0_  = ~n3384 ;
  assign \g37897/_0_  = ~n3392 ;
  assign \g37899/_0_  = ~n3400 ;
  assign \g37900/_0_  = ~n3408 ;
  assign \g37907/_0_  = n3420 ;
  assign \g37925/_0_  = ~n3467 ;
  assign \g37927/_0_  = ~n3633 ;
  assign \g37928/_0_  = ~n3648 ;
  assign \g37929/_0_  = n3657 ;
  assign \g37930/_0_  = ~n3668 ;
  assign \g37932/_0_  = ~n3688 ;
  assign \g37933/_0_  = ~n3701 ;
  assign \g37934/_0_  = ~n3717 ;
  assign \g37935/_0_  = ~n3730 ;
  assign \g37936/_0_  = ~n3742 ;
  assign \g37937/_0_  = ~n3755 ;
  assign \g37938/_0_  = ~n3768 ;
  assign \g37939/_0_  = ~n3785 ;
  assign \g37941/_0_  = ~n3797 ;
  assign \g37942/_0_  = ~n3805 ;
  assign \g37943/_0_  = ~n3813 ;
  assign \g37944/_0_  = ~n3821 ;
  assign \g37945/_0_  = ~n3829 ;
  assign \g38030/_3_  = ~n4017 ;
  assign \g38035/_0_  = n4030 ;
  assign \g38036/_0_  = n4041 ;
  assign \g38054/_0_  = n4052 ;
  assign \g38129/_0_  = n4058 ;
  assign \g38130/_0_  = ~n4119 ;
  assign \g38148/_3_  = ~n4135 ;
  assign \g38149/_3_  = ~n4163 ;
  assign \g38150/_3_  = ~n4179 ;
  assign \g38166/_0_  = n4193 ;
  assign \g38198/_0_  = ~n4200 ;
  assign \g38201/_0_  = ~n4235 ;
  assign \g38257/_0_  = ~n4243 ;
  assign \g38286/_0_  = ~n4266 ;
  assign \g38294/_3_  = ~n4283 ;
  assign \g38295/_3_  = ~n4293 ;
  assign \g38296/_3_  = ~n4307 ;
  assign \g38297/_3_  = ~n4319 ;
  assign \g38332/_0_  = n4320 ;
  assign \g38350/_0_  = n4321 ;
  assign \g38365/_3_  = ~n4333 ;
  assign \g38366/_3_  = ~n4345 ;
  assign \g38367/_3_  = ~n4353 ;
  assign \g38389/_0_  = n4354 ;
  assign \g38397/_0_  = n4365 ;
  assign \g38398/_0_  = n4376 ;
  assign \g38399/_0_  = n4387 ;
  assign \g38400/_0_  = n4398 ;
  assign \g38417/_3_  = ~n4413 ;
  assign \g38418/_3_  = n4432 ;
  assign \g38422/_0_  = ~n4487 ;
  assign \g38440/_0_  = n4500 ;
  assign \g38443/_0_  = ~n4520 ;
  assign \g38448/_3_  = ~n4523 ;
  assign \g38449/_0_  = ~n4529 ;
  assign \g38450/_0_  = n4554 ;
  assign \g38460/_0_  = ~n4770 ;
  assign \g38466/_0_  = ~n4775 ;
  assign \g38467/_0_  = ~n4782 ;
  assign \g38468/_0_  = ~n4787 ;
  assign \g38469/_0_  = ~n4792 ;
  assign \g38470/_0_  = ~n4799 ;
  assign \g38471/_0_  = ~n4804 ;
  assign \g38472/_0_  = ~n4811 ;
  assign \g38473/_0_  = ~n4816 ;
  assign \g38474/_0_  = ~n4821 ;
  assign \g38475/_0_  = ~n4828 ;
  assign \g38476/_0_  = ~n4833 ;
  assign \g38477/_0_  = ~n4838 ;
  assign \g38478/_0_  = ~n4847 ;
  assign \g38479/_0_  = ~n4852 ;
  assign \g38528/_0_  = n4858 ;
  assign \g38533/_0_  = ~n4866 ;
  assign \g38534/_0_  = n4868 ;
  assign \g38536/_0_  = n4879 ;
  assign \g38545/_0_  = ~n4890 ;
  assign \g38551/_0_  = ~n4489 ;
  assign \g38554/_0_  = ~n4897 ;
  assign \g38555/_0_  = ~n4905 ;
  assign \g38556/_0_  = ~n5121 ;
  assign \g38575/_0_  = n5124 ;
  assign \g38616/_0_  = ~n5125 ;
  assign \g38653/_0_  = ~n5201 ;
  assign \g38656/_0_  = ~n5250 ;
  assign \g38657/_0_  = ~n5299 ;
  assign \g38658/_0_  = ~n5348 ;
  assign \g38660/_0_  = ~n5397 ;
  assign \g38706/_0_  = n5415 ;
  assign \g38716/_0_  = n5435 ;
  assign \g38717/_0_  = ~n5444 ;
  assign \g38738/_1_  = ~n1750 ;
  assign \g38763/_0_  = ~n5448 ;
  assign \g38790/_0_  = n5452 ;
  assign \g38792/_0_  = n5456 ;
  assign \g38801/_0_  = n5460 ;
  assign \g38803/_0_  = n5464 ;
  assign \g38804/_0_  = ~n5475 ;
  assign \g38805/_0_  = ~n5484 ;
  assign \g38806/_0_  = ~n5505 ;
  assign \g38807/_0_  = ~n5517 ;
  assign \g38808/_0_  = ~n5529 ;
  assign \g38809/_0_  = ~n5541 ;
  assign \g38810/_0_  = ~n5553 ;
  assign \g38814/_0_  = ~n5575 ;
  assign \g38833/_0_  = n5589 ;
  assign \g38834/_0_  = n5594 ;
  assign \g38839/_0_  = ~n5601 ;
  assign \g38840/_0_  = ~n5608 ;
  assign \g38841/_0_  = ~n5615 ;
  assign \g38842/_0_  = ~n5622 ;
  assign \g38846/_0_  = ~n5631 ;
  assign \g38847/_0_  = ~n5637 ;
  assign \g38848/_0_  = n5646 ;
  assign \g38849/_0_  = n5654 ;
  assign \g38853/_0_  = ~n5665 ;
  assign \g38857/_0_  = n5668 ;
  assign \g38872/_0_  = ~n5733 ;
  assign \g38882/_0_  = ~n5775 ;
  assign \g38884/_0_  = ~n5813 ;
  assign \g38885/_0_  = ~n5851 ;
  assign \g38886/_0_  = ~n5889 ;
  assign \g38887/_0_  = ~n5927 ;
  assign \g38931/_0_  = n5934 ;
  assign \g38952/_0_  = n5943 ;
  assign \g38960/_0_  = n5979 ;
  assign \g38971/_0_  = n5986 ;
  assign \g38973/_0_  = n5989 ;
  assign \g38974/_0_  = n5992 ;
  assign \g38975/_0_  = n5997 ;
  assign \g38976/_0_  = ~n6004 ;
  assign \g38978/_0_  = n6007 ;
  assign \g38981/_0_  = n6010 ;
  assign \g38986/_0_  = n6013 ;
  assign \g38987/_0_  = n6022 ;
  assign \g39001/_3_  = ~n6024 ;
  assign \g39003/_3_  = n6025 ;
  assign \g39009/_3_  = ~n6027 ;
  assign \g39011/_3_  = ~n6029 ;
  assign \g39013/_3_  = ~n6031 ;
  assign \g39015/_2_  = ~n6033 ;
  assign \g39017/_2_  = ~n6035 ;
  assign \g39019/_2_  = ~n6037 ;
  assign \g39021/_2_  = ~n6039 ;
  assign \g39060/_0_  = ~n6045 ;
  assign \g39061/_3_  = ~n6048 ;
  assign \g39062/_0_  = ~n6051 ;
  assign \g39063/_0_  = ~n6062 ;
  assign \g39065/_0_  = ~n6072 ;
  assign \g39066/_0_  = ~n6081 ;
  assign \g39093/_0_  = n6129 ;
  assign \g39099/_2_  = n6211 ;
  assign \g39118/_0_  = ~n6227 ;
  assign \g39123/_0_  = ~n6241 ;
  assign \g39174/_0_  = ~n6299 ;
  assign \g39175/_0_  = ~n6356 ;
  assign \g39176/_0_  = ~n6414 ;
  assign \g39177/_0_  = n6476 ;
  assign \g39178/_0_  = n6482 ;
  assign \g39185/_0_  = n6486 ;
  assign \g39186/_0_  = n6491 ;
  assign \g39187/_0_  = ~n6498 ;
  assign \g39188/_0_  = n6500 ;
  assign \g39194/_0_  = n6504 ;
  assign \g39195/_0_  = n6508 ;
  assign \g39196/_0_  = n6512 ;
  assign \g39197/_0_  = n6516 ;
  assign \g39198/_0_  = n6520 ;
  assign \g39199/_0_  = n6524 ;
  assign \g39200/_0_  = n6528 ;
  assign \g39201/_0_  = n6532 ;
  assign \g39202/_0_  = n6536 ;
  assign \g39203/_0_  = n6540 ;
  assign \g39204/_0_  = n6544 ;
  assign \g39216/_3_  = ~n6547 ;
  assign \g39217/_3_  = ~n6550 ;
  assign \g39218/_0_  = ~n6553 ;
  assign \g39219/_0_  = ~n6556 ;
  assign \g39220/_0_  = ~n6562 ;
  assign \g39221/_0_  = n6570 ;
  assign \g39299/_0_  = ~n6604 ;
  assign \g39300/_0_  = ~n6638 ;
  assign \g39301/_0_  = n6666 ;
  assign \g39302/_0_  = n6694 ;
  assign \g39303/_0_  = n6705 ;
  assign \g39304/_0_  = n6708 ;
  assign \g39305/_0_  = n6720 ;
  assign \g39306/_0_  = n6728 ;
  assign \g39307/_0_  = n6735 ;
  assign \g39308/_0_  = n6799 ;
  assign \g39309/_0_  = n6863 ;
  assign \g39310/_0_  = n6927 ;
  assign \g39311/_0_  = n6992 ;
  assign \g39315/_0_  = n6994 ;
  assign \g39318/_0_  = n7002 ;
  assign \g39321/_0_  = n7007 ;
  assign \g39322/_0_  = n7009 ;
  assign \g39323/_0_  = n7024 ;
  assign \g39333/_0_  = n7030 ;
  assign \g39334/_0_  = n7037 ;
  assign \g39336/_0_  = n7045 ;
  assign \g39338/_0_  = n7052 ;
  assign \g39339/_0_  = n7060 ;
  assign \g39340/_0_  = n7070 ;
  assign \g39341/_0_  = n7077 ;
  assign \g39342/_0_  = n7085 ;
  assign \g39343/_0_  = n7090 ;
  assign \g39344/_0_  = n7097 ;
  assign \g39345/_0_  = n7103 ;
  assign \g39346/_0_  = n7109 ;
  assign \g39349/_0_  = n7117 ;
  assign \g39352/_3_  = n7122 ;
  assign \g39354/_3_  = n7171 ;
  assign \g39371/_3_  = ~n7174 ;
  assign \g39372/_3_  = ~n7177 ;
  assign \g39373/_3_  = ~n7180 ;
  assign \g39374/_3_  = ~n7183 ;
  assign \g39376/_0_  = ~n7191 ;
  assign \g39377/_0_  = ~n7197 ;
  assign \g39471/_0_  = n7215 ;
  assign \g39472/_0_  = n7236 ;
  assign \g39473/_0_  = n7257 ;
  assign \g39474/_0_  = n7283 ;
  assign \g39475/_0_  = ~n7300 ;
  assign \g39476/_0_  = ~n7331 ;
  assign \g39477/_0_  = n7350 ;
  assign \g39478/_0_  = ~n7381 ;
  assign \g39479/_0_  = n7400 ;
  assign \g39480/_0_  = ~n7431 ;
  assign \g39481/_0_  = n7450 ;
  assign \g39482/_0_  = ~n7481 ;
  assign \g39483/_0_  = n7500 ;
  assign \g39484/_0_  = n7531 ;
  assign \g39485/_0_  = n7561 ;
  assign \g39486/_0_  = ~n7577 ;
  assign \g39487/_0_  = n7589 ;
  assign \g39488/_0_  = n7597 ;
  assign \g39492/_0_  = n7600 ;
  assign \g39497/_0_  = n7604 ;
  assign \g39501/_0_  = n7609 ;
  assign \g39502/_0_  = n7615 ;
  assign \g39503/_0_  = n7623 ;
  assign \g39504/_0_  = n7628 ;
  assign \g39505/_0_  = n7635 ;
  assign \g39506/_0_  = n7643 ;
  assign \g39539/_0_  = ~n7653 ;
  assign \g39541/_0_  = n7659 ;
  assign \g39542/_0_  = ~n7664 ;
  assign \g39543/_0_  = n7668 ;
  assign \g39544/_0_  = ~n7673 ;
  assign \g39545/_0_  = n7679 ;
  assign \g39546/_0_  = n7682 ;
  assign \g39547/_0_  = ~n7687 ;
  assign \g39550/_0_  = n7694 ;
  assign \g39551/_0_  = ~n7700 ;
  assign \g39563/_0_  = n7702 ;
  assign \g39568/_00_  = ~n7760 ;
  assign \g39617/_0_  = ~n7763 ;
  assign \g39618/_0_  = ~n7766 ;
  assign \g39621/_0_  = ~n7774 ;
  assign \g39622/_0_  = ~n7783 ;
  assign \g39623/_0_  = ~n7793 ;
  assign \g39624/_00_  = n7805 ;
  assign \g39685/_0_  = ~n7813 ;
  assign \g39690/_0_  = n7877 ;
  assign \g39693/_0_  = n7942 ;
  assign \g39695/_0_  = n7951 ;
  assign \g39697/_0_  = n7952 ;
  assign \g39706/_0_  = ~n7962 ;
  assign \g39749/_0_  = ~n7971 ;
  assign \g39750/_0_  = ~n7978 ;
  assign \g39751/_0_  = ~n7985 ;
  assign \g39752/_0_  = ~n7992 ;
  assign \g39753/_0_  = ~n7999 ;
  assign \g39754/_0_  = ~n8006 ;
  assign \g39755/_0_  = ~n8015 ;
  assign \g39756/_0_  = ~n8023 ;
  assign \g39757/_0_  = ~n8030 ;
  assign \g39758/_0_  = ~n8038 ;
  assign \g39759/_0_  = ~n8044 ;
  assign \g39760/_0_  = ~n8050 ;
  assign \g39761/_0_  = ~n8056 ;
  assign \g39762/_0_  = ~n8062 ;
  assign \g39763/_0_  = ~n8071 ;
  assign \g39764/_0_  = ~n8077 ;
  assign \g39765/_0_  = ~n8083 ;
  assign \g39766/_0_  = ~n8090 ;
  assign \g39767/_0_  = ~n8096 ;
  assign \g39768/_0_  = ~n8102 ;
  assign \g39769/_0_  = ~n8108 ;
  assign \g39770/_0_  = ~n8114 ;
  assign \g39772/_0_  = ~n8120 ;
  assign \g39773/_0_  = ~n8126 ;
  assign \g39775/_3_  = ~n8134 ;
  assign \g39776/_3_  = ~n8140 ;
  assign \g39777/_3_  = ~n8146 ;
  assign \g39778/_3_  = ~n8153 ;
  assign \g39779/_3_  = ~n8159 ;
  assign \g39780/_3_  = ~n8165 ;
  assign \g39781/_3_  = ~n8171 ;
  assign \g39782/_3_  = ~n8177 ;
  assign \g39788/_3_  = n8195 ;
  assign \g39799/_0_  = ~n8203 ;
  assign \g39800/_0_  = ~n8214 ;
  assign \g39801/_0_  = n8226 ;
  assign \g39802/_0_  = n8237 ;
  assign \g39927/_0_  = ~n8252 ;
  assign \g39928/_0_  = n8276 ;
  assign \g39929/_0_  = n8300 ;
  assign \g39930/_0_  = n8323 ;
  assign \g39931/_0_  = n8350 ;
  assign \g39932/_0_  = n8374 ;
  assign \g39933/_0_  = ~n8398 ;
  assign \g39934/_0_  = n8422 ;
  assign \g39935/_0_  = ~n8446 ;
  assign \g39936/_0_  = n8461 ;
  assign \g39937/_0_  = n8476 ;
  assign \g39938/_0_  = n8491 ;
  assign \g39939/_0_  = n8506 ;
  assign \g39940/_0_  = n8517 ;
  assign \g39942/_0_  = ~n8542 ;
  assign \g39943/_0_  = ~n8569 ;
  assign \g39944/_0_  = n8593 ;
  assign \g39945/_0_  = n8617 ;
  assign \g39956/_0_  = n8622 ;
  assign \g39957/_0_  = n8627 ;
  assign \g39958/_0_  = ~n8634 ;
  assign \g39959/_0_  = n8640 ;
  assign \g39960/_0_  = n8643 ;
  assign \g39961/_0_  = ~n8648 ;
  assign \g39962/_0_  = n8654 ;
  assign \g39963/_0_  = ~n8659 ;
  assign \g39964/_0_  = n8680 ;
  assign \g39969/_0_  = n8743 ;
  assign \g39974/_0_  = n8807 ;
  assign \g39975/_0_  = n8808 ;
  assign \g39993/_0_  = n8811 ;
  assign \g39994/_0_  = n8814 ;
  assign \g40003/_0_  = ~n8876 ;
  assign \g40004/_0_  = ~n8930 ;
  assign \g40005/_0_  = ~n8984 ;
  assign \g40006/_0_  = ~n9038 ;
  assign \g40016/_0_  = ~n9047 ;
  assign \g40023/_3_  = ~n9050 ;
  assign \g40033/_0_  = ~n9055 ;
  assign \g40034/_0_  = n9060 ;
  assign \g40035/_0_  = ~n9109 ;
  assign \g40036/_0_  = ~n9158 ;
  assign \g40037/_0_  = ~n9207 ;
  assign \g40038/_0_  = ~n9256 ;
  assign \g40199/_0_  = n9276 ;
  assign \g40200/_0_  = ~n9301 ;
  assign \g40201/_0_  = n9321 ;
  assign \g40202/_0_  = ~n9346 ;
  assign \g40203/_0_  = ~n9369 ;
  assign \g40204/_0_  = ~n9394 ;
  assign \g40205/_0_  = n9415 ;
  assign \g40206/_0_  = n9439 ;
  assign \g40207/_0_  = n9462 ;
  assign \g40208/_0_  = n9485 ;
  assign \g40209/_0_  = n9510 ;
  assign \g40210/_0_  = n9535 ;
  assign \g40224/_0_  = n9560 ;
  assign \g40225/_0_  = n9585 ;
  assign \g40226/_0_  = n9610 ;
  assign \g40227/_0_  = n9635 ;
  assign \g40234/_0_  = ~n9644 ;
  assign \g40235/_0_  = ~n9653 ;
  assign \g40236/_0_  = ~n9662 ;
  assign \g40237/_0_  = ~n9671 ;
  assign \g40238/_0_  = ~n9680 ;
  assign \g40239/_0_  = ~n9689 ;
  assign \g40240/_0_  = ~n9698 ;
  assign \g40241/_0_  = ~n9707 ;
  assign \g40242/_0_  = ~n9716 ;
  assign \g40243/_0_  = ~n9725 ;
  assign \g40244/_0_  = ~n9734 ;
  assign \g40246/_0_  = ~n9743 ;
  assign \g40247/_0_  = ~n9752 ;
  assign \g40248/_0_  = ~n9761 ;
  assign \g40249/_0_  = ~n9770 ;
  assign \g40250/_0_  = ~n9779 ;
  assign \g40251/_0_  = ~n9788 ;
  assign \g40252/_0_  = ~n9797 ;
  assign \g40253/_0_  = ~n9806 ;
  assign \g40254/_0_  = ~n9815 ;
  assign \g40255/_0_  = ~n9824 ;
  assign \g40257/_0_  = ~n9833 ;
  assign \g40258/_0_  = ~n9842 ;
  assign \g40262/_0_  = ~n9854 ;
  assign \g40264/_0_  = ~n9855 ;
  assign \g40265/_0_  = n9864 ;
  assign \g40266/_0_  = ~n9872 ;
  assign \g40267/_0_  = ~n9880 ;
  assign \g40268/_0_  = ~n9888 ;
  assign \g40269/_0_  = ~n9896 ;
  assign \g40270/_0_  = ~n9904 ;
  assign \g40271/_0_  = ~n9912 ;
  assign \g40272/_0_  = ~n9920 ;
  assign \g40273/_0_  = ~n9928 ;
  assign \g40274/_0_  = ~n9936 ;
  assign \g40275/_0_  = ~n9944 ;
  assign \g40276/_0_  = ~n9952 ;
  assign \g40277/_0_  = ~n9960 ;
  assign \g40278/_0_  = ~n9968 ;
  assign \g40280/_2_  = ~n10015 ;
  assign \g40281/_0_  = ~n10023 ;
  assign \g40282/_0_  = ~n10031 ;
  assign \g40283/_0_  = ~n10039 ;
  assign \g40284/_0_  = ~n10047 ;
  assign \g40285/_0_  = ~n10055 ;
  assign \g40286/_0_  = ~n10063 ;
  assign \g40287/_0_  = ~n10071 ;
  assign \g40288/_0_  = ~n10079 ;
  assign \g40289/_0_  = ~n10087 ;
  assign \g40290/_0_  = ~n10095 ;
  assign \g40291/_0_  = n10101 ;
  assign \g40297/_0_  = ~n10109 ;
  assign \g40298/_0_  = ~n10117 ;
  assign \g40299/_0_  = ~n10125 ;
  assign \g40300/_0_  = ~n10133 ;
  assign \g40301/_0_  = ~n10141 ;
  assign \g40302/_0_  = ~n10149 ;
  assign \g40303/_0_  = ~n10157 ;
  assign \g40304/_0_  = ~n10165 ;
  assign \g40306/_0_  = ~n10173 ;
  assign \g40307/_0_  = ~n10181 ;
  assign \g40308/_0_  = ~n10189 ;
  assign \g40309/_0_  = ~n10197 ;
  assign \g40310/_0_  = ~n10205 ;
  assign \g40311/_0_  = ~n10213 ;
  assign \g40312/_0_  = ~n10221 ;
  assign \g40313/_0_  = ~n10229 ;
  assign \g40314/_0_  = ~n10237 ;
  assign \g40315/_0_  = ~n10245 ;
  assign \g40316/_0_  = ~n10253 ;
  assign \g40317/_0_  = ~n10261 ;
  assign \g40318/_0_  = ~n10269 ;
  assign \g40319/_0_  = ~n10277 ;
  assign \g40320/_0_  = ~n10285 ;
  assign \g40324/_0_  = n6499 ;
  assign \g40325/_0_  = ~n10293 ;
  assign \g40326/_0_  = ~n10301 ;
  assign \g40327/_0_  = ~n10309 ;
  assign \g40328/_0_  = ~n10317 ;
  assign \g40329/_0_  = ~n10325 ;
  assign \g40330/_0_  = ~n10333 ;
  assign \g40331/_0_  = ~n10341 ;
  assign \g40332/_0_  = ~n10349 ;
  assign \g40333/_0_  = ~n10357 ;
  assign \g40334/_0_  = ~n10365 ;
  assign \g40335/_0_  = ~n10373 ;
  assign \g40336/_0_  = ~n10381 ;
  assign \g40337/_0_  = ~n10389 ;
  assign \g40338/_0_  = ~n10397 ;
  assign \g40339/_0_  = ~n10405 ;
  assign \g40340/_0_  = ~n10413 ;
  assign \g40341/_0_  = ~n10421 ;
  assign \g40342/_0_  = ~n10429 ;
  assign \g40343/_0_  = ~n10437 ;
  assign \g40344/_0_  = ~n10445 ;
  assign \g40345/_0_  = ~n10453 ;
  assign \g40346/_0_  = ~n10461 ;
  assign \g40347/_0_  = ~n10469 ;
  assign \g40350/_0_  = ~n10482 ;
  assign \g40353/_0_  = ~n10560 ;
  assign \g40354/_0_  = ~n10619 ;
  assign \g40355/_0_  = ~n10633 ;
  assign \g40374/_0_  = n10638 ;
  assign \g40457/_0_  = n10642 ;
  assign \g40458/_0_  = n10650 ;
  assign \g40549/_0_  = ~n10671 ;
  assign \g40550/_0_  = ~n10692 ;
  assign \g40551/_0_  = ~n10702 ;
  assign \g40552/_0_  = ~n10712 ;
  assign \g40553/_0_  = ~n10722 ;
  assign \g40554/_0_  = ~n10732 ;
  assign \g40556/_0_  = n10749 ;
  assign \g40557/_0_  = n10769 ;
  assign \g40558/_0_  = ~n10790 ;
  assign \g40559/_0_  = n10801 ;
  assign \g40561/_0_  = n10818 ;
  assign \g40562/_0_  = n10839 ;
  assign \g40563/_0_  = ~n10859 ;
  assign \g40565/_0_  = n10876 ;
  assign \g40566/_0_  = n10896 ;
  assign \g40567/_0_  = ~n10917 ;
  assign \g40569/_0_  = n10934 ;
  assign \g40570/_0_  = n10954 ;
  assign \g40571/_0_  = ~n10974 ;
  assign \g40572/_0_  = n10993 ;
  assign \g40573/_0_  = ~n11014 ;
  assign \g40574/_0_  = ~n11037 ;
  assign \g40575/_0_  = n11056 ;
  assign \g40576/_0_  = ~n11076 ;
  assign \g40577/_0_  = ~n11099 ;
  assign \g40578/_0_  = n11119 ;
  assign \g40579/_0_  = ~n11140 ;
  assign \g40580/_0_  = ~n11163 ;
  assign \g40581/_0_  = n11183 ;
  assign \g40582/_0_  = ~n11203 ;
  assign \g40583/_0_  = ~n11226 ;
  assign \g40584/_0_  = n11235 ;
  assign \g40586/_0_  = n11252 ;
  assign \g40587/_0_  = n11269 ;
  assign \g40588/_0_  = n11286 ;
  assign \g40589/_0_  = n11303 ;
  assign \g40591/_0_  = ~n11313 ;
  assign \g40592/_0_  = ~n11324 ;
  assign \g40593/_0_  = ~n11335 ;
  assign \g40594/_0_  = ~n11346 ;
  assign \g40595/_0_  = ~n11357 ;
  assign \g40596/_0_  = ~n11368 ;
  assign \g40597/_0_  = ~n11379 ;
  assign \g40598/_0_  = ~n11390 ;
  assign \g40599/_0_  = ~n11401 ;
  assign \g40600/_0_  = ~n11412 ;
  assign \g40601/_0_  = ~n11423 ;
  assign \g40602/_0_  = ~n11434 ;
  assign \g40603/_0_  = ~n11445 ;
  assign \g40604/_0_  = ~n11456 ;
  assign \g40605/_0_  = ~n11467 ;
  assign \g40606/_0_  = ~n11478 ;
  assign \g40607/_0_  = ~n11489 ;
  assign \g40608/_0_  = ~n11500 ;
  assign \g40609/_0_  = ~n11511 ;
  assign \g40610/_0_  = ~n11522 ;
  assign \g40611/_0_  = ~n11533 ;
  assign \g40612/_0_  = ~n11544 ;
  assign \g40613/_0_  = ~n11555 ;
  assign \g40614/_0_  = ~n11566 ;
  assign \g40617/_0_  = ~n11570 ;
  assign \g40629/_0_  = n11578 ;
  assign \g40632/_0_  = ~n11588 ;
  assign \g40633/_0_  = ~n11598 ;
  assign \g40634/_0_  = ~n11608 ;
  assign \g40635/_0_  = ~n11618 ;
  assign \g40636/_0_  = ~n11628 ;
  assign \g40637/_0_  = ~n11638 ;
  assign \g40638/_0_  = ~n11648 ;
  assign \g40639/_0_  = ~n11658 ;
  assign \g40640/_0_  = ~n11668 ;
  assign \g40641/_0_  = ~n11678 ;
  assign \g40642/_0_  = ~n11688 ;
  assign \g40643/_0_  = ~n11698 ;
  assign \g40644/_0_  = ~n11708 ;
  assign \g40645/_0_  = ~n11718 ;
  assign \g40646/_0_  = ~n11728 ;
  assign \g40647/_0_  = ~n11738 ;
  assign \g40648/_0_  = ~n11748 ;
  assign \g40649/_0_  = ~n11758 ;
  assign \g40650/_0_  = ~n11768 ;
  assign \g40651/_0_  = ~n11778 ;
  assign \g40652/_0_  = ~n11788 ;
  assign \g40653/_0_  = ~n11798 ;
  assign \g40654/_0_  = ~n11808 ;
  assign \g40655/_0_  = n11814 ;
  assign \g40661/_0_  = ~n11818 ;
  assign \g40663/_0_  = ~n11828 ;
  assign \g40664/_0_  = ~n11838 ;
  assign \g40665/_0_  = ~n11848 ;
  assign \g40666/_0_  = ~n11858 ;
  assign \g40667/_0_  = ~n11868 ;
  assign \g40668/_0_  = ~n11878 ;
  assign \g40669/_0_  = ~n11888 ;
  assign \g40670/_0_  = ~n11898 ;
  assign \g40671/_0_  = ~n11908 ;
  assign \g40672/_0_  = ~n11918 ;
  assign \g40673/_0_  = ~n11928 ;
  assign \g40674/_0_  = ~n11938 ;
  assign \g40675/_0_  = ~n11948 ;
  assign \g40676/_0_  = ~n11958 ;
  assign \g40677/_0_  = ~n11968 ;
  assign \g40678/_0_  = ~n11978 ;
  assign \g40679/_0_  = ~n11988 ;
  assign \g40680/_0_  = ~n11998 ;
  assign \g40681/_0_  = ~n12008 ;
  assign \g40682/_0_  = ~n12018 ;
  assign \g40683/_0_  = ~n12028 ;
  assign \g40684/_0_  = ~n12038 ;
  assign \g40685/_0_  = ~n12048 ;
  assign \g40689/_0_  = ~n12052 ;
  assign \g40690/_0_  = ~n12062 ;
  assign \g40691/_0_  = ~n12072 ;
  assign \g40692/_0_  = ~n12082 ;
  assign \g40693/_0_  = ~n12092 ;
  assign \g40694/_0_  = ~n12102 ;
  assign \g40695/_0_  = ~n12112 ;
  assign \g40696/_0_  = ~n12122 ;
  assign \g40697/_0_  = ~n12132 ;
  assign \g40698/_0_  = ~n12142 ;
  assign \g40699/_0_  = ~n12152 ;
  assign \g40700/_0_  = ~n12162 ;
  assign \g40701/_0_  = ~n12172 ;
  assign \g40702/_0_  = ~n12182 ;
  assign \g40703/_0_  = ~n12192 ;
  assign \g40704/_0_  = ~n12202 ;
  assign \g40705/_0_  = ~n12212 ;
  assign \g40706/_0_  = ~n12222 ;
  assign \g40707/_0_  = ~n12232 ;
  assign \g40708/_0_  = ~n12242 ;
  assign \g40709/_0_  = ~n12252 ;
  assign \g40710/_0_  = ~n12262 ;
  assign \g40711/_0_  = ~n12272 ;
  assign \g40712/_0_  = ~n12282 ;
  assign \g40758/_00_  = n12285 ;
  assign \g40759/_0_  = n12288 ;
  assign \g40812/_0_  = ~n12325 ;
  assign \g40816/_0_  = n12329 ;
  assign \g40817/_0_  = n12333 ;
  assign \g40818/_0_  = ~n12376 ;
  assign \g40819/_0_  = n12380 ;
  assign \g40820/_0_  = n12384 ;
  assign \g40822/_3_  = ~n12387 ;
  assign \g40823/_3_  = ~n12390 ;
  assign \g40824/_3_  = ~n12393 ;
  assign \g40825/_3_  = ~n12396 ;
  assign \g40849/_3_  = ~n12399 ;
  assign \g40915/_0_  = n12408 ;
  assign \g40916/_0_  = n12422 ;
  assign \g40917/_0_  = n12426 ;
  assign \g40920/_0_  = n12435 ;
  assign \g40923/_0_  = ~n12452 ;
  assign \g40926/_0_  = n12461 ;
  assign \g40927/_0_  = n12475 ;
  assign \g40930/_0_  = n12484 ;
  assign \g40931/_0_  = n12498 ;
  assign \g41138/_0_  = ~n12505 ;
  assign \g41152/_0_  = n12513 ;
  assign \g41180/_0_  = n12520 ;
  assign \g41185/_0_  = ~n12537 ;
  assign \g41186/_0_  = n12540 ;
  assign \g41187/_0_  = n12543 ;
  assign \g41189/_0_  = n12549 ;
  assign \g41190/_0_  = n12555 ;
  assign \g41191/_0_  = n12561 ;
  assign \g41192/_0_  = n12567 ;
  assign \g41193/_0_  = n12573 ;
  assign \g41195/_0_  = n12583 ;
  assign \g41199/_0_  = n12590 ;
  assign \g41207/_0_  = ~n12605 ;
  assign \g41221/_0_  = n12609 ;
  assign \g41226/_0_  = n12615 ;
  assign \g41227/_0_  = n12622 ;
  assign \g41230/_0_  = n12629 ;
  assign \g41231/_0_  = ~n12637 ;
  assign \g41234/_0_  = n12662 ;
  assign \g41238/_0_  = ~n12670 ;
  assign \g41239/_0_  = n12677 ;
  assign \g41275/_0_  = ~n12710 ;
  assign \g41277/_0_  = ~n12718 ;
  assign \g41278/_0_  = ~n12726 ;
  assign \g41279/_0_  = ~n12734 ;
  assign \g41280/_0_  = ~n12742 ;
  assign \g41281/_0_  = ~n12750 ;
  assign \g41282/_0_  = ~n12757 ;
  assign \g41283/_0_  = ~n12771 ;
  assign \g41284/_0_  = ~n12779 ;
  assign \g41285/_0_  = ~n12798 ;
  assign \g41286/_0_  = ~n12809 ;
  assign \g41287/_0_  = ~n12823 ;
  assign \g41288/_0_  = ~n12836 ;
  assign \g41289/_0_  = ~n12850 ;
  assign \g41291/_3_  = ~n12897 ;
  assign \g41330/_0_  = ~n12903 ;
  assign \g41332/_0_  = n12919 ;
  assign \g41334/_0_  = ~n12922 ;
  assign \g41340/_0_  = n12938 ;
  assign \g41343/_0_  = ~n12941 ;
  assign \g41345/_0_  = n12957 ;
  assign \g41348/_0_  = ~n12960 ;
  assign \g41349/_0_  = n12977 ;
  assign \g41350/_0_  = ~n12997 ;
  assign \g41351/_0_  = ~n13005 ;
  assign \g41356/_0_  = ~n13033 ;
  assign \g41394/_0_  = n13038 ;
  assign \g41423/_0_  = ~n13042 ;
  assign \g41426/_3_  = ~n13045 ;
  assign \g41427/_3_  = ~n13048 ;
  assign \g41428/_3_  = ~n13051 ;
  assign \g41429/_3_  = ~n13054 ;
  assign \g41430/_3_  = ~n13057 ;
  assign \g41431/_3_  = ~n13060 ;
  assign \g41432/_3_  = ~n13063 ;
  assign \g41433/_3_  = ~n13066 ;
  assign \g41434/_3_  = ~n13069 ;
  assign \g41435/_3_  = ~n13072 ;
  assign \g41436/_3_  = ~n13075 ;
  assign \g41437/_3_  = ~n13078 ;
  assign \g41438/_3_  = ~n13081 ;
  assign \g41439/_3_  = ~n13084 ;
  assign \g41440/_3_  = ~n13087 ;
  assign \g41441/_3_  = ~n13090 ;
  assign \g41442/_0_  = ~n13096 ;
  assign \g41445/_3_  = ~n13099 ;
  assign \g41446/_0_  = ~n13103 ;
  assign \g41449/_0_  = ~n13107 ;
  assign \g41464/_0_  = ~n13110 ;
  assign \g41466/_0_  = ~n13113 ;
  assign \g41468/_0_  = ~n13116 ;
  assign \g41469/_0_  = ~n13121 ;
  assign \g41471/_0_  = ~n13124 ;
  assign \g41795/_0_  = n13131 ;
  assign \g41799/_0_  = n13140 ;
  assign \g41800/_0_  = ~n13150 ;
  assign \g41801/_0_  = ~n13160 ;
  assign \g41802/_0_  = ~n13170 ;
  assign \g41803/_0_  = ~n13180 ;
  assign \g41804/_0_  = ~n13190 ;
  assign \g41805/_0_  = ~n13200 ;
  assign \g41806/_0_  = ~n13210 ;
  assign \g41807/_0_  = ~n13220 ;
  assign \g41808/_0_  = ~n13230 ;
  assign \g41809/_0_  = ~n13240 ;
  assign \g41810/_0_  = ~n13250 ;
  assign \g41811/_0_  = ~n13260 ;
  assign \g41812/_0_  = ~n13270 ;
  assign \g41814/_0_  = ~n13280 ;
  assign \g41815/_0_  = ~n13290 ;
  assign \g41816/_0_  = ~n13300 ;
  assign \g41817/_0_  = ~n13310 ;
  assign \g41818/_0_  = ~n13320 ;
  assign \g41819/_0_  = ~n13330 ;
  assign \g41820/_0_  = ~n13340 ;
  assign \g41821/_0_  = ~n13350 ;
  assign \g41822/_0_  = ~n13360 ;
  assign \g41823/_0_  = ~n13370 ;
  assign \g41825/_0_  = ~n13380 ;
  assign \g41826/_0_  = ~n13390 ;
  assign \g41827/_0_  = ~n13400 ;
  assign \g41828/_0_  = ~n13410 ;
  assign \g41829/_0_  = ~n13420 ;
  assign \g41830/_0_  = ~n13430 ;
  assign \g41831/_0_  = ~n13440 ;
  assign \g41832/_0_  = ~n13450 ;
  assign \g41833/_0_  = ~n13460 ;
  assign \g41834/_0_  = ~n13470 ;
  assign \g41835/_0_  = ~n13480 ;
  assign \g41836/_0_  = ~n13490 ;
  assign \g41837/_0_  = ~n13500 ;
  assign \g41838/_0_  = ~n13510 ;
  assign \g41839/_0_  = ~n13520 ;
  assign \g41840/_0_  = ~n13530 ;
  assign \g41841/_0_  = ~n13540 ;
  assign \g41842/_0_  = ~n13550 ;
  assign \g41843/_0_  = ~n13560 ;
  assign \g41844/_0_  = ~n13570 ;
  assign \g41845/_0_  = ~n13580 ;
  assign \g41846/_0_  = ~n13590 ;
  assign \g41847/_0_  = ~n13600 ;
  assign \g41848/_0_  = ~n13610 ;
  assign \g41849/_0_  = ~n13620 ;
  assign \g41850/_0_  = ~n13630 ;
  assign \g41851/_0_  = ~n13640 ;
  assign \g41852/_0_  = ~n13650 ;
  assign \g41853/_0_  = ~n13660 ;
  assign \g41854/_0_  = ~n13670 ;
  assign \g41855/_0_  = ~n13680 ;
  assign \g41856/_0_  = ~n13690 ;
  assign \g41857/_0_  = ~n13700 ;
  assign \g41858/_0_  = ~n13710 ;
  assign \g41859/_0_  = ~n13720 ;
  assign \g41860/_0_  = ~n13730 ;
  assign \g41861/_0_  = ~n13740 ;
  assign \g41862/_0_  = ~n13750 ;
  assign \g41863/_0_  = ~n13760 ;
  assign \g41864/_0_  = ~n13770 ;
  assign \g41865/_0_  = ~n13780 ;
  assign \g41866/_0_  = ~n13790 ;
  assign \g41867/_0_  = ~n13800 ;
  assign \g41868/_0_  = ~n13810 ;
  assign \g41869/_0_  = ~n13820 ;
  assign \g41870/_0_  = ~n13830 ;
  assign \g41871/_0_  = ~n13840 ;
  assign \g41872/_0_  = ~n13850 ;
  assign \g41873/_0_  = ~n13860 ;
  assign \g41874/_0_  = ~n13870 ;
  assign \g41875/_0_  = ~n13880 ;
  assign \g41876/_0_  = ~n13890 ;
  assign \g41877/_0_  = ~n13900 ;
  assign \g41878/_0_  = ~n13910 ;
  assign \g41879/_0_  = ~n13920 ;
  assign \g41880/_0_  = ~n13930 ;
  assign \g41881/_0_  = ~n13940 ;
  assign \g41882/_0_  = ~n13950 ;
  assign \g41883/_0_  = ~n13960 ;
  assign \g41884/_0_  = ~n13970 ;
  assign \g41885/_0_  = ~n13980 ;
  assign \g41886/_0_  = ~n13990 ;
  assign \g41887/_0_  = ~n14000 ;
  assign \g41888/_0_  = ~n14010 ;
  assign \g41889/_0_  = ~n14020 ;
  assign \g41890/_0_  = ~n14030 ;
  assign \g41891/_0_  = ~n14040 ;
  assign \g41902/_0_  = n14048 ;
  assign \g41904/_0_  = n14051 ;
  assign \g41906/_0_  = n14057 ;
  assign \g41907/_0_  = ~n14063 ;
  assign \g41954/_0_  = n14076 ;
  assign \g41955/_0_  = n14082 ;
  assign \g41956/_0_  = n14088 ;
  assign \g41957/_0_  = n14094 ;
  assign \g41958/_0_  = n14100 ;
  assign \g41959/_0_  = n14106 ;
  assign \g41960/_0_  = n14112 ;
  assign \g41962/_0_  = n14119 ;
  assign \g41963/_0_  = n14124 ;
  assign \g41964/_0_  = n14129 ;
  assign \g41965/_0_  = n14134 ;
  assign \g41966/_0_  = n14139 ;
  assign \g41967/_0_  = n14144 ;
  assign \g41968/_0_  = n14149 ;
  assign \g41969/_0_  = n14155 ;
  assign \g41970/_0_  = n14161 ;
  assign \g41971/_0_  = n14167 ;
  assign \g41972/_0_  = n14173 ;
  assign \g41973/_0_  = n14179 ;
  assign \g41974/_0_  = n14185 ;
  assign \g41975/_0_  = n14191 ;
  assign \g41976/_0_  = n14197 ;
  assign \g41977/_0_  = n14203 ;
  assign \g41978/_0_  = n14209 ;
  assign \g41979/_0_  = n14215 ;
  assign \g42062/_0_  = ~n14225 ;
  assign \g42079/_0_  = ~n14235 ;
  assign \g42142/_0_  = n14237 ;
  assign \g42143/_0_  = n14239 ;
  assign \g42144/_0_  = n14241 ;
  assign \g42154/_0_  = n14261 ;
  assign \g42157/_0_  = ~n14273 ;
  assign \g42160/_0_  = n14276 ;
  assign \g42181/_0_  = ~n14291 ;
  assign \g42203/_0_  = ~n14304 ;
  assign \g42204/_3_  = ~n14307 ;
  assign \g42205/_3_  = ~n14310 ;
  assign \g42206/_3_  = ~n14313 ;
  assign \g42208/_0_  = ~n14318 ;
  assign \g42220/_0_  = ~n14331 ;
  assign \g42225/_0_  = ~n14346 ;
  assign \g42251/_0_  = n14355 ;
  assign \g42273/_0_  = n14364 ;
  assign \g42335/_0_  = n14373 ;
  assign \g42357/_0_  = n14382 ;
  assign \g42380/_0_  = n14384 ;
  assign \g42381/_0_  = ~n14387 ;
  assign \g42383/_0_  = ~n14390 ;
  assign \g42386/_0_  = ~n14393 ;
  assign \g42388/_0_  = ~n14396 ;
  assign \g42475/_0_  = n14403 ;
  assign \g42476/_0_  = n14408 ;
  assign \g42477/_0_  = n14413 ;
  assign \g42478/_0_  = n14418 ;
  assign \g42479/_0_  = n14423 ;
  assign \g42480/_0_  = n14428 ;
  assign \g42481/_0_  = n14433 ;
  assign \g42482/_0_  = n14438 ;
  assign \g42483/_0_  = n14443 ;
  assign \g42484/_0_  = n14448 ;
  assign \g42485/_0_  = n14453 ;
  assign \g42486/_0_  = n14458 ;
  assign \g42487/_0_  = ~n14464 ;
  assign \g42488/_0_  = n14471 ;
  assign \g42490/_0_  = ~n14473 ;
  assign \g42491/_0_  = ~n14475 ;
  assign \g42493/_0_  = ~n14477 ;
  assign \g42494/_0_  = ~n14479 ;
  assign \g42495/_0_  = ~n14481 ;
  assign \g42496/_0_  = ~n14483 ;
  assign \g42497/_0_  = ~n14485 ;
  assign \g42498/_0_  = ~n14487 ;
  assign \g42499/_0_  = ~n14489 ;
  assign \g42500/_0_  = ~n14491 ;
  assign \g42501/_0_  = ~n14493 ;
  assign \g42502/_0_  = ~n14495 ;
  assign \g42503/_0_  = ~n14497 ;
  assign \g42504/_0_  = ~n14499 ;
  assign \g42505/_0_  = ~n14501 ;
  assign \g42506/_0_  = ~n14503 ;
  assign \g42507/_0_  = ~n14505 ;
  assign \g42508/_0_  = ~n14507 ;
  assign \g42509/_0_  = ~n14509 ;
  assign \g42510/_0_  = ~n14511 ;
  assign \g42511/_0_  = ~n14513 ;
  assign \g42512/_0_  = ~n14515 ;
  assign \g42513/_0_  = ~n14517 ;
  assign \g42514/_0_  = ~n14519 ;
  assign \g42515/_0_  = ~n14521 ;
  assign \g42516/_0_  = ~n14523 ;
  assign \g42517/_0_  = ~n14525 ;
  assign \g42518/_0_  = ~n14527 ;
  assign \g42519/_0_  = ~n14529 ;
  assign \g42521/_0_  = n14534 ;
  assign \g42522/_0_  = n14540 ;
  assign \g42523/_0_  = n14545 ;
  assign \g42524/_0_  = n14550 ;
  assign \g42525/_0_  = n14555 ;
  assign \g42526/_0_  = n14560 ;
  assign \g42527/_0_  = n14565 ;
  assign \g42528/_0_  = n14570 ;
  assign \g42529/_0_  = n14575 ;
  assign \g42530/_0_  = n14580 ;
  assign \g42531/_0_  = n14585 ;
  assign \g42532/_0_  = n14590 ;
  assign \g42533/_0_  = n14595 ;
  assign \g42534/_0_  = n14600 ;
  assign \g42535/_0_  = n14604 ;
  assign \g42536/_0_  = n14609 ;
  assign \g42537/_0_  = n14614 ;
  assign \g42538/_0_  = n14619 ;
  assign \g42539/_0_  = n14624 ;
  assign \g42540/_0_  = n14629 ;
  assign \g42541/_0_  = n14634 ;
  assign \g42542/_0_  = n14639 ;
  assign \g42543/_0_  = n14644 ;
  assign \g42544/_0_  = n14649 ;
  assign \g42545/_0_  = n14654 ;
  assign \g42548/_0_  = ~n14656 ;
  assign \g42557/_0_  = ~n14693 ;
  assign \g42564/_0_  = ~n14695 ;
  assign \g42565/_0_  = n14700 ;
  assign \g42566/_0_  = n14704 ;
  assign \g42567/_0_  = n14708 ;
  assign \g42568/_0_  = n14712 ;
  assign \g42569/_0_  = n14716 ;
  assign \g42570/_0_  = n14720 ;
  assign \g42571/_0_  = n14724 ;
  assign \g42572/_0_  = n14728 ;
  assign \g42573/_0_  = n14732 ;
  assign \g42574/_0_  = n14736 ;
  assign \g42575/_0_  = n14740 ;
  assign \g42576/_0_  = n14744 ;
  assign \g42577/_0_  = ~n14750 ;
  assign \g42578/_0_  = n14754 ;
  assign \g42581/_0_  = ~n14791 ;
  assign \g42589/_0_  = ~n14793 ;
  assign \g42590/_0_  = ~n14795 ;
  assign \g42591/_0_  = ~n14797 ;
  assign \g42592/_0_  = ~n14799 ;
  assign \g42593/_0_  = ~n14801 ;
  assign \g42594/_0_  = ~n14803 ;
  assign \g42595/_0_  = ~n14805 ;
  assign \g42596/_0_  = ~n14807 ;
  assign \g42597/_0_  = ~n14809 ;
  assign \g42598/_0_  = ~n14811 ;
  assign \g42599/_0_  = ~n14813 ;
  assign \g42600/_0_  = ~n14815 ;
  assign \g42601/_0_  = ~n14817 ;
  assign \g42602/_0_  = ~n14819 ;
  assign \g42603/_0_  = ~n14821 ;
  assign \g42604/_0_  = ~n14823 ;
  assign \g42605/_0_  = ~n14825 ;
  assign \g42606/_0_  = ~n14827 ;
  assign \g42607/_0_  = ~n14829 ;
  assign \g42608/_0_  = ~n14831 ;
  assign \g42609/_0_  = ~n14833 ;
  assign \g42610/_0_  = ~n14835 ;
  assign \g42611/_0_  = ~n14837 ;
  assign \g42612/_0_  = ~n14839 ;
  assign \g42613/_0_  = ~n14841 ;
  assign \g42614/_0_  = ~n14843 ;
  assign \g42615/_0_  = ~n14845 ;
  assign \g42616/_0_  = ~n14847 ;
  assign \g42617/_0_  = ~n14849 ;
  assign \g42618/_0_  = ~n14851 ;
  assign \g42619/_0_  = ~n14853 ;
  assign \g42620/_0_  = ~n14855 ;
  assign \g42622/_0_  = ~n14892 ;
  assign \g42623/_0_  = n14895 ;
  assign \g42627/_0_  = n14900 ;
  assign \g42628/_0_  = n14904 ;
  assign \g42629/_0_  = n14908 ;
  assign \g42630/_0_  = n14912 ;
  assign \g42631/_0_  = n14916 ;
  assign \g42632/_0_  = n14920 ;
  assign \g42633/_0_  = n14924 ;
  assign \g42634/_0_  = n14928 ;
  assign \g42635/_0_  = n14932 ;
  assign \g42636/_0_  = n14936 ;
  assign \g42637/_0_  = n14940 ;
  assign \g42638/_0_  = n14944 ;
  assign \g42639/_0_  = n14948 ;
  assign \g42640/_0_  = n14952 ;
  assign \g42641/_0_  = n14956 ;
  assign \g42642/_0_  = n14960 ;
  assign \g42643/_0_  = n14964 ;
  assign \g42644/_0_  = n14968 ;
  assign \g42645/_0_  = n14972 ;
  assign \g42646/_0_  = n14976 ;
  assign \g42647/_0_  = n14980 ;
  assign \g42648/_0_  = n14984 ;
  assign \g42649/_0_  = n14988 ;
  assign \g42650/_0_  = n14992 ;
  assign \g42666/_0_  = ~n14994 ;
  assign \g42667/_0_  = n14999 ;
  assign \g42668/_0_  = n15003 ;
  assign \g42669/_0_  = n15007 ;
  assign \g42670/_0_  = n15011 ;
  assign \g42671/_0_  = n15015 ;
  assign \g42672/_0_  = n15019 ;
  assign \g42673/_0_  = n15023 ;
  assign \g42674/_0_  = n15027 ;
  assign \g42675/_0_  = n15031 ;
  assign \g42676/_0_  = n15035 ;
  assign \g42677/_0_  = n15039 ;
  assign \g42678/_0_  = n15043 ;
  assign \g42680/_0_  = ~n15049 ;
  assign \g42681/_0_  = n15053 ;
  assign \g42685/_0_  = ~n15055 ;
  assign \g42686/_0_  = ~n15057 ;
  assign \g42688/_0_  = ~n15059 ;
  assign \g42689/_0_  = ~n15061 ;
  assign \g42690/_0_  = ~n15063 ;
  assign \g42691/_0_  = ~n15065 ;
  assign \g42692/_0_  = ~n15067 ;
  assign \g42693/_0_  = ~n15069 ;
  assign \g42694/_0_  = ~n15071 ;
  assign \g42695/_0_  = ~n15073 ;
  assign \g42696/_0_  = ~n15075 ;
  assign \g42697/_0_  = ~n15077 ;
  assign \g42698/_0_  = ~n15079 ;
  assign \g42699/_0_  = ~n15081 ;
  assign \g42700/_0_  = ~n15083 ;
  assign \g42701/_0_  = ~n15085 ;
  assign \g42702/_0_  = ~n15087 ;
  assign \g42703/_0_  = ~n15089 ;
  assign \g42704/_0_  = ~n15091 ;
  assign \g42705/_0_  = ~n15093 ;
  assign \g42706/_0_  = ~n15095 ;
  assign \g42707/_0_  = ~n15097 ;
  assign \g42708/_0_  = ~n15099 ;
  assign \g42709/_0_  = ~n15101 ;
  assign \g42710/_0_  = ~n15103 ;
  assign \g42711/_0_  = ~n15105 ;
  assign \g42712/_0_  = ~n15107 ;
  assign \g42713/_0_  = ~n15109 ;
  assign \g42715/_0_  = ~n15111 ;
  assign \g42716/_0_  = ~n15113 ;
  assign \g42717/_0_  = ~n15115 ;
  assign \g42718/_0_  = ~n15117 ;
  assign \g42723/_1_  = ~n15118 ;
  assign \g42727/_0_  = n15123 ;
  assign \g42728/_0_  = n15127 ;
  assign \g42729/_0_  = n15131 ;
  assign \g42730/_0_  = n15135 ;
  assign \g42731/_0_  = n15139 ;
  assign \g42732/_0_  = n15143 ;
  assign \g42733/_0_  = n15147 ;
  assign \g42734/_0_  = n15151 ;
  assign \g42735/_0_  = n15155 ;
  assign \g42736/_0_  = n15159 ;
  assign \g42737/_0_  = n15163 ;
  assign \g42738/_0_  = n15167 ;
  assign \g42739/_0_  = n15171 ;
  assign \g42740/_0_  = n15175 ;
  assign \g42741/_0_  = n15179 ;
  assign \g42742/_0_  = n15183 ;
  assign \g42743/_0_  = n15187 ;
  assign \g42744/_0_  = n15191 ;
  assign \g42745/_0_  = n15195 ;
  assign \g42746/_0_  = n15199 ;
  assign \g42747/_0_  = n15203 ;
  assign \g42748/_0_  = n15207 ;
  assign \g42749/_0_  = n15211 ;
  assign \g42750/_0_  = n15215 ;
  assign \g42751/_0_  = n15219 ;
  assign \g42754/_0_  = n15224 ;
  assign \g42767/_0_  = n15228 ;
  assign \g42768/_0_  = n15244 ;
  assign \g42772/_0_  = n15249 ;
  assign \g42773/_0_  = n15253 ;
  assign \g42774/_0_  = n15257 ;
  assign \g42775/_0_  = n15261 ;
  assign \g42776/_0_  = n15265 ;
  assign \g42777/_0_  = n15269 ;
  assign \g42778/_0_  = n15273 ;
  assign \g42779/_0_  = n15277 ;
  assign \g42780/_0_  = n15281 ;
  assign \g42781/_0_  = n15285 ;
  assign \g42782/_0_  = n15289 ;
  assign \g42783/_0_  = n15293 ;
  assign \g42784/_0_  = ~n15299 ;
  assign \g42785/_0_  = n15303 ;
  assign \g42790/_0_  = ~n15305 ;
  assign \g42791/_0_  = ~n15307 ;
  assign \g42792/_0_  = ~n15309 ;
  assign \g42793/_0_  = ~n15311 ;
  assign \g42794/_0_  = ~n15313 ;
  assign \g42795/_0_  = ~n15315 ;
  assign \g42796/_0_  = ~n15317 ;
  assign \g42797/_0_  = ~n15319 ;
  assign \g42798/_0_  = ~n15321 ;
  assign \g42799/_0_  = ~n15323 ;
  assign \g42800/_0_  = ~n15325 ;
  assign \g42801/_0_  = ~n15327 ;
  assign \g42802/_0_  = ~n15329 ;
  assign \g42803/_0_  = ~n15331 ;
  assign \g42804/_0_  = ~n15333 ;
  assign \g42805/_0_  = ~n15335 ;
  assign \g42806/_0_  = ~n15337 ;
  assign \g42807/_0_  = ~n15339 ;
  assign \g42808/_0_  = ~n15341 ;
  assign \g42809/_0_  = ~n15343 ;
  assign \g42810/_0_  = ~n15345 ;
  assign \g42811/_0_  = ~n15347 ;
  assign \g42812/_0_  = ~n15349 ;
  assign \g42813/_0_  = ~n15351 ;
  assign \g42814/_0_  = ~n15353 ;
  assign \g42815/_0_  = ~n15355 ;
  assign \g42816/_0_  = ~n15357 ;
  assign \g42817/_0_  = ~n15359 ;
  assign \g42818/_0_  = ~n15361 ;
  assign \g42819/_0_  = ~n15363 ;
  assign \g42820/_0_  = ~n15365 ;
  assign \g42821/_0_  = ~n15367 ;
  assign \g42824/_0_  = n15371 ;
  assign \g42825/_0_  = n15375 ;
  assign \g42826/_0_  = n15379 ;
  assign \g42827/_0_  = n15383 ;
  assign \g42828/_0_  = n15387 ;
  assign \g42829/_0_  = n15391 ;
  assign \g42830/_0_  = n15395 ;
  assign \g42831/_0_  = n15399 ;
  assign \g42832/_0_  = n15403 ;
  assign \g42833/_0_  = n15407 ;
  assign \g42834/_0_  = n15411 ;
  assign \g42835/_0_  = n15415 ;
  assign \g42836/_0_  = n15419 ;
  assign \g42837/_0_  = n15423 ;
  assign \g42838/_0_  = n15427 ;
  assign \g42839/_0_  = n15431 ;
  assign \g42840/_0_  = n15435 ;
  assign \g42841/_0_  = n15439 ;
  assign \g42842/_0_  = n15443 ;
  assign \g42843/_0_  = n15447 ;
  assign \g42844/_0_  = n15451 ;
  assign \g42845/_0_  = n15455 ;
  assign \g42846/_0_  = n15459 ;
  assign \g42907/_0_  = n15471 ;
  assign \g42914/_0_  = n15479 ;
  assign \g42924/_0_  = n15482 ;
  assign \g42925/_0_  = n15485 ;
  assign \g42926/_0_  = n15488 ;
  assign \g42927/_0_  = ~n15497 ;
  assign \g42928/_0_  = ~n15510 ;
  assign \g42929/_0_  = ~n15517 ;
  assign \g42930/_0_  = ~n15568 ;
  assign \g42931/_0_  = ~n15575 ;
  assign \g42933/_0_  = n15584 ;
  assign \g42941/_0_  = ~n15591 ;
  assign \g42947/_0_  = ~n15598 ;
  assign \g42950/_0_  = ~n15603 ;
  assign \g42955/_0_  = ~n15608 ;
  assign \g42956/_0_  = ~n15613 ;
  assign \g42972/_3_  = ~n15616 ;
  assign \g42973/_3_  = ~n15619 ;
  assign \g42974/_3_  = ~n15622 ;
  assign \g43178/_0_  = ~n15628 ;
  assign \g43179/_0_  = n15636 ;
  assign \g43184/_0_  = ~n15667 ;
  assign \g43186/_0_  = ~n15698 ;
  assign \g43187/_0_  = ~n15737 ;
  assign \g43190/_0_  = ~n15743 ;
  assign \g43191/_0_  = ~n15748 ;
  assign \g43192/_0_  = ~n15753 ;
  assign \g43202/_0_  = ~n15792 ;
  assign \g43205/_0_  = ~n15797 ;
  assign \g43206/_0_  = ~n15801 ;
  assign \g43207/_0_  = ~n15806 ;
  assign \g43209/_2_  = ~n15840 ;
  assign \g43228/_0_  = ~n15844 ;
  assign \g43233/_0_  = ~n15848 ;
  assign \g43235/_0_  = ~n15853 ;
  assign \g43236/_0_  = ~n15857 ;
  assign \g43237/_0_  = ~n15861 ;
  assign \g43238/_0_  = ~n15865 ;
  assign \g43280/_0_  = ~n15875 ;
  assign \g43287/_0_  = ~n15879 ;
  assign \g43289/_0_  = ~n15884 ;
  assign \g43290/_0_  = ~n15888 ;
  assign \g43291/_0_  = ~n15892 ;
  assign \g43292/_0_  = ~n15896 ;
  assign \g43303/_0_  = ~n15898 ;
  assign \g43311/_0_  = n15906 ;
  assign \g43312/_0_  = n15909 ;
  assign \g43363/_0_  = ~n15951 ;
  assign \g43364/_0_  = ~n15993 ;
  assign \g43366/_0_  = ~n16035 ;
  assign \g43367/_0_  = ~n16077 ;
  assign \g43370/_0_  = ~n16119 ;
  assign \g43371/_0_  = ~n16161 ;
  assign \g43374/_0_  = ~n16203 ;
  assign \g43413/_0_  = ~n16248 ;
  assign \g43414/_0_  = ~n16293 ;
  assign \g43415/_0_  = ~n16338 ;
  assign \g43416/_0_  = n16341 ;
  assign \g43422/_0_  = ~n16351 ;
  assign \g43427/_0_  = ~n16399 ;
  assign \g43428/_0_  = ~n16447 ;
  assign \g43528/_1__syn_2  = n10521 ;
  assign \g43630/_0_  = n16451 ;
  assign \g43633/_3_  = ~n16454 ;
  assign \g43647/_0_  = n16464 ;
  assign \g43648/_0_  = n16474 ;
  assign \g43656/_0_  = n16484 ;
  assign \g43657/_0_  = n16494 ;
  assign \g43667/_0_  = n16504 ;
  assign \g43668/_0_  = n16514 ;
  assign \g43675/_0_  = n16524 ;
  assign \g43678/_0_  = n16534 ;
  assign \g43787/_0_  = ~n16541 ;
  assign \g44055/_0_  = n16544 ;
  assign \g44092/_0_  = ~n16575 ;
  assign \g44093/_0_  = ~n16606 ;
  assign \g44176/_0_  = ~n16637 ;
  assign \g44181/_0_  = n16642 ;
  assign \g44433/_0_  = n16647 ;
  assign \g44510/_0_  = n16654 ;
  assign \g44515/_2_  = ~n16657 ;
  assign \g44522/_0_  = n16662 ;
  assign \g44529/_2_  = ~n16665 ;
  assign \g44537/_2_  = ~n16668 ;
  assign \g44544/_2_  = ~n16671 ;
  assign \g44594/_0_  = n16674 ;
  assign \g44695/_0_  = n16680 ;
  assign \g44697/_0_  = n16686 ;
  assign \g44699/_0_  = n16692 ;
  assign \g44700/_0_  = n16698 ;
  assign \g44843/_0_  = ~n16715 ;
  assign \g44844/_0_  = ~n16732 ;
  assign \g44879/_0_  = n16740 ;
  assign \g44880/_0_  = n16745 ;
  assign \g44881/_0_  = n16750 ;
  assign \g44882/_0_  = n16755 ;
  assign \g44906/_2_  = ~n16782 ;
  assign \g44910/_0_  = ~n16809 ;
  assign \g44912/_0_  = ~n16836 ;
  assign \g44954/_0_  = n16840 ;
  assign \g45000/_0_  = ~n16846 ;
  assign \g45001/_0_  = ~n16851 ;
  assign \g45002/_0_  = ~n16856 ;
  assign \g45003/_0_  = ~n16861 ;
  assign \g45021/_1_  = n7206 ;
  assign \g45025/_0_  = ~n16863 ;
  assign \g45051/_0_  = n16866 ;
  assign \g45104/_0_  = ~n16872 ;
  assign \g45111/_0_  = ~n16878 ;
  assign \g45112/_0_  = n16882 ;
  assign \g45116/_0_  = n16883 ;
  assign \g45155/_0_  = ~n5198 ;
  assign \g45238/_0_  = ~n16884 ;
  assign \g45239/_0_  = ~n16885 ;
  assign \g45240/_0_  = ~n16886 ;
  assign \g45241/_0_  = ~n16887 ;
  assign \g45249/_0_  = n16888 ;
  assign \g45257/_0_  = n16894 ;
  assign \g45332/_0_  = ~n16897 ;
  assign \g45334/_0_  = ~n16900 ;
  assign \g45336/_0_  = ~n16903 ;
  assign \g45337/_0_  = ~n16907 ;
  assign \g45342/_0_  = ~n16910 ;
  assign \g45459/_0_  = ~n16915 ;
  assign \g45460/_0_  = n16921 ;
  assign \g45466/_0_  = ~n16923 ;
  assign \g45469/_0_  = ~n16925 ;
  assign \g45470/_0_  = ~n16927 ;
  assign \g45474/_0_  = ~n16932 ;
  assign \g45475/_0_  = n16938 ;
  assign \g45477/_0_  = ~n16940 ;
  assign \g45481/_0_  = ~n16945 ;
  assign \g45482/_0_  = n16951 ;
  assign \g45487/_0_  = ~n16956 ;
  assign \g45488/_0_  = n16962 ;
  assign \g45518/_3_  = ~n16970 ;
  assign \g45519/_3_  = ~n16977 ;
  assign \g45520/_3_  = ~n16984 ;
  assign \g45521/_3_  = ~n16991 ;
  assign \g45522/_3_  = ~n16998 ;
  assign \g45523/_3_  = ~n17005 ;
  assign \g45524/_3_  = ~n17012 ;
  assign \g45525/_3_  = ~n17019 ;
  assign \g45526/_3_  = ~n17026 ;
  assign \g45530/_3_  = ~n17033 ;
  assign \g45531/_3_  = ~n17040 ;
  assign \g45532/_3_  = ~n17047 ;
  assign \g45533/_3_  = ~n17054 ;
  assign \g45534/_3_  = ~n17061 ;
  assign \g45535/_3_  = ~n17068 ;
  assign \g45536/_3_  = ~n17075 ;
  assign \g45559/_3_  = ~n17082 ;
  assign \g45596/_0_  = n17088 ;
  assign \g45605/_0_  = n17093 ;
  assign \g45622/_0_  = n17105 ;
  assign \g45623/_0_  = n17117 ;
  assign \g45630/_0_  = n17123 ;
  assign \g45747/_0_  = n17124 ;
  assign \g45753/_0_  = n17125 ;
  assign \g45796/_0_  = ~n17130 ;
  assign \g45837/_0_  = ~n17149 ;
  assign \g45882/_0_  = ~n17153 ;
  assign \g45903/_0_  = n17154 ;
  assign \g45912/_0_  = n16731 ;
  assign \g45946/_0_  = n16714 ;
  assign \g45999/_0_  = ~n17157 ;
  assign \g46000/_0_  = ~n17160 ;
  assign \g46001/_0_  = ~n17163 ;
  assign \g46002/_0_  = ~n17165 ;
  assign \g46012/_0_  = ~n17167 ;
  assign \g46014/_0_  = ~n17169 ;
  assign \g46017/_0_  = ~n17172 ;
  assign \g46018/_0_  = ~n17174 ;
  assign \g46021/_0_  = ~n17176 ;
  assign \g46024/_0_  = ~n17178 ;
  assign \g46026/_0_  = ~n17180 ;
  assign \g46029/_0_  = ~n17182 ;
  assign \g46053/_0_  = n17185 ;
  assign \g46083/_0_  = n17189 ;
  assign \g46093/_0_  = n17152 ;
  assign \g46142/_0_  = n17193 ;
  assign \g46154/_1__syn_2  = n10624 ;
  assign \g46265/_0_  = ~n17205 ;
  assign \g46266/_0_  = ~n17216 ;
  assign \g46268/_0_  = ~n17228 ;
  assign \g46270/_0_  = ~n17239 ;
  assign \g46273/_0_  = ~n17251 ;
  assign \g46274/_0_  = ~n17262 ;
  assign \g46275/_0_  = ~n17274 ;
  assign \g46276/_0_  = ~n17285 ;
  assign \g46278/_0_  = n17291 ;
  assign \g46385/_0_  = n17296 ;
  assign \g46411/_0_  = n17302 ;
  assign \g46414/_0_  = n17305 ;
  assign \g46479/_0_  = n17307 ;
  assign \g46520/_0_  = n17309 ;
  assign \g46521/_0_  = n17311 ;
  assign \g46530/_0_  = n17313 ;
  assign \g46531/_0_  = n17318 ;
  assign \g46597/_0_  = n17319 ;
  assign \g46610/_0_  = ~n17323 ;
  assign \g46617/_0_  = ~n17327 ;
  assign \g46632/_0_  = ~n17331 ;
  assign \g46637/_0_  = ~n17335 ;
  assign \g46722/_0_  = n17338 ;
  assign \g46723/_0_  = n17341 ;
  assign \g46724/_0_  = n17344 ;
  assign \g46725/_0_  = n17347 ;
  assign \g46813/_0_  = n5140 ;
  assign \g46842/_0_  = n5171 ;
  assign \g46888/_0_  = n4936 ;
  assign \g46891/_0_  = n17350 ;
  assign \g46894/_0_  = ~n15631 ;
  assign \g46905/_0_  = n17353 ;
  assign \g46940/_0_  = n17354 ;
  assign \g46992/_0_  = n5155 ;
  assign \g46995/_0_  = n5193 ;
  assign \g47037/_3_  = n17356 ;
  assign \g47053/_0_  = n17357 ;
  assign \g47140/_0_  = ~n17372 ;
  assign \g47155/_3_  = ~n17375 ;
  assign \g47209/_0_  = n17378 ;
  assign \g47211/_0_  = n17381 ;
  assign \g47213/_0_  = n17384 ;
  assign \g47215/_0_  = n17387 ;
  assign \g47337/_0_  = n17388 ;
  assign \g47433/_0_  = n17389 ;
  assign \g47972/_0_  = n17391 ;
  assign \g47976/_0_  = n17392 ;
  assign \g48081/_0_  = ~n17393 ;
  assign \g48171/_0_  = n17394 ;
  assign \g48227/_0_  = n17395 ;
  assign \g48234/_1_  = n3447 ;
  assign \g48257/_1_  = n5016 ;
  assign \g48266/_0_  = n2355 ;
  assign \g48281/_0_  = n17396 ;
  assign \g48291/_1_  = n17397 ;
  assign \g48322/_0_  = ~n17398 ;
  assign \g48345/_0_  = n17400 ;
  assign \g48429/_0_  = n17401 ;
  assign \g48495/_1_  = n5759 ;
  assign \g48549/_0_  = n5767 ;
  assign \g48589/_0_  = n2352 ;
  assign \g48642/_0_  = n5765 ;
  assign \g48722/_0_  = ~n17402 ;
  assign \g48748/_0_  = ~n17403 ;
  assign \g48749/_0_  = ~n17404 ;
  assign \g48763/_0_  = ~n17405 ;
  assign \g48867/_0_  = n17407 ;
  assign \g48876/_0_  = n17409 ;
  assign \g48880/_0_  = n17411 ;
  assign \g49023/_0_  = ~n5748 ;
  assign \g49205/_0_  = n17412 ;
  assign \g49314/_0_  = n17413 ;
  assign \g49432/_0__syn_2  = n17414 ;
  assign \g49512/_0_  = n17415 ;
  assign \g49707/_0_  = n17416 ;
  assign \g49737/_0_  = n17417 ;
  assign \g49831/_0_  = n17418 ;
  assign \g49922/_1_  = n17419 ;
  assign \g50132/_0_  = ~n5753 ;
  assign \g51376/_0_  = ~\u4_u2_buf0_orig_reg[19]/P0001  ;
  assign \g51412/_0_  = ~\u4_u0_buf0_orig_reg[19]/P0001  ;
  assign \g51822/_0_  = ~\u4_u3_buf0_orig_reg[19]/P0001  ;
  assign \g52114/_0_  = ~\u4_u1_buf0_orig_reg[19]/P0001  ;
  assign \g52156/_0_  = ~\u0_u0_idle_cnt1_reg[0]/P0001  ;
  assign \g54427/_0_  = n3460 ;
  assign \g54557/_0_  = ~n17428 ;
  assign \g54561/_3_  = ~n5497 ;
  assign \g55079/_0_  = ~n17430 ;
  assign \sram_adr_o[0]_pad  = ~n17439 ;
  assign \sram_adr_o[10]_pad  = ~n17444 ;
  assign \sram_adr_o[11]_pad  = ~n17449 ;
  assign \sram_adr_o[12]_pad  = ~n17454 ;
  assign \sram_adr_o[13]_pad  = ~n17459 ;
  assign \sram_adr_o[14]_pad  = ~n17464 ;
  assign \sram_adr_o[1]_pad  = ~n17469 ;
  assign \sram_adr_o[2]_pad  = ~n17474 ;
  assign \sram_adr_o[3]_pad  = ~n17479 ;
  assign \sram_adr_o[4]_pad  = ~n17484 ;
  assign \sram_adr_o[5]_pad  = ~n17489 ;
  assign \sram_adr_o[6]_pad  = ~n17494 ;
  assign \sram_adr_o[7]_pad  = ~n17499 ;
  assign \sram_adr_o[8]_pad  = ~n17504 ;
  assign \sram_adr_o[9]_pad  = ~n17509 ;
  assign \sram_data_o[0]_pad  = ~n17514 ;
  assign \sram_data_o[10]_pad  = ~n17519 ;
  assign \sram_data_o[11]_pad  = ~n17524 ;
  assign \sram_data_o[12]_pad  = ~n17529 ;
  assign \sram_data_o[13]_pad  = ~n17534 ;
  assign \sram_data_o[14]_pad  = ~n17539 ;
  assign \sram_data_o[15]_pad  = ~n17544 ;
  assign \sram_data_o[16]_pad  = ~n17549 ;
  assign \sram_data_o[17]_pad  = ~n17554 ;
  assign \sram_data_o[18]_pad  = ~n17559 ;
  assign \sram_data_o[19]_pad  = ~n17564 ;
  assign \sram_data_o[1]_pad  = ~n17569 ;
  assign \sram_data_o[20]_pad  = ~n17574 ;
  assign \sram_data_o[21]_pad  = ~n17579 ;
  assign \sram_data_o[22]_pad  = ~n17584 ;
  assign \sram_data_o[23]_pad  = ~n17589 ;
  assign \sram_data_o[24]_pad  = ~n17594 ;
  assign \sram_data_o[25]_pad  = ~n17599 ;
  assign \sram_data_o[26]_pad  = ~n17604 ;
  assign \sram_data_o[27]_pad  = ~n17609 ;
  assign \sram_data_o[28]_pad  = ~n17614 ;
  assign \sram_data_o[29]_pad  = ~n17619 ;
  assign \sram_data_o[2]_pad  = ~n17624 ;
  assign \sram_data_o[30]_pad  = ~n17629 ;
  assign \sram_data_o[31]_pad  = ~n17634 ;
  assign \sram_data_o[3]_pad  = ~n17639 ;
  assign \sram_data_o[4]_pad  = ~n17644 ;
  assign \sram_data_o[5]_pad  = ~n17649 ;
  assign \sram_data_o[6]_pad  = ~n17654 ;
  assign \sram_data_o[7]_pad  = ~n17659 ;
  assign \sram_data_o[8]_pad  = ~n17664 ;
  assign \sram_data_o[9]_pad  = ~n17669 ;
  assign sram_re_o_pad = ~1'b0 ;
  assign sram_we_o_pad = ~n17678 ;
  assign \u4_utmi_vend_ctrl_r_reg[0]/P0001_reg_syn_3  = ~n17684 ;
  assign \u4_utmi_vend_ctrl_r_reg[1]/P0001_reg_syn_3  = ~n17688 ;
  assign \u4_utmi_vend_ctrl_r_reg[2]/P0001_reg_syn_3  = ~n17692 ;
  assign \u4_utmi_vend_ctrl_r_reg[3]/P0001_reg_syn_3  = ~n17697 ;
endmodule
