module top (\C_0_pad , \C_10_pad , \C_11_pad , \C_12_pad , \C_13_pad , \C_14_pad , \C_15_pad , \C_16_pad , \C_17_pad , \C_18_pad , \C_19_pad , \C_1_pad , \C_20_pad , \C_21_pad , \C_22_pad , \C_23_pad , \C_24_pad , \C_25_pad , \C_26_pad , \C_27_pad , \C_28_pad , \C_29_pad , \C_2_pad , \C_30_pad , \C_31_pad , \C_32_pad , \C_3_pad , \C_4_pad , \C_5_pad , \C_6_pad , \C_7_pad , \C_8_pad , \C_9_pad , \P_0_pad , \X_10_reg/NET0131 , \X_11_reg/NET0131 , \X_12_reg/NET0131 , \X_13_reg/NET0131 , \X_14_reg/NET0131 , \X_15_reg/NET0131 , \X_16_reg/NET0131 , \X_17_reg/NET0131 , \X_18_reg/NET0131 , \X_19_reg/NET0131 , \X_1_reg/NET0131 , \X_20_reg/NET0131 , \X_21_reg/NET0131 , \X_22_reg/NET0131 , \X_23_reg/NET0131 , \X_24_reg/NET0131 , \X_25_reg/NET0131 , \X_26_reg/NET0131 , \X_27_reg/NET0131 , \X_28_reg/NET0131 , \X_29_reg/NET0131 , \X_2_reg/NET0131 , \X_30_reg/P0002 , \X_31_reg/P0002 , \X_32_reg/P0002 , \X_3_reg/NET0131 , \X_4_reg/NET0131 , \X_5_reg/NET0131 , \X_6_reg/NET0131 , \X_7_reg/NET0131 , \X_8_reg/NET0131 , \X_9_reg/NET0131 , \X_30_reg/P0000 , \X_31_reg/P0000 , \X_32_reg/P0000 , Z_pad, \_al_n0 , \_al_n1 , \g1375/_1_ , \g1387/_0_ , \g1398/_0_ , \g1400/_0_ , \g1419/_0_ , \g1433/_0_ , \g1443/_0_ , \g1457/_0_ , \g1458/_0_ , \g1468/_0_ , \g1483/_0_ , \g1486/_0_ , \g1493/_0_ , \g1504/_0_ , \g1505/_0_ , \g1512/_0_ , \g1525/_0_ , \g1535/_0_ , \g1544/_0_ , \g1565/_0_ , \g1871/_0_ , \g1900/_0_ , \g1955/_0_ , \g1961/_0_ , \g1991/_0_ , \g2026/_0_ , \g2040/_0_ , \g2046/_0_ , \g2051/_1_ , \g2098/_0_ , \g21/_0_ , \g2101/_0_ );
	input \C_0_pad  ;
	input \C_10_pad  ;
	input \C_11_pad  ;
	input \C_12_pad  ;
	input \C_13_pad  ;
	input \C_14_pad  ;
	input \C_15_pad  ;
	input \C_16_pad  ;
	input \C_17_pad  ;
	input \C_18_pad  ;
	input \C_19_pad  ;
	input \C_1_pad  ;
	input \C_20_pad  ;
	input \C_21_pad  ;
	input \C_22_pad  ;
	input \C_23_pad  ;
	input \C_24_pad  ;
	input \C_25_pad  ;
	input \C_26_pad  ;
	input \C_27_pad  ;
	input \C_28_pad  ;
	input \C_29_pad  ;
	input \C_2_pad  ;
	input \C_30_pad  ;
	input \C_31_pad  ;
	input \C_32_pad  ;
	input \C_3_pad  ;
	input \C_4_pad  ;
	input \C_5_pad  ;
	input \C_6_pad  ;
	input \C_7_pad  ;
	input \C_8_pad  ;
	input \C_9_pad  ;
	input \P_0_pad  ;
	input \X_10_reg/NET0131  ;
	input \X_11_reg/NET0131  ;
	input \X_12_reg/NET0131  ;
	input \X_13_reg/NET0131  ;
	input \X_14_reg/NET0131  ;
	input \X_15_reg/NET0131  ;
	input \X_16_reg/NET0131  ;
	input \X_17_reg/NET0131  ;
	input \X_18_reg/NET0131  ;
	input \X_19_reg/NET0131  ;
	input \X_1_reg/NET0131  ;
	input \X_20_reg/NET0131  ;
	input \X_21_reg/NET0131  ;
	input \X_22_reg/NET0131  ;
	input \X_23_reg/NET0131  ;
	input \X_24_reg/NET0131  ;
	input \X_25_reg/NET0131  ;
	input \X_26_reg/NET0131  ;
	input \X_27_reg/NET0131  ;
	input \X_28_reg/NET0131  ;
	input \X_29_reg/NET0131  ;
	input \X_2_reg/NET0131  ;
	input \X_30_reg/P0002  ;
	input \X_31_reg/P0002  ;
	input \X_32_reg/P0002  ;
	input \X_3_reg/NET0131  ;
	input \X_4_reg/NET0131  ;
	input \X_5_reg/NET0131  ;
	input \X_6_reg/NET0131  ;
	input \X_7_reg/NET0131  ;
	input \X_8_reg/NET0131  ;
	input \X_9_reg/NET0131  ;
	output \X_30_reg/P0000  ;
	output \X_31_reg/P0000  ;
	output \X_32_reg/P0000  ;
	output Z_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1375/_1_  ;
	output \g1387/_0_  ;
	output \g1398/_0_  ;
	output \g1400/_0_  ;
	output \g1419/_0_  ;
	output \g1433/_0_  ;
	output \g1443/_0_  ;
	output \g1457/_0_  ;
	output \g1458/_0_  ;
	output \g1468/_0_  ;
	output \g1483/_0_  ;
	output \g1486/_0_  ;
	output \g1493/_0_  ;
	output \g1504/_0_  ;
	output \g1505/_0_  ;
	output \g1512/_0_  ;
	output \g1525/_0_  ;
	output \g1535/_0_  ;
	output \g1544/_0_  ;
	output \g1565/_0_  ;
	output \g1871/_0_  ;
	output \g1900/_0_  ;
	output \g1955/_0_  ;
	output \g1961/_0_  ;
	output \g1991/_0_  ;
	output \g2026/_0_  ;
	output \g2040/_0_  ;
	output \g2046/_0_  ;
	output \g2051/_1_  ;
	output \g2098/_0_  ;
	output \g21/_0_  ;
	output \g2101/_0_  ;
	wire _w324_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\X_10_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\X_11_reg/NET0131 ,
		\X_12_reg/NET0131 ,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\X_3_reg/NET0131 ,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\X_4_reg/NET0131 ,
		\X_5_reg/NET0131 ,
		_w73_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		\X_6_reg/NET0131 ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w72_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w71_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\C_14_pad ,
		\X_14_reg/NET0131 ,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\C_16_pad ,
		\X_14_reg/NET0131 ,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		\X_15_reg/NET0131 ,
		\X_16_reg/NET0131 ,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w77_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		\X_13_reg/NET0131 ,
		_w69_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w81_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		_w76_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\X_4_reg/NET0131 ,
		_w71_,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\C_5_pad ,
		\X_5_reg/NET0131 ,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w85_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\X_13_reg/NET0131 ,
		\X_14_reg/NET0131 ,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\X_15_reg/NET0131 ,
		\X_16_reg/NET0131 ,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w88_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\X_17_reg/NET0131 ,
		\X_18_reg/NET0131 ,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\X_19_reg/NET0131 ,
		\X_1_reg/NET0131 ,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\X_20_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		\X_3_reg/NET0131 ,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w91_,
		_w92_,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w69_,
		_w90_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w75_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		\C_21_pad ,
		\X_21_reg/NET0131 ,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\C_22_pad ,
		\X_22_reg/NET0131 ,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		\C_23_pad ,
		\X_22_reg/NET0131 ,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		\X_23_reg/NET0131 ,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\X_21_reg/NET0131 ,
		_w101_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		_w103_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w100_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w99_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\C_0_pad ,
		_w87_,
		_w108_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w84_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w107_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\P_0_pad ,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\C_17_pad ,
		\X_17_reg/NET0131 ,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\C_19_pad ,
		\X_19_reg/NET0131 ,
		_w113_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		\C_20_pad ,
		\X_19_reg/NET0131 ,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\X_20_reg/NET0131 ,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w113_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		_w91_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w112_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		_w90_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\C_13_pad ,
		\X_13_reg/NET0131 ,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\C_15_pad ,
		\X_15_reg/NET0131 ,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w88_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\C_18_pad ,
		\X_17_reg/NET0131 ,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\X_18_reg/NET0131 ,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w90_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w120_,
		_w122_,
		_w126_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w119_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\P_0_pad ,
		_w76_,
		_w129_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w69_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w128_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\C_11_pad ,
		\X_11_reg/NET0131 ,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\C_12_pad ,
		\X_11_reg/NET0131 ,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\X_12_reg/NET0131 ,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w132_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		_w67_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\C_9_pad ,
		\X_9_reg/NET0131 ,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\C_10_pad ,
		\X_10_reg/NET0131 ,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		\X_9_reg/NET0131 ,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w137_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		_w136_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		_w129_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\C_2_pad ,
		\X_2_reg/NET0131 ,
		_w144_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		\C_4_pad ,
		\X_2_reg/NET0131 ,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\X_3_reg/NET0131 ,
		\X_4_reg/NET0131 ,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w144_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		_w143_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\C_1_pad ,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\C_3_pad ,
		\X_2_reg/NET0131 ,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		\X_3_reg/NET0131 ,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w143_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		\C_6_pad ,
		\X_6_reg/NET0131 ,
		_w155_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\C_8_pad ,
		\X_7_reg/NET0131 ,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\X_8_reg/NET0131 ,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\C_7_pad ,
		\X_7_reg/NET0131 ,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\X_6_reg/NET0131 ,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w157_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		\P_0_pad ,
		\X_5_reg/NET0131 ,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w155_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w85_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w160_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		\X_21_reg/NET0131 ,
		\X_22_reg/NET0131 ,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w99_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\C_24_pad ,
		\P_0_pad ,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		\X_23_reg/NET0131 ,
		\X_24_reg/NET0131 ,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w167_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w166_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		\C_25_pad ,
		\X_25_reg/NET0131 ,
		_w171_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		\C_26_pad ,
		\X_26_reg/NET0131 ,
		_w172_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		\C_28_pad ,
		\X_27_reg/NET0131 ,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\X_28_reg/NET0131 ,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\C_27_pad ,
		\X_27_reg/NET0131 ,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\X_26_reg/NET0131 ,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w174_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\X_25_reg/NET0131 ,
		_w172_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w171_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		\P_0_pad ,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\C_30_pad ,
		\X_30_reg/P0002 ,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		\C_31_pad ,
		\X_31_reg/P0002 ,
		_w183_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\C_32_pad ,
		\X_31_reg/P0002 ,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\X_32_reg/P0002 ,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w183_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		\X_30_reg/P0002 ,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\X_29_reg/NET0131 ,
		_w182_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		_w187_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		\C_29_pad ,
		\X_29_reg/NET0131 ,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		\P_0_pad ,
		\X_25_reg/NET0131 ,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\X_26_reg/NET0131 ,
		\X_27_reg/NET0131 ,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		\X_28_reg/NET0131 ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		_w190_,
		_w191_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w193_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w189_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w181_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\X_23_reg/NET0131 ,
		\X_24_reg/NET0131 ,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w166_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		_w197_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w151_,
		_w154_,
		_w201_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w149_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w164_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		_w142_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		_w170_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		_w111_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		_w131_,
		_w200_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		\X_10_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w209_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\X_11_reg/NET0131 ,
		\X_12_reg/NET0131 ,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w212_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		_w211_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		\X_14_reg/NET0131 ,
		\X_15_reg/NET0131 ,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		\X_16_reg/NET0131 ,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\X_17_reg/NET0131 ,
		\X_18_reg/NET0131 ,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\X_19_reg/NET0131 ,
		\X_1_reg/NET0131 ,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		\X_20_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\X_4_reg/NET0131 ,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		_w218_,
		_w219_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w221_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		_w217_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w215_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\P_0_pad ,
		\X_13_reg/NET0131 ,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\X_2_reg/NET0131 ,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\X_21_reg/NET0131 ,
		\X_22_reg/NET0131 ,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		\X_23_reg/NET0131 ,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\X_24_reg/NET0131 ,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\X_25_reg/NET0131 ,
		_w227_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w230_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		_w225_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		\X_26_reg/NET0131 ,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\X_27_reg/NET0131 ,
		\X_28_reg/NET0131 ,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w234_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\X_29_reg/NET0131 ,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		\X_30_reg/P0002 ,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\X_31_reg/P0002 ,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		\X_26_reg/NET0131 ,
		_w233_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w234_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w225_,
		_w227_,
		_w242_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		\X_21_reg/NET0131 ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\X_22_reg/NET0131 ,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w228_,
		_w242_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w244_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		\X_27_reg/NET0131 ,
		_w234_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		\X_27_reg/NET0131 ,
		_w234_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w247_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\X_23_reg/NET0131 ,
		_w245_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w229_,
		_w242_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\X_21_reg/NET0131 ,
		_w242_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w243_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		\X_2_reg/NET0131 ,
		_w150_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		\X_3_reg/NET0131 ,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\X_4_reg/NET0131 ,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		_w215_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\X_13_reg/NET0131 ,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w217_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w218_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\X_19_reg/NET0131 ,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		\X_19_reg/NET0131 ,
		_w261_,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w262_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\X_5_reg/NET0131 ,
		_w257_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		\X_6_reg/NET0131 ,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w211_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		\X_11_reg/NET0131 ,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\X_12_reg/NET0131 ,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w258_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		\X_17_reg/NET0131 ,
		_w260_,
		_w271_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		\X_17_reg/NET0131 ,
		_w260_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\X_14_reg/NET0131 ,
		_w259_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		\X_15_reg/NET0131 ,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		\X_15_reg/NET0131 ,
		_w274_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		\X_13_reg/NET0131 ,
		_w258_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w259_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		\X_6_reg/NET0131 ,
		_w265_,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w266_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\X_11_reg/NET0131 ,
		_w267_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w268_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		\X_4_reg/NET0131 ,
		_w256_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w257_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w209_,
		_w266_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\X_9_reg/NET0131 ,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		\X_9_reg/NET0131 ,
		_w286_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		_w287_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name223 (
		\X_7_reg/NET0131 ,
		_w266_,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		\X_7_reg/NET0131 ,
		_w266_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w290_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		\X_5_reg/NET0131 ,
		_w257_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w265_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		\X_3_reg/NET0131 ,
		_w255_,
		_w295_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w256_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		\X_2_reg/NET0131 ,
		_w150_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w255_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w143_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		\X_20_reg/NET0131 ,
		_w262_,
		_w301_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		\X_20_reg/NET0131 ,
		_w262_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w301_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		\X_14_reg/NET0131 ,
		_w259_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w274_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		\X_18_reg/NET0131 ,
		_w271_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w261_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\X_24_reg/NET0131 ,
		_w251_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w230_,
		_w242_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		\X_25_reg/NET0131 ,
		_w309_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		_w233_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		\X_29_reg/NET0131 ,
		_w236_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w237_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		_w72_,
		_w209_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		_w291_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		_w291_,
		_w315_,
		_w317_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w316_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		\X_28_reg/NET0131 ,
		_w247_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w236_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		\X_16_reg/NET0131 ,
		_w276_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w260_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		\X_10_reg/NET0131 ,
		_w287_,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w267_,
		_w323_,
		_w324_
	);
	assign \X_30_reg/P0000  = \X_30_reg/P0002 ;
	assign \X_31_reg/P0000  = \X_31_reg/P0002 ;
	assign \X_32_reg/P0000  = \X_32_reg/P0002 ;
	assign Z_pad = _w208_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1375/_1_  = _w239_ ;
	assign \g1387/_0_  = _w241_ ;
	assign \g1398/_0_  = _w246_ ;
	assign \g1400/_0_  = _w249_ ;
	assign \g1419/_0_  = _w252_ ;
	assign \g1433/_0_  = _w254_ ;
	assign \g1443/_0_  = _w264_ ;
	assign \g1457/_0_  = _w270_ ;
	assign \g1458/_0_  = _w273_ ;
	assign \g1468/_0_  = _w277_ ;
	assign \g1483/_0_  = _w279_ ;
	assign \g1486/_0_  = _w281_ ;
	assign \g1493/_0_  = _w283_ ;
	assign \g1504/_0_  = _w285_ ;
	assign \g1505/_0_  = _w289_ ;
	assign \g1512/_0_  = _w292_ ;
	assign \g1525/_0_  = _w294_ ;
	assign \g1535/_0_  = _w296_ ;
	assign \g1544/_0_  = _w298_ ;
	assign \g1565/_0_  = _w300_ ;
	assign \g1871/_0_  = _w303_ ;
	assign \g1900/_0_  = _w305_ ;
	assign \g1955/_0_  = _w307_ ;
	assign \g1961/_0_  = _w310_ ;
	assign \g1991/_0_  = _w312_ ;
	assign \g2026/_0_  = _w314_ ;
	assign \g2040/_0_  = _w318_ ;
	assign \g2046/_0_  = _w238_ ;
	assign \g2051/_1_  = _w237_ ;
	assign \g2098/_0_  = _w320_ ;
	assign \g21/_0_  = _w322_ ;
	assign \g2101/_0_  = _w324_ ;
endmodule;