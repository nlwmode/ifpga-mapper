module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G18_pad , \G1_pad , \G2_pad , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G4_pad , \G5_pad , \G6_pad , \G7_pad , \G8_pad , \G9_pad , \G288_pad , \G290_pad , \G296_pad , \G302_pad , \G315_pad , \G325_pad , \G327_pad , \G45_pad , \G47_pad , \G49_pad , \G53_pad , \G55_pad , \_al_n0 , \_al_n1 , \g1404/_0_ , \g1412/_0_ , \g1416/_0_ , \g1451/_2_ , \g1459/_3_ , \g1511/_3_ , \g1527/_3_ , \g1529/_3_ , \g31/_0_ , \g33/_1_ , \g56/_3_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G18_pad  ;
	input \G1_pad  ;
	input \G2_pad  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G6_pad  ;
	input \G7_pad  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G288_pad  ;
	output \G290_pad  ;
	output \G296_pad  ;
	output \G302_pad  ;
	output \G315_pad  ;
	output \G325_pad  ;
	output \G327_pad  ;
	output \G45_pad  ;
	output \G47_pad  ;
	output \G49_pad  ;
	output \G53_pad  ;
	output \G55_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1404/_0_  ;
	output \g1412/_0_  ;
	output \g1416/_0_  ;
	output \g1451/_2_  ;
	output \g1459/_3_  ;
	output \g1511/_3_  ;
	output \g1527/_3_  ;
	output \g1529/_3_  ;
	output \g31/_0_  ;
	output \g33/_1_  ;
	output \g56/_3_  ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w25_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w26_
	);
	LUT3 #(
		.INIT('h01)
	) name2 (
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w27_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w25_,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\G15_pad ,
		\G39_reg/NET0131 ,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w30_
	);
	LUT3 #(
		.INIT('h01)
	) name6 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w29_,
		_w31_,
		_w32_
	);
	LUT3 #(
		.INIT('h08)
	) name8 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w33_
	);
	LUT4 #(
		.INIT('h0040)
	) name9 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\G39_reg/NET0131 ,
		_w34_,
		_w35_
	);
	LUT4 #(
		.INIT('hccc4)
	) name11 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w37_
	);
	LUT3 #(
		.INIT('h15)
	) name13 (
		\G16_pad ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w38_
	);
	LUT4 #(
		.INIT('h0111)
	) name14 (
		\G16_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w39_
	);
	LUT4 #(
		.INIT('haa08)
	) name15 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w36_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\G16_pad ,
		\G4_pad ,
		_w41_
	);
	LUT3 #(
		.INIT('h80)
	) name17 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w42_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name18 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w43_
	);
	LUT3 #(
		.INIT('h15)
	) name19 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w44_
	);
	LUT4 #(
		.INIT('h5444)
	) name20 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w45_
	);
	LUT3 #(
		.INIT('h10)
	) name21 (
		_w41_,
		_w43_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w47_
	);
	LUT4 #(
		.INIT('h0001)
	) name23 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\G16_pad ,
		\G38_reg/NET0131 ,
		_w49_
	);
	LUT3 #(
		.INIT('h02)
	) name25 (
		\G16_pad ,
		\G1_pad ,
		\G38_reg/NET0131 ,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w48_,
		_w50_,
		_w51_
	);
	LUT3 #(
		.INIT('hfe)
	) name27 (
		_w46_,
		_w40_,
		_w51_,
		_w52_
	);
	LUT4 #(
		.INIT('h8000)
	) name28 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w53_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name29 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\G38_reg/NET0131 ,
		_w54_,
		_w55_
	);
	LUT3 #(
		.INIT('h80)
	) name31 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w26_,
		_w56_,
		_w57_
	);
	LUT3 #(
		.INIT('h80)
	) name33 (
		\G15_pad ,
		\G39_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w30_,
		_w58_,
		_w59_
	);
	LUT3 #(
		.INIT('h08)
	) name35 (
		\G15_pad ,
		\G16_pad ,
		\G38_reg/NET0131 ,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w61_
	);
	LUT4 #(
		.INIT('h000e)
	) name37 (
		\G10_pad ,
		\G11_pad ,
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w62_
	);
	LUT3 #(
		.INIT('h07)
	) name38 (
		\G10_pad ,
		\G11_pad ,
		\G12_pad ,
		_w63_
	);
	LUT4 #(
		.INIT('h2000)
	) name39 (
		_w33_,
		_w63_,
		_w60_,
		_w62_,
		_w64_
	);
	LUT3 #(
		.INIT('h40)
	) name40 (
		\G5_pad ,
		_w25_,
		_w27_,
		_w65_
	);
	LUT4 #(
		.INIT('h01ab)
	) name41 (
		\G39_reg/NET0131 ,
		_w43_,
		_w44_,
		_w36_,
		_w66_
	);
	LUT3 #(
		.INIT('h04)
	) name42 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT3 #(
		.INIT('h80)
	) name45 (
		\G5_pad ,
		_w25_,
		_w27_,
		_w70_
	);
	LUT3 #(
		.INIT('h80)
	) name46 (
		\G13_pad ,
		\G15_pad ,
		\G42_reg/NET0131 ,
		_w71_
	);
	LUT3 #(
		.INIT('hc4)
	) name47 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w72_
	);
	LUT4 #(
		.INIT('hf020)
	) name48 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w73_
	);
	LUT3 #(
		.INIT('h45)
	) name49 (
		\G39_reg/NET0131 ,
		_w71_,
		_w73_,
		_w74_
	);
	LUT4 #(
		.INIT('h8000)
	) name50 (
		\G6_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		_w77_
	);
	LUT3 #(
		.INIT('he0)
	) name53 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w78_
	);
	LUT4 #(
		.INIT('h1f00)
	) name54 (
		\G40_reg/NET0131 ,
		_w75_,
		_w76_,
		_w78_,
		_w79_
	);
	LUT3 #(
		.INIT('h01)
	) name55 (
		\G1_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w80_
	);
	LUT3 #(
		.INIT('h10)
	) name56 (
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w81_
	);
	LUT4 #(
		.INIT('h0800)
	) name57 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		\G6_pad ,
		_w82_
	);
	LUT4 #(
		.INIT('ha888)
	) name58 (
		_w68_,
		_w80_,
		_w81_,
		_w82_,
		_w83_
	);
	LUT3 #(
		.INIT('h45)
	) name59 (
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w84_
	);
	LUT4 #(
		.INIT('h070a)
	) name60 (
		\G15_pad ,
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w85_
	);
	LUT4 #(
		.INIT('h0100)
	) name61 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w86_
	);
	LUT3 #(
		.INIT('h0b)
	) name62 (
		_w84_,
		_w85_,
		_w86_,
		_w87_
	);
	LUT4 #(
		.INIT('h0b00)
	) name63 (
		_w74_,
		_w79_,
		_w83_,
		_w87_,
		_w88_
	);
	LUT3 #(
		.INIT('h23)
	) name64 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		\G5_pad ,
		_w89_
	);
	LUT4 #(
		.INIT('h0100)
	) name65 (
		\G1_pad ,
		\G3_pad ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w90_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name66 (
		\G2_pad ,
		_w25_,
		_w89_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		\G15_pad ,
		\G39_reg/NET0131 ,
		_w92_
	);
	LUT3 #(
		.INIT('h08)
	) name68 (
		\G14_pad ,
		\G15_pad ,
		\G39_reg/NET0131 ,
		_w93_
	);
	LUT4 #(
		.INIT('hea00)
	) name69 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		\G4_pad ,
		_w94_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name70 (
		\G39_reg/NET0131 ,
		_w67_,
		_w93_,
		_w94_,
		_w95_
	);
	LUT3 #(
		.INIT('h45)
	) name71 (
		\G38_reg/NET0131 ,
		_w91_,
		_w95_,
		_w96_
	);
	LUT3 #(
		.INIT('h08)
	) name72 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w36_,
		_w97_
	);
	LUT4 #(
		.INIT('h4c40)
	) name73 (
		\G0_pad ,
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w42_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w97_,
		_w99_,
		_w100_
	);
	LUT4 #(
		.INIT('h0d00)
	) name76 (
		\G16_pad ,
		_w88_,
		_w96_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\G18_pad ,
		_w101_,
		_w102_
	);
	LUT3 #(
		.INIT('h01)
	) name78 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		\G4_pad ,
		_w103_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name79 (
		\G0_pad ,
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w103_,
		_w104_,
		_w105_
	);
	LUT4 #(
		.INIT('hccc8)
	) name81 (
		\G38_reg/NET0131 ,
		_w25_,
		_w89_,
		_w90_,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		_w108_
	);
	LUT3 #(
		.INIT('h2a)
	) name84 (
		\G16_pad ,
		_w75_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w110_
	);
	LUT3 #(
		.INIT('h02)
	) name86 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G4_pad ,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w37_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w109_,
		_w112_,
		_w113_
	);
	LUT3 #(
		.INIT('h02)
	) name89 (
		\G16_pad ,
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w114_
	);
	LUT3 #(
		.INIT('h10)
	) name90 (
		_w44_,
		_w77_,
		_w114_,
		_w115_
	);
	LUT3 #(
		.INIT('h0e)
	) name91 (
		\G10_pad ,
		\G11_pad ,
		\G42_reg/NET0131 ,
		_w116_
	);
	LUT3 #(
		.INIT('h80)
	) name92 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w117_
	);
	LUT3 #(
		.INIT('h45)
	) name93 (
		_w43_,
		_w116_,
		_w117_,
		_w118_
	);
	LUT4 #(
		.INIT('h0010)
	) name94 (
		\G16_pad ,
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		\G41_reg/NET0131 ,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w121_
	);
	LUT3 #(
		.INIT('hb0)
	) name97 (
		\G14_pad ,
		\G15_pad ,
		\G41_reg/NET0131 ,
		_w122_
	);
	LUT3 #(
		.INIT('h08)
	) name98 (
		_w68_,
		_w121_,
		_w122_,
		_w123_
	);
	LUT4 #(
		.INIT('h7077)
	) name99 (
		_w115_,
		_w118_,
		_w120_,
		_w123_,
		_w124_
	);
	LUT4 #(
		.INIT('h5455)
	) name100 (
		\G18_pad ,
		_w107_,
		_w113_,
		_w124_,
		_w125_
	);
	LUT4 #(
		.INIT('haa2a)
	) name101 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w126_
	);
	LUT4 #(
		.INIT('h62ea)
	) name102 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w126_,
		_w127_,
		_w128_
	);
	LUT3 #(
		.INIT('h13)
	) name104 (
		\G10_pad ,
		\G11_pad ,
		\G12_pad ,
		_w129_
	);
	LUT3 #(
		.INIT('h08)
	) name105 (
		_w34_,
		_w92_,
		_w129_,
		_w130_
	);
	LUT3 #(
		.INIT('ha8)
	) name106 (
		_w41_,
		_w128_,
		_w130_,
		_w131_
	);
	LUT3 #(
		.INIT('h01)
	) name107 (
		\G16_pad ,
		\G1_pad ,
		\G38_reg/NET0131 ,
		_w132_
	);
	LUT4 #(
		.INIT('h5f01)
	) name108 (
		\G16_pad ,
		\G1_pad ,
		\G38_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w133_
	);
	LUT3 #(
		.INIT('h08)
	) name109 (
		\G0_pad ,
		\G38_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w134_
	);
	LUT3 #(
		.INIT('h01)
	) name110 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w135_
	);
	LUT3 #(
		.INIT('h10)
	) name111 (
		_w134_,
		_w133_,
		_w135_,
		_w136_
	);
	LUT3 #(
		.INIT('h40)
	) name112 (
		\G0_pad ,
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w137_
	);
	LUT3 #(
		.INIT('h08)
	) name113 (
		\G1_pad ,
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w138_
	);
	LUT4 #(
		.INIT('hc400)
	) name114 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w139_
	);
	LUT3 #(
		.INIT('he0)
	) name115 (
		_w137_,
		_w138_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w136_,
		_w140_,
		_w141_
	);
	LUT3 #(
		.INIT('h45)
	) name117 (
		\G18_pad ,
		_w131_,
		_w141_,
		_w142_
	);
	LUT3 #(
		.INIT('h7e)
	) name118 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w143_
	);
	LUT3 #(
		.INIT('h02)
	) name119 (
		\G1_pad ,
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w143_,
		_w144_,
		_w145_
	);
	LUT3 #(
		.INIT('h80)
	) name121 (
		\G3_pad ,
		_w48_,
		_w132_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w49_,
		_w53_,
		_w147_
	);
	LUT3 #(
		.INIT('h80)
	) name123 (
		\G15_pad ,
		_w67_,
		_w68_,
		_w148_
	);
	LUT3 #(
		.INIT('h40)
	) name124 (
		\G38_reg/NET0131 ,
		_w67_,
		_w93_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\G39_reg/NET0131 ,
		_w94_,
		_w150_
	);
	LUT4 #(
		.INIT('h0800)
	) name126 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w151_
	);
	LUT4 #(
		.INIT('hf3d1)
	) name127 (
		\G16_pad ,
		_w121_,
		_w122_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		\G41_reg/NET0131 ,
		\G4_pad ,
		_w153_
	);
	LUT4 #(
		.INIT('h5173)
	) name129 (
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G4_pad ,
		\G5_pad ,
		_w154_
	);
	LUT4 #(
		.INIT('h40cc)
	) name130 (
		\G16_pad ,
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w155_
	);
	LUT4 #(
		.INIT('h3efe)
	) name131 (
		\G16_pad ,
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w156_
	);
	LUT4 #(
		.INIT('h0004)
	) name132 (
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		\G41_reg/NET0131 ,
		_w157_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name133 (
		_w154_,
		_w155_,
		_w156_,
		_w157_,
		_w158_
	);
	LUT4 #(
		.INIT('h4055)
	) name134 (
		\G38_reg/NET0131 ,
		_w150_,
		_w152_,
		_w158_,
		_w159_
	);
	LUT3 #(
		.INIT('h0e)
	) name135 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w160_
	);
	LUT3 #(
		.INIT('h04)
	) name136 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		\G4_pad ,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		_w160_,
		_w161_,
		_w162_
	);
	LUT3 #(
		.INIT('h80)
	) name138 (
		\G13_pad ,
		\G15_pad ,
		\G16_pad ,
		_w163_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name139 (
		_w42_,
		_w61_,
		_w137_,
		_w163_,
		_w164_
	);
	LUT4 #(
		.INIT('h444c)
	) name140 (
		\G15_pad ,
		\G16_pad ,
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w165_
	);
	LUT3 #(
		.INIT('h08)
	) name141 (
		_w44_,
		_w110_,
		_w165_,
		_w166_
	);
	LUT4 #(
		.INIT('h0103)
	) name142 (
		_w109_,
		_w164_,
		_w166_,
		_w162_,
		_w167_
	);
	LUT3 #(
		.INIT('h45)
	) name143 (
		\G18_pad ,
		_w159_,
		_w167_,
		_w168_
	);
	LUT4 #(
		.INIT('h0006)
	) name144 (
		\G10_pad ,
		\G11_pad ,
		\G12_pad ,
		\G42_reg/NET0131 ,
		_w169_
	);
	LUT3 #(
		.INIT('h08)
	) name145 (
		\G15_pad ,
		\G16_pad ,
		\G39_reg/NET0131 ,
		_w170_
	);
	LUT4 #(
		.INIT('h0800)
	) name146 (
		_w72_,
		_w153_,
		_w169_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		_w38_,
		_w111_,
		_w172_
	);
	LUT3 #(
		.INIT('h80)
	) name148 (
		_w27_,
		_w47_,
		_w119_,
		_w173_
	);
	LUT3 #(
		.INIT('h01)
	) name149 (
		_w172_,
		_w171_,
		_w173_,
		_w174_
	);
	LUT3 #(
		.INIT('h45)
	) name150 (
		\G18_pad ,
		_w107_,
		_w174_,
		_w175_
	);
	assign \G288_pad  = _w28_ ;
	assign \G290_pad  = _w32_ ;
	assign \G296_pad  = _w35_ ;
	assign \G302_pad  = _w52_ ;
	assign \G315_pad  = _w55_ ;
	assign \G325_pad  = _w57_ ;
	assign \G327_pad  = _w59_ ;
	assign \G45_pad  = _w64_ ;
	assign \G47_pad  = _w65_ ;
	assign \G49_pad  = _w66_ ;
	assign \G53_pad  = _w69_ ;
	assign \G55_pad  = _w70_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1404/_0_  = _w102_ ;
	assign \g1412/_0_  = _w125_ ;
	assign \g1416/_0_  = _w142_ ;
	assign \g1451/_2_  = _w145_ ;
	assign \g1459/_3_  = _w146_ ;
	assign \g1511/_3_  = _w147_ ;
	assign \g1527/_3_  = _w148_ ;
	assign \g1529/_3_  = _w149_ ;
	assign \g31/_0_  = _w168_ ;
	assign \g33/_1_  = _w175_ ;
	assign \g56/_3_  = _w113_ ;
endmodule;