module top( \address_reg[0]/NET0131  , \address_reg[1]/NET0131  , \address_reg[2]/NET0131  , \address_reg[3]/NET0131  , \address_reg[4]/NET0131  , \count_reg[0]/NET0131  , \count_reg[0]1198/NET0131  , \count_reg[1]/NET0131  , \count_reg[1]1200/NET0131  , \count_reg[2]/NET0131  , \count_reg[3]/NET0131  , \count_reg[4]/NET0131  , \count_reg[5]/NET0131  , \counter_reg[0]/NET0131  , \counter_reg[1]/NET0131  , \counter_reg[2]/NET0131  , \data_in_reg[0]/NET0131  , \data_in_reg[1]/NET0131  , \data_out_reg[0]/NET0131  , \data_out_reg[1]/NET0131  , \gamma_reg[0]/NET0131  , \gamma_reg[1]/NET0131  , \gamma_reg[2]/NET0131  , \gamma_reg[3]/NET0131  , \gamma_reg[4]/NET0131  , \ind_reg[0]/NET0131  , \ind_reg[1]/NET0131  , \k[0]_pad  , \k[1]_pad  , \k[2]_pad  , \k[3]_pad  , \max_reg[0]/NET0131  , \max_reg[1]/NET0131  , \max_reg[2]/NET0131  , \max_reg[3]/NET0131  , \max_reg[4]/NET0131  , \memory_reg[0][0]/NET0131  , \memory_reg[0][1]/NET0131  , \memory_reg[10][0]/NET0131  , \memory_reg[10][1]/NET0131  , \memory_reg[11][0]/NET0131  , \memory_reg[11][1]/NET0131  , \memory_reg[12][0]/NET0131  , \memory_reg[12][1]/NET0131  , \memory_reg[13][0]/NET0131  , \memory_reg[13][1]/NET0131  , \memory_reg[14][0]/NET0131  , \memory_reg[14][1]/NET0131  , \memory_reg[15][0]/NET0131  , \memory_reg[15][1]/NET0131  , \memory_reg[16][0]/NET0131  , \memory_reg[16][1]/NET0131  , \memory_reg[17][0]/NET0131  , \memory_reg[17][1]/NET0131  , \memory_reg[18][0]/NET0131  , \memory_reg[18][1]/NET0131  , \memory_reg[19][0]/NET0131  , \memory_reg[19][1]/NET0131  , \memory_reg[1][0]/NET0131  , \memory_reg[1][1]/NET0131  , \memory_reg[20][0]/NET0131  , \memory_reg[20][1]/NET0131  , \memory_reg[21][0]/NET0131  , \memory_reg[21][1]/NET0131  , \memory_reg[22][0]/NET0131  , \memory_reg[22][1]/NET0131  , \memory_reg[23][0]/NET0131  , \memory_reg[23][1]/NET0131  , \memory_reg[24][0]/NET0131  , \memory_reg[24][1]/NET0131  , \memory_reg[25][0]/NET0131  , \memory_reg[25][1]/NET0131  , \memory_reg[26][0]/NET0131  , \memory_reg[26][1]/NET0131  , \memory_reg[27][0]/NET0131  , \memory_reg[27][1]/NET0131  , \memory_reg[28][0]/NET0131  , \memory_reg[28][1]/NET0131  , \memory_reg[29][0]/NET0131  , \memory_reg[29][1]/NET0131  , \memory_reg[2][0]/NET0131  , \memory_reg[2][1]/NET0131  , \memory_reg[30][0]/NET0131  , \memory_reg[30][1]/NET0131  , \memory_reg[31][0]/NET0131  , \memory_reg[31][1]/NET0131  , \memory_reg[3][0]/NET0131  , \memory_reg[3][1]/NET0131  , \memory_reg[4][0]/NET0131  , \memory_reg[4][1]/NET0131  , \memory_reg[5][0]/NET0131  , \memory_reg[5][1]/NET0131  , \memory_reg[6][0]/NET0131  , \memory_reg[6][1]/NET0131  , \memory_reg[7][0]/NET0131  , \memory_reg[7][1]/NET0131  , \memory_reg[8][0]/NET0131  , \memory_reg[8][1]/NET0131  , \memory_reg[9][0]/NET0131  , \memory_reg[9][1]/NET0131  , \nl[0]_pad  , \nl[2]_pad  , \nl[3]_pad  , \nl_reg[1]/NET0131  , nloss_pad , \play_reg/NET0131  , \s_reg/NET0131  , \scan_reg[0]/NET0131  , \scan_reg[1]/NET0131  , \scan_reg[2]/NET0131  , \scan_reg[3]/NET0131  , \scan_reg[4]/NET0131  , \sound_reg[0]/NET0131  , \sound_reg[1]/NET0131  , \sound_reg[2]/NET0131  , speaker_pad , start_pad , \timebase_reg[0]/NET0131  , \timebase_reg[1]/NET0131  , \timebase_reg[2]/NET0131  , \timebase_reg[3]/NET0131  , \timebase_reg[4]/NET0131  , \timebase_reg[5]/NET0131  , \wr_reg/NET0131  , \_al_n0  , \_al_n1  , \count_reg[0]/P0001  , \g10376/_0_  , \g11078/_0_  , \g11102/_0_  , \g11126/_0_  , \g11156/_0_  , \g11299/_0_  , \g11308/_0_  , \g11318/_0_  , \g11346/_0_  , \g11378/_0_  , \g11516/_0_  , \g63/_0_  , \g8501/_0_  , \g8516/_0_  , \g8517/_0_  , \g8519/_0_  , \g8520/_0_  , \g8522/_0_  , \g8526/_0_  , \g8529/_2_  , \g8545/_0_  , \g8546/_0_  , \g8547/_0_  , \g8555/_0_  , \g8556/_0_  , \g8557/_0_  , \g8558/_0_  , \g8559/_0_  , \g8560/_0_  , \g8562/_0_  , \g8563/_0_  , \g8581/_0_  , \g8586/_0_  , \g8591/_0_  , \g8594/_0_  , \g8606/_0_  , \g8608/_0_  , \g8647/_0_  , \g8659/_0_  , \g8695/_0_  , \g8784/_0_  , \g8797/_0_  , \g8854/_2_  , \g8869/_0_  , \g8871/_0_  , \g8889/_0_  , \g8891/_0_  , \g8892/_0_  , \g8894/_0_  , \g8970/_0_  , \g8975/_0_  , \g8992/_0_  , \g9180/_0_  , \g9183/_0_  , \g9511/u3_syn_4  , \g9513/u3_syn_4  , \g9515/u3_syn_4  , \g9517/u3_syn_4  , \g9519/u3_syn_4  , \g9521/u3_syn_4  , \g9523/u3_syn_4  , \g9525/u3_syn_4  , \g9527/u3_syn_4  , \g9529/u3_syn_4  , \g9531/u3_syn_4  , \g9533/u3_syn_4  , \g9535/u3_syn_4  , \g9537/u3_syn_4  , \g9539/u3_syn_4  , \g9541/u3_syn_4  , \g9543/u3_syn_4  , \g9545/u3_syn_4  , \g9547/u3_syn_4  , \g9549/u3_syn_4  , \g9551/u3_syn_4  , \g9553/u3_syn_4  , \g9555/u3_syn_4  , \g9557/u3_syn_4  , \g9559/u3_syn_4  , \g9560/u3_syn_4  , \g9562/u3_syn_4  , \g9564/u3_syn_4  , \g9566/u3_syn_4  , \g9568/u3_syn_4  , \g9570/u3_syn_4  , \g9572/u3_syn_4  );
  input \address_reg[0]/NET0131  ;
  input \address_reg[1]/NET0131  ;
  input \address_reg[2]/NET0131  ;
  input \address_reg[3]/NET0131  ;
  input \address_reg[4]/NET0131  ;
  input \count_reg[0]/NET0131  ;
  input \count_reg[0]1198/NET0131  ;
  input \count_reg[1]/NET0131  ;
  input \count_reg[1]1200/NET0131  ;
  input \count_reg[2]/NET0131  ;
  input \count_reg[3]/NET0131  ;
  input \count_reg[4]/NET0131  ;
  input \count_reg[5]/NET0131  ;
  input \counter_reg[0]/NET0131  ;
  input \counter_reg[1]/NET0131  ;
  input \counter_reg[2]/NET0131  ;
  input \data_in_reg[0]/NET0131  ;
  input \data_in_reg[1]/NET0131  ;
  input \data_out_reg[0]/NET0131  ;
  input \data_out_reg[1]/NET0131  ;
  input \gamma_reg[0]/NET0131  ;
  input \gamma_reg[1]/NET0131  ;
  input \gamma_reg[2]/NET0131  ;
  input \gamma_reg[3]/NET0131  ;
  input \gamma_reg[4]/NET0131  ;
  input \ind_reg[0]/NET0131  ;
  input \ind_reg[1]/NET0131  ;
  input \k[0]_pad  ;
  input \k[1]_pad  ;
  input \k[2]_pad  ;
  input \k[3]_pad  ;
  input \max_reg[0]/NET0131  ;
  input \max_reg[1]/NET0131  ;
  input \max_reg[2]/NET0131  ;
  input \max_reg[3]/NET0131  ;
  input \max_reg[4]/NET0131  ;
  input \memory_reg[0][0]/NET0131  ;
  input \memory_reg[0][1]/NET0131  ;
  input \memory_reg[10][0]/NET0131  ;
  input \memory_reg[10][1]/NET0131  ;
  input \memory_reg[11][0]/NET0131  ;
  input \memory_reg[11][1]/NET0131  ;
  input \memory_reg[12][0]/NET0131  ;
  input \memory_reg[12][1]/NET0131  ;
  input \memory_reg[13][0]/NET0131  ;
  input \memory_reg[13][1]/NET0131  ;
  input \memory_reg[14][0]/NET0131  ;
  input \memory_reg[14][1]/NET0131  ;
  input \memory_reg[15][0]/NET0131  ;
  input \memory_reg[15][1]/NET0131  ;
  input \memory_reg[16][0]/NET0131  ;
  input \memory_reg[16][1]/NET0131  ;
  input \memory_reg[17][0]/NET0131  ;
  input \memory_reg[17][1]/NET0131  ;
  input \memory_reg[18][0]/NET0131  ;
  input \memory_reg[18][1]/NET0131  ;
  input \memory_reg[19][0]/NET0131  ;
  input \memory_reg[19][1]/NET0131  ;
  input \memory_reg[1][0]/NET0131  ;
  input \memory_reg[1][1]/NET0131  ;
  input \memory_reg[20][0]/NET0131  ;
  input \memory_reg[20][1]/NET0131  ;
  input \memory_reg[21][0]/NET0131  ;
  input \memory_reg[21][1]/NET0131  ;
  input \memory_reg[22][0]/NET0131  ;
  input \memory_reg[22][1]/NET0131  ;
  input \memory_reg[23][0]/NET0131  ;
  input \memory_reg[23][1]/NET0131  ;
  input \memory_reg[24][0]/NET0131  ;
  input \memory_reg[24][1]/NET0131  ;
  input \memory_reg[25][0]/NET0131  ;
  input \memory_reg[25][1]/NET0131  ;
  input \memory_reg[26][0]/NET0131  ;
  input \memory_reg[26][1]/NET0131  ;
  input \memory_reg[27][0]/NET0131  ;
  input \memory_reg[27][1]/NET0131  ;
  input \memory_reg[28][0]/NET0131  ;
  input \memory_reg[28][1]/NET0131  ;
  input \memory_reg[29][0]/NET0131  ;
  input \memory_reg[29][1]/NET0131  ;
  input \memory_reg[2][0]/NET0131  ;
  input \memory_reg[2][1]/NET0131  ;
  input \memory_reg[30][0]/NET0131  ;
  input \memory_reg[30][1]/NET0131  ;
  input \memory_reg[31][0]/NET0131  ;
  input \memory_reg[31][1]/NET0131  ;
  input \memory_reg[3][0]/NET0131  ;
  input \memory_reg[3][1]/NET0131  ;
  input \memory_reg[4][0]/NET0131  ;
  input \memory_reg[4][1]/NET0131  ;
  input \memory_reg[5][0]/NET0131  ;
  input \memory_reg[5][1]/NET0131  ;
  input \memory_reg[6][0]/NET0131  ;
  input \memory_reg[6][1]/NET0131  ;
  input \memory_reg[7][0]/NET0131  ;
  input \memory_reg[7][1]/NET0131  ;
  input \memory_reg[8][0]/NET0131  ;
  input \memory_reg[8][1]/NET0131  ;
  input \memory_reg[9][0]/NET0131  ;
  input \memory_reg[9][1]/NET0131  ;
  input \nl[0]_pad  ;
  input \nl[2]_pad  ;
  input \nl[3]_pad  ;
  input \nl_reg[1]/NET0131  ;
  input nloss_pad ;
  input \play_reg/NET0131  ;
  input \s_reg/NET0131  ;
  input \scan_reg[0]/NET0131  ;
  input \scan_reg[1]/NET0131  ;
  input \scan_reg[2]/NET0131  ;
  input \scan_reg[3]/NET0131  ;
  input \scan_reg[4]/NET0131  ;
  input \sound_reg[0]/NET0131  ;
  input \sound_reg[1]/NET0131  ;
  input \sound_reg[2]/NET0131  ;
  input speaker_pad ;
  input start_pad ;
  input \timebase_reg[0]/NET0131  ;
  input \timebase_reg[1]/NET0131  ;
  input \timebase_reg[2]/NET0131  ;
  input \timebase_reg[3]/NET0131  ;
  input \timebase_reg[4]/NET0131  ;
  input \timebase_reg[5]/NET0131  ;
  input \wr_reg/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \count_reg[0]/P0001  ;
  output \g10376/_0_  ;
  output \g11078/_0_  ;
  output \g11102/_0_  ;
  output \g11126/_0_  ;
  output \g11156/_0_  ;
  output \g11299/_0_  ;
  output \g11308/_0_  ;
  output \g11318/_0_  ;
  output \g11346/_0_  ;
  output \g11378/_0_  ;
  output \g11516/_0_  ;
  output \g63/_0_  ;
  output \g8501/_0_  ;
  output \g8516/_0_  ;
  output \g8517/_0_  ;
  output \g8519/_0_  ;
  output \g8520/_0_  ;
  output \g8522/_0_  ;
  output \g8526/_0_  ;
  output \g8529/_2_  ;
  output \g8545/_0_  ;
  output \g8546/_0_  ;
  output \g8547/_0_  ;
  output \g8555/_0_  ;
  output \g8556/_0_  ;
  output \g8557/_0_  ;
  output \g8558/_0_  ;
  output \g8559/_0_  ;
  output \g8560/_0_  ;
  output \g8562/_0_  ;
  output \g8563/_0_  ;
  output \g8581/_0_  ;
  output \g8586/_0_  ;
  output \g8591/_0_  ;
  output \g8594/_0_  ;
  output \g8606/_0_  ;
  output \g8608/_0_  ;
  output \g8647/_0_  ;
  output \g8659/_0_  ;
  output \g8695/_0_  ;
  output \g8784/_0_  ;
  output \g8797/_0_  ;
  output \g8854/_2_  ;
  output \g8869/_0_  ;
  output \g8871/_0_  ;
  output \g8889/_0_  ;
  output \g8891/_0_  ;
  output \g8892/_0_  ;
  output \g8894/_0_  ;
  output \g8970/_0_  ;
  output \g8975/_0_  ;
  output \g8992/_0_  ;
  output \g9180/_0_  ;
  output \g9183/_0_  ;
  output \g9511/u3_syn_4  ;
  output \g9513/u3_syn_4  ;
  output \g9515/u3_syn_4  ;
  output \g9517/u3_syn_4  ;
  output \g9519/u3_syn_4  ;
  output \g9521/u3_syn_4  ;
  output \g9523/u3_syn_4  ;
  output \g9525/u3_syn_4  ;
  output \g9527/u3_syn_4  ;
  output \g9529/u3_syn_4  ;
  output \g9531/u3_syn_4  ;
  output \g9533/u3_syn_4  ;
  output \g9535/u3_syn_4  ;
  output \g9537/u3_syn_4  ;
  output \g9539/u3_syn_4  ;
  output \g9541/u3_syn_4  ;
  output \g9543/u3_syn_4  ;
  output \g9545/u3_syn_4  ;
  output \g9547/u3_syn_4  ;
  output \g9549/u3_syn_4  ;
  output \g9551/u3_syn_4  ;
  output \g9553/u3_syn_4  ;
  output \g9555/u3_syn_4  ;
  output \g9557/u3_syn_4  ;
  output \g9559/u3_syn_4  ;
  output \g9560/u3_syn_4  ;
  output \g9562/u3_syn_4  ;
  output \g9564/u3_syn_4  ;
  output \g9566/u3_syn_4  ;
  output \g9568/u3_syn_4  ;
  output \g9570/u3_syn_4  ;
  output \g9572/u3_syn_4  ;
  wire n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 ;
  assign n125 = \count_reg[0]/NET0131  & ~\count_reg[1]/NET0131  ;
  assign n126 = ~\count_reg[0]/NET0131  & \count_reg[1]/NET0131  ;
  assign n127 = ~n125 & ~n126 ;
  assign n152 = ~\gamma_reg[0]/NET0131  & ~start_pad ;
  assign n153 = \gamma_reg[2]/NET0131  & ~start_pad ;
  assign n154 = \gamma_reg[1]/NET0131  & ~start_pad ;
  assign n155 = n153 & ~n154 ;
  assign n156 = \gamma_reg[4]/NET0131  & ~start_pad ;
  assign n157 = \gamma_reg[3]/NET0131  & ~start_pad ;
  assign n158 = ~n156 & n157 ;
  assign n159 = n155 & n158 ;
  assign n160 = ~n152 & n159 ;
  assign n161 = ~\count_reg[0]1198/NET0131  & ~\count_reg[1]1200/NET0131  ;
  assign n162 = ~\count_reg[2]/NET0131  & n161 ;
  assign n163 = ~\count_reg[3]/NET0131  & ~\count_reg[4]/NET0131  ;
  assign n164 = n162 & n163 ;
  assign n165 = ~\count_reg[5]/NET0131  & n164 ;
  assign n181 = n160 & ~n165 ;
  assign n175 = ~n153 & n154 ;
  assign n176 = n158 & n175 ;
  assign n177 = ~n152 & n176 ;
  assign n169 = ~n156 & ~n157 ;
  assign n172 = n153 & n154 ;
  assign n178 = n169 & n172 ;
  assign n179 = ~\gamma_reg[0]/NET0131  & n178 ;
  assign n180 = ~n177 & ~n179 ;
  assign n170 = n155 & n169 ;
  assign n171 = n156 & ~n157 ;
  assign n173 = n171 & n172 ;
  assign n174 = ~n170 & ~n173 ;
  assign n182 = n169 & n175 ;
  assign n183 = ~n152 & n182 ;
  assign n184 = n174 & ~n183 ;
  assign n185 = n180 & n184 ;
  assign n186 = ~n181 & n185 ;
  assign n193 = ~\gamma_reg[0]/NET0131  & n171 ;
  assign n194 = n155 & n193 ;
  assign n190 = n158 & n172 ;
  assign n195 = \gamma_reg[0]/NET0131  & n190 ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = \gamma_reg[0]/NET0131  & n171 ;
  assign n198 = ~n153 & n197 ;
  assign n199 = n196 & ~n198 ;
  assign n187 = ~n153 & ~n154 ;
  assign n188 = ~n171 & n187 ;
  assign n189 = n152 & n159 ;
  assign n191 = ~\gamma_reg[0]/NET0131  & n190 ;
  assign n192 = ~n189 & ~n191 ;
  assign n206 = ~n188 & n192 ;
  assign n200 = n175 & n193 ;
  assign n201 = n155 & n197 ;
  assign n202 = ~n200 & ~n201 ;
  assign n203 = n152 & n176 ;
  assign n204 = n187 & n193 ;
  assign n205 = ~n203 & ~n204 ;
  assign n207 = n202 & n205 ;
  assign n208 = n206 & n207 ;
  assign n209 = n199 & n208 ;
  assign n210 = n186 & n209 ;
  assign n211 = \scan_reg[1]/NET0131  & ~n210 ;
  assign n128 = \max_reg[3]/NET0131  & \scan_reg[3]/NET0131  ;
  assign n129 = ~\max_reg[3]/NET0131  & ~\scan_reg[3]/NET0131  ;
  assign n130 = ~n128 & ~n129 ;
  assign n133 = ~\max_reg[4]/NET0131  & ~\scan_reg[4]/NET0131  ;
  assign n134 = \max_reg[4]/NET0131  & \scan_reg[4]/NET0131  ;
  assign n135 = ~n133 & ~n134 ;
  assign n131 = \max_reg[1]/NET0131  & ~\scan_reg[1]/NET0131  ;
  assign n132 = ~\max_reg[1]/NET0131  & \scan_reg[1]/NET0131  ;
  assign n142 = ~n131 & ~n132 ;
  assign n143 = ~n135 & n142 ;
  assign n136 = ~\max_reg[2]/NET0131  & ~\scan_reg[2]/NET0131  ;
  assign n137 = \max_reg[2]/NET0131  & \scan_reg[2]/NET0131  ;
  assign n138 = ~n136 & ~n137 ;
  assign n139 = ~\max_reg[0]/NET0131  & ~\scan_reg[0]/NET0131  ;
  assign n140 = \max_reg[0]/NET0131  & \scan_reg[0]/NET0131  ;
  assign n141 = ~n139 & ~n140 ;
  assign n144 = ~n138 & ~n141 ;
  assign n145 = n143 & n144 ;
  assign n146 = ~n130 & n145 ;
  assign n148 = \scan_reg[0]/NET0131  & \scan_reg[1]/NET0131  ;
  assign n149 = ~\scan_reg[0]/NET0131  & ~\scan_reg[1]/NET0131  ;
  assign n150 = ~n148 & ~n149 ;
  assign n151 = ~n146 & ~n150 ;
  assign n147 = ~\scan_reg[1]/NET0131  & n146 ;
  assign n166 = n160 & n165 ;
  assign n167 = ~n147 & n166 ;
  assign n168 = ~n151 & n167 ;
  assign n212 = \scan_reg[1]/NET0131  & ~n165 ;
  assign n213 = ~n146 & n165 ;
  assign n214 = n150 & n213 ;
  assign n215 = ~n212 & ~n214 ;
  assign n216 = \gamma_reg[0]/NET0131  & n178 ;
  assign n217 = ~n215 & n216 ;
  assign n218 = ~n168 & ~n217 ;
  assign n219 = ~n211 & n218 ;
  assign n244 = \gamma_reg[0]/NET0131  & n170 ;
  assign n220 = n158 & n187 ;
  assign n245 = ~n152 & n220 ;
  assign n246 = ~n244 & ~n245 ;
  assign n232 = ~n153 & n193 ;
  assign n233 = ~n160 & ~n232 ;
  assign n234 = ~n190 & ~n216 ;
  assign n254 = n233 & n234 ;
  assign n255 = n246 & n254 ;
  assign n235 = \gamma_reg[3]/NET0131  & n156 ;
  assign n236 = n187 & n235 ;
  assign n237 = n152 & n236 ;
  assign n238 = ~n201 & ~n203 ;
  assign n239 = ~n237 & n238 ;
  assign n231 = n175 & n197 ;
  assign n228 = n169 & n187 ;
  assign n229 = ~n152 & n228 ;
  assign n230 = n152 & n170 ;
  assign n252 = ~n229 & ~n230 ;
  assign n253 = ~n231 & n252 ;
  assign n256 = n239 & n253 ;
  assign n240 = ~n179 & ~n189 ;
  assign n241 = n152 & n228 ;
  assign n242 = ~n177 & ~n241 ;
  assign n243 = n240 & n242 ;
  assign n247 = n152 & n173 ;
  assign n248 = ~n194 & ~n247 ;
  assign n249 = ~n173 & ~n236 ;
  assign n250 = ~n152 & ~n249 ;
  assign n251 = n248 & ~n250 ;
  assign n257 = n243 & n251 ;
  assign n258 = n256 & n257 ;
  assign n259 = n255 & n258 ;
  assign n260 = \address_reg[0]/NET0131  & ~n259 ;
  assign n221 = n152 & n220 ;
  assign n222 = ~n183 & ~n221 ;
  assign n223 = \scan_reg[0]/NET0131  & ~n222 ;
  assign n224 = n187 & n197 ;
  assign n225 = n152 & n182 ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = \max_reg[0]/NET0131  & ~n226 ;
  assign n261 = ~n223 & ~n227 ;
  assign n262 = ~n260 & n261 ;
  assign n263 = ~\count_reg[5]/NET0131  & n163 ;
  assign n264 = \count_reg[3]/NET0131  & ~n162 ;
  assign n265 = ~\count_reg[3]/NET0131  & n162 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = ~n263 & ~n266 ;
  assign n268 = n146 & n165 ;
  assign n269 = \max_reg[0]/NET0131  & \max_reg[1]/NET0131  ;
  assign n270 = \max_reg[2]/NET0131  & n269 ;
  assign n271 = \max_reg[3]/NET0131  & n270 ;
  assign n272 = \max_reg[4]/NET0131  & n271 ;
  assign n273 = ~\count_reg[3]/NET0131  & ~n272 ;
  assign n274 = n268 & ~n273 ;
  assign n275 = ~n267 & ~n274 ;
  assign n276 = n160 & ~n275 ;
  assign n292 = ~n225 & ~n241 ;
  assign n293 = ~n224 & n292 ;
  assign n294 = \count_reg[3]/NET0131  & ~n293 ;
  assign n290 = ~n231 & ~n244 ;
  assign n291 = \timebase_reg[3]/NET0131  & ~n290 ;
  assign n295 = n165 & n201 ;
  assign n296 = n146 & n295 ;
  assign n309 = ~n291 & ~n296 ;
  assign n310 = ~n294 & n309 ;
  assign n297 = \timebase_reg[3]/NET0131  & n165 ;
  assign n298 = ~n267 & ~n297 ;
  assign n299 = n196 & n240 ;
  assign n300 = ~n298 & ~n299 ;
  assign n302 = ~\k[0]_pad  & ~\k[1]_pad  ;
  assign n303 = ~\k[2]_pad  & ~\k[3]_pad  ;
  assign n304 = n302 & n303 ;
  assign n306 = n266 & n304 ;
  assign n301 = ~n165 & n203 ;
  assign n305 = ~\timebase_reg[3]/NET0131  & ~n304 ;
  assign n307 = n301 & ~n305 ;
  assign n308 = ~n306 & n307 ;
  assign n311 = ~n300 & ~n308 ;
  assign n312 = n310 & n311 ;
  assign n278 = ~n183 & ~n229 ;
  assign n279 = ~n200 & ~n230 ;
  assign n280 = n278 & n279 ;
  assign n277 = ~n177 & ~n191 ;
  assign n281 = ~n245 & n277 ;
  assign n282 = n280 & n281 ;
  assign n283 = \count_reg[3]/NET0131  & ~n282 ;
  assign n285 = ~n201 & ~n204 ;
  assign n286 = ~n263 & ~n285 ;
  assign n284 = ~n165 & n216 ;
  assign n287 = n249 & ~n284 ;
  assign n288 = ~n286 & n287 ;
  assign n289 = ~n266 & ~n288 ;
  assign n313 = ~n283 & ~n289 ;
  assign n314 = n312 & n313 ;
  assign n315 = ~n276 & n314 ;
  assign n320 = ~n195 & ~n203 ;
  assign n321 = ~n165 & ~n320 ;
  assign n322 = ~n173 & ~n191 ;
  assign n323 = ~n200 & n322 ;
  assign n326 = ~n296 & n323 ;
  assign n327 = ~n321 & n326 ;
  assign n317 = n146 & ~n272 ;
  assign n318 = n166 & n317 ;
  assign n316 = n216 & ~n268 ;
  assign n319 = ~n179 & ~n229 ;
  assign n324 = n226 & n246 ;
  assign n325 = n319 & n324 ;
  assign n328 = ~n316 & n325 ;
  assign n329 = ~n318 & n328 ;
  assign n330 = n327 & n329 ;
  assign n358 = n128 & n145 ;
  assign n359 = n270 & n358 ;
  assign n360 = \max_reg[4]/NET0131  & n359 ;
  assign n361 = n166 & ~n360 ;
  assign n362 = ~n182 & n319 ;
  assign n355 = ~n189 & ~n224 ;
  assign n356 = ~n190 & ~n194 ;
  assign n357 = n355 & n356 ;
  assign n341 = ~n152 & n173 ;
  assign n363 = ~n216 & ~n220 ;
  assign n364 = ~n341 & n363 ;
  assign n365 = n357 & n364 ;
  assign n366 = n362 & n365 ;
  assign n367 = ~n361 & n366 ;
  assign n368 = \sound_reg[0]/NET0131  & ~n367 ;
  assign n349 = ~n177 & ~n201 ;
  assign n350 = ~n247 & n349 ;
  assign n351 = ~n181 & n350 ;
  assign n344 = ~n204 & ~n237 ;
  assign n345 = n279 & n344 ;
  assign n346 = ~n152 & n236 ;
  assign n347 = ~n165 & n346 ;
  assign n348 = ~n241 & ~n347 ;
  assign n352 = n345 & n348 ;
  assign n353 = n351 & n352 ;
  assign n354 = \sound_reg[0]/NET0131  & ~n353 ;
  assign n331 = ~\k[0]_pad  & ~\k[2]_pad  ;
  assign n332 = ~n165 & ~n331 ;
  assign n333 = \k[3]_pad  & ~n165 ;
  assign n334 = ~\sound_reg[0]/NET0131  & ~n333 ;
  assign n335 = ~n332 & ~n334 ;
  assign n336 = ~\k[0]_pad  & \k[1]_pad  ;
  assign n337 = ~n165 & n336 ;
  assign n338 = ~n335 & ~n337 ;
  assign n339 = n203 & ~n338 ;
  assign n340 = \data_out_reg[0]/NET0131  & ~n290 ;
  assign n342 = n165 & n341 ;
  assign n343 = ~n296 & ~n342 ;
  assign n369 = ~n340 & n343 ;
  assign n370 = ~n339 & n369 ;
  assign n371 = ~n354 & n370 ;
  assign n372 = ~n368 & n371 ;
  assign n375 = \count_reg[4]/NET0131  & ~n265 ;
  assign n376 = ~n164 & ~n375 ;
  assign n377 = ~n165 & ~n376 ;
  assign n378 = n165 & ~n299 ;
  assign n379 = \timebase_reg[4]/NET0131  & n378 ;
  assign n380 = ~n377 & ~n379 ;
  assign n382 = ~n160 & ~n341 ;
  assign n381 = ~n201 & ~n216 ;
  assign n383 = ~n237 & n381 ;
  assign n384 = n382 & n383 ;
  assign n385 = ~n204 & n384 ;
  assign n386 = ~n247 & ~n346 ;
  assign n387 = n240 & n386 ;
  assign n388 = n196 & n387 ;
  assign n389 = n385 & n388 ;
  assign n390 = ~n380 & ~n389 ;
  assign n373 = n282 & n293 ;
  assign n374 = \count_reg[4]/NET0131  & ~n373 ;
  assign n391 = n301 & n304 ;
  assign n392 = ~n376 & n391 ;
  assign n393 = n301 & ~n304 ;
  assign n394 = n290 & ~n393 ;
  assign n395 = \timebase_reg[4]/NET0131  & ~n394 ;
  assign n396 = ~n392 & ~n395 ;
  assign n397 = ~n374 & n396 ;
  assign n398 = ~n390 & n397 ;
  assign n405 = \count_reg[5]/NET0131  & ~n164 ;
  assign n406 = n385 & ~n391 ;
  assign n407 = n405 & ~n406 ;
  assign n399 = ~n164 & ~n386 ;
  assign n400 = ~n220 & n277 ;
  assign n401 = n280 & n400 ;
  assign n402 = n293 & n401 ;
  assign n403 = ~n399 & n402 ;
  assign n404 = \count_reg[5]/NET0131  & ~n403 ;
  assign n408 = ~n378 & n394 ;
  assign n409 = \timebase_reg[5]/NET0131  & ~n408 ;
  assign n410 = ~n299 & n405 ;
  assign n411 = ~n221 & ~n410 ;
  assign n412 = ~n409 & n411 ;
  assign n413 = ~n404 & n412 ;
  assign n414 = ~n407 & n413 ;
  assign n415 = ~n165 & ~n388 ;
  assign n416 = ~n224 & ~n415 ;
  assign n418 = ~n165 & n201 ;
  assign n419 = ~n200 & ~n418 ;
  assign n417 = n205 & ~n341 ;
  assign n420 = n292 & n417 ;
  assign n421 = n419 & n420 ;
  assign n422 = n416 & n421 ;
  assign n423 = \nl_reg[1]/NET0131  & ~n422 ;
  assign n430 = \data_out_reg[0]/NET0131  & ~\data_out_reg[1]/NET0131  ;
  assign n431 = n290 & n343 ;
  assign n432 = n430 & ~n431 ;
  assign n433 = ~n183 & ~n230 ;
  assign n434 = n363 & n433 ;
  assign n435 = n290 & ~n295 ;
  assign n436 = n434 & n435 ;
  assign n437 = \nl_reg[1]/NET0131  & ~n436 ;
  assign n424 = ~n160 & n277 ;
  assign n425 = ~n237 & n424 ;
  assign n426 = \ind_reg[0]/NET0131  & ~\ind_reg[1]/NET0131  ;
  assign n427 = ~n277 & n426 ;
  assign n428 = ~\nl_reg[1]/NET0131  & ~n427 ;
  assign n429 = ~n425 & ~n428 ;
  assign n438 = n165 & n237 ;
  assign n439 = ~n429 & ~n438 ;
  assign n440 = ~n437 & n439 ;
  assign n441 = ~n432 & n440 ;
  assign n442 = ~n423 & n441 ;
  assign n445 = n268 & ~n272 ;
  assign n446 = n160 & ~n445 ;
  assign n443 = n216 & n268 ;
  assign n444 = n157 & n187 ;
  assign n447 = ~n189 & ~n444 ;
  assign n448 = n277 & n447 ;
  assign n449 = ~n321 & n448 ;
  assign n450 = ~n443 & n449 ;
  assign n451 = ~n446 & n450 ;
  assign n457 = n242 & ~n341 ;
  assign n458 = ~n160 & n386 ;
  assign n459 = n357 & n458 ;
  assign n460 = n457 & n459 ;
  assign n452 = ~n165 & ~n303 ;
  assign n453 = ~n165 & ~n302 ;
  assign n454 = n203 & ~n453 ;
  assign n455 = ~n452 & n454 ;
  assign n456 = ~n221 & n345 ;
  assign n461 = ~n455 & n456 ;
  assign n462 = n460 & n461 ;
  assign n463 = \sound_reg[2]/NET0131  & ~n462 ;
  assign n466 = ~\sound_reg[2]/NET0131  & ~n296 ;
  assign n467 = ~n245 & n362 ;
  assign n468 = n381 & n467 ;
  assign n469 = ~n466 & ~n468 ;
  assign n464 = n166 & n360 ;
  assign n465 = n165 & n250 ;
  assign n470 = ~n464 & ~n465 ;
  assign n471 = ~n469 & n470 ;
  assign n472 = ~n463 & n471 ;
  assign n475 = ~\gamma_reg[4]/NET0131  & n155 ;
  assign n476 = ~n190 & ~n475 ;
  assign n477 = ~n198 & n476 ;
  assign n478 = n180 & n477 ;
  assign n479 = n363 & n478 ;
  assign n480 = n251 & n479 ;
  assign n473 = n202 & ~n241 ;
  assign n474 = n344 & n473 ;
  assign n481 = ~n182 & n474 ;
  assign n482 = n480 & n481 ;
  assign n483 = nloss_pad & ~n482 ;
  assign n484 = \k[1]_pad  & ~n430 ;
  assign n487 = \data_out_reg[0]/NET0131  & \data_out_reg[1]/NET0131  ;
  assign n488 = ~\k[2]_pad  & n487 ;
  assign n485 = ~\data_out_reg[0]/NET0131  & \data_out_reg[1]/NET0131  ;
  assign n486 = \k[2]_pad  & n485 ;
  assign n489 = ~\k[1]_pad  & ~n303 ;
  assign n490 = ~n486 & n489 ;
  assign n491 = ~n488 & n490 ;
  assign n492 = ~n484 & ~n491 ;
  assign n493 = ~\k[0]_pad  & ~n492 ;
  assign n494 = ~\data_out_reg[0]/NET0131  & ~\data_out_reg[1]/NET0131  ;
  assign n495 = \k[0]_pad  & ~n494 ;
  assign n496 = ~n493 & ~n495 ;
  assign n497 = ~nloss_pad & ~n165 ;
  assign n498 = n496 & n497 ;
  assign n499 = n203 & ~n498 ;
  assign n500 = ~n483 & ~n499 ;
  assign n515 = n201 & ~n268 ;
  assign n501 = \k[3]_pad  & n488 ;
  assign n502 = ~n486 & ~n501 ;
  assign n503 = n302 & ~n502 ;
  assign n504 = ~\k[0]_pad  & ~n430 ;
  assign n505 = ~n302 & ~n495 ;
  assign n506 = ~n504 & n505 ;
  assign n507 = ~n503 & ~n506 ;
  assign n508 = n203 & ~n507 ;
  assign n522 = ~n316 & ~n508 ;
  assign n523 = ~n515 & n522 ;
  assign n509 = ~n203 & n240 ;
  assign n510 = n248 & n344 ;
  assign n511 = n509 & n510 ;
  assign n512 = n165 & ~n511 ;
  assign n513 = ~n165 & n195 ;
  assign n518 = n279 & ~n347 ;
  assign n519 = ~n513 & n518 ;
  assign n514 = ~n165 & ~n382 ;
  assign n516 = ~n191 & ~n221 ;
  assign n517 = ~n225 & n516 ;
  assign n520 = ~n514 & n517 ;
  assign n521 = n519 & n520 ;
  assign n524 = ~n512 & n521 ;
  assign n525 = n523 & n524 ;
  assign n527 = n301 & ~n496 ;
  assign n528 = n201 & ~n213 ;
  assign n529 = n192 & ~n284 ;
  assign n526 = ~n194 & ~n231 ;
  assign n530 = ~n513 & n526 ;
  assign n531 = n529 & n530 ;
  assign n532 = n186 & n531 ;
  assign n533 = ~n528 & n532 ;
  assign n534 = ~n527 & n533 ;
  assign n537 = ~n237 & n434 ;
  assign n538 = n202 & n292 ;
  assign n539 = n537 & n538 ;
  assign n540 = n417 & n539 ;
  assign n541 = \nl[0]_pad  & ~n540 ;
  assign n535 = n290 & ~n415 ;
  assign n536 = \nl[0]_pad  & ~n535 ;
  assign n542 = ~n431 & n494 ;
  assign n543 = ~\ind_reg[0]/NET0131  & ~\ind_reg[1]/NET0131  ;
  assign n544 = ~n277 & n543 ;
  assign n545 = ~\nl[0]_pad  & ~n544 ;
  assign n546 = ~n224 & n424 ;
  assign n547 = ~n545 & ~n546 ;
  assign n548 = ~n438 & ~n547 ;
  assign n549 = ~n542 & n548 ;
  assign n550 = ~n536 & n549 ;
  assign n551 = ~n541 & n550 ;
  assign n563 = ~n160 & n205 ;
  assign n564 = n293 & n563 ;
  assign n565 = n419 & n564 ;
  assign n566 = n537 & n565 ;
  assign n567 = ~n415 & n566 ;
  assign n568 = \nl[2]_pad  & ~n567 ;
  assign n558 = ~\nl[2]_pad  & ~n485 ;
  assign n559 = ~\nl[2]_pad  & ~n165 ;
  assign n560 = n341 & ~n559 ;
  assign n561 = n290 & ~n560 ;
  assign n562 = ~n558 & ~n561 ;
  assign n552 = n146 & n485 ;
  assign n553 = ~\nl[2]_pad  & ~n552 ;
  assign n554 = n295 & ~n553 ;
  assign n555 = ~\ind_reg[0]/NET0131  & \ind_reg[1]/NET0131  ;
  assign n556 = ~\nl[2]_pad  & ~n555 ;
  assign n557 = ~n277 & ~n556 ;
  assign n569 = ~n438 & ~n557 ;
  assign n570 = ~n554 & n569 ;
  assign n571 = ~n562 & n570 ;
  assign n572 = ~n568 & n571 ;
  assign n573 = n416 & n539 ;
  assign n574 = \nl[3]_pad  & ~n573 ;
  assign n575 = \nl[3]_pad  & ~n290 ;
  assign n576 = ~n487 & ~n575 ;
  assign n577 = ~n431 & ~n576 ;
  assign n578 = n417 & n424 ;
  assign n579 = \ind_reg[0]/NET0131  & \ind_reg[1]/NET0131  ;
  assign n580 = ~n277 & n579 ;
  assign n581 = ~\nl[3]_pad  & ~n580 ;
  assign n582 = ~n578 & ~n581 ;
  assign n583 = ~n438 & ~n582 ;
  assign n584 = ~n577 & n583 ;
  assign n585 = ~n574 & n584 ;
  assign n590 = ~n183 & ~n236 ;
  assign n591 = ~n244 & n590 ;
  assign n592 = ~n181 & n192 ;
  assign n593 = n279 & ~n301 ;
  assign n597 = n592 & n593 ;
  assign n598 = n591 & n597 ;
  assign n586 = ~n173 & ~n195 ;
  assign n587 = n180 & n586 ;
  assign n588 = n293 & n587 ;
  assign n594 = n363 & ~n418 ;
  assign n589 = ~n165 & n204 ;
  assign n595 = n526 & ~n589 ;
  assign n596 = n594 & n595 ;
  assign n599 = n588 & n596 ;
  assign n600 = n598 & n599 ;
  assign n601 = \max_reg[4]/NET0131  & ~n600 ;
  assign n602 = ~\max_reg[4]/NET0131  & ~n359 ;
  assign n603 = n166 & ~n602 ;
  assign n604 = \scan_reg[4]/NET0131  & n146 ;
  assign n605 = ~\max_reg[4]/NET0131  & ~n271 ;
  assign n606 = ~n272 & ~n605 ;
  assign n607 = ~n146 & n606 ;
  assign n608 = ~n604 & ~n607 ;
  assign n609 = n295 & ~n608 ;
  assign n610 = ~n603 & ~n609 ;
  assign n611 = ~n601 & n610 ;
  assign n612 = n165 & n360 ;
  assign n613 = ~\play_reg/NET0131  & ~n612 ;
  assign n614 = n160 & ~n613 ;
  assign n615 = ~n165 & ~n299 ;
  assign n616 = n226 & ~n615 ;
  assign n617 = \play_reg/NET0131  & ~n616 ;
  assign n624 = ~n165 & n247 ;
  assign n625 = ~n191 & ~n346 ;
  assign n626 = ~n624 & n625 ;
  assign n627 = n457 & n626 ;
  assign n628 = \play_reg/NET0131  & ~n627 ;
  assign n618 = ~\play_reg/NET0131  & ~n296 ;
  assign n619 = ~n232 & n238 ;
  assign n620 = n434 & n619 ;
  assign n621 = ~n618 & ~n620 ;
  assign n622 = \play_reg/NET0131  & ~n165 ;
  assign n623 = n237 & n622 ;
  assign n629 = ~n465 & ~n623 ;
  assign n630 = n394 & n629 ;
  assign n631 = ~n621 & n630 ;
  assign n632 = ~n628 & n631 ;
  assign n633 = ~n617 & n632 ;
  assign n634 = ~n614 & n633 ;
  assign n635 = n385 & n387 ;
  assign n636 = ~\count_reg[0]1198/NET0131  & ~n165 ;
  assign n637 = ~n635 & n636 ;
  assign n641 = \count_reg[0]1198/NET0131  & ~n402 ;
  assign n638 = n165 & ~n240 ;
  assign n639 = n290 & ~n638 ;
  assign n640 = \timebase_reg[0]/NET0131  & ~n639 ;
  assign n646 = \timebase_reg[0]/NET0131  & n165 ;
  assign n647 = ~n636 & ~n646 ;
  assign n648 = ~n196 & ~n647 ;
  assign n642 = ~\timebase_reg[0]/NET0131  & ~n304 ;
  assign n643 = \count_reg[0]1198/NET0131  & n304 ;
  assign n644 = ~n642 & ~n643 ;
  assign n645 = n301 & n644 ;
  assign n649 = ~n221 & ~n645 ;
  assign n650 = ~n648 & n649 ;
  assign n651 = ~n640 & n650 ;
  assign n652 = ~n641 & n651 ;
  assign n653 = ~n637 & n652 ;
  assign n655 = \count_reg[2]/NET0131  & ~n161 ;
  assign n656 = ~n162 & ~n655 ;
  assign n657 = ~n165 & ~n656 ;
  assign n658 = \timebase_reg[2]/NET0131  & n378 ;
  assign n659 = ~n657 & ~n658 ;
  assign n660 = n384 & n388 ;
  assign n661 = ~n659 & ~n660 ;
  assign n654 = \count_reg[2]/NET0131  & ~n373 ;
  assign n662 = \timebase_reg[2]/NET0131  & ~n394 ;
  assign n663 = ~n391 & ~n589 ;
  assign n664 = ~n656 & ~n663 ;
  assign n665 = ~n662 & ~n664 ;
  assign n666 = ~n654 & n665 ;
  assign n667 = ~n661 & n666 ;
  assign n668 = ~\timebase_reg[0]/NET0131  & ~\timebase_reg[1]/NET0131  ;
  assign n669 = ~n272 & n668 ;
  assign n670 = ~\timebase_reg[2]/NET0131  & n669 ;
  assign n671 = n268 & n670 ;
  assign n672 = ~\timebase_reg[3]/NET0131  & n671 ;
  assign n673 = ~\timebase_reg[4]/NET0131  & n672 ;
  assign n674 = ~\timebase_reg[5]/NET0131  & ~n673 ;
  assign n675 = ~\timebase_reg[4]/NET0131  & \timebase_reg[5]/NET0131  ;
  assign n676 = n672 & n675 ;
  assign n677 = n160 & ~n676 ;
  assign n678 = ~n674 & n677 ;
  assign n680 = n239 & n363 ;
  assign n679 = ~n172 & n193 ;
  assign n681 = n192 & ~n679 ;
  assign n682 = n433 & n681 ;
  assign n683 = n588 & n682 ;
  assign n684 = n680 & n683 ;
  assign n685 = \timebase_reg[5]/NET0131  & ~n684 ;
  assign n686 = n290 & ~n346 ;
  assign n687 = \timebase_reg[5]/NET0131  & ~n686 ;
  assign n688 = ~n229 & ~n687 ;
  assign n689 = ~n685 & n688 ;
  assign n690 = ~n678 & n689 ;
  assign n691 = \max_reg[3]/NET0131  & ~n600 ;
  assign n692 = \max_reg[3]/NET0131  & ~n317 ;
  assign n693 = ~\max_reg[3]/NET0131  & ~n270 ;
  assign n694 = ~n271 & ~n693 ;
  assign n695 = n146 & n694 ;
  assign n696 = ~n692 & ~n695 ;
  assign n697 = n166 & ~n696 ;
  assign n698 = ~n146 & n694 ;
  assign n699 = ~n358 & ~n698 ;
  assign n700 = n295 & ~n699 ;
  assign n701 = ~n697 & ~n700 ;
  assign n702 = ~n691 & n701 ;
  assign n703 = \timebase_reg[3]/NET0131  & ~n671 ;
  assign n704 = ~n672 & ~n703 ;
  assign n705 = n160 & ~n704 ;
  assign n706 = n684 & n686 ;
  assign n707 = \timebase_reg[3]/NET0131  & ~n706 ;
  assign n708 = ~n705 & ~n707 ;
  assign n710 = \count_reg[0]1198/NET0131  & \count_reg[1]1200/NET0131  ;
  assign n711 = ~n161 & ~n710 ;
  assign n712 = ~n165 & ~n711 ;
  assign n713 = \timebase_reg[1]/NET0131  & n378 ;
  assign n714 = ~n712 & ~n713 ;
  assign n715 = ~n389 & ~n714 ;
  assign n709 = \count_reg[1]1200/NET0131  & ~n373 ;
  assign n716 = n391 & ~n711 ;
  assign n717 = \timebase_reg[1]/NET0131  & ~n394 ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = ~n709 & n718 ;
  assign n720 = ~n715 & n719 ;
  assign n729 = \scan_reg[3]/NET0131  & ~n210 ;
  assign n721 = \scan_reg[3]/NET0131  & ~n165 ;
  assign n722 = \scan_reg[2]/NET0131  & n148 ;
  assign n723 = \scan_reg[3]/NET0131  & n722 ;
  assign n724 = ~\scan_reg[3]/NET0131  & ~n722 ;
  assign n725 = ~n723 & ~n724 ;
  assign n726 = n213 & n725 ;
  assign n727 = ~n721 & ~n726 ;
  assign n728 = n216 & ~n727 ;
  assign n730 = ~n146 & n725 ;
  assign n731 = ~n358 & ~n730 ;
  assign n732 = n166 & ~n731 ;
  assign n733 = ~n728 & ~n732 ;
  assign n734 = ~n729 & n733 ;
  assign n742 = \scan_reg[4]/NET0131  & ~n210 ;
  assign n735 = \scan_reg[4]/NET0131  & ~n165 ;
  assign n736 = \scan_reg[4]/NET0131  & ~n723 ;
  assign n737 = ~\scan_reg[4]/NET0131  & n723 ;
  assign n738 = ~n736 & ~n737 ;
  assign n739 = n213 & ~n738 ;
  assign n740 = ~n735 & ~n739 ;
  assign n741 = n216 & ~n740 ;
  assign n743 = ~n146 & ~n738 ;
  assign n744 = ~n604 & ~n743 ;
  assign n745 = n166 & ~n744 ;
  assign n746 = ~n741 & ~n745 ;
  assign n747 = ~n742 & n746 ;
  assign n758 = n234 & n456 ;
  assign n759 = ~n361 & n758 ;
  assign n760 = \sound_reg[1]/NET0131  & ~n759 ;
  assign n754 = ~n177 & n355 ;
  assign n755 = n467 & n754 ;
  assign n756 = ~n515 & n755 ;
  assign n757 = \sound_reg[1]/NET0131  & ~n756 ;
  assign n751 = n248 & n348 ;
  assign n752 = ~n514 & n751 ;
  assign n753 = \sound_reg[1]/NET0131  & ~n752 ;
  assign n748 = ~\sound_reg[1]/NET0131  & ~n452 ;
  assign n749 = n454 & ~n748 ;
  assign n750 = \data_out_reg[1]/NET0131  & ~n290 ;
  assign n761 = ~n749 & ~n750 ;
  assign n762 = ~n753 & n761 ;
  assign n763 = ~n757 & n762 ;
  assign n764 = ~n760 & n763 ;
  assign n765 = \timebase_reg[1]/NET0131  & ~n706 ;
  assign n766 = ~\timebase_reg[0]/NET0131  & n445 ;
  assign n767 = \timebase_reg[1]/NET0131  & ~n766 ;
  assign n768 = n268 & n669 ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = n160 & ~n769 ;
  assign n771 = ~n765 & ~n770 ;
  assign n772 = \timebase_reg[2]/NET0131  & ~n768 ;
  assign n773 = ~n671 & ~n772 ;
  assign n774 = n160 & ~n773 ;
  assign n775 = \timebase_reg[2]/NET0131  & ~n706 ;
  assign n776 = ~n774 & ~n775 ;
  assign n777 = \timebase_reg[4]/NET0131  & ~n706 ;
  assign n778 = \timebase_reg[4]/NET0131  & ~n672 ;
  assign n779 = ~n673 & ~n778 ;
  assign n780 = n160 & ~n779 ;
  assign n781 = ~n777 & ~n780 ;
  assign n785 = \timebase_reg[0]/NET0131  & ~n684 ;
  assign n782 = \timebase_reg[0]/NET0131  & ~n445 ;
  assign n783 = ~n766 & ~n782 ;
  assign n784 = n160 & ~n783 ;
  assign n786 = \timebase_reg[0]/NET0131  & ~n686 ;
  assign n787 = ~n229 & ~n786 ;
  assign n788 = ~n784 & n787 ;
  assign n789 = ~n785 & n788 ;
  assign n790 = \max_reg[2]/NET0131  & ~n600 ;
  assign n794 = ~\max_reg[2]/NET0131  & ~n317 ;
  assign n791 = ~\max_reg[2]/NET0131  & ~n269 ;
  assign n792 = ~n270 & ~n791 ;
  assign n793 = n317 & ~n792 ;
  assign n795 = n166 & ~n793 ;
  assign n796 = ~n794 & n795 ;
  assign n798 = ~\max_reg[2]/NET0131  & n146 ;
  assign n797 = ~n146 & ~n792 ;
  assign n799 = n295 & ~n797 ;
  assign n800 = ~n798 & n799 ;
  assign n801 = ~n796 & ~n800 ;
  assign n802 = ~n790 & n801 ;
  assign n803 = \max_reg[0]/NET0131  & ~n600 ;
  assign n804 = ~\max_reg[0]/NET0131  & ~n146 ;
  assign n805 = \max_reg[0]/NET0131  & n146 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = ~n360 & ~n806 ;
  assign n808 = n166 & ~n807 ;
  assign n809 = n295 & ~n806 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = ~n803 & n810 ;
  assign n812 = \max_reg[1]/NET0131  & ~n600 ;
  assign n816 = ~\max_reg[1]/NET0131  & ~n317 ;
  assign n813 = ~\max_reg[0]/NET0131  & ~\max_reg[1]/NET0131  ;
  assign n814 = ~n269 & ~n813 ;
  assign n815 = n317 & ~n814 ;
  assign n817 = n166 & ~n815 ;
  assign n818 = ~n816 & n817 ;
  assign n820 = ~\max_reg[1]/NET0131  & n146 ;
  assign n819 = ~n146 & ~n814 ;
  assign n821 = n295 & ~n819 ;
  assign n822 = ~n820 & n821 ;
  assign n823 = ~n818 & ~n822 ;
  assign n824 = ~n812 & n823 ;
  assign n825 = n146 & n166 ;
  assign n826 = ~n284 & ~n825 ;
  assign n827 = n210 & n826 ;
  assign n828 = \scan_reg[0]/NET0131  & ~n827 ;
  assign n829 = ~n160 & ~n216 ;
  assign n830 = ~\scan_reg[0]/NET0131  & ~n829 ;
  assign n831 = n213 & n830 ;
  assign n832 = ~n828 & ~n831 ;
  assign n840 = \scan_reg[2]/NET0131  & ~n210 ;
  assign n834 = ~\scan_reg[2]/NET0131  & ~n148 ;
  assign n835 = ~n722 & ~n834 ;
  assign n836 = ~n146 & n835 ;
  assign n837 = n165 & ~n836 ;
  assign n833 = ~\scan_reg[2]/NET0131  & ~n165 ;
  assign n838 = n216 & ~n833 ;
  assign n839 = ~n837 & n838 ;
  assign n841 = \scan_reg[2]/NET0131  & n146 ;
  assign n842 = ~n836 & ~n841 ;
  assign n843 = n166 & ~n842 ;
  assign n844 = ~n839 & ~n843 ;
  assign n845 = ~n840 & n844 ;
  assign n846 = n165 & ~n320 ;
  assign n847 = ~n171 & ~n236 ;
  assign n848 = ~n846 & n847 ;
  assign n849 = ~n464 & n848 ;
  assign n850 = ~n229 & n482 ;
  assign n851 = \ind_reg[0]/NET0131  & ~n850 ;
  assign n853 = ~\ind_reg[0]/NET0131  & ~\k[3]_pad  ;
  assign n854 = n331 & ~n853 ;
  assign n855 = ~n165 & n854 ;
  assign n852 = \ind_reg[0]/NET0131  & n165 ;
  assign n856 = ~n337 & ~n852 ;
  assign n857 = ~n855 & n856 ;
  assign n858 = n203 & ~n857 ;
  assign n859 = ~n851 & ~n858 ;
  assign n860 = \ind_reg[1]/NET0131  & ~n850 ;
  assign n861 = ~\ind_reg[1]/NET0131  & ~n452 ;
  assign n862 = n454 & ~n861 ;
  assign n863 = ~n860 & ~n862 ;
  assign n878 = ~\sound_reg[1]/NET0131  & ~\sound_reg[2]/NET0131  ;
  assign n864 = ~\sound_reg[1]/NET0131  & \sound_reg[2]/NET0131  ;
  assign n875 = \sound_reg[1]/NET0131  & ~\sound_reg[2]/NET0131  ;
  assign n893 = ~n864 & ~n875 ;
  assign n894 = ~n878 & n893 ;
  assign n884 = ~\sound_reg[0]/NET0131  & n878 ;
  assign n885 = \counter_reg[0]/NET0131  & \counter_reg[1]/NET0131  ;
  assign n886 = ~\counter_reg[2]/NET0131  & ~n885 ;
  assign n895 = n884 & n886 ;
  assign n888 = ~\sound_reg[0]/NET0131  & n864 ;
  assign n889 = \counter_reg[2]/NET0131  & n885 ;
  assign n896 = n888 & ~n889 ;
  assign n897 = ~n895 & ~n896 ;
  assign n898 = ~n894 & n897 ;
  assign n899 = speaker_pad & ~n898 ;
  assign n871 = \counter_reg[1]/NET0131  & \counter_reg[2]/NET0131  ;
  assign n872 = speaker_pad & ~n871 ;
  assign n873 = ~\s_reg/NET0131  & n871 ;
  assign n874 = ~n872 & ~n873 ;
  assign n876 = \sound_reg[0]/NET0131  & n875 ;
  assign n877 = ~n874 & n876 ;
  assign n865 = \sound_reg[0]/NET0131  & n864 ;
  assign n866 = ~\counter_reg[1]/NET0131  & ~\counter_reg[2]/NET0131  ;
  assign n867 = ~\s_reg/NET0131  & ~n866 ;
  assign n868 = speaker_pad & n866 ;
  assign n869 = ~n867 & ~n868 ;
  assign n870 = n865 & ~n869 ;
  assign n879 = \sound_reg[0]/NET0131  & n878 ;
  assign n880 = ~\counter_reg[2]/NET0131  & speaker_pad ;
  assign n881 = \counter_reg[2]/NET0131  & ~\s_reg/NET0131  ;
  assign n882 = ~n880 & ~n881 ;
  assign n883 = n879 & ~n882 ;
  assign n907 = ~n870 & ~n883 ;
  assign n908 = ~n877 & n907 ;
  assign n887 = n884 & ~n886 ;
  assign n890 = n888 & n889 ;
  assign n891 = ~n887 & ~n890 ;
  assign n892 = ~\s_reg/NET0131  & ~n891 ;
  assign n900 = ~\sound_reg[0]/NET0131  & n875 ;
  assign n901 = ~\counter_reg[0]/NET0131  & ~\counter_reg[1]/NET0131  ;
  assign n902 = \counter_reg[2]/NET0131  & ~n901 ;
  assign n903 = speaker_pad & ~n902 ;
  assign n904 = n881 & ~n901 ;
  assign n905 = ~n903 & ~n904 ;
  assign n906 = n900 & ~n905 ;
  assign n909 = ~n892 & ~n906 ;
  assign n910 = n908 & n909 ;
  assign n911 = ~n899 & n910 ;
  assign n912 = \play_reg/NET0131  & ~n911 ;
  assign n913 = ~n203 & n474 ;
  assign n914 = n480 & n913 ;
  assign n915 = \wr_reg/NET0131  & ~n914 ;
  assign n916 = ~n225 & ~n915 ;
  assign n924 = n900 & ~n902 ;
  assign n925 = n865 & n866 ;
  assign n926 = ~n924 & ~n925 ;
  assign n927 = n897 & n926 ;
  assign n928 = \s_reg/NET0131  & ~n894 ;
  assign n929 = n927 & n928 ;
  assign n930 = n885 & n888 ;
  assign n931 = n900 & ~n901 ;
  assign n932 = ~n930 & ~n931 ;
  assign n933 = \counter_reg[2]/NET0131  & ~n932 ;
  assign n934 = ~\s_reg/NET0131  & ~n887 ;
  assign n935 = ~n933 & n934 ;
  assign n936 = ~n929 & ~n935 ;
  assign n921 = \s_reg/NET0131  & ~n871 ;
  assign n922 = ~n873 & ~n921 ;
  assign n923 = n876 & ~n922 ;
  assign n917 = n865 & n867 ;
  assign n918 = ~\counter_reg[2]/NET0131  & \s_reg/NET0131  ;
  assign n919 = ~n881 & ~n918 ;
  assign n920 = n879 & ~n919 ;
  assign n937 = ~n917 & ~n920 ;
  assign n938 = ~n923 & n937 ;
  assign n939 = ~n936 & n938 ;
  assign n940 = \count_reg[0]/NET0131  & n225 ;
  assign n941 = n174 & n233 ;
  assign n942 = n278 & n625 ;
  assign n943 = n941 & n942 ;
  assign n944 = n199 & n243 ;
  assign n945 = n943 & n944 ;
  assign n946 = n680 & n945 ;
  assign n947 = \data_in_reg[0]/NET0131  & ~n946 ;
  assign n948 = ~n940 & ~n947 ;
  assign n949 = \count_reg[1]/NET0131  & n225 ;
  assign n950 = \data_in_reg[1]/NET0131  & ~n946 ;
  assign n951 = ~n949 & ~n950 ;
  assign n954 = \address_reg[2]/NET0131  & ~n259 ;
  assign n952 = \scan_reg[2]/NET0131  & ~n222 ;
  assign n953 = \max_reg[2]/NET0131  & ~n226 ;
  assign n955 = ~n952 & ~n953 ;
  assign n956 = ~n954 & n955 ;
  assign n959 = \address_reg[3]/NET0131  & ~n259 ;
  assign n957 = \scan_reg[3]/NET0131  & ~n222 ;
  assign n958 = \max_reg[3]/NET0131  & ~n226 ;
  assign n960 = ~n957 & ~n958 ;
  assign n961 = ~n959 & n960 ;
  assign n964 = \address_reg[4]/NET0131  & ~n259 ;
  assign n962 = \scan_reg[4]/NET0131  & ~n222 ;
  assign n963 = \max_reg[4]/NET0131  & ~n226 ;
  assign n965 = ~n962 & ~n963 ;
  assign n966 = ~n964 & n965 ;
  assign n969 = \address_reg[1]/NET0131  & ~n259 ;
  assign n967 = \scan_reg[1]/NET0131  & ~n222 ;
  assign n968 = \max_reg[1]/NET0131  & ~n226 ;
  assign n970 = ~n967 & ~n968 ;
  assign n971 = ~n969 & n970 ;
  assign n972 = ~\counter_reg[2]/NET0131  & n879 ;
  assign n973 = ~n876 & ~n972 ;
  assign n974 = ~n871 & ~n973 ;
  assign n975 = n927 & ~n974 ;
  assign n976 = \play_reg/NET0131  & ~n975 ;
  assign n977 = ~n886 & ~n889 ;
  assign n978 = n976 & n977 ;
  assign n979 = ~n885 & ~n901 ;
  assign n980 = n976 & n979 ;
  assign n981 = ~\counter_reg[0]/NET0131  & n976 ;
  assign n986 = ~\address_reg[2]/NET0131  & \address_reg[3]/NET0131  ;
  assign n990 = \address_reg[1]/NET0131  & ~\address_reg[4]/NET0131  ;
  assign n1008 = n986 & n990 ;
  assign n1009 = \memory_reg[10][0]/NET0131  & n1008 ;
  assign n983 = ~\address_reg[1]/NET0131  & \address_reg[4]/NET0131  ;
  assign n1002 = \address_reg[2]/NET0131  & \address_reg[3]/NET0131  ;
  assign n1003 = n983 & n1002 ;
  assign n1004 = \memory_reg[28][0]/NET0131  & n1003 ;
  assign n1005 = \address_reg[1]/NET0131  & \address_reg[4]/NET0131  ;
  assign n1006 = n986 & n1005 ;
  assign n1007 = \memory_reg[26][0]/NET0131  & n1006 ;
  assign n1014 = ~n1004 & ~n1007 ;
  assign n1015 = ~n1009 & n1014 ;
  assign n993 = ~\address_reg[2]/NET0131  & ~\address_reg[3]/NET0131  ;
  assign n994 = n990 & n993 ;
  assign n995 = \memory_reg[2][0]/NET0131  & n994 ;
  assign n996 = n983 & n986 ;
  assign n997 = \memory_reg[24][0]/NET0131  & n996 ;
  assign n1012 = ~n995 & ~n997 ;
  assign n982 = \address_reg[2]/NET0131  & ~\address_reg[3]/NET0131  ;
  assign n987 = ~\address_reg[1]/NET0131  & ~\address_reg[4]/NET0131  ;
  assign n998 = n982 & n987 ;
  assign n999 = \memory_reg[4][0]/NET0131  & n998 ;
  assign n1000 = n983 & n993 ;
  assign n1001 = \memory_reg[16][0]/NET0131  & n1000 ;
  assign n1013 = ~n999 & ~n1001 ;
  assign n1016 = n1012 & n1013 ;
  assign n984 = n982 & n983 ;
  assign n985 = \memory_reg[20][0]/NET0131  & n984 ;
  assign n1010 = ~\address_reg[0]/NET0131  & ~n985 ;
  assign n988 = n986 & n987 ;
  assign n989 = \memory_reg[8][0]/NET0131  & n988 ;
  assign n991 = n982 & n990 ;
  assign n992 = \memory_reg[6][0]/NET0131  & n991 ;
  assign n1011 = ~n989 & ~n992 ;
  assign n1017 = n1010 & n1011 ;
  assign n1018 = n1016 & n1017 ;
  assign n1019 = n1015 & n1018 ;
  assign n1029 = \memory_reg[27][0]/NET0131  & n1006 ;
  assign n1026 = n993 & n1005 ;
  assign n1027 = \memory_reg[19][0]/NET0131  & n1026 ;
  assign n1028 = \memory_reg[17][0]/NET0131  & n1000 ;
  assign n1033 = ~n1027 & ~n1028 ;
  assign n1034 = ~n1029 & n1033 ;
  assign n1020 = n990 & n1002 ;
  assign n1021 = \memory_reg[15][0]/NET0131  & n1020 ;
  assign n1030 = \address_reg[0]/NET0131  & ~n1021 ;
  assign n1022 = \memory_reg[5][0]/NET0131  & n998 ;
  assign n1023 = \memory_reg[9][0]/NET0131  & n988 ;
  assign n1031 = ~n1022 & ~n1023 ;
  assign n1024 = \memory_reg[21][0]/NET0131  & n984 ;
  assign n1025 = \memory_reg[25][0]/NET0131  & n996 ;
  assign n1032 = ~n1024 & ~n1025 ;
  assign n1035 = n1031 & n1032 ;
  assign n1036 = n1030 & n1035 ;
  assign n1037 = n1034 & n1036 ;
  assign n1038 = ~n1019 & ~n1037 ;
  assign n1057 = \memory_reg[14][0]/NET0131  & n1020 ;
  assign n1056 = \memory_reg[18][0]/NET0131  & n1026 ;
  assign n1058 = ~\address_reg[0]/NET0131  & ~n1056 ;
  assign n1059 = ~n1057 & n1058 ;
  assign n1061 = \memory_reg[11][0]/NET0131  & n1008 ;
  assign n1060 = \memory_reg[3][0]/NET0131  & n994 ;
  assign n1062 = \address_reg[0]/NET0131  & ~n1060 ;
  assign n1063 = ~n1061 & n1062 ;
  assign n1064 = ~n1059 & ~n1063 ;
  assign n1069 = n987 & n993 ;
  assign n1070 = ~\address_reg[0]/NET0131  & ~\memory_reg[0][0]/NET0131  ;
  assign n1071 = \address_reg[0]/NET0131  & ~\memory_reg[1][0]/NET0131  ;
  assign n1072 = ~n1070 & ~n1071 ;
  assign n1073 = n1069 & n1072 ;
  assign n1051 = n987 & n1002 ;
  assign n1052 = ~\address_reg[0]/NET0131  & ~\memory_reg[12][0]/NET0131  ;
  assign n1053 = \address_reg[0]/NET0131  & ~\memory_reg[13][0]/NET0131  ;
  assign n1054 = ~n1052 & ~n1053 ;
  assign n1055 = n1051 & n1054 ;
  assign n1065 = \address_reg[0]/NET0131  & ~\address_reg[3]/NET0131  ;
  assign n1066 = \address_reg[2]/NET0131  & n1065 ;
  assign n1067 = \memory_reg[7][0]/NET0131  & n990 ;
  assign n1068 = n1066 & n1067 ;
  assign n1075 = ~n1055 & ~n1068 ;
  assign n1076 = ~n1073 & n1075 ;
  assign n1039 = \address_reg[0]/NET0131  & n1003 ;
  assign n1040 = \memory_reg[29][0]/NET0131  & n1039 ;
  assign n1041 = n982 & n1005 ;
  assign n1042 = ~\address_reg[0]/NET0131  & ~\memory_reg[22][0]/NET0131  ;
  assign n1043 = \address_reg[0]/NET0131  & ~\memory_reg[23][0]/NET0131  ;
  assign n1044 = ~n1042 & ~n1043 ;
  assign n1045 = n1041 & n1044 ;
  assign n1046 = n1002 & n1005 ;
  assign n1047 = ~\address_reg[0]/NET0131  & ~\memory_reg[30][0]/NET0131  ;
  assign n1048 = \address_reg[0]/NET0131  & ~\memory_reg[31][0]/NET0131  ;
  assign n1049 = ~n1047 & ~n1048 ;
  assign n1050 = n1046 & n1049 ;
  assign n1074 = ~n1045 & ~n1050 ;
  assign n1077 = ~n1040 & n1074 ;
  assign n1078 = n1076 & n1077 ;
  assign n1079 = ~n1064 & n1078 ;
  assign n1080 = ~n1038 & n1079 ;
  assign n1128 = \memory_reg[17][1]/NET0131  & n1000 ;
  assign n1132 = \address_reg[0]/NET0131  & ~n1128 ;
  assign n1131 = \memory_reg[5][1]/NET0131  & n998 ;
  assign n1129 = \memory_reg[1][1]/NET0131  & n1069 ;
  assign n1130 = \memory_reg[15][1]/NET0131  & n1020 ;
  assign n1133 = ~n1129 & ~n1130 ;
  assign n1134 = ~n1131 & n1133 ;
  assign n1135 = n1132 & n1134 ;
  assign n1136 = \memory_reg[12][1]/NET0131  & n1051 ;
  assign n1141 = ~\address_reg[0]/NET0131  & ~n1136 ;
  assign n1137 = \memory_reg[28][1]/NET0131  & n1003 ;
  assign n1138 = \memory_reg[20][1]/NET0131  & n984 ;
  assign n1142 = ~n1137 & ~n1138 ;
  assign n1139 = \memory_reg[26][1]/NET0131  & n1006 ;
  assign n1140 = \memory_reg[24][1]/NET0131  & n996 ;
  assign n1143 = ~n1139 & ~n1140 ;
  assign n1144 = n1142 & n1143 ;
  assign n1145 = n1141 & n1144 ;
  assign n1146 = ~n1135 & ~n1145 ;
  assign n1086 = \memory_reg[4][1]/NET0131  & n998 ;
  assign n1084 = \memory_reg[8][1]/NET0131  & n988 ;
  assign n1085 = \memory_reg[16][1]/NET0131  & n1000 ;
  assign n1089 = ~n1084 & ~n1085 ;
  assign n1090 = ~n1086 & n1089 ;
  assign n1081 = \memory_reg[14][1]/NET0131  & n1020 ;
  assign n1087 = ~\address_reg[0]/NET0131  & ~n1081 ;
  assign n1082 = \memory_reg[2][1]/NET0131  & n994 ;
  assign n1083 = \memory_reg[6][1]/NET0131  & n991 ;
  assign n1088 = ~n1082 & ~n1083 ;
  assign n1091 = n1087 & n1088 ;
  assign n1092 = n1090 & n1091 ;
  assign n1098 = \memory_reg[9][1]/NET0131  & n988 ;
  assign n1096 = \memory_reg[13][1]/NET0131  & n1051 ;
  assign n1097 = \memory_reg[25][1]/NET0131  & n996 ;
  assign n1101 = ~n1096 & ~n1097 ;
  assign n1102 = ~n1098 & n1101 ;
  assign n1093 = \memory_reg[27][1]/NET0131  & n1006 ;
  assign n1099 = \address_reg[0]/NET0131  & ~n1093 ;
  assign n1094 = \memory_reg[19][1]/NET0131  & n1026 ;
  assign n1095 = \memory_reg[3][1]/NET0131  & n994 ;
  assign n1100 = ~n1094 & ~n1095 ;
  assign n1103 = n1099 & n1100 ;
  assign n1104 = n1102 & n1103 ;
  assign n1105 = ~n1092 & ~n1104 ;
  assign n1108 = \memory_reg[18][1]/NET0131  & n1026 ;
  assign n1107 = \memory_reg[0][1]/NET0131  & n1069 ;
  assign n1109 = ~\address_reg[0]/NET0131  & ~n1107 ;
  assign n1110 = ~n1108 & n1109 ;
  assign n1112 = \memory_reg[7][1]/NET0131  & n991 ;
  assign n1111 = \memory_reg[21][1]/NET0131  & n984 ;
  assign n1113 = \address_reg[0]/NET0131  & ~n1111 ;
  assign n1114 = ~n1112 & n1113 ;
  assign n1115 = ~n1110 & ~n1114 ;
  assign n1106 = \memory_reg[29][1]/NET0131  & n1039 ;
  assign n1124 = ~\address_reg[0]/NET0131  & ~\memory_reg[10][1]/NET0131  ;
  assign n1125 = \address_reg[0]/NET0131  & ~\memory_reg[11][1]/NET0131  ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = n1008 & n1126 ;
  assign n1116 = ~\address_reg[0]/NET0131  & ~\memory_reg[22][1]/NET0131  ;
  assign n1117 = \address_reg[0]/NET0131  & ~\memory_reg[23][1]/NET0131  ;
  assign n1118 = ~n1116 & ~n1117 ;
  assign n1119 = n1041 & n1118 ;
  assign n1120 = ~\address_reg[0]/NET0131  & ~\memory_reg[30][1]/NET0131  ;
  assign n1121 = \address_reg[0]/NET0131  & ~\memory_reg[31][1]/NET0131  ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = n1046 & n1122 ;
  assign n1147 = ~n1119 & ~n1123 ;
  assign n1148 = ~n1127 & n1147 ;
  assign n1149 = ~n1106 & n1148 ;
  assign n1150 = ~n1115 & n1149 ;
  assign n1151 = ~n1105 & n1150 ;
  assign n1152 = ~n1146 & n1151 ;
  assign n1153 = ~\address_reg[0]/NET0131  & ~\address_reg[3]/NET0131  ;
  assign n1154 = ~\address_reg[2]/NET0131  & n1153 ;
  assign n1155 = \wr_reg/NET0131  & n987 ;
  assign n1156 = n1154 & n1155 ;
  assign n1157 = ~\address_reg[0]/NET0131  & \address_reg[3]/NET0131  ;
  assign n1158 = ~\address_reg[2]/NET0131  & n1157 ;
  assign n1159 = \wr_reg/NET0131  & n990 ;
  assign n1160 = n1158 & n1159 ;
  assign n1161 = \address_reg[0]/NET0131  & \address_reg[3]/NET0131  ;
  assign n1162 = ~\address_reg[2]/NET0131  & n1161 ;
  assign n1163 = n1159 & n1162 ;
  assign n1164 = \address_reg[2]/NET0131  & n1157 ;
  assign n1165 = n1155 & n1164 ;
  assign n1166 = \address_reg[2]/NET0131  & n1161 ;
  assign n1167 = n1155 & n1166 ;
  assign n1168 = n1159 & n1164 ;
  assign n1169 = n1159 & n1166 ;
  assign n1170 = \wr_reg/NET0131  & n983 ;
  assign n1171 = n1154 & n1170 ;
  assign n1172 = ~\address_reg[2]/NET0131  & n1065 ;
  assign n1173 = n1170 & n1172 ;
  assign n1174 = \wr_reg/NET0131  & n1005 ;
  assign n1175 = n1154 & n1174 ;
  assign n1176 = n1172 & n1174 ;
  assign n1177 = n1155 & n1172 ;
  assign n1178 = \address_reg[2]/NET0131  & n1153 ;
  assign n1179 = n1170 & n1178 ;
  assign n1180 = n1066 & n1170 ;
  assign n1181 = n1174 & n1178 ;
  assign n1182 = n1066 & n1174 ;
  assign n1183 = n1158 & n1170 ;
  assign n1184 = n1162 & n1170 ;
  assign n1185 = n1158 & n1174 ;
  assign n1186 = n1162 & n1174 ;
  assign n1187 = n1164 & n1170 ;
  assign n1188 = \wr_reg/NET0131  & n1039 ;
  assign n1189 = n1154 & n1159 ;
  assign n1190 = n1164 & n1174 ;
  assign n1191 = n1166 & n1174 ;
  assign n1192 = n1159 & n1172 ;
  assign n1193 = n1155 & n1178 ;
  assign n1194 = n1066 & n1155 ;
  assign n1195 = n1159 & n1178 ;
  assign n1196 = n1066 & n1159 ;
  assign n1197 = n1155 & n1158 ;
  assign n1198 = n1155 & n1162 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \count_reg[0]/P0001  = ~\count_reg[0]/NET0131  ;
  assign \g10376/_0_  = ~n127 ;
  assign \g11078/_0_  = ~n219 ;
  assign \g11102/_0_  = ~n262 ;
  assign \g11126/_0_  = ~n315 ;
  assign \g11156/_0_  = ~n330 ;
  assign \g11299/_0_  = ~n372 ;
  assign \g11308/_0_  = ~n398 ;
  assign \g11318/_0_  = ~n414 ;
  assign \g11346/_0_  = ~n442 ;
  assign \g11378/_0_  = ~n451 ;
  assign \g11516/_0_  = ~n472 ;
  assign \g63/_0_  = ~n500 ;
  assign \g8501/_0_  = ~n525 ;
  assign \g8516/_0_  = ~n534 ;
  assign \g8517/_0_  = ~n551 ;
  assign \g8519/_0_  = ~n572 ;
  assign \g8520/_0_  = ~n585 ;
  assign \g8522/_0_  = ~n611 ;
  assign \g8526/_0_  = ~n634 ;
  assign \g8529/_2_  = ~n653 ;
  assign \g8545/_0_  = ~n667 ;
  assign \g8546/_0_  = ~n690 ;
  assign \g8547/_0_  = ~n702 ;
  assign \g8555/_0_  = ~n708 ;
  assign \g8556/_0_  = ~n720 ;
  assign \g8557/_0_  = ~n734 ;
  assign \g8558/_0_  = ~n747 ;
  assign \g8559/_0_  = ~n764 ;
  assign \g8560/_0_  = ~n771 ;
  assign \g8562/_0_  = ~n776 ;
  assign \g8563/_0_  = ~n781 ;
  assign \g8581/_0_  = ~n789 ;
  assign \g8586/_0_  = ~n802 ;
  assign \g8591/_0_  = ~n811 ;
  assign \g8594/_0_  = ~n824 ;
  assign \g8606/_0_  = ~n832 ;
  assign \g8608/_0_  = ~n845 ;
  assign \g8647/_0_  = ~n849 ;
  assign \g8659/_0_  = ~n859 ;
  assign \g8695/_0_  = ~n863 ;
  assign \g8784/_0_  = n912 ;
  assign \g8797/_0_  = ~n916 ;
  assign \g8854/_2_  = ~n939 ;
  assign \g8869/_0_  = ~n948 ;
  assign \g8871/_0_  = ~n951 ;
  assign \g8889/_0_  = ~n956 ;
  assign \g8891/_0_  = ~n961 ;
  assign \g8892/_0_  = ~n966 ;
  assign \g8894/_0_  = ~n971 ;
  assign \g8970/_0_  = n978 ;
  assign \g8975/_0_  = n980 ;
  assign \g8992/_0_  = n981 ;
  assign \g9180/_0_  = ~n1080 ;
  assign \g9183/_0_  = ~n1152 ;
  assign \g9511/u3_syn_4  = n1156 ;
  assign \g9513/u3_syn_4  = n1160 ;
  assign \g9515/u3_syn_4  = n1163 ;
  assign \g9517/u3_syn_4  = n1165 ;
  assign \g9519/u3_syn_4  = n1167 ;
  assign \g9521/u3_syn_4  = n1168 ;
  assign \g9523/u3_syn_4  = n1169 ;
  assign \g9525/u3_syn_4  = n1171 ;
  assign \g9527/u3_syn_4  = n1173 ;
  assign \g9529/u3_syn_4  = n1175 ;
  assign \g9531/u3_syn_4  = n1176 ;
  assign \g9533/u3_syn_4  = n1177 ;
  assign \g9535/u3_syn_4  = n1179 ;
  assign \g9537/u3_syn_4  = n1180 ;
  assign \g9539/u3_syn_4  = n1181 ;
  assign \g9541/u3_syn_4  = n1182 ;
  assign \g9543/u3_syn_4  = n1183 ;
  assign \g9545/u3_syn_4  = n1184 ;
  assign \g9547/u3_syn_4  = n1185 ;
  assign \g9549/u3_syn_4  = n1186 ;
  assign \g9551/u3_syn_4  = n1187 ;
  assign \g9553/u3_syn_4  = n1188 ;
  assign \g9555/u3_syn_4  = n1189 ;
  assign \g9557/u3_syn_4  = n1190 ;
  assign \g9559/u3_syn_4  = n1191 ;
  assign \g9560/u3_syn_4  = n1192 ;
  assign \g9562/u3_syn_4  = n1193 ;
  assign \g9564/u3_syn_4  = n1194 ;
  assign \g9566/u3_syn_4  = n1195 ;
  assign \g9568/u3_syn_4  = n1196 ;
  assign \g9570/u3_syn_4  = n1197 ;
  assign \g9572/u3_syn_4  = n1198 ;
endmodule
