module top (\data_i[0]_pad , \data_i[10]_pad , \data_i[11]_pad , \data_i[12]_pad , \data_i[13]_pad , \data_i[14]_pad , \data_i[15]_pad , \data_i[16]_pad , \data_i[17]_pad , \data_i[18]_pad , \data_i[19]_pad , \data_i[1]_pad , \data_i[20]_pad , \data_i[21]_pad , \data_i[22]_pad , \data_i[23]_pad , \data_i[24]_pad , \data_i[25]_pad , \data_i[26]_pad , \data_i[27]_pad , \data_i[28]_pad , \data_i[29]_pad , \data_i[2]_pad , \data_i[30]_pad , \data_i[31]_pad , \data_i[32]_pad , \data_i[33]_pad , \data_i[34]_pad , \data_i[35]_pad , \data_i[36]_pad , \data_i[37]_pad , \data_i[38]_pad , \data_i[39]_pad , \data_i[3]_pad , \data_i[40]_pad , \data_i[41]_pad , \data_i[42]_pad , \data_i[43]_pad , \data_i[44]_pad , \data_i[45]_pad , \data_i[46]_pad , \data_i[47]_pad , \data_i[48]_pad , \data_i[49]_pad , \data_i[4]_pad , \data_i[50]_pad , \data_i[51]_pad , \data_i[52]_pad , \data_i[53]_pad , \data_i[54]_pad , \data_i[55]_pad , \data_i[56]_pad , \data_i[57]_pad , \data_i[58]_pad , \data_i[59]_pad , \data_i[5]_pad , \data_i[60]_pad , \data_i[61]_pad , \data_i[62]_pad , \data_i[63]_pad , \data_i[6]_pad , \data_i[7]_pad , \data_i[8]_pad , \data_i[9]_pad , \data_ready_reg/NET0131 , decrypt_i_pad, \key_i[10]_pad , \key_i[11]_pad , \key_i[12]_pad , \key_i[13]_pad , \key_i[14]_pad , \key_i[15]_pad , \key_i[17]_pad , \key_i[18]_pad , \key_i[19]_pad , \key_i[1]_pad , \key_i[20]_pad , \key_i[21]_pad , \key_i[22]_pad , \key_i[23]_pad , \key_i[25]_pad , \key_i[26]_pad , \key_i[27]_pad , \key_i[28]_pad , \key_i[29]_pad , \key_i[2]_pad , \key_i[30]_pad , \key_i[31]_pad , \key_i[33]_pad , \key_i[34]_pad , \key_i[35]_pad , \key_i[36]_pad , \key_i[37]_pad , \key_i[38]_pad , \key_i[39]_pad , \key_i[3]_pad , \key_i[41]_pad , \key_i[42]_pad , \key_i[43]_pad , \key_i[44]_pad , \key_i[45]_pad , \key_i[46]_pad , \key_i[47]_pad , \key_i[49]_pad , \key_i[4]_pad , \key_i[50]_pad , \key_i[51]_pad , \key_i[52]_pad , \key_i[53]_pad , \key_i[54]_pad , \key_i[55]_pad , \key_i[57]_pad , \key_i[58]_pad , \key_i[59]_pad , \key_i[5]_pad , \key_i[60]_pad , \key_i[61]_pad , \key_i[62]_pad , \key_i[63]_pad , \key_i[6]_pad , \key_i[7]_pad , \key_i[9]_pad , load_i_pad, \rd1_Key_o_reg[0]/NET0131 , \rd1_Key_o_reg[10]/NET0131 , \rd1_Key_o_reg[11]/NET0131 , \rd1_Key_o_reg[12]/NET0131 , \rd1_Key_o_reg[13]/NET0131 , \rd1_Key_o_reg[14]/NET0131 , \rd1_Key_o_reg[15]/NET0131 , \rd1_Key_o_reg[16]/NET0131 , \rd1_Key_o_reg[17]/NET0131 , \rd1_Key_o_reg[18]/NET0131 , \rd1_Key_o_reg[19]/NET0131 , \rd1_Key_o_reg[1]/NET0131 , \rd1_Key_o_reg[20]/NET0131 , \rd1_Key_o_reg[21]/NET0131 , \rd1_Key_o_reg[22]/NET0131 , \rd1_Key_o_reg[23]/NET0131 , \rd1_Key_o_reg[24]/NET0131 , \rd1_Key_o_reg[25]/NET0131 , \rd1_Key_o_reg[26]/NET0131 , \rd1_Key_o_reg[27]/NET0131 , \rd1_Key_o_reg[28]/NET0131 , \rd1_Key_o_reg[29]/NET0131 , \rd1_Key_o_reg[2]/NET0131 , \rd1_Key_o_reg[30]/NET0131 , \rd1_Key_o_reg[31]/NET0131 , \rd1_Key_o_reg[32]/NET0131 , \rd1_Key_o_reg[33]/NET0131 , \rd1_Key_o_reg[34]/NET0131 , \rd1_Key_o_reg[35]/NET0131 , \rd1_Key_o_reg[36]/NET0131 , \rd1_Key_o_reg[37]/NET0131 , \rd1_Key_o_reg[38]/NET0131 , \rd1_Key_o_reg[39]/NET0131 , \rd1_Key_o_reg[3]/NET0131 , \rd1_Key_o_reg[40]/NET0131 , \rd1_Key_o_reg[41]/NET0131 , \rd1_Key_o_reg[42]/NET0131 , \rd1_Key_o_reg[43]/NET0131 , \rd1_Key_o_reg[44]/NET0131 , \rd1_Key_o_reg[45]/NET0131 , \rd1_Key_o_reg[46]/NET0131 , \rd1_Key_o_reg[47]/NET0131 , \rd1_Key_o_reg[48]/NET0131 , \rd1_Key_o_reg[49]/NET0131 , \rd1_Key_o_reg[4]/NET0131 , \rd1_Key_o_reg[50]/NET0131 , \rd1_Key_o_reg[51]/NET0131 , \rd1_Key_o_reg[52]/NET0131 , \rd1_Key_o_reg[53]/NET0131 , \rd1_Key_o_reg[54]/NET0131 , \rd1_Key_o_reg[55]/NET0131 , \rd1_Key_o_reg[5]/NET0131 , \rd1_Key_o_reg[6]/NET0131 , \rd1_Key_o_reg[7]/NET0131 , \rd1_Key_o_reg[8]/NET0131 , \rd1_Key_o_reg[9]/NET0131 , \rd1_L_o_reg[0]/NET0131 , \rd1_L_o_reg[10]/NET0131 , \rd1_L_o_reg[11]/NET0131 , \rd1_L_o_reg[12]/NET0131 , \rd1_L_o_reg[13]/NET0131 , \rd1_L_o_reg[14]/NET0131 , \rd1_L_o_reg[15]/NET0131 , \rd1_L_o_reg[16]/NET0131 , \rd1_L_o_reg[17]/NET0131 , \rd1_L_o_reg[18]/NET0131 , \rd1_L_o_reg[19]/NET0131 , \rd1_L_o_reg[1]/NET0131 , \rd1_L_o_reg[20]/NET0131 , \rd1_L_o_reg[21]/NET0131 , \rd1_L_o_reg[22]/NET0131 , \rd1_L_o_reg[23]/NET0131 , \rd1_L_o_reg[24]/NET0131 , \rd1_L_o_reg[25]/NET0131 , \rd1_L_o_reg[26]/NET0131 , \rd1_L_o_reg[27]/NET0131 , \rd1_L_o_reg[28]/NET0131 , \rd1_L_o_reg[29]/NET0131 , \rd1_L_o_reg[2]/NET0131 , \rd1_L_o_reg[30]/NET0131 , \rd1_L_o_reg[31]/NET0131 , \rd1_L_o_reg[3]/NET0131 , \rd1_L_o_reg[4]/NET0131 , \rd1_L_o_reg[5]/NET0131 , \rd1_L_o_reg[6]/NET0131 , \rd1_L_o_reg[7]/NET0131 , \rd1_L_o_reg[8]/NET0131 , \rd1_L_o_reg[9]/NET0131 , \rd1_R_o_reg[0]/NET0131 , \rd1_R_o_reg[10]/NET0131 , \rd1_R_o_reg[11]/NET0131 , \rd1_R_o_reg[12]/NET0131 , \rd1_R_o_reg[13]/NET0131 , \rd1_R_o_reg[14]/NET0131 , \rd1_R_o_reg[15]/NET0131 , \rd1_R_o_reg[16]/NET0131 , \rd1_R_o_reg[17]/NET0131 , \rd1_R_o_reg[18]/NET0131 , \rd1_R_o_reg[19]/NET0131 , \rd1_R_o_reg[1]/NET0131 , \rd1_R_o_reg[20]/NET0131 , \rd1_R_o_reg[21]/NET0131 , \rd1_R_o_reg[22]/NET0131 , \rd1_R_o_reg[23]/NET0131 , \rd1_R_o_reg[24]/NET0131 , \rd1_R_o_reg[25]/NET0131 , \rd1_R_o_reg[26]/NET0131 , \rd1_R_o_reg[27]/NET0131 , \rd1_R_o_reg[28]/NET0131 , \rd1_R_o_reg[29]/NET0131 , \rd1_R_o_reg[2]/NET0131 , \rd1_R_o_reg[30]/NET0131 , \rd1_R_o_reg[31]/NET0131 , \rd1_R_o_reg[3]/NET0131 , \rd1_R_o_reg[4]/NET0131 , \rd1_R_o_reg[5]/NET0131 , \rd1_R_o_reg[6]/NET0131 , \rd1_R_o_reg[7]/NET0131 , \rd1_R_o_reg[8]/NET0131 , \rd1_R_o_reg[9]/NET0131 , \stage1_iter_reg[0]/NET0131 , \stage1_iter_reg[1]/NET0131 , \stage1_iter_reg[2]/NET0131 , \stage1_iter_reg[3]/NET0131 , \_al_n0 , \_al_n1 , \g10087/_0_ , \g10220/_1_ , \g11117/_0_ , \g11124/_0_ , \g11125/_0_ , \g11170/_0_ , \g11182/_0_ , \g11184/_0_ , \g11378/_0_ , \g11393/_0_ , \g11415/_0_ , \g11432/_0_ , \g11433/_0_ , \g11453/_0_ , \g11500/_0_ , \g11588/_0_ , \g11607/_0_ , \g11616/_0_ , \g11625/_0_ , \g11641_dup/_0_ , \g11648/_0_ , \g11655/_0_ , \g11683/_0_ , \g11689/_2_ , \g11694/_0_ , \g11748/_0_ , \g11880/_0_ , \g11962/_1_ , \g12016/_0_ , \g12038/_0_ , \g12039/_0_ , \g12094/_0_ , \g12100/_0_ , \g12132/_0_ , \g12151/_0_ , \g12251/_0_ , \g12279/_0_ , \g12288/_0_ , \g12290/_0_ , \g12311/_0_ , \g12313/_0_ , \g12356/_0_ , \g12357/_0_ , \g12427/_0_ , \g12441/_0_ , \g12442/_0_ , \g12480/_0_ , \g12485/_0_ , \g12506/_0_ , \g12544/_0_ , \g12549/_2_ , \g12614/_0_ , \g12678/_0_ , \g12680/_0_ , \g12748/_0_ , \g15/_0_ , \g25/_0_ , \g31/_0_ , \g6843/_0_ , \g6861/_0_ , \g6863/_0_ , \g6865/_0_ , \g6887/_0_ , \g6888/_0_ , \g6889/_0_ , \g6890/_0_ , \g6891/_0_ , \g6892/_0_ , \g6893/_0_ , \g6894/_0_ , \g6922/_0_ , \g6923/_0_ , \g6924/_3_ , \g6926/_0_ , \g6927/_0_ , \g6928/_0_ , \g6931/_0_ , \g6933/_0_ , \g6967/_0_ , \g6968/_0_ , \g6969/_0_ , \g6974/_0_ , \g6975/_0_ , \g6976/_3_ , \g7006/_3_ , \g8882/_0_ , \g8883/_0_ , \g8884/_0_ , \g8895/_0_ , \g8896/_0_ , \g8898/_0_ , \g8900/_2_ , \g8902/_0_ , \g8907/_0_ , \g8911/_0_ , \g8924/_0_ , \g8927/_0_ , \g8929/_2_ , \g8967/_0_ , \g8969/_0_ , \g8973/_2_ , \g8987/_0_ , \g8989/_0_ , \g8991/_0_ , \g8996/_0_ , \g9099/_0_ , \g9543/_1_ , \g9751/_1_ , \g9755/_0_ , \g9786/_0_ , \g9794/_0_ , \g9817/_0_ , \g9836/_0_ , \g9859/_0_ , \g9862/_0_ , \g9867/_0_ , \g9869/_0_ , \g9876/_0_ , \g9887/_0_ , \g9895/_0_ , \g9897/_0_ , \g9908/_0_ , \g9910/_0_ , \g9915/_0_ , \g9938/_0_ , \g9970/_0_ );
	input \data_i[0]_pad  ;
	input \data_i[10]_pad  ;
	input \data_i[11]_pad  ;
	input \data_i[12]_pad  ;
	input \data_i[13]_pad  ;
	input \data_i[14]_pad  ;
	input \data_i[15]_pad  ;
	input \data_i[16]_pad  ;
	input \data_i[17]_pad  ;
	input \data_i[18]_pad  ;
	input \data_i[19]_pad  ;
	input \data_i[1]_pad  ;
	input \data_i[20]_pad  ;
	input \data_i[21]_pad  ;
	input \data_i[22]_pad  ;
	input \data_i[23]_pad  ;
	input \data_i[24]_pad  ;
	input \data_i[25]_pad  ;
	input \data_i[26]_pad  ;
	input \data_i[27]_pad  ;
	input \data_i[28]_pad  ;
	input \data_i[29]_pad  ;
	input \data_i[2]_pad  ;
	input \data_i[30]_pad  ;
	input \data_i[31]_pad  ;
	input \data_i[32]_pad  ;
	input \data_i[33]_pad  ;
	input \data_i[34]_pad  ;
	input \data_i[35]_pad  ;
	input \data_i[36]_pad  ;
	input \data_i[37]_pad  ;
	input \data_i[38]_pad  ;
	input \data_i[39]_pad  ;
	input \data_i[3]_pad  ;
	input \data_i[40]_pad  ;
	input \data_i[41]_pad  ;
	input \data_i[42]_pad  ;
	input \data_i[43]_pad  ;
	input \data_i[44]_pad  ;
	input \data_i[45]_pad  ;
	input \data_i[46]_pad  ;
	input \data_i[47]_pad  ;
	input \data_i[48]_pad  ;
	input \data_i[49]_pad  ;
	input \data_i[4]_pad  ;
	input \data_i[50]_pad  ;
	input \data_i[51]_pad  ;
	input \data_i[52]_pad  ;
	input \data_i[53]_pad  ;
	input \data_i[54]_pad  ;
	input \data_i[55]_pad  ;
	input \data_i[56]_pad  ;
	input \data_i[57]_pad  ;
	input \data_i[58]_pad  ;
	input \data_i[59]_pad  ;
	input \data_i[5]_pad  ;
	input \data_i[60]_pad  ;
	input \data_i[61]_pad  ;
	input \data_i[62]_pad  ;
	input \data_i[63]_pad  ;
	input \data_i[6]_pad  ;
	input \data_i[7]_pad  ;
	input \data_i[8]_pad  ;
	input \data_i[9]_pad  ;
	input \data_ready_reg/NET0131  ;
	input decrypt_i_pad ;
	input \key_i[10]_pad  ;
	input \key_i[11]_pad  ;
	input \key_i[12]_pad  ;
	input \key_i[13]_pad  ;
	input \key_i[14]_pad  ;
	input \key_i[15]_pad  ;
	input \key_i[17]_pad  ;
	input \key_i[18]_pad  ;
	input \key_i[19]_pad  ;
	input \key_i[1]_pad  ;
	input \key_i[20]_pad  ;
	input \key_i[21]_pad  ;
	input \key_i[22]_pad  ;
	input \key_i[23]_pad  ;
	input \key_i[25]_pad  ;
	input \key_i[26]_pad  ;
	input \key_i[27]_pad  ;
	input \key_i[28]_pad  ;
	input \key_i[29]_pad  ;
	input \key_i[2]_pad  ;
	input \key_i[30]_pad  ;
	input \key_i[31]_pad  ;
	input \key_i[33]_pad  ;
	input \key_i[34]_pad  ;
	input \key_i[35]_pad  ;
	input \key_i[36]_pad  ;
	input \key_i[37]_pad  ;
	input \key_i[38]_pad  ;
	input \key_i[39]_pad  ;
	input \key_i[3]_pad  ;
	input \key_i[41]_pad  ;
	input \key_i[42]_pad  ;
	input \key_i[43]_pad  ;
	input \key_i[44]_pad  ;
	input \key_i[45]_pad  ;
	input \key_i[46]_pad  ;
	input \key_i[47]_pad  ;
	input \key_i[49]_pad  ;
	input \key_i[4]_pad  ;
	input \key_i[50]_pad  ;
	input \key_i[51]_pad  ;
	input \key_i[52]_pad  ;
	input \key_i[53]_pad  ;
	input \key_i[54]_pad  ;
	input \key_i[55]_pad  ;
	input \key_i[57]_pad  ;
	input \key_i[58]_pad  ;
	input \key_i[59]_pad  ;
	input \key_i[5]_pad  ;
	input \key_i[60]_pad  ;
	input \key_i[61]_pad  ;
	input \key_i[62]_pad  ;
	input \key_i[63]_pad  ;
	input \key_i[6]_pad  ;
	input \key_i[7]_pad  ;
	input \key_i[9]_pad  ;
	input load_i_pad ;
	input \rd1_Key_o_reg[0]/NET0131  ;
	input \rd1_Key_o_reg[10]/NET0131  ;
	input \rd1_Key_o_reg[11]/NET0131  ;
	input \rd1_Key_o_reg[12]/NET0131  ;
	input \rd1_Key_o_reg[13]/NET0131  ;
	input \rd1_Key_o_reg[14]/NET0131  ;
	input \rd1_Key_o_reg[15]/NET0131  ;
	input \rd1_Key_o_reg[16]/NET0131  ;
	input \rd1_Key_o_reg[17]/NET0131  ;
	input \rd1_Key_o_reg[18]/NET0131  ;
	input \rd1_Key_o_reg[19]/NET0131  ;
	input \rd1_Key_o_reg[1]/NET0131  ;
	input \rd1_Key_o_reg[20]/NET0131  ;
	input \rd1_Key_o_reg[21]/NET0131  ;
	input \rd1_Key_o_reg[22]/NET0131  ;
	input \rd1_Key_o_reg[23]/NET0131  ;
	input \rd1_Key_o_reg[24]/NET0131  ;
	input \rd1_Key_o_reg[25]/NET0131  ;
	input \rd1_Key_o_reg[26]/NET0131  ;
	input \rd1_Key_o_reg[27]/NET0131  ;
	input \rd1_Key_o_reg[28]/NET0131  ;
	input \rd1_Key_o_reg[29]/NET0131  ;
	input \rd1_Key_o_reg[2]/NET0131  ;
	input \rd1_Key_o_reg[30]/NET0131  ;
	input \rd1_Key_o_reg[31]/NET0131  ;
	input \rd1_Key_o_reg[32]/NET0131  ;
	input \rd1_Key_o_reg[33]/NET0131  ;
	input \rd1_Key_o_reg[34]/NET0131  ;
	input \rd1_Key_o_reg[35]/NET0131  ;
	input \rd1_Key_o_reg[36]/NET0131  ;
	input \rd1_Key_o_reg[37]/NET0131  ;
	input \rd1_Key_o_reg[38]/NET0131  ;
	input \rd1_Key_o_reg[39]/NET0131  ;
	input \rd1_Key_o_reg[3]/NET0131  ;
	input \rd1_Key_o_reg[40]/NET0131  ;
	input \rd1_Key_o_reg[41]/NET0131  ;
	input \rd1_Key_o_reg[42]/NET0131  ;
	input \rd1_Key_o_reg[43]/NET0131  ;
	input \rd1_Key_o_reg[44]/NET0131  ;
	input \rd1_Key_o_reg[45]/NET0131  ;
	input \rd1_Key_o_reg[46]/NET0131  ;
	input \rd1_Key_o_reg[47]/NET0131  ;
	input \rd1_Key_o_reg[48]/NET0131  ;
	input \rd1_Key_o_reg[49]/NET0131  ;
	input \rd1_Key_o_reg[4]/NET0131  ;
	input \rd1_Key_o_reg[50]/NET0131  ;
	input \rd1_Key_o_reg[51]/NET0131  ;
	input \rd1_Key_o_reg[52]/NET0131  ;
	input \rd1_Key_o_reg[53]/NET0131  ;
	input \rd1_Key_o_reg[54]/NET0131  ;
	input \rd1_Key_o_reg[55]/NET0131  ;
	input \rd1_Key_o_reg[5]/NET0131  ;
	input \rd1_Key_o_reg[6]/NET0131  ;
	input \rd1_Key_o_reg[7]/NET0131  ;
	input \rd1_Key_o_reg[8]/NET0131  ;
	input \rd1_Key_o_reg[9]/NET0131  ;
	input \rd1_L_o_reg[0]/NET0131  ;
	input \rd1_L_o_reg[10]/NET0131  ;
	input \rd1_L_o_reg[11]/NET0131  ;
	input \rd1_L_o_reg[12]/NET0131  ;
	input \rd1_L_o_reg[13]/NET0131  ;
	input \rd1_L_o_reg[14]/NET0131  ;
	input \rd1_L_o_reg[15]/NET0131  ;
	input \rd1_L_o_reg[16]/NET0131  ;
	input \rd1_L_o_reg[17]/NET0131  ;
	input \rd1_L_o_reg[18]/NET0131  ;
	input \rd1_L_o_reg[19]/NET0131  ;
	input \rd1_L_o_reg[1]/NET0131  ;
	input \rd1_L_o_reg[20]/NET0131  ;
	input \rd1_L_o_reg[21]/NET0131  ;
	input \rd1_L_o_reg[22]/NET0131  ;
	input \rd1_L_o_reg[23]/NET0131  ;
	input \rd1_L_o_reg[24]/NET0131  ;
	input \rd1_L_o_reg[25]/NET0131  ;
	input \rd1_L_o_reg[26]/NET0131  ;
	input \rd1_L_o_reg[27]/NET0131  ;
	input \rd1_L_o_reg[28]/NET0131  ;
	input \rd1_L_o_reg[29]/NET0131  ;
	input \rd1_L_o_reg[2]/NET0131  ;
	input \rd1_L_o_reg[30]/NET0131  ;
	input \rd1_L_o_reg[31]/NET0131  ;
	input \rd1_L_o_reg[3]/NET0131  ;
	input \rd1_L_o_reg[4]/NET0131  ;
	input \rd1_L_o_reg[5]/NET0131  ;
	input \rd1_L_o_reg[6]/NET0131  ;
	input \rd1_L_o_reg[7]/NET0131  ;
	input \rd1_L_o_reg[8]/NET0131  ;
	input \rd1_L_o_reg[9]/NET0131  ;
	input \rd1_R_o_reg[0]/NET0131  ;
	input \rd1_R_o_reg[10]/NET0131  ;
	input \rd1_R_o_reg[11]/NET0131  ;
	input \rd1_R_o_reg[12]/NET0131  ;
	input \rd1_R_o_reg[13]/NET0131  ;
	input \rd1_R_o_reg[14]/NET0131  ;
	input \rd1_R_o_reg[15]/NET0131  ;
	input \rd1_R_o_reg[16]/NET0131  ;
	input \rd1_R_o_reg[17]/NET0131  ;
	input \rd1_R_o_reg[18]/NET0131  ;
	input \rd1_R_o_reg[19]/NET0131  ;
	input \rd1_R_o_reg[1]/NET0131  ;
	input \rd1_R_o_reg[20]/NET0131  ;
	input \rd1_R_o_reg[21]/NET0131  ;
	input \rd1_R_o_reg[22]/NET0131  ;
	input \rd1_R_o_reg[23]/NET0131  ;
	input \rd1_R_o_reg[24]/NET0131  ;
	input \rd1_R_o_reg[25]/NET0131  ;
	input \rd1_R_o_reg[26]/NET0131  ;
	input \rd1_R_o_reg[27]/NET0131  ;
	input \rd1_R_o_reg[28]/NET0131  ;
	input \rd1_R_o_reg[29]/NET0131  ;
	input \rd1_R_o_reg[2]/NET0131  ;
	input \rd1_R_o_reg[30]/NET0131  ;
	input \rd1_R_o_reg[31]/NET0131  ;
	input \rd1_R_o_reg[3]/NET0131  ;
	input \rd1_R_o_reg[4]/NET0131  ;
	input \rd1_R_o_reg[5]/NET0131  ;
	input \rd1_R_o_reg[6]/NET0131  ;
	input \rd1_R_o_reg[7]/NET0131  ;
	input \rd1_R_o_reg[8]/NET0131  ;
	input \rd1_R_o_reg[9]/NET0131  ;
	input \stage1_iter_reg[0]/NET0131  ;
	input \stage1_iter_reg[1]/NET0131  ;
	input \stage1_iter_reg[2]/NET0131  ;
	input \stage1_iter_reg[3]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g10087/_0_  ;
	output \g10220/_1_  ;
	output \g11117/_0_  ;
	output \g11124/_0_  ;
	output \g11125/_0_  ;
	output \g11170/_0_  ;
	output \g11182/_0_  ;
	output \g11184/_0_  ;
	output \g11378/_0_  ;
	output \g11393/_0_  ;
	output \g11415/_0_  ;
	output \g11432/_0_  ;
	output \g11433/_0_  ;
	output \g11453/_0_  ;
	output \g11500/_0_  ;
	output \g11588/_0_  ;
	output \g11607/_0_  ;
	output \g11616/_0_  ;
	output \g11625/_0_  ;
	output \g11641_dup/_0_  ;
	output \g11648/_0_  ;
	output \g11655/_0_  ;
	output \g11683/_0_  ;
	output \g11689/_2_  ;
	output \g11694/_0_  ;
	output \g11748/_0_  ;
	output \g11880/_0_  ;
	output \g11962/_1_  ;
	output \g12016/_0_  ;
	output \g12038/_0_  ;
	output \g12039/_0_  ;
	output \g12094/_0_  ;
	output \g12100/_0_  ;
	output \g12132/_0_  ;
	output \g12151/_0_  ;
	output \g12251/_0_  ;
	output \g12279/_0_  ;
	output \g12288/_0_  ;
	output \g12290/_0_  ;
	output \g12311/_0_  ;
	output \g12313/_0_  ;
	output \g12356/_0_  ;
	output \g12357/_0_  ;
	output \g12427/_0_  ;
	output \g12441/_0_  ;
	output \g12442/_0_  ;
	output \g12480/_0_  ;
	output \g12485/_0_  ;
	output \g12506/_0_  ;
	output \g12544/_0_  ;
	output \g12549/_2_  ;
	output \g12614/_0_  ;
	output \g12678/_0_  ;
	output \g12680/_0_  ;
	output \g12748/_0_  ;
	output \g15/_0_  ;
	output \g25/_0_  ;
	output \g31/_0_  ;
	output \g6843/_0_  ;
	output \g6861/_0_  ;
	output \g6863/_0_  ;
	output \g6865/_0_  ;
	output \g6887/_0_  ;
	output \g6888/_0_  ;
	output \g6889/_0_  ;
	output \g6890/_0_  ;
	output \g6891/_0_  ;
	output \g6892/_0_  ;
	output \g6893/_0_  ;
	output \g6894/_0_  ;
	output \g6922/_0_  ;
	output \g6923/_0_  ;
	output \g6924/_3_  ;
	output \g6926/_0_  ;
	output \g6927/_0_  ;
	output \g6928/_0_  ;
	output \g6931/_0_  ;
	output \g6933/_0_  ;
	output \g6967/_0_  ;
	output \g6968/_0_  ;
	output \g6969/_0_  ;
	output \g6974/_0_  ;
	output \g6975/_0_  ;
	output \g6976/_3_  ;
	output \g7006/_3_  ;
	output \g8882/_0_  ;
	output \g8883/_0_  ;
	output \g8884/_0_  ;
	output \g8895/_0_  ;
	output \g8896/_0_  ;
	output \g8898/_0_  ;
	output \g8900/_2_  ;
	output \g8902/_0_  ;
	output \g8907/_0_  ;
	output \g8911/_0_  ;
	output \g8924/_0_  ;
	output \g8927/_0_  ;
	output \g8929/_2_  ;
	output \g8967/_0_  ;
	output \g8969/_0_  ;
	output \g8973/_2_  ;
	output \g8987/_0_  ;
	output \g8989/_0_  ;
	output \g8991/_0_  ;
	output \g8996/_0_  ;
	output \g9099/_0_  ;
	output \g9543/_1_  ;
	output \g9751/_1_  ;
	output \g9755/_0_  ;
	output \g9786/_0_  ;
	output \g9794/_0_  ;
	output \g9817/_0_  ;
	output \g9836/_0_  ;
	output \g9859/_0_  ;
	output \g9862/_0_  ;
	output \g9867/_0_  ;
	output \g9869/_0_  ;
	output \g9876/_0_  ;
	output \g9887/_0_  ;
	output \g9895/_0_  ;
	output \g9897/_0_  ;
	output \g9908/_0_  ;
	output \g9910/_0_  ;
	output \g9915/_0_  ;
	output \g9938/_0_  ;
	output \g9970/_0_  ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[3]/NET0131 ,
		_w249_
	);
	LUT4 #(
		.INIT('h0001)
	) name1 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[1]/NET0131 ,
		\stage1_iter_reg[2]/NET0131 ,
		\stage1_iter_reg[3]/NET0131 ,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\data_ready_reg/NET0131 ,
		load_i_pad,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h6)
	) name4 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[1]/NET0131 ,
		_w253_
	);
	LUT3 #(
		.INIT('hb8)
	) name5 (
		\key_i[9]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[26]/NET0131 ,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w250_,
		_w254_,
		_w255_
	);
	LUT4 #(
		.INIT('h7efc)
	) name7 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[1]/NET0131 ,
		\stage1_iter_reg[2]/NET0131 ,
		\stage1_iter_reg[3]/NET0131 ,
		_w256_
	);
	LUT4 #(
		.INIT('h00e2)
	) name8 (
		\rd1_Key_o_reg[26]/NET0131 ,
		_w250_,
		_w254_,
		_w256_,
		_w257_
	);
	LUT3 #(
		.INIT('hb8)
	) name9 (
		\key_i[17]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[25]/NET0131 ,
		_w258_
	);
	LUT4 #(
		.INIT('he020)
	) name10 (
		\rd1_Key_o_reg[25]/NET0131 ,
		_w250_,
		_w256_,
		_w258_,
		_w259_
	);
	LUT3 #(
		.INIT('h54)
	) name11 (
		decrypt_i_pad,
		_w257_,
		_w259_,
		_w260_
	);
	LUT3 #(
		.INIT('hb8)
	) name12 (
		\key_i[60]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[0]/NET0131 ,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w250_,
		_w261_,
		_w262_
	);
	LUT4 #(
		.INIT('h8102)
	) name14 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[1]/NET0131 ,
		\stage1_iter_reg[2]/NET0131 ,
		\stage1_iter_reg[3]/NET0131 ,
		_w263_
	);
	LUT4 #(
		.INIT('he200)
	) name15 (
		\rd1_Key_o_reg[0]/NET0131 ,
		_w250_,
		_w261_,
		_w263_,
		_w264_
	);
	LUT3 #(
		.INIT('hb8)
	) name16 (
		\key_i[1]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[27]/NET0131 ,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		_w250_,
		_w265_,
		_w266_
	);
	LUT4 #(
		.INIT('h470f)
	) name18 (
		\key_i[52]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[1]/NET0131 ,
		_w250_,
		_w267_
	);
	LUT4 #(
		.INIT('h0031)
	) name19 (
		_w256_,
		_w266_,
		_w267_,
		_w264_,
		_w268_
	);
	LUT3 #(
		.INIT('hce)
	) name20 (
		decrypt_i_pad,
		_w260_,
		_w268_,
		_w269_
	);
	LUT4 #(
		.INIT('h470f)
	) name21 (
		\data_i[43]_pad ,
		load_i_pad,
		\rd1_R_o_reg[10]/NET0131 ,
		_w250_,
		_w270_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name22 (
		\data_i[43]_pad ,
		load_i_pad,
		\rd1_R_o_reg[10]/NET0131 ,
		_w250_,
		_w271_
	);
	LUT4 #(
		.INIT('h470f)
	) name23 (
		\key_i[36]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[3]/NET0131 ,
		_w250_,
		_w272_
	);
	LUT3 #(
		.INIT('hb8)
	) name24 (
		\key_i[59]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[4]/NET0131 ,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		_w250_,
		_w273_,
		_w274_
	);
	LUT3 #(
		.INIT('h1d)
	) name26 (
		\rd1_Key_o_reg[4]/NET0131 ,
		_w250_,
		_w273_,
		_w275_
	);
	LUT4 #(
		.INIT('h0415)
	) name27 (
		decrypt_i_pad,
		_w256_,
		_w272_,
		_w275_,
		_w276_
	);
	LUT3 #(
		.INIT('hb8)
	) name28 (
		\key_i[43]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[6]/NET0131 ,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w250_,
		_w277_,
		_w278_
	);
	LUT3 #(
		.INIT('h1d)
	) name30 (
		\rd1_Key_o_reg[6]/NET0131 ,
		_w250_,
		_w277_,
		_w279_
	);
	LUT4 #(
		.INIT('he020)
	) name31 (
		\rd1_Key_o_reg[6]/NET0131 ,
		_w250_,
		_w263_,
		_w277_,
		_w280_
	);
	LUT4 #(
		.INIT('h470f)
	) name32 (
		\key_i[51]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[5]/NET0131 ,
		_w250_,
		_w281_
	);
	LUT4 #(
		.INIT('hb800)
	) name33 (
		\key_i[51]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[5]/NET0131 ,
		_w250_,
		_w282_
	);
	LUT3 #(
		.INIT('hb8)
	) name34 (
		\key_i[35]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[7]/NET0131 ,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w250_,
		_w283_,
		_w284_
	);
	LUT4 #(
		.INIT('he020)
	) name36 (
		\rd1_Key_o_reg[7]/NET0131 ,
		_w250_,
		_w256_,
		_w283_,
		_w285_
	);
	LUT4 #(
		.INIT('haaa8)
	) name37 (
		decrypt_i_pad,
		_w282_,
		_w285_,
		_w280_,
		_w286_
	);
	LUT2 #(
		.INIT('he)
	) name38 (
		_w276_,
		_w286_,
		_w287_
	);
	LUT3 #(
		.INIT('hb8)
	) name39 (
		\key_i[28]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[28]/NET0131 ,
		_w288_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w250_,
		_w288_,
		_w289_
	);
	LUT4 #(
		.INIT('h0e02)
	) name41 (
		\rd1_Key_o_reg[28]/NET0131 ,
		_w250_,
		_w256_,
		_w288_,
		_w290_
	);
	LUT3 #(
		.INIT('hb8)
	) name42 (
		\key_i[7]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[55]/NET0131 ,
		_w291_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w250_,
		_w291_,
		_w292_
	);
	LUT3 #(
		.INIT('h1d)
	) name44 (
		\rd1_Key_o_reg[55]/NET0131 ,
		_w250_,
		_w291_,
		_w293_
	);
	LUT4 #(
		.INIT('he020)
	) name45 (
		\rd1_Key_o_reg[55]/NET0131 ,
		_w250_,
		_w256_,
		_w291_,
		_w294_
	);
	LUT3 #(
		.INIT('h54)
	) name46 (
		decrypt_i_pad,
		_w290_,
		_w294_,
		_w295_
	);
	LUT3 #(
		.INIT('hb8)
	) name47 (
		\key_i[12]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[30]/NET0131 ,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w250_,
		_w296_,
		_w297_
	);
	LUT4 #(
		.INIT('he020)
	) name49 (
		\rd1_Key_o_reg[30]/NET0131 ,
		_w250_,
		_w263_,
		_w296_,
		_w298_
	);
	LUT3 #(
		.INIT('hb8)
	) name50 (
		\key_i[20]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[29]/NET0131 ,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w250_,
		_w299_,
		_w300_
	);
	LUT3 #(
		.INIT('hb8)
	) name52 (
		\key_i[4]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[31]/NET0131 ,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w250_,
		_w301_,
		_w302_
	);
	LUT4 #(
		.INIT('he020)
	) name54 (
		\rd1_Key_o_reg[31]/NET0131 ,
		_w250_,
		_w256_,
		_w301_,
		_w303_
	);
	LUT4 #(
		.INIT('haaa8)
	) name55 (
		decrypt_i_pad,
		_w300_,
		_w303_,
		_w298_,
		_w304_
	);
	LUT2 #(
		.INIT('he)
	) name56 (
		_w295_,
		_w304_,
		_w305_
	);
	LUT4 #(
		.INIT('h470f)
	) name57 (
		\data_i[25]_pad ,
		load_i_pad,
		\rd1_R_o_reg[4]/NET0131 ,
		_w250_,
		_w306_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name58 (
		\data_i[25]_pad ,
		load_i_pad,
		\rd1_R_o_reg[4]/NET0131 ,
		_w250_,
		_w307_
	);
	LUT3 #(
		.INIT('hb8)
	) name59 (
		\key_i[49]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[21]/NET0131 ,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w250_,
		_w308_,
		_w309_
	);
	LUT4 #(
		.INIT('h0e02)
	) name61 (
		\rd1_Key_o_reg[21]/NET0131 ,
		_w250_,
		_w256_,
		_w308_,
		_w310_
	);
	LUT3 #(
		.INIT('hb8)
	) name62 (
		\key_i[57]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[20]/NET0131 ,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w250_,
		_w311_,
		_w312_
	);
	LUT3 #(
		.INIT('h1d)
	) name64 (
		\rd1_Key_o_reg[20]/NET0131 ,
		_w250_,
		_w311_,
		_w313_
	);
	LUT4 #(
		.INIT('he020)
	) name65 (
		\rd1_Key_o_reg[20]/NET0131 ,
		_w250_,
		_w256_,
		_w311_,
		_w314_
	);
	LUT3 #(
		.INIT('h54)
	) name66 (
		decrypt_i_pad,
		_w310_,
		_w314_,
		_w315_
	);
	LUT4 #(
		.INIT('h470f)
	) name67 (
		\key_i[33]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[23]/NET0131 ,
		_w250_,
		_w316_
	);
	LUT3 #(
		.INIT('hb8)
	) name68 (
		\key_i[25]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[24]/NET0131 ,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w250_,
		_w317_,
		_w318_
	);
	LUT3 #(
		.INIT('h1d)
	) name70 (
		\rd1_Key_o_reg[24]/NET0131 ,
		_w250_,
		_w317_,
		_w319_
	);
	LUT4 #(
		.INIT('he020)
	) name71 (
		\rd1_Key_o_reg[24]/NET0131 ,
		_w250_,
		_w256_,
		_w317_,
		_w320_
	);
	LUT3 #(
		.INIT('hb8)
	) name72 (
		\key_i[41]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[22]/NET0131 ,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w250_,
		_w321_,
		_w322_
	);
	LUT4 #(
		.INIT('h0031)
	) name74 (
		_w263_,
		_w320_,
		_w316_,
		_w322_,
		_w323_
	);
	LUT3 #(
		.INIT('hce)
	) name75 (
		decrypt_i_pad,
		_w315_,
		_w323_,
		_w324_
	);
	LUT4 #(
		.INIT('h0415)
	) name76 (
		decrypt_i_pad,
		_w256_,
		_w281_,
		_w279_,
		_w325_
	);
	LUT4 #(
		.INIT('h470f)
	) name77 (
		\key_i[27]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[8]/NET0131 ,
		_w250_,
		_w326_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		_w263_,
		_w326_,
		_w327_
	);
	LUT4 #(
		.INIT('h470f)
	) name79 (
		\key_i[19]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[9]/NET0131 ,
		_w250_,
		_w328_
	);
	LUT3 #(
		.INIT('h31)
	) name80 (
		_w256_,
		_w284_,
		_w328_,
		_w329_
	);
	LUT4 #(
		.INIT('h1311)
	) name81 (
		decrypt_i_pad,
		_w325_,
		_w327_,
		_w329_,
		_w330_
	);
	LUT4 #(
		.INIT('hecee)
	) name82 (
		decrypt_i_pad,
		_w325_,
		_w327_,
		_w329_,
		_w331_
	);
	LUT3 #(
		.INIT('hb8)
	) name83 (
		\key_i[11]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[10]/NET0131 ,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w250_,
		_w332_,
		_w333_
	);
	LUT3 #(
		.INIT('h1d)
	) name85 (
		\rd1_Key_o_reg[10]/NET0131 ,
		_w250_,
		_w332_,
		_w334_
	);
	LUT4 #(
		.INIT('h0415)
	) name86 (
		decrypt_i_pad,
		_w256_,
		_w328_,
		_w334_,
		_w335_
	);
	LUT4 #(
		.INIT('h470f)
	) name87 (
		\key_i[50]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[13]/NET0131 ,
		_w250_,
		_w336_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w256_,
		_w336_,
		_w337_
	);
	LUT4 #(
		.INIT('h470f)
	) name89 (
		\key_i[58]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[12]/NET0131 ,
		_w250_,
		_w338_
	);
	LUT3 #(
		.INIT('hb8)
	) name90 (
		\key_i[3]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[11]/NET0131 ,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w250_,
		_w339_,
		_w340_
	);
	LUT3 #(
		.INIT('h0d)
	) name92 (
		_w263_,
		_w338_,
		_w340_,
		_w341_
	);
	LUT4 #(
		.INIT('h1311)
	) name93 (
		decrypt_i_pad,
		_w335_,
		_w337_,
		_w341_,
		_w342_
	);
	LUT4 #(
		.INIT('hecee)
	) name94 (
		decrypt_i_pad,
		_w335_,
		_w337_,
		_w341_,
		_w343_
	);
	LUT4 #(
		.INIT('h0e02)
	) name95 (
		\rd1_Key_o_reg[29]/NET0131 ,
		_w250_,
		_w256_,
		_w299_,
		_w344_
	);
	LUT4 #(
		.INIT('he020)
	) name96 (
		\rd1_Key_o_reg[28]/NET0131 ,
		_w250_,
		_w256_,
		_w288_,
		_w345_
	);
	LUT3 #(
		.INIT('h54)
	) name97 (
		decrypt_i_pad,
		_w344_,
		_w345_,
		_w346_
	);
	LUT4 #(
		.INIT('he020)
	) name98 (
		\rd1_Key_o_reg[31]/NET0131 ,
		_w250_,
		_w263_,
		_w301_,
		_w347_
	);
	LUT3 #(
		.INIT('hb8)
	) name99 (
		\key_i[61]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[32]/NET0131 ,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w250_,
		_w348_,
		_w349_
	);
	LUT4 #(
		.INIT('he020)
	) name101 (
		\rd1_Key_o_reg[32]/NET0131 ,
		_w250_,
		_w256_,
		_w348_,
		_w350_
	);
	LUT4 #(
		.INIT('haaa8)
	) name102 (
		decrypt_i_pad,
		_w297_,
		_w350_,
		_w347_,
		_w351_
	);
	LUT2 #(
		.INIT('he)
	) name103 (
		_w346_,
		_w351_,
		_w352_
	);
	LUT4 #(
		.INIT('h0e02)
	) name104 (
		\rd1_Key_o_reg[31]/NET0131 ,
		_w250_,
		_w256_,
		_w301_,
		_w353_
	);
	LUT4 #(
		.INIT('he020)
	) name105 (
		\rd1_Key_o_reg[30]/NET0131 ,
		_w250_,
		_w256_,
		_w296_,
		_w354_
	);
	LUT3 #(
		.INIT('h54)
	) name106 (
		decrypt_i_pad,
		_w353_,
		_w354_,
		_w355_
	);
	LUT4 #(
		.INIT('h470f)
	) name107 (
		\key_i[53]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[33]/NET0131 ,
		_w250_,
		_w356_
	);
	LUT3 #(
		.INIT('hb8)
	) name108 (
		\key_i[45]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[34]/NET0131 ,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w250_,
		_w357_,
		_w358_
	);
	LUT3 #(
		.INIT('h1d)
	) name110 (
		\rd1_Key_o_reg[34]/NET0131 ,
		_w250_,
		_w357_,
		_w359_
	);
	LUT4 #(
		.INIT('he020)
	) name111 (
		\rd1_Key_o_reg[34]/NET0131 ,
		_w250_,
		_w256_,
		_w357_,
		_w360_
	);
	LUT4 #(
		.INIT('h0301)
	) name112 (
		_w263_,
		_w349_,
		_w360_,
		_w356_,
		_w361_
	);
	LUT3 #(
		.INIT('hce)
	) name113 (
		decrypt_i_pad,
		_w355_,
		_w361_,
		_w362_
	);
	LUT4 #(
		.INIT('h470f)
	) name114 (
		\data_i[23]_pad ,
		load_i_pad,
		\rd1_R_o_reg[29]/NET0131 ,
		_w250_,
		_w363_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name115 (
		\data_i[23]_pad ,
		load_i_pad,
		\rd1_R_o_reg[29]/NET0131 ,
		_w250_,
		_w364_
	);
	LUT4 #(
		.INIT('hb800)
	) name116 (
		\key_i[19]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[9]/NET0131 ,
		_w250_,
		_w365_
	);
	LUT4 #(
		.INIT('hfe32)
	) name117 (
		_w249_,
		_w256_,
		_w328_,
		_w326_,
		_w366_
	);
	LUT4 #(
		.INIT('he020)
	) name118 (
		\rd1_Key_o_reg[11]/NET0131 ,
		_w250_,
		_w263_,
		_w339_,
		_w367_
	);
	LUT4 #(
		.INIT('h0031)
	) name119 (
		_w256_,
		_w333_,
		_w338_,
		_w367_,
		_w368_
	);
	LUT4 #(
		.INIT('hba10)
	) name120 (
		decrypt_i_pad,
		_w365_,
		_w366_,
		_w368_,
		_w369_
	);
	LUT4 #(
		.INIT('h45ef)
	) name121 (
		decrypt_i_pad,
		_w365_,
		_w366_,
		_w368_,
		_w370_
	);
	LUT4 #(
		.INIT('h0e02)
	) name122 (
		\rd1_Key_o_reg[32]/NET0131 ,
		_w250_,
		_w256_,
		_w348_,
		_w371_
	);
	LUT3 #(
		.INIT('h54)
	) name123 (
		decrypt_i_pad,
		_w303_,
		_w371_,
		_w372_
	);
	LUT4 #(
		.INIT('he020)
	) name124 (
		\rd1_Key_o_reg[34]/NET0131 ,
		_w250_,
		_w263_,
		_w357_,
		_w373_
	);
	LUT4 #(
		.INIT('hb800)
	) name125 (
		\key_i[53]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[33]/NET0131 ,
		_w250_,
		_w374_
	);
	LUT3 #(
		.INIT('hb8)
	) name126 (
		\key_i[37]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[35]/NET0131 ,
		_w375_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w250_,
		_w375_,
		_w376_
	);
	LUT4 #(
		.INIT('he020)
	) name128 (
		\rd1_Key_o_reg[35]/NET0131 ,
		_w250_,
		_w256_,
		_w375_,
		_w377_
	);
	LUT4 #(
		.INIT('haaa8)
	) name129 (
		decrypt_i_pad,
		_w374_,
		_w377_,
		_w373_,
		_w378_
	);
	LUT2 #(
		.INIT('he)
	) name130 (
		_w372_,
		_w378_,
		_w379_
	);
	LUT4 #(
		.INIT('h0e02)
	) name131 (
		\rd1_Key_o_reg[22]/NET0131 ,
		_w250_,
		_w256_,
		_w321_,
		_w380_
	);
	LUT4 #(
		.INIT('he020)
	) name132 (
		\rd1_Key_o_reg[21]/NET0131 ,
		_w250_,
		_w256_,
		_w308_,
		_w381_
	);
	LUT3 #(
		.INIT('h54)
	) name133 (
		decrypt_i_pad,
		_w380_,
		_w381_,
		_w382_
	);
	LUT4 #(
		.INIT('he020)
	) name134 (
		\rd1_Key_o_reg[24]/NET0131 ,
		_w250_,
		_w263_,
		_w317_,
		_w383_
	);
	LUT4 #(
		.INIT('hb800)
	) name135 (
		\key_i[33]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[23]/NET0131 ,
		_w250_,
		_w384_
	);
	LUT4 #(
		.INIT('haaa8)
	) name136 (
		decrypt_i_pad,
		_w259_,
		_w384_,
		_w383_,
		_w385_
	);
	LUT2 #(
		.INIT('he)
	) name137 (
		_w382_,
		_w385_,
		_w386_
	);
	LUT4 #(
		.INIT('h0e02)
	) name138 (
		\rd1_Key_o_reg[0]/NET0131 ,
		_w250_,
		_w256_,
		_w261_,
		_w387_
	);
	LUT3 #(
		.INIT('h20)
	) name139 (
		\rd1_Key_o_reg[27]/NET0131 ,
		_w250_,
		_w256_,
		_w388_
	);
	LUT3 #(
		.INIT('h54)
	) name140 (
		decrypt_i_pad,
		_w387_,
		_w388_,
		_w389_
	);
	LUT3 #(
		.INIT('hb8)
	) name141 (
		\key_i[44]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[2]/NET0131 ,
		_w390_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w250_,
		_w390_,
		_w391_
	);
	LUT3 #(
		.INIT('h1d)
	) name143 (
		\rd1_Key_o_reg[2]/NET0131 ,
		_w250_,
		_w390_,
		_w392_
	);
	LUT4 #(
		.INIT('he020)
	) name144 (
		\rd1_Key_o_reg[2]/NET0131 ,
		_w250_,
		_w263_,
		_w390_,
		_w393_
	);
	LUT4 #(
		.INIT('hb800)
	) name145 (
		\key_i[52]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[1]/NET0131 ,
		_w250_,
		_w394_
	);
	LUT4 #(
		.INIT('h000d)
	) name146 (
		_w256_,
		_w272_,
		_w394_,
		_w393_,
		_w395_
	);
	LUT3 #(
		.INIT('hce)
	) name147 (
		decrypt_i_pad,
		_w389_,
		_w395_,
		_w396_
	);
	LUT3 #(
		.INIT('hb8)
	) name148 (
		\key_i[55]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[49]/NET0131 ,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w250_,
		_w397_,
		_w398_
	);
	LUT4 #(
		.INIT('he020)
	) name150 (
		\rd1_Key_o_reg[49]/NET0131 ,
		_w250_,
		_w263_,
		_w397_,
		_w399_
	);
	LUT3 #(
		.INIT('hb8)
	) name151 (
		\key_i[63]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[48]/NET0131 ,
		_w400_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w250_,
		_w400_,
		_w401_
	);
	LUT3 #(
		.INIT('hb8)
	) name153 (
		\key_i[47]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[50]/NET0131 ,
		_w402_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		_w250_,
		_w402_,
		_w403_
	);
	LUT4 #(
		.INIT('he020)
	) name155 (
		\rd1_Key_o_reg[50]/NET0131 ,
		_w250_,
		_w256_,
		_w402_,
		_w404_
	);
	LUT4 #(
		.INIT('haaa8)
	) name156 (
		decrypt_i_pad,
		_w401_,
		_w404_,
		_w399_,
		_w405_
	);
	LUT4 #(
		.INIT('h470f)
	) name157 (
		\key_i[6]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[47]/NET0131 ,
		_w250_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		_w263_,
		_w406_,
		_w407_
	);
	LUT4 #(
		.INIT('hb800)
	) name159 (
		\key_i[6]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[47]/NET0131 ,
		_w250_,
		_w408_
	);
	LUT4 #(
		.INIT('h470f)
	) name160 (
		\key_i[14]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[46]/NET0131 ,
		_w250_,
		_w409_
	);
	LUT3 #(
		.INIT('h31)
	) name161 (
		_w256_,
		_w408_,
		_w409_,
		_w410_
	);
	LUT4 #(
		.INIT('h2322)
	) name162 (
		decrypt_i_pad,
		_w405_,
		_w407_,
		_w410_,
		_w411_
	);
	LUT4 #(
		.INIT('hdcdd)
	) name163 (
		decrypt_i_pad,
		_w405_,
		_w407_,
		_w410_,
		_w412_
	);
	LUT4 #(
		.INIT('h470f)
	) name164 (
		\data_i[19]_pad ,
		load_i_pad,
		\rd1_R_o_reg[13]/NET0131 ,
		_w250_,
		_w413_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name165 (
		\data_i[19]_pad ,
		load_i_pad,
		\rd1_R_o_reg[13]/NET0131 ,
		_w250_,
		_w414_
	);
	LUT4 #(
		.INIT('h0e02)
	) name166 (
		\rd1_Key_o_reg[35]/NET0131 ,
		_w250_,
		_w256_,
		_w375_,
		_w415_
	);
	LUT3 #(
		.INIT('h54)
	) name167 (
		decrypt_i_pad,
		_w360_,
		_w415_,
		_w416_
	);
	LUT3 #(
		.INIT('hb8)
	) name168 (
		\key_i[21]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[37]/NET0131 ,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w250_,
		_w417_,
		_w418_
	);
	LUT4 #(
		.INIT('he020)
	) name170 (
		\rd1_Key_o_reg[37]/NET0131 ,
		_w250_,
		_w263_,
		_w417_,
		_w419_
	);
	LUT3 #(
		.INIT('hb8)
	) name171 (
		\key_i[29]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[36]/NET0131 ,
		_w420_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w250_,
		_w420_,
		_w421_
	);
	LUT4 #(
		.INIT('h470f)
	) name173 (
		\key_i[13]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[38]/NET0131 ,
		_w250_,
		_w422_
	);
	LUT4 #(
		.INIT('h0031)
	) name174 (
		_w256_,
		_w421_,
		_w422_,
		_w419_,
		_w423_
	);
	LUT3 #(
		.INIT('hce)
	) name175 (
		decrypt_i_pad,
		_w416_,
		_w423_,
		_w424_
	);
	LUT3 #(
		.INIT('h1d)
	) name176 (
		\rd1_Key_o_reg[48]/NET0131 ,
		_w250_,
		_w400_,
		_w425_
	);
	LUT4 #(
		.INIT('h0415)
	) name177 (
		decrypt_i_pad,
		_w256_,
		_w406_,
		_w425_,
		_w426_
	);
	LUT4 #(
		.INIT('he020)
	) name178 (
		\rd1_Key_o_reg[50]/NET0131 ,
		_w250_,
		_w263_,
		_w402_,
		_w427_
	);
	LUT3 #(
		.INIT('hb8)
	) name179 (
		\key_i[39]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[51]/NET0131 ,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w250_,
		_w428_,
		_w429_
	);
	LUT4 #(
		.INIT('he020)
	) name181 (
		\rd1_Key_o_reg[51]/NET0131 ,
		_w250_,
		_w256_,
		_w428_,
		_w430_
	);
	LUT4 #(
		.INIT('haaa8)
	) name182 (
		decrypt_i_pad,
		_w398_,
		_w430_,
		_w427_,
		_w431_
	);
	LUT2 #(
		.INIT('he)
	) name183 (
		_w426_,
		_w431_,
		_w432_
	);
	LUT3 #(
		.INIT('hb8)
	) name184 (
		\key_i[34]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[15]/NET0131 ,
		_w433_
	);
	LUT4 #(
		.INIT('he020)
	) name185 (
		\rd1_Key_o_reg[15]/NET0131 ,
		_w250_,
		_w256_,
		_w433_,
		_w434_
	);
	LUT3 #(
		.INIT('hb8)
	) name186 (
		\key_i[26]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[16]/NET0131 ,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w250_,
		_w435_,
		_w436_
	);
	LUT4 #(
		.INIT('h0e02)
	) name188 (
		\rd1_Key_o_reg[16]/NET0131 ,
		_w250_,
		_w256_,
		_w435_,
		_w437_
	);
	LUT3 #(
		.INIT('h54)
	) name189 (
		decrypt_i_pad,
		_w434_,
		_w437_,
		_w438_
	);
	LUT3 #(
		.INIT('hb8)
	) name190 (
		\key_i[10]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[18]/NET0131 ,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		_w250_,
		_w439_,
		_w440_
	);
	LUT4 #(
		.INIT('he020)
	) name192 (
		\rd1_Key_o_reg[18]/NET0131 ,
		_w250_,
		_w263_,
		_w439_,
		_w441_
	);
	LUT3 #(
		.INIT('hb8)
	) name193 (
		\key_i[18]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[17]/NET0131 ,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w250_,
		_w442_,
		_w443_
	);
	LUT4 #(
		.INIT('h470f)
	) name195 (
		\key_i[2]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[19]/NET0131 ,
		_w250_,
		_w444_
	);
	LUT4 #(
		.INIT('h0031)
	) name196 (
		_w256_,
		_w443_,
		_w444_,
		_w441_,
		_w445_
	);
	LUT3 #(
		.INIT('hce)
	) name197 (
		decrypt_i_pad,
		_w438_,
		_w445_,
		_w446_
	);
	LUT4 #(
		.INIT('h470f)
	) name198 (
		\data_i[57]_pad ,
		load_i_pad,
		\rd1_R_o_reg[0]/NET0131 ,
		_w250_,
		_w447_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name199 (
		\data_i[57]_pad ,
		load_i_pad,
		\rd1_R_o_reg[0]/NET0131 ,
		_w250_,
		_w448_
	);
	LUT4 #(
		.INIT('h470f)
	) name200 (
		\data_i[61]_pad ,
		load_i_pad,
		\rd1_R_o_reg[16]/NET0131 ,
		_w250_,
		_w449_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name201 (
		\data_i[61]_pad ,
		load_i_pad,
		\rd1_R_o_reg[16]/NET0131 ,
		_w250_,
		_w450_
	);
	LUT3 #(
		.INIT('hb8)
	) name202 (
		\key_i[42]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[14]/NET0131 ,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		_w250_,
		_w451_,
		_w452_
	);
	LUT3 #(
		.INIT('h1d)
	) name204 (
		\rd1_Key_o_reg[14]/NET0131 ,
		_w250_,
		_w451_,
		_w453_
	);
	LUT4 #(
		.INIT('h0415)
	) name205 (
		decrypt_i_pad,
		_w256_,
		_w336_,
		_w453_,
		_w454_
	);
	LUT4 #(
		.INIT('he020)
	) name206 (
		\rd1_Key_o_reg[16]/NET0131 ,
		_w250_,
		_w263_,
		_w435_,
		_w455_
	);
	LUT3 #(
		.INIT('h20)
	) name207 (
		\rd1_Key_o_reg[17]/NET0131 ,
		_w250_,
		_w256_,
		_w456_
	);
	LUT4 #(
		.INIT('h13df)
	) name208 (
		\rd1_Key_o_reg[17]/NET0131 ,
		_w250_,
		_w256_,
		_w433_,
		_w457_
	);
	LUT3 #(
		.INIT('h8a)
	) name209 (
		decrypt_i_pad,
		_w455_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('he)
	) name210 (
		_w454_,
		_w458_,
		_w459_
	);
	LUT4 #(
		.INIT('h470f)
	) name211 (
		\data_i[1]_pad ,
		load_i_pad,
		\rd1_R_o_reg[7]/NET0131 ,
		_w250_,
		_w460_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name212 (
		\data_i[1]_pad ,
		load_i_pad,
		\rd1_R_o_reg[7]/NET0131 ,
		_w250_,
		_w461_
	);
	LUT4 #(
		.INIT('he020)
	) name213 (
		\rd1_Key_o_reg[28]/NET0131 ,
		_w250_,
		_w263_,
		_w288_,
		_w462_
	);
	LUT4 #(
		.INIT('he020)
	) name214 (
		\rd1_Key_o_reg[29]/NET0131 ,
		_w250_,
		_w256_,
		_w299_,
		_w463_
	);
	LUT4 #(
		.INIT('haaa8)
	) name215 (
		decrypt_i_pad,
		_w292_,
		_w463_,
		_w462_,
		_w464_
	);
	LUT4 #(
		.INIT('h470f)
	) name216 (
		\key_i[15]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[54]/NET0131 ,
		_w250_,
		_w465_
	);
	LUT4 #(
		.INIT('hb800)
	) name217 (
		\key_i[15]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[54]/NET0131 ,
		_w250_,
		_w466_
	);
	LUT3 #(
		.INIT('hb8)
	) name218 (
		\key_i[23]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[53]/NET0131 ,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w250_,
		_w467_,
		_w468_
	);
	LUT4 #(
		.INIT('he020)
	) name220 (
		\rd1_Key_o_reg[53]/NET0131 ,
		_w250_,
		_w256_,
		_w467_,
		_w469_
	);
	LUT4 #(
		.INIT('h00f1)
	) name221 (
		_w250_,
		_w263_,
		_w465_,
		_w469_,
		_w470_
	);
	LUT3 #(
		.INIT('hcd)
	) name222 (
		decrypt_i_pad,
		_w464_,
		_w470_,
		_w471_
	);
	LUT3 #(
		.INIT('hb8)
	) name223 (
		\key_i[22]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[45]/NET0131 ,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w250_,
		_w472_,
		_w473_
	);
	LUT4 #(
		.INIT('h0e02)
	) name225 (
		\rd1_Key_o_reg[45]/NET0131 ,
		_w250_,
		_w256_,
		_w472_,
		_w474_
	);
	LUT3 #(
		.INIT('hb8)
	) name226 (
		\key_i[30]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[44]/NET0131 ,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w250_,
		_w475_,
		_w476_
	);
	LUT4 #(
		.INIT('he020)
	) name228 (
		\rd1_Key_o_reg[44]/NET0131 ,
		_w250_,
		_w256_,
		_w475_,
		_w477_
	);
	LUT3 #(
		.INIT('h01)
	) name229 (
		decrypt_i_pad,
		_w477_,
		_w474_,
		_w478_
	);
	LUT4 #(
		.INIT('hb800)
	) name230 (
		\key_i[14]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[46]/NET0131 ,
		_w250_,
		_w479_
	);
	LUT4 #(
		.INIT('he020)
	) name231 (
		\rd1_Key_o_reg[48]/NET0131 ,
		_w250_,
		_w256_,
		_w400_,
		_w480_
	);
	LUT4 #(
		.INIT('h00a2)
	) name232 (
		decrypt_i_pad,
		_w263_,
		_w406_,
		_w480_,
		_w481_
	);
	LUT3 #(
		.INIT('h45)
	) name233 (
		_w478_,
		_w479_,
		_w481_,
		_w482_
	);
	LUT4 #(
		.INIT('h0e02)
	) name234 (
		\rd1_Key_o_reg[36]/NET0131 ,
		_w250_,
		_w256_,
		_w420_,
		_w483_
	);
	LUT3 #(
		.INIT('h54)
	) name235 (
		decrypt_i_pad,
		_w377_,
		_w483_,
		_w484_
	);
	LUT3 #(
		.INIT('hb8)
	) name236 (
		\key_i[5]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[39]/NET0131 ,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w250_,
		_w485_,
		_w486_
	);
	LUT3 #(
		.INIT('h1d)
	) name238 (
		\rd1_Key_o_reg[39]/NET0131 ,
		_w250_,
		_w485_,
		_w487_
	);
	LUT4 #(
		.INIT('he020)
	) name239 (
		\rd1_Key_o_reg[39]/NET0131 ,
		_w250_,
		_w256_,
		_w485_,
		_w488_
	);
	LUT4 #(
		.INIT('h000d)
	) name240 (
		_w263_,
		_w422_,
		_w418_,
		_w488_,
		_w489_
	);
	LUT3 #(
		.INIT('hce)
	) name241 (
		decrypt_i_pad,
		_w484_,
		_w489_,
		_w490_
	);
	LUT4 #(
		.INIT('h470f)
	) name242 (
		\data_i[15]_pad ,
		load_i_pad,
		\rd1_R_o_reg[30]/NET0131 ,
		_w250_,
		_w491_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name243 (
		\data_i[15]_pad ,
		load_i_pad,
		\rd1_R_o_reg[30]/NET0131 ,
		_w250_,
		_w492_
	);
	LUT4 #(
		.INIT('h0e02)
	) name244 (
		\rd1_Key_o_reg[44]/NET0131 ,
		_w250_,
		_w256_,
		_w475_,
		_w493_
	);
	LUT3 #(
		.INIT('hb8)
	) name245 (
		\key_i[38]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[43]/NET0131 ,
		_w494_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w250_,
		_w494_,
		_w495_
	);
	LUT3 #(
		.INIT('h1d)
	) name247 (
		\rd1_Key_o_reg[43]/NET0131 ,
		_w250_,
		_w494_,
		_w496_
	);
	LUT4 #(
		.INIT('he020)
	) name248 (
		\rd1_Key_o_reg[43]/NET0131 ,
		_w250_,
		_w256_,
		_w494_,
		_w497_
	);
	LUT3 #(
		.INIT('h54)
	) name249 (
		decrypt_i_pad,
		_w493_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		_w263_,
		_w409_,
		_w499_
	);
	LUT3 #(
		.INIT('h0d)
	) name251 (
		_w256_,
		_w406_,
		_w473_,
		_w500_
	);
	LUT4 #(
		.INIT('h1311)
	) name252 (
		decrypt_i_pad,
		_w498_,
		_w499_,
		_w500_,
		_w501_
	);
	LUT4 #(
		.INIT('hecee)
	) name253 (
		decrypt_i_pad,
		_w498_,
		_w499_,
		_w500_,
		_w502_
	);
	LUT4 #(
		.INIT('he020)
	) name254 (
		\rd1_Key_o_reg[15]/NET0131 ,
		_w250_,
		_w263_,
		_w433_,
		_w503_
	);
	LUT4 #(
		.INIT('he020)
	) name255 (
		\rd1_Key_o_reg[16]/NET0131 ,
		_w250_,
		_w256_,
		_w435_,
		_w504_
	);
	LUT4 #(
		.INIT('haaa8)
	) name256 (
		decrypt_i_pad,
		_w452_,
		_w504_,
		_w503_,
		_w505_
	);
	LUT4 #(
		.INIT('hb800)
	) name257 (
		\key_i[50]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[13]/NET0131 ,
		_w250_,
		_w506_
	);
	LUT4 #(
		.INIT('hf3e2)
	) name258 (
		_w249_,
		_w256_,
		_w338_,
		_w336_,
		_w507_
	);
	LUT4 #(
		.INIT('h2322)
	) name259 (
		decrypt_i_pad,
		_w505_,
		_w506_,
		_w507_,
		_w508_
	);
	LUT4 #(
		.INIT('hdcdd)
	) name260 (
		decrypt_i_pad,
		_w505_,
		_w506_,
		_w507_,
		_w509_
	);
	LUT4 #(
		.INIT('h470f)
	) name261 (
		\data_i[33]_pad ,
		load_i_pad,
		\rd1_R_o_reg[3]/NET0131 ,
		_w250_,
		_w510_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name262 (
		\data_i[33]_pad ,
		load_i_pad,
		\rd1_R_o_reg[3]/NET0131 ,
		_w250_,
		_w511_
	);
	LUT2 #(
		.INIT('h9)
	) name263 (
		_w508_,
		_w510_,
		_w512_
	);
	LUT4 #(
		.INIT('he020)
	) name264 (
		\rd1_Key_o_reg[7]/NET0131 ,
		_w250_,
		_w263_,
		_w283_,
		_w513_
	);
	LUT4 #(
		.INIT('h0031)
	) name265 (
		_w256_,
		_w278_,
		_w326_,
		_w513_,
		_w514_
	);
	LUT4 #(
		.INIT('he020)
	) name266 (
		\rd1_Key_o_reg[4]/NET0131 ,
		_w250_,
		_w256_,
		_w273_,
		_w515_
	);
	LUT4 #(
		.INIT('h00f1)
	) name267 (
		_w250_,
		_w263_,
		_w281_,
		_w515_,
		_w516_
	);
	LUT3 #(
		.INIT('h27)
	) name268 (
		decrypt_i_pad,
		_w514_,
		_w516_,
		_w517_
	);
	LUT4 #(
		.INIT('h470f)
	) name269 (
		\data_i[41]_pad ,
		load_i_pad,
		\rd1_R_o_reg[2]/NET0131 ,
		_w250_,
		_w518_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name270 (
		\data_i[41]_pad ,
		load_i_pad,
		\rd1_R_o_reg[2]/NET0131 ,
		_w250_,
		_w519_
	);
	LUT4 #(
		.INIT('hd827)
	) name271 (
		decrypt_i_pad,
		_w514_,
		_w516_,
		_w518_,
		_w520_
	);
	LUT3 #(
		.INIT('h06)
	) name272 (
		_w508_,
		_w510_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h9)
	) name273 (
		_w306_,
		_w369_,
		_w522_
	);
	LUT4 #(
		.INIT('he020)
	) name274 (
		\rd1_Key_o_reg[21]/NET0131 ,
		_w250_,
		_w263_,
		_w308_,
		_w523_
	);
	LUT4 #(
		.INIT('he020)
	) name275 (
		\rd1_Key_o_reg[22]/NET0131 ,
		_w250_,
		_w256_,
		_w321_,
		_w524_
	);
	LUT4 #(
		.INIT('haaa8)
	) name276 (
		decrypt_i_pad,
		_w312_,
		_w524_,
		_w523_,
		_w525_
	);
	LUT4 #(
		.INIT('hb800)
	) name277 (
		\key_i[2]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[19]/NET0131 ,
		_w250_,
		_w526_
	);
	LUT4 #(
		.INIT('he020)
	) name278 (
		\rd1_Key_o_reg[18]/NET0131 ,
		_w250_,
		_w256_,
		_w439_,
		_w527_
	);
	LUT4 #(
		.INIT('h00f1)
	) name279 (
		_w250_,
		_w263_,
		_w444_,
		_w527_,
		_w528_
	);
	LUT3 #(
		.INIT('hcd)
	) name280 (
		decrypt_i_pad,
		_w525_,
		_w528_,
		_w529_
	);
	LUT4 #(
		.INIT('h470f)
	) name281 (
		\data_i[49]_pad ,
		load_i_pad,
		\rd1_R_o_reg[1]/NET0131 ,
		_w250_,
		_w530_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name282 (
		\data_i[49]_pad ,
		load_i_pad,
		\rd1_R_o_reg[1]/NET0131 ,
		_w250_,
		_w531_
	);
	LUT4 #(
		.INIT('h32cd)
	) name283 (
		decrypt_i_pad,
		_w525_,
		_w528_,
		_w530_,
		_w532_
	);
	LUT4 #(
		.INIT('h6006)
	) name284 (
		_w306_,
		_w369_,
		_w508_,
		_w510_,
		_w533_
	);
	LUT3 #(
		.INIT('h20)
	) name285 (
		_w520_,
		_w532_,
		_w533_,
		_w534_
	);
	LUT4 #(
		.INIT('hfff6)
	) name286 (
		_w512_,
		_w520_,
		_w522_,
		_w532_,
		_w535_
	);
	LUT3 #(
		.INIT('h09)
	) name287 (
		_w306_,
		_w369_,
		_w520_,
		_w536_
	);
	LUT3 #(
		.INIT('h90)
	) name288 (
		_w508_,
		_w510_,
		_w532_,
		_w537_
	);
	LUT4 #(
		.INIT('h0900)
	) name289 (
		_w508_,
		_w510_,
		_w520_,
		_w532_,
		_w538_
	);
	LUT4 #(
		.INIT('h0990)
	) name290 (
		_w306_,
		_w369_,
		_w508_,
		_w510_,
		_w539_
	);
	LUT3 #(
		.INIT('h54)
	) name291 (
		_w536_,
		_w538_,
		_w539_,
		_w540_
	);
	LUT4 #(
		.INIT('h31ce)
	) name292 (
		decrypt_i_pad,
		_w260_,
		_w268_,
		_w447_,
		_w541_
	);
	LUT3 #(
		.INIT('hd0)
	) name293 (
		_w535_,
		_w540_,
		_w541_,
		_w542_
	);
	LUT3 #(
		.INIT('h90)
	) name294 (
		_w306_,
		_w369_,
		_w520_,
		_w543_
	);
	LUT4 #(
		.INIT('h0090)
	) name295 (
		_w306_,
		_w369_,
		_w520_,
		_w541_,
		_w544_
	);
	LUT3 #(
		.INIT('h8c)
	) name296 (
		_w520_,
		_w532_,
		_w541_,
		_w545_
	);
	LUT3 #(
		.INIT('hd0)
	) name297 (
		_w512_,
		_w544_,
		_w545_,
		_w546_
	);
	LUT4 #(
		.INIT('h090f)
	) name298 (
		_w306_,
		_w369_,
		_w532_,
		_w541_,
		_w547_
	);
	LUT4 #(
		.INIT('h000d)
	) name299 (
		_w263_,
		_w316_,
		_w384_,
		_w524_,
		_w548_
	);
	LUT4 #(
		.INIT('he200)
	) name300 (
		\rd1_Key_o_reg[25]/NET0131 ,
		_w250_,
		_w258_,
		_w263_,
		_w549_
	);
	LUT4 #(
		.INIT('he200)
	) name301 (
		\rd1_Key_o_reg[26]/NET0131 ,
		_w250_,
		_w254_,
		_w256_,
		_w550_
	);
	LUT4 #(
		.INIT('haaa8)
	) name302 (
		decrypt_i_pad,
		_w318_,
		_w550_,
		_w549_,
		_w551_
	);
	LUT3 #(
		.INIT('hf1)
	) name303 (
		decrypt_i_pad,
		_w548_,
		_w551_,
		_w552_
	);
	LUT4 #(
		.INIT('h470f)
	) name304 (
		\data_i[7]_pad ,
		load_i_pad,
		\rd1_R_o_reg[31]/NET0131 ,
		_w250_,
		_w553_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name305 (
		\data_i[7]_pad ,
		load_i_pad,
		\rd1_R_o_reg[31]/NET0131 ,
		_w250_,
		_w554_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name306 (
		decrypt_i_pad,
		_w548_,
		_w551_,
		_w553_,
		_w555_
	);
	LUT4 #(
		.INIT('h00df)
	) name307 (
		_w512_,
		_w544_,
		_w547_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		_w546_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w542_,
		_w557_,
		_w558_
	);
	LUT3 #(
		.INIT('h70)
	) name310 (
		_w520_,
		_w533_,
		_w541_,
		_w559_
	);
	LUT4 #(
		.INIT('h4ee4)
	) name311 (
		_w512_,
		_w520_,
		_w522_,
		_w532_,
		_w560_
	);
	LUT3 #(
		.INIT('h80)
	) name312 (
		_w535_,
		_w559_,
		_w560_,
		_w561_
	);
	LUT3 #(
		.INIT('h90)
	) name313 (
		_w306_,
		_w369_,
		_w532_,
		_w562_
	);
	LUT3 #(
		.INIT('h02)
	) name314 (
		_w520_,
		_w533_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w538_,
		_w541_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		_w563_,
		_w564_,
		_w565_
	);
	LUT4 #(
		.INIT('h0009)
	) name317 (
		_w306_,
		_w369_,
		_w520_,
		_w532_,
		_w566_
	);
	LUT3 #(
		.INIT('h8c)
	) name318 (
		_w512_,
		_w555_,
		_w566_,
		_w567_
	);
	LUT3 #(
		.INIT('he0)
	) name319 (
		_w561_,
		_w565_,
		_w567_,
		_w568_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name320 (
		\data_i[16]_pad ,
		load_i_pad,
		\rd1_L_o_reg[5]/NET0131 ,
		_w250_,
		_w569_
	);
	LUT3 #(
		.INIT('he1)
	) name321 (
		_w558_,
		_w568_,
		_w569_,
		_w570_
	);
	LUT4 #(
		.INIT('h470f)
	) name322 (
		\key_i[46]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[42]/NET0131 ,
		_w250_,
		_w571_
	);
	LUT4 #(
		.INIT('hb800)
	) name323 (
		\key_i[46]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[42]/NET0131 ,
		_w250_,
		_w572_
	);
	LUT3 #(
		.INIT('hb8)
	) name324 (
		\key_i[54]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[41]/NET0131 ,
		_w573_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w250_,
		_w573_,
		_w574_
	);
	LUT4 #(
		.INIT('he020)
	) name326 (
		\rd1_Key_o_reg[41]/NET0131 ,
		_w250_,
		_w256_,
		_w573_,
		_w575_
	);
	LUT4 #(
		.INIT('h000d)
	) name327 (
		_w263_,
		_w571_,
		_w572_,
		_w575_,
		_w576_
	);
	LUT4 #(
		.INIT('he020)
	) name328 (
		\rd1_Key_o_reg[44]/NET0131 ,
		_w250_,
		_w263_,
		_w475_,
		_w577_
	);
	LUT4 #(
		.INIT('he020)
	) name329 (
		\rd1_Key_o_reg[45]/NET0131 ,
		_w250_,
		_w256_,
		_w472_,
		_w578_
	);
	LUT4 #(
		.INIT('haaa8)
	) name330 (
		decrypt_i_pad,
		_w495_,
		_w578_,
		_w577_,
		_w579_
	);
	LUT3 #(
		.INIT('hf1)
	) name331 (
		decrypt_i_pad,
		_w576_,
		_w579_,
		_w580_
	);
	LUT4 #(
		.INIT('h33c9)
	) name332 (
		decrypt_i_pad,
		_w449_,
		_w576_,
		_w579_,
		_w581_
	);
	LUT4 #(
		.INIT('h470f)
	) name333 (
		\data_i[53]_pad ,
		load_i_pad,
		\rd1_R_o_reg[17]/NET0131 ,
		_w250_,
		_w582_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name334 (
		\data_i[53]_pad ,
		load_i_pad,
		\rd1_R_o_reg[17]/NET0131 ,
		_w250_,
		_w583_
	);
	LUT4 #(
		.INIT('h31ce)
	) name335 (
		decrypt_i_pad,
		_w416_,
		_w423_,
		_w582_,
		_w584_
	);
	LUT4 #(
		.INIT('h470f)
	) name336 (
		\data_i[37]_pad ,
		load_i_pad,
		\rd1_R_o_reg[19]/NET0131 ,
		_w250_,
		_w585_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name337 (
		\data_i[37]_pad ,
		load_i_pad,
		\rd1_R_o_reg[19]/NET0131 ,
		_w250_,
		_w586_
	);
	LUT3 #(
		.INIT('h1e)
	) name338 (
		_w426_,
		_w431_,
		_w585_,
		_w587_
	);
	LUT4 #(
		.INIT('h0415)
	) name339 (
		decrypt_i_pad,
		_w256_,
		_w422_,
		_w487_,
		_w588_
	);
	LUT4 #(
		.INIT('he020)
	) name340 (
		\rd1_Key_o_reg[41]/NET0131 ,
		_w250_,
		_w263_,
		_w573_,
		_w589_
	);
	LUT3 #(
		.INIT('hb8)
	) name341 (
		\key_i[62]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[40]/NET0131 ,
		_w590_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		_w250_,
		_w590_,
		_w591_
	);
	LUT4 #(
		.INIT('h0031)
	) name343 (
		_w256_,
		_w591_,
		_w571_,
		_w589_,
		_w592_
	);
	LUT3 #(
		.INIT('hce)
	) name344 (
		decrypt_i_pad,
		_w588_,
		_w592_,
		_w593_
	);
	LUT4 #(
		.INIT('h470f)
	) name345 (
		\data_i[29]_pad ,
		load_i_pad,
		\rd1_R_o_reg[20]/NET0131 ,
		_w250_,
		_w594_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name346 (
		\data_i[29]_pad ,
		load_i_pad,
		\rd1_R_o_reg[20]/NET0131 ,
		_w250_,
		_w595_
	);
	LUT4 #(
		.INIT('h31ce)
	) name347 (
		decrypt_i_pad,
		_w588_,
		_w592_,
		_w594_,
		_w596_
	);
	LUT4 #(
		.INIT('h470f)
	) name348 (
		\data_i[45]_pad ,
		load_i_pad,
		\rd1_R_o_reg[18]/NET0131 ,
		_w250_,
		_w597_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name349 (
		\data_i[45]_pad ,
		load_i_pad,
		\rd1_R_o_reg[18]/NET0131 ,
		_w250_,
		_w598_
	);
	LUT3 #(
		.INIT('h1e)
	) name350 (
		_w295_,
		_w304_,
		_w597_,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w599_,
		_w584_,
		_w600_
	);
	LUT4 #(
		.INIT('h3eef)
	) name352 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w601_
	);
	LUT4 #(
		.INIT('h4004)
	) name353 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w602_
	);
	LUT3 #(
		.INIT('hd6)
	) name354 (
		_w599_,
		_w587_,
		_w596_,
		_w603_
	);
	LUT4 #(
		.INIT('h5404)
	) name355 (
		_w602_,
		_w603_,
		_w581_,
		_w601_,
		_w604_
	);
	LUT4 #(
		.INIT('h0e02)
	) name356 (
		\rd1_Key_o_reg[53]/NET0131 ,
		_w250_,
		_w256_,
		_w467_,
		_w605_
	);
	LUT3 #(
		.INIT('hb8)
	) name357 (
		\key_i[31]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[52]/NET0131 ,
		_w606_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		_w250_,
		_w606_,
		_w607_
	);
	LUT4 #(
		.INIT('he020)
	) name359 (
		\rd1_Key_o_reg[52]/NET0131 ,
		_w250_,
		_w256_,
		_w606_,
		_w608_
	);
	LUT3 #(
		.INIT('h54)
	) name360 (
		decrypt_i_pad,
		_w605_,
		_w608_,
		_w609_
	);
	LUT4 #(
		.INIT('he020)
	) name361 (
		\rd1_Key_o_reg[55]/NET0131 ,
		_w250_,
		_w263_,
		_w291_,
		_w610_
	);
	LUT4 #(
		.INIT('haaa8)
	) name362 (
		decrypt_i_pad,
		_w345_,
		_w466_,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('he)
	) name363 (
		_w609_,
		_w611_,
		_w612_
	);
	LUT4 #(
		.INIT('h470f)
	) name364 (
		\data_i[3]_pad ,
		load_i_pad,
		\rd1_R_o_reg[15]/NET0131 ,
		_w250_,
		_w613_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name365 (
		\data_i[3]_pad ,
		load_i_pad,
		\rd1_R_o_reg[15]/NET0131 ,
		_w250_,
		_w614_
	);
	LUT3 #(
		.INIT('h1e)
	) name366 (
		_w609_,
		_w611_,
		_w613_,
		_w615_
	);
	LUT2 #(
		.INIT('h4)
	) name367 (
		_w604_,
		_w615_,
		_w616_
	);
	LUT4 #(
		.INIT('hf15c)
	) name368 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w617_
	);
	LUT3 #(
		.INIT('h04)
	) name369 (
		_w599_,
		_w584_,
		_w596_,
		_w618_
	);
	LUT4 #(
		.INIT('h1000)
	) name370 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w619_
	);
	LUT4 #(
		.INIT('h00b1)
	) name371 (
		_w581_,
		_w618_,
		_w617_,
		_w619_,
		_w620_
	);
	LUT4 #(
		.INIT('haffc)
	) name372 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w621_
	);
	LUT3 #(
		.INIT('h02)
	) name373 (
		_w581_,
		_w600_,
		_w621_,
		_w622_
	);
	LUT4 #(
		.INIT('h0800)
	) name374 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w623_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		_w599_,
		_w584_,
		_w624_
	);
	LUT4 #(
		.INIT('hdfd3)
	) name376 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w625_
	);
	LUT3 #(
		.INIT('h32)
	) name377 (
		_w581_,
		_w623_,
		_w625_,
		_w626_
	);
	LUT4 #(
		.INIT('h0e00)
	) name378 (
		_w615_,
		_w620_,
		_w622_,
		_w626_,
		_w627_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name379 (
		\data_i[8]_pad ,
		load_i_pad,
		\rd1_L_o_reg[6]/NET0131 ,
		_w250_,
		_w628_
	);
	LUT3 #(
		.INIT('hb4)
	) name380 (
		_w616_,
		_w627_,
		_w628_,
		_w629_
	);
	LUT4 #(
		.INIT('h0e02)
	) name381 (
		\rd1_Key_o_reg[25]/NET0131 ,
		_w250_,
		_w256_,
		_w258_,
		_w630_
	);
	LUT3 #(
		.INIT('h54)
	) name382 (
		decrypt_i_pad,
		_w320_,
		_w630_,
		_w631_
	);
	LUT4 #(
		.INIT('he200)
	) name383 (
		\rd1_Key_o_reg[27]/NET0131 ,
		_w250_,
		_w265_,
		_w263_,
		_w632_
	);
	LUT4 #(
		.INIT('he020)
	) name384 (
		\rd1_Key_o_reg[0]/NET0131 ,
		_w250_,
		_w256_,
		_w261_,
		_w633_
	);
	LUT4 #(
		.INIT('haaa8)
	) name385 (
		decrypt_i_pad,
		_w255_,
		_w633_,
		_w632_,
		_w634_
	);
	LUT2 #(
		.INIT('he)
	) name386 (
		_w631_,
		_w634_,
		_w635_
	);
	LUT4 #(
		.INIT('h0e02)
	) name387 (
		\rd1_Key_o_reg[50]/NET0131 ,
		_w250_,
		_w256_,
		_w402_,
		_w636_
	);
	LUT4 #(
		.INIT('he020)
	) name388 (
		\rd1_Key_o_reg[49]/NET0131 ,
		_w250_,
		_w256_,
		_w397_,
		_w637_
	);
	LUT3 #(
		.INIT('h54)
	) name389 (
		decrypt_i_pad,
		_w636_,
		_w637_,
		_w638_
	);
	LUT4 #(
		.INIT('he020)
	) name390 (
		\rd1_Key_o_reg[52]/NET0131 ,
		_w250_,
		_w263_,
		_w606_,
		_w639_
	);
	LUT4 #(
		.INIT('haaa8)
	) name391 (
		decrypt_i_pad,
		_w429_,
		_w469_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('he)
	) name392 (
		_w638_,
		_w640_,
		_w641_
	);
	LUT4 #(
		.INIT('h0e02)
	) name393 (
		\rd1_Key_o_reg[18]/NET0131 ,
		_w250_,
		_w256_,
		_w439_,
		_w642_
	);
	LUT3 #(
		.INIT('h54)
	) name394 (
		decrypt_i_pad,
		_w456_,
		_w642_,
		_w643_
	);
	LUT4 #(
		.INIT('he020)
	) name395 (
		\rd1_Key_o_reg[20]/NET0131 ,
		_w250_,
		_w263_,
		_w311_,
		_w644_
	);
	LUT4 #(
		.INIT('haaa8)
	) name396 (
		decrypt_i_pad,
		_w381_,
		_w526_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('he)
	) name397 (
		_w643_,
		_w645_,
		_w646_
	);
	LUT4 #(
		.INIT('he020)
	) name398 (
		\rd1_Key_o_reg[6]/NET0131 ,
		_w250_,
		_w256_,
		_w277_,
		_w647_
	);
	LUT4 #(
		.INIT('h0031)
	) name399 (
		_w263_,
		_w274_,
		_w281_,
		_w647_,
		_w648_
	);
	LUT4 #(
		.INIT('hb800)
	) name400 (
		\key_i[36]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[3]/NET0131 ,
		_w250_,
		_w649_
	);
	LUT4 #(
		.INIT('he020)
	) name401 (
		\rd1_Key_o_reg[2]/NET0131 ,
		_w250_,
		_w256_,
		_w390_,
		_w650_
	);
	LUT4 #(
		.INIT('h00f1)
	) name402 (
		_w250_,
		_w263_,
		_w272_,
		_w650_,
		_w651_
	);
	LUT3 #(
		.INIT('h27)
	) name403 (
		decrypt_i_pad,
		_w648_,
		_w651_,
		_w652_
	);
	LUT4 #(
		.INIT('h470f)
	) name404 (
		\data_i[31]_pad ,
		load_i_pad,
		\rd1_R_o_reg[28]/NET0131 ,
		_w250_,
		_w653_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name405 (
		\data_i[31]_pad ,
		load_i_pad,
		\rd1_R_o_reg[28]/NET0131 ,
		_w250_,
		_w654_
	);
	LUT4 #(
		.INIT('h0e02)
	) name406 (
		\rd1_Key_o_reg[52]/NET0131 ,
		_w250_,
		_w256_,
		_w606_,
		_w655_
	);
	LUT3 #(
		.INIT('h54)
	) name407 (
		decrypt_i_pad,
		_w430_,
		_w655_,
		_w656_
	);
	LUT4 #(
		.INIT('h0031)
	) name408 (
		_w263_,
		_w294_,
		_w465_,
		_w468_,
		_w657_
	);
	LUT3 #(
		.INIT('hce)
	) name409 (
		decrypt_i_pad,
		_w656_,
		_w657_,
		_w658_
	);
	LUT4 #(
		.INIT('h0e02)
	) name410 (
		\rd1_Key_o_reg[40]/NET0131 ,
		_w250_,
		_w256_,
		_w590_,
		_w659_
	);
	LUT3 #(
		.INIT('h54)
	) name411 (
		decrypt_i_pad,
		_w488_,
		_w659_,
		_w660_
	);
	LUT4 #(
		.INIT('h0031)
	) name412 (
		_w263_,
		_w497_,
		_w571_,
		_w574_,
		_w661_
	);
	LUT3 #(
		.INIT('hce)
	) name413 (
		decrypt_i_pad,
		_w660_,
		_w661_,
		_w662_
	);
	LUT4 #(
		.INIT('h470f)
	) name414 (
		\data_i[47]_pad ,
		load_i_pad,
		\rd1_R_o_reg[26]/NET0131 ,
		_w250_,
		_w663_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name415 (
		\data_i[47]_pad ,
		load_i_pad,
		\rd1_R_o_reg[26]/NET0131 ,
		_w250_,
		_w664_
	);
	LUT3 #(
		.INIT('h56)
	) name416 (
		_w449_,
		_w454_,
		_w458_,
		_w665_
	);
	LUT4 #(
		.INIT('hc693)
	) name417 (
		decrypt_i_pad,
		_w613_,
		_w648_,
		_w651_,
		_w666_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		_w665_,
		_w666_,
		_w667_
	);
	LUT3 #(
		.INIT('h56)
	) name419 (
		_w413_,
		_w643_,
		_w645_,
		_w668_
	);
	LUT4 #(
		.INIT('h0145)
	) name420 (
		decrypt_i_pad,
		_w256_,
		_w319_,
		_w316_,
		_w669_
	);
	LUT4 #(
		.INIT('he200)
	) name421 (
		\rd1_Key_o_reg[26]/NET0131 ,
		_w250_,
		_w254_,
		_w263_,
		_w670_
	);
	LUT4 #(
		.INIT('h13df)
	) name422 (
		\rd1_Key_o_reg[27]/NET0131 ,
		_w250_,
		_w256_,
		_w258_,
		_w671_
	);
	LUT3 #(
		.INIT('h8a)
	) name423 (
		decrypt_i_pad,
		_w670_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('he)
	) name424 (
		_w669_,
		_w672_,
		_w673_
	);
	LUT4 #(
		.INIT('h470f)
	) name425 (
		\data_i[11]_pad ,
		load_i_pad,
		\rd1_R_o_reg[14]/NET0131 ,
		_w250_,
		_w674_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name426 (
		\data_i[11]_pad ,
		load_i_pad,
		\rd1_R_o_reg[14]/NET0131 ,
		_w250_,
		_w675_
	);
	LUT3 #(
		.INIT('h1e)
	) name427 (
		_w669_,
		_w672_,
		_w674_,
		_w676_
	);
	LUT4 #(
		.INIT('h0046)
	) name428 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w677_
	);
	LUT3 #(
		.INIT('h20)
	) name429 (
		_w666_,
		_w668_,
		_w676_,
		_w678_
	);
	LUT4 #(
		.INIT('hb800)
	) name430 (
		\key_i[27]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[8]/NET0131 ,
		_w250_,
		_w679_
	);
	LUT4 #(
		.INIT('h0031)
	) name431 (
		_w263_,
		_w285_,
		_w326_,
		_w679_,
		_w680_
	);
	LUT4 #(
		.INIT('he020)
	) name432 (
		\rd1_Key_o_reg[10]/NET0131 ,
		_w250_,
		_w263_,
		_w332_,
		_w681_
	);
	LUT4 #(
		.INIT('he020)
	) name433 (
		\rd1_Key_o_reg[11]/NET0131 ,
		_w250_,
		_w256_,
		_w339_,
		_w682_
	);
	LUT4 #(
		.INIT('haaa8)
	) name434 (
		decrypt_i_pad,
		_w365_,
		_w682_,
		_w681_,
		_w683_
	);
	LUT3 #(
		.INIT('hf1)
	) name435 (
		decrypt_i_pad,
		_w680_,
		_w683_,
		_w684_
	);
	LUT4 #(
		.INIT('h470f)
	) name436 (
		\data_i[27]_pad ,
		load_i_pad,
		\rd1_R_o_reg[12]/NET0131 ,
		_w250_,
		_w685_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name437 (
		\data_i[27]_pad ,
		load_i_pad,
		\rd1_R_o_reg[12]/NET0131 ,
		_w250_,
		_w686_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name438 (
		decrypt_i_pad,
		_w680_,
		_w683_,
		_w685_,
		_w687_
	);
	LUT4 #(
		.INIT('h5455)
	) name439 (
		_w687_,
		_w665_,
		_w666_,
		_w668_,
		_w688_
	);
	LUT3 #(
		.INIT('h10)
	) name440 (
		_w677_,
		_w678_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h4)
	) name441 (
		_w666_,
		_w676_,
		_w690_
	);
	LUT4 #(
		.INIT('ha280)
	) name442 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w691_
	);
	LUT4 #(
		.INIT('haa2a)
	) name443 (
		_w687_,
		_w665_,
		_w666_,
		_w676_,
		_w692_
	);
	LUT4 #(
		.INIT('h0001)
	) name444 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w693_
	);
	LUT3 #(
		.INIT('h02)
	) name445 (
		_w692_,
		_w691_,
		_w693_,
		_w694_
	);
	LUT4 #(
		.INIT('hfb7f)
	) name446 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w695_
	);
	LUT4 #(
		.INIT('h470f)
	) name447 (
		\data_i[35]_pad ,
		load_i_pad,
		\rd1_R_o_reg[11]/NET0131 ,
		_w250_,
		_w696_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name448 (
		\data_i[35]_pad ,
		load_i_pad,
		\rd1_R_o_reg[11]/NET0131 ,
		_w250_,
		_w697_
	);
	LUT4 #(
		.INIT('h31ce)
	) name449 (
		decrypt_i_pad,
		_w389_,
		_w395_,
		_w696_,
		_w698_
	);
	LUT4 #(
		.INIT('h001f)
	) name450 (
		_w689_,
		_w694_,
		_w695_,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w665_,
		_w676_,
		_w700_
	);
	LUT4 #(
		.INIT('h0008)
	) name452 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w701_
	);
	LUT4 #(
		.INIT('h5cf6)
	) name453 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w702_
	);
	LUT4 #(
		.INIT('h0040)
	) name454 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w703_
	);
	LUT4 #(
		.INIT('h5504)
	) name455 (
		_w687_,
		_w698_,
		_w702_,
		_w703_,
		_w704_
	);
	LUT4 #(
		.INIT('ha020)
	) name456 (
		_w687_,
		_w666_,
		_w668_,
		_w676_,
		_w705_
	);
	LUT4 #(
		.INIT('h082e)
	) name457 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w706_
	);
	LUT4 #(
		.INIT('h23af)
	) name458 (
		_w665_,
		_w692_,
		_w705_,
		_w706_,
		_w707_
	);
	LUT3 #(
		.INIT('h80)
	) name459 (
		_w665_,
		_w666_,
		_w668_,
		_w708_
	);
	LUT2 #(
		.INIT('h2)
	) name460 (
		_w687_,
		_w676_,
		_w709_
	);
	LUT3 #(
		.INIT('h47)
	) name461 (
		_w687_,
		_w668_,
		_w698_,
		_w710_
	);
	LUT3 #(
		.INIT('h10)
	) name462 (
		_w665_,
		_w666_,
		_w676_,
		_w711_
	);
	LUT4 #(
		.INIT('h7077)
	) name463 (
		_w708_,
		_w709_,
		_w710_,
		_w711_,
		_w712_
	);
	LUT4 #(
		.INIT('h3100)
	) name464 (
		_w698_,
		_w704_,
		_w707_,
		_w712_,
		_w713_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name465 (
		\data_i[44]_pad ,
		load_i_pad,
		\rd1_L_o_reg[18]/NET0131 ,
		_w250_,
		_w714_
	);
	LUT3 #(
		.INIT('h4b)
	) name466 (
		_w699_,
		_w713_,
		_w714_,
		_w715_
	);
	LUT4 #(
		.INIT('h470f)
	) name467 (
		\data_i[59]_pad ,
		load_i_pad,
		\rd1_R_o_reg[8]/NET0131 ,
		_w250_,
		_w716_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name468 (
		\data_i[59]_pad ,
		load_i_pad,
		\rd1_R_o_reg[8]/NET0131 ,
		_w250_,
		_w717_
	);
	LUT4 #(
		.INIT('h0e02)
	) name469 (
		\rd1_Key_o_reg[11]/NET0131 ,
		_w250_,
		_w256_,
		_w339_,
		_w718_
	);
	LUT4 #(
		.INIT('he020)
	) name470 (
		\rd1_Key_o_reg[10]/NET0131 ,
		_w250_,
		_w256_,
		_w332_,
		_w719_
	);
	LUT3 #(
		.INIT('h54)
	) name471 (
		decrypt_i_pad,
		_w718_,
		_w719_,
		_w720_
	);
	LUT4 #(
		.INIT('hb800)
	) name472 (
		\key_i[58]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[12]/NET0131 ,
		_w250_,
		_w721_
	);
	LUT4 #(
		.INIT('he020)
	) name473 (
		\rd1_Key_o_reg[14]/NET0131 ,
		_w250_,
		_w256_,
		_w451_,
		_w722_
	);
	LUT4 #(
		.INIT('h000d)
	) name474 (
		_w263_,
		_w336_,
		_w721_,
		_w722_,
		_w723_
	);
	LUT3 #(
		.INIT('hce)
	) name475 (
		decrypt_i_pad,
		_w720_,
		_w723_,
		_w724_
	);
	LUT4 #(
		.INIT('h0e02)
	) name476 (
		\rd1_Key_o_reg[15]/NET0131 ,
		_w250_,
		_w256_,
		_w433_,
		_w725_
	);
	LUT3 #(
		.INIT('h54)
	) name477 (
		decrypt_i_pad,
		_w722_,
		_w725_,
		_w726_
	);
	LUT4 #(
		.INIT('he020)
	) name478 (
		\rd1_Key_o_reg[17]/NET0131 ,
		_w250_,
		_w263_,
		_w442_,
		_w727_
	);
	LUT4 #(
		.INIT('haaa8)
	) name479 (
		decrypt_i_pad,
		_w436_,
		_w527_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('he)
	) name480 (
		_w726_,
		_w728_,
		_w729_
	);
	LUT4 #(
		.INIT('h0e02)
	) name481 (
		\rd1_Key_o_reg[7]/NET0131 ,
		_w250_,
		_w256_,
		_w283_,
		_w730_
	);
	LUT3 #(
		.INIT('h54)
	) name482 (
		decrypt_i_pad,
		_w647_,
		_w730_,
		_w731_
	);
	LUT4 #(
		.INIT('h000d)
	) name483 (
		_w263_,
		_w328_,
		_w679_,
		_w719_,
		_w732_
	);
	LUT3 #(
		.INIT('hce)
	) name484 (
		decrypt_i_pad,
		_w731_,
		_w732_,
		_w733_
	);
	LUT4 #(
		.INIT('h470f)
	) name485 (
		\data_i[5]_pad ,
		load_i_pad,
		\rd1_R_o_reg[23]/NET0131 ,
		_w250_,
		_w734_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name486 (
		\data_i[5]_pad ,
		load_i_pad,
		\rd1_R_o_reg[23]/NET0131 ,
		_w250_,
		_w735_
	);
	LUT4 #(
		.INIT('hba45)
	) name487 (
		_w478_,
		_w479_,
		_w481_,
		_w734_,
		_w736_
	);
	LUT4 #(
		.INIT('h3c36)
	) name488 (
		decrypt_i_pad,
		_w653_,
		_w656_,
		_w657_,
		_w737_
	);
	LUT4 #(
		.INIT('h31ce)
	) name489 (
		decrypt_i_pad,
		_w660_,
		_w661_,
		_w663_,
		_w738_
	);
	LUT4 #(
		.INIT('h0145)
	) name490 (
		decrypt_i_pad,
		_w256_,
		_w293_,
		_w465_,
		_w739_
	);
	LUT4 #(
		.INIT('he020)
	) name491 (
		\rd1_Key_o_reg[29]/NET0131 ,
		_w250_,
		_w263_,
		_w299_,
		_w740_
	);
	LUT4 #(
		.INIT('haaa8)
	) name492 (
		decrypt_i_pad,
		_w289_,
		_w354_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('he)
	) name493 (
		_w739_,
		_w741_,
		_w742_
	);
	LUT4 #(
		.INIT('h470f)
	) name494 (
		\data_i[39]_pad ,
		load_i_pad,
		\rd1_R_o_reg[27]/NET0131 ,
		_w250_,
		_w743_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name495 (
		\data_i[39]_pad ,
		load_i_pad,
		\rd1_R_o_reg[27]/NET0131 ,
		_w250_,
		_w744_
	);
	LUT3 #(
		.INIT('h1e)
	) name496 (
		_w739_,
		_w741_,
		_w743_,
		_w745_
	);
	LUT4 #(
		.INIT('h0e02)
	) name497 (
		\rd1_Key_o_reg[49]/NET0131 ,
		_w250_,
		_w256_,
		_w397_,
		_w746_
	);
	LUT3 #(
		.INIT('h54)
	) name498 (
		decrypt_i_pad,
		_w480_,
		_w746_,
		_w747_
	);
	LUT4 #(
		.INIT('he020)
	) name499 (
		\rd1_Key_o_reg[51]/NET0131 ,
		_w250_,
		_w263_,
		_w428_,
		_w748_
	);
	LUT4 #(
		.INIT('haaa8)
	) name500 (
		decrypt_i_pad,
		_w403_,
		_w608_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('he)
	) name501 (
		_w747_,
		_w749_,
		_w750_
	);
	LUT4 #(
		.INIT('h470f)
	) name502 (
		\data_i[55]_pad ,
		load_i_pad,
		\rd1_R_o_reg[25]/NET0131 ,
		_w250_,
		_w751_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name503 (
		\data_i[55]_pad ,
		load_i_pad,
		\rd1_R_o_reg[25]/NET0131 ,
		_w250_,
		_w752_
	);
	LUT3 #(
		.INIT('h1e)
	) name504 (
		_w747_,
		_w749_,
		_w751_,
		_w753_
	);
	LUT4 #(
		.INIT('hfe3e)
	) name505 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w754_
	);
	LUT3 #(
		.INIT('h08)
	) name506 (
		_w753_,
		_w738_,
		_w737_,
		_w755_
	);
	LUT4 #(
		.INIT('hf638)
	) name507 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w756_
	);
	LUT3 #(
		.INIT('h80)
	) name508 (
		_w738_,
		_w745_,
		_w737_,
		_w757_
	);
	LUT4 #(
		.INIT('h4000)
	) name509 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w758_
	);
	LUT4 #(
		.INIT('h0145)
	) name510 (
		decrypt_i_pad,
		_w256_,
		_w359_,
		_w356_,
		_w759_
	);
	LUT4 #(
		.INIT('he020)
	) name511 (
		\rd1_Key_o_reg[36]/NET0131 ,
		_w250_,
		_w263_,
		_w420_,
		_w760_
	);
	LUT4 #(
		.INIT('he020)
	) name512 (
		\rd1_Key_o_reg[37]/NET0131 ,
		_w250_,
		_w256_,
		_w417_,
		_w761_
	);
	LUT4 #(
		.INIT('haaa8)
	) name513 (
		decrypt_i_pad,
		_w376_,
		_w761_,
		_w760_,
		_w762_
	);
	LUT2 #(
		.INIT('he)
	) name514 (
		_w759_,
		_w762_,
		_w763_
	);
	LUT4 #(
		.INIT('h470f)
	) name515 (
		\data_i[63]_pad ,
		load_i_pad,
		\rd1_R_o_reg[24]/NET0131 ,
		_w250_,
		_w764_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name516 (
		\data_i[63]_pad ,
		load_i_pad,
		\rd1_R_o_reg[24]/NET0131 ,
		_w250_,
		_w765_
	);
	LUT3 #(
		.INIT('h1e)
	) name517 (
		_w759_,
		_w762_,
		_w764_,
		_w766_
	);
	LUT4 #(
		.INIT('h00f2)
	) name518 (
		_w736_,
		_w756_,
		_w758_,
		_w766_,
		_w767_
	);
	LUT3 #(
		.INIT('h07)
	) name519 (
		_w753_,
		_w738_,
		_w766_,
		_w768_
	);
	LUT3 #(
		.INIT('he4)
	) name520 (
		_w738_,
		_w745_,
		_w737_,
		_w769_
	);
	LUT4 #(
		.INIT('h0008)
	) name521 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w770_
	);
	LUT4 #(
		.INIT('h1200)
	) name522 (
		_w738_,
		_w745_,
		_w737_,
		_w766_,
		_w771_
	);
	LUT4 #(
		.INIT('h0111)
	) name523 (
		_w770_,
		_w771_,
		_w768_,
		_w769_,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w736_,
		_w772_,
		_w773_
	);
	LUT4 #(
		.INIT('h0040)
	) name525 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w774_
	);
	LUT4 #(
		.INIT('h5f9e)
	) name526 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w775_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		_w766_,
		_w775_,
		_w776_
	);
	LUT4 #(
		.INIT('h2000)
	) name528 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w777_
	);
	LUT4 #(
		.INIT('h4000)
	) name529 (
		_w738_,
		_w745_,
		_w737_,
		_w766_,
		_w778_
	);
	LUT4 #(
		.INIT('h1000)
	) name530 (
		_w753_,
		_w745_,
		_w737_,
		_w766_,
		_w779_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name531 (
		_w738_,
		_w736_,
		_w778_,
		_w779_,
		_w780_
	);
	LUT3 #(
		.INIT('h01)
	) name532 (
		_w777_,
		_w780_,
		_w776_,
		_w781_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name533 (
		\data_i[14]_pad ,
		load_i_pad,
		\rd1_L_o_reg[30]/NET0131 ,
		_w250_,
		_w782_
	);
	LUT4 #(
		.INIT('h10ef)
	) name534 (
		_w767_,
		_w773_,
		_w781_,
		_w782_,
		_w783_
	);
	LUT4 #(
		.INIT('he020)
	) name535 (
		\rd1_Key_o_reg[40]/NET0131 ,
		_w250_,
		_w256_,
		_w590_,
		_w784_
	);
	LUT4 #(
		.INIT('h0e02)
	) name536 (
		\rd1_Key_o_reg[41]/NET0131 ,
		_w250_,
		_w256_,
		_w573_,
		_w785_
	);
	LUT3 #(
		.INIT('h54)
	) name537 (
		decrypt_i_pad,
		_w784_,
		_w785_,
		_w786_
	);
	LUT4 #(
		.INIT('he020)
	) name538 (
		\rd1_Key_o_reg[43]/NET0131 ,
		_w250_,
		_w263_,
		_w494_,
		_w787_
	);
	LUT4 #(
		.INIT('haaa8)
	) name539 (
		decrypt_i_pad,
		_w477_,
		_w572_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('he)
	) name540 (
		_w786_,
		_w788_,
		_w789_
	);
	LUT4 #(
		.INIT('h0e02)
	) name541 (
		\rd1_Key_o_reg[27]/NET0131 ,
		_w250_,
		_w256_,
		_w265_,
		_w790_
	);
	LUT3 #(
		.INIT('h54)
	) name542 (
		decrypt_i_pad,
		_w550_,
		_w790_,
		_w791_
	);
	LUT4 #(
		.INIT('h0023)
	) name543 (
		_w267_,
		_w262_,
		_w263_,
		_w650_,
		_w792_
	);
	LUT3 #(
		.INIT('hce)
	) name544 (
		decrypt_i_pad,
		_w791_,
		_w792_,
		_w793_
	);
	LUT4 #(
		.INIT('hf35f)
	) name545 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w794_
	);
	LUT4 #(
		.INIT('h0001)
	) name546 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w795_
	);
	LUT3 #(
		.INIT('h0e)
	) name547 (
		_w581_,
		_w794_,
		_w795_,
		_w796_
	);
	LUT3 #(
		.INIT('hd0)
	) name548 (
		_w584_,
		_w587_,
		_w581_,
		_w797_
	);
	LUT4 #(
		.INIT('h1800)
	) name549 (
		_w584_,
		_w587_,
		_w596_,
		_w581_,
		_w798_
	);
	LUT4 #(
		.INIT('h4000)
	) name550 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w799_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		_w798_,
		_w799_,
		_w800_
	);
	LUT3 #(
		.INIT('h15)
	) name552 (
		_w615_,
		_w796_,
		_w800_,
		_w801_
	);
	LUT4 #(
		.INIT('h2000)
	) name553 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w802_
	);
	LUT4 #(
		.INIT('h5145)
	) name554 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w803_
	);
	LUT4 #(
		.INIT('hd700)
	) name555 (
		_w599_,
		_w587_,
		_w596_,
		_w581_,
		_w804_
	);
	LUT4 #(
		.INIT('h8a88)
	) name556 (
		_w615_,
		_w802_,
		_w803_,
		_w804_,
		_w805_
	);
	LUT4 #(
		.INIT('ha7fb)
	) name557 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w806_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		_w581_,
		_w806_,
		_w807_
	);
	LUT4 #(
		.INIT('h2000)
	) name559 (
		_w599_,
		_w584_,
		_w596_,
		_w581_,
		_w808_
	);
	LUT4 #(
		.INIT('h0080)
	) name560 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w809_
	);
	LUT3 #(
		.INIT('ha8)
	) name561 (
		_w587_,
		_w808_,
		_w809_,
		_w810_
	);
	LUT3 #(
		.INIT('h01)
	) name562 (
		_w587_,
		_w596_,
		_w581_,
		_w811_
	);
	LUT4 #(
		.INIT('hee0e)
	) name563 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w812_
	);
	LUT4 #(
		.INIT('h0e00)
	) name564 (
		_w584_,
		_w596_,
		_w581_,
		_w615_,
		_w813_
	);
	LUT4 #(
		.INIT('h7077)
	) name565 (
		_w624_,
		_w811_,
		_w812_,
		_w813_,
		_w814_
	);
	LUT4 #(
		.INIT('h0100)
	) name566 (
		_w805_,
		_w810_,
		_w807_,
		_w814_,
		_w815_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name567 (
		\data_i[12]_pad ,
		load_i_pad,
		\rd1_L_o_reg[22]/NET0131 ,
		_w250_,
		_w816_
	);
	LUT3 #(
		.INIT('h4b)
	) name568 (
		_w801_,
		_w815_,
		_w816_,
		_w817_
	);
	LUT4 #(
		.INIT('h0415)
	) name569 (
		decrypt_i_pad,
		_w256_,
		_w267_,
		_w392_,
		_w818_
	);
	LUT4 #(
		.INIT('he020)
	) name570 (
		\rd1_Key_o_reg[4]/NET0131 ,
		_w250_,
		_w263_,
		_w273_,
		_w819_
	);
	LUT4 #(
		.INIT('h000d)
	) name571 (
		_w256_,
		_w281_,
		_w649_,
		_w819_,
		_w820_
	);
	LUT3 #(
		.INIT('hce)
	) name572 (
		decrypt_i_pad,
		_w818_,
		_w820_,
		_w821_
	);
	LUT4 #(
		.INIT('h3c36)
	) name573 (
		decrypt_i_pad,
		_w510_,
		_w818_,
		_w820_,
		_w822_
	);
	LUT4 #(
		.INIT('h3c36)
	) name574 (
		decrypt_i_pad,
		_w306_,
		_w315_,
		_w323_,
		_w823_
	);
	LUT4 #(
		.INIT('h3c36)
	) name575 (
		decrypt_i_pad,
		_w716_,
		_w720_,
		_w723_,
		_w824_
	);
	LUT4 #(
		.INIT('h470f)
	) name576 (
		\data_i[9]_pad ,
		load_i_pad,
		\rd1_R_o_reg[6]/NET0131 ,
		_w250_,
		_w825_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name577 (
		\data_i[9]_pad ,
		load_i_pad,
		\rd1_R_o_reg[6]/NET0131 ,
		_w250_,
		_w826_
	);
	LUT4 #(
		.INIT('h31ce)
	) name578 (
		decrypt_i_pad,
		_w438_,
		_w445_,
		_w825_,
		_w827_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w824_,
		_w827_,
		_w828_
	);
	LUT3 #(
		.INIT('h06)
	) name580 (
		_w330_,
		_w460_,
		_w824_,
		_w829_
	);
	LUT4 #(
		.INIT('h470f)
	) name581 (
		\data_i[17]_pad ,
		load_i_pad,
		\rd1_R_o_reg[5]/NET0131 ,
		_w250_,
		_w830_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name582 (
		\data_i[17]_pad ,
		load_i_pad,
		\rd1_R_o_reg[5]/NET0131 ,
		_w250_,
		_w831_
	);
	LUT4 #(
		.INIT('h31ce)
	) name583 (
		decrypt_i_pad,
		_w791_,
		_w792_,
		_w830_,
		_w832_
	);
	LUT4 #(
		.INIT('h0900)
	) name584 (
		_w330_,
		_w460_,
		_w827_,
		_w832_,
		_w833_
	);
	LUT3 #(
		.INIT('h32)
	) name585 (
		_w829_,
		_w828_,
		_w833_,
		_w834_
	);
	LUT3 #(
		.INIT('h90)
	) name586 (
		_w330_,
		_w460_,
		_w824_,
		_w835_
	);
	LUT3 #(
		.INIT('h69)
	) name587 (
		_w330_,
		_w460_,
		_w824_,
		_w836_
	);
	LUT3 #(
		.INIT('h07)
	) name588 (
		_w824_,
		_w827_,
		_w832_,
		_w837_
	);
	LUT2 #(
		.INIT('h8)
	) name589 (
		_w836_,
		_w837_,
		_w838_
	);
	LUT3 #(
		.INIT('h60)
	) name590 (
		_w330_,
		_w460_,
		_w832_,
		_w839_
	);
	LUT4 #(
		.INIT('h0600)
	) name591 (
		_w330_,
		_w460_,
		_w824_,
		_w832_,
		_w840_
	);
	LUT2 #(
		.INIT('h4)
	) name592 (
		_w824_,
		_w827_,
		_w841_
	);
	LUT2 #(
		.INIT('h9)
	) name593 (
		_w824_,
		_w827_,
		_w842_
	);
	LUT4 #(
		.INIT('h090f)
	) name594 (
		_w330_,
		_w460_,
		_w823_,
		_w832_,
		_w843_
	);
	LUT4 #(
		.INIT('h26bf)
	) name595 (
		_w824_,
		_w827_,
		_w839_,
		_w843_,
		_w844_
	);
	LUT4 #(
		.INIT('h5700)
	) name596 (
		_w823_,
		_w834_,
		_w838_,
		_w844_,
		_w845_
	);
	LUT4 #(
		.INIT('h0006)
	) name597 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w846_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		_w823_,
		_w846_,
		_w847_
	);
	LUT4 #(
		.INIT('h0600)
	) name599 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w848_
	);
	LUT4 #(
		.INIT('h9099)
	) name600 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w849_
	);
	LUT3 #(
		.INIT('h02)
	) name601 (
		_w832_,
		_w849_,
		_w848_,
		_w850_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		_w847_,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w822_,
		_w823_,
		_w852_
	);
	LUT4 #(
		.INIT('h0060)
	) name604 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w853_
	);
	LUT3 #(
		.INIT('h09)
	) name605 (
		_w330_,
		_w460_,
		_w832_,
		_w854_
	);
	LUT4 #(
		.INIT('h0090)
	) name606 (
		_w330_,
		_w460_,
		_w824_,
		_w832_,
		_w855_
	);
	LUT4 #(
		.INIT('h000b)
	) name607 (
		_w832_,
		_w848_,
		_w853_,
		_w855_,
		_w856_
	);
	LUT3 #(
		.INIT('h96)
	) name608 (
		_w330_,
		_w460_,
		_w832_,
		_w857_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w823_,
		_w832_,
		_w858_
	);
	LUT4 #(
		.INIT('h80c0)
	) name610 (
		_w823_,
		_w824_,
		_w827_,
		_w832_,
		_w859_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		_w857_,
		_w859_,
		_w860_
	);
	LUT4 #(
		.INIT('h0777)
	) name612 (
		_w853_,
		_w858_,
		_w854_,
		_w828_,
		_w861_
	);
	LUT4 #(
		.INIT('h5100)
	) name613 (
		_w860_,
		_w852_,
		_w856_,
		_w861_,
		_w862_
	);
	LUT4 #(
		.INIT('he400)
	) name614 (
		_w822_,
		_w851_,
		_w845_,
		_w862_,
		_w863_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name615 (
		\data_i[42]_pad ,
		load_i_pad,
		\rd1_L_o_reg[10]/NET0131 ,
		_w250_,
		_w864_
	);
	LUT2 #(
		.INIT('h9)
	) name616 (
		_w863_,
		_w864_,
		_w865_
	);
	LUT4 #(
		.INIT('h9000)
	) name617 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w866_
	);
	LUT4 #(
		.INIT('h5400)
	) name618 (
		_w823_,
		_w824_,
		_w827_,
		_w832_,
		_w867_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		_w866_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h2)
	) name620 (
		_w823_,
		_w832_,
		_w869_
	);
	LUT4 #(
		.INIT('h5d04)
	) name621 (
		_w823_,
		_w824_,
		_w827_,
		_w832_,
		_w870_
	);
	LUT3 #(
		.INIT('hb0)
	) name622 (
		_w866_,
		_w867_,
		_w870_,
		_w871_
	);
	LUT4 #(
		.INIT('h6900)
	) name623 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w872_
	);
	LUT3 #(
		.INIT('h09)
	) name624 (
		_w330_,
		_w460_,
		_w824_,
		_w873_
	);
	LUT4 #(
		.INIT('h4d4f)
	) name625 (
		_w823_,
		_w832_,
		_w872_,
		_w873_,
		_w874_
	);
	LUT3 #(
		.INIT('h8a)
	) name626 (
		_w822_,
		_w871_,
		_w874_,
		_w875_
	);
	LUT4 #(
		.INIT('h008a)
	) name627 (
		_w823_,
		_w824_,
		_w833_,
		_w866_,
		_w876_
	);
	LUT4 #(
		.INIT('h0111)
	) name628 (
		_w823_,
		_w848_,
		_w854_,
		_w828_,
		_w877_
	);
	LUT4 #(
		.INIT('h131f)
	) name629 (
		_w823_,
		_w827_,
		_w855_,
		_w840_,
		_w878_
	);
	LUT4 #(
		.INIT('h0e00)
	) name630 (
		_w876_,
		_w877_,
		_w868_,
		_w878_,
		_w879_
	);
	LUT3 #(
		.INIT('h40)
	) name631 (
		_w823_,
		_w827_,
		_w840_,
		_w880_
	);
	LUT4 #(
		.INIT('h96f9)
	) name632 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w881_
	);
	LUT2 #(
		.INIT('h2)
	) name633 (
		_w869_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		_w880_,
		_w882_,
		_w883_
	);
	LUT4 #(
		.INIT('h0e00)
	) name635 (
		_w822_,
		_w879_,
		_w875_,
		_w883_,
		_w884_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name636 (
		\data_i[54]_pad ,
		load_i_pad,
		\rd1_L_o_reg[25]/NET0131 ,
		_w250_,
		_w885_
	);
	LUT2 #(
		.INIT('h9)
	) name637 (
		_w884_,
		_w885_,
		_w886_
	);
	LUT3 #(
		.INIT('h1e)
	) name638 (
		_w638_,
		_w640_,
		_w743_,
		_w887_
	);
	LUT4 #(
		.INIT('h32cd)
	) name639 (
		decrypt_i_pad,
		_w464_,
		_w470_,
		_w653_,
		_w888_
	);
	LUT2 #(
		.INIT('h9)
	) name640 (
		_w491_,
		_w501_,
		_w889_
	);
	LUT4 #(
		.INIT('hb800)
	) name641 (
		\key_i[13]_pad ,
		load_i_pad,
		\rd1_Key_o_reg[38]/NET0131 ,
		_w250_,
		_w890_
	);
	LUT4 #(
		.INIT('h000d)
	) name642 (
		_w263_,
		_w422_,
		_w761_,
		_w890_,
		_w891_
	);
	LUT4 #(
		.INIT('he020)
	) name643 (
		\rd1_Key_o_reg[40]/NET0131 ,
		_w250_,
		_w263_,
		_w590_,
		_w892_
	);
	LUT4 #(
		.INIT('haaa8)
	) name644 (
		decrypt_i_pad,
		_w486_,
		_w575_,
		_w892_,
		_w893_
	);
	LUT3 #(
		.INIT('hf1)
	) name645 (
		decrypt_i_pad,
		_w891_,
		_w893_,
		_w894_
	);
	LUT4 #(
		.INIT('h33c9)
	) name646 (
		decrypt_i_pad,
		_w553_,
		_w891_,
		_w893_,
		_w895_
	);
	LUT3 #(
		.INIT('h56)
	) name647 (
		_w447_,
		_w786_,
		_w788_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name648 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT4 #(
		.INIT('h6000)
	) name649 (
		_w491_,
		_w501_,
		_w895_,
		_w896_,
		_w898_
	);
	LUT4 #(
		.INIT('h96ff)
	) name650 (
		_w491_,
		_w501_,
		_w895_,
		_w896_,
		_w899_
	);
	LUT4 #(
		.INIT('h31ce)
	) name651 (
		decrypt_i_pad,
		_w355_,
		_w361_,
		_w363_,
		_w900_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		_w895_,
		_w896_,
		_w901_
	);
	LUT3 #(
		.INIT('h08)
	) name653 (
		_w900_,
		_w895_,
		_w896_,
		_w902_
	);
	LUT3 #(
		.INIT('h20)
	) name654 (
		_w900_,
		_w895_,
		_w896_,
		_w903_
	);
	LUT3 #(
		.INIT('h86)
	) name655 (
		_w900_,
		_w895_,
		_w896_,
		_w904_
	);
	LUT3 #(
		.INIT('ha2)
	) name656 (
		_w888_,
		_w899_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w895_,
		_w896_,
		_w906_
	);
	LUT3 #(
		.INIT('h60)
	) name658 (
		_w491_,
		_w501_,
		_w900_,
		_w907_
	);
	LUT2 #(
		.INIT('h8)
	) name659 (
		_w906_,
		_w907_,
		_w908_
	);
	LUT3 #(
		.INIT('ha8)
	) name660 (
		_w887_,
		_w905_,
		_w908_,
		_w909_
	);
	LUT4 #(
		.INIT('h0006)
	) name661 (
		_w491_,
		_w501_,
		_w900_,
		_w895_,
		_w910_
	);
	LUT3 #(
		.INIT('h40)
	) name662 (
		_w900_,
		_w895_,
		_w896_,
		_w911_
	);
	LUT3 #(
		.INIT('hb7)
	) name663 (
		_w900_,
		_w895_,
		_w896_,
		_w912_
	);
	LUT4 #(
		.INIT('hce00)
	) name664 (
		_w889_,
		_w910_,
		_w912_,
		_w888_,
		_w913_
	);
	LUT3 #(
		.INIT('h09)
	) name665 (
		_w491_,
		_w501_,
		_w895_,
		_w914_
	);
	LUT4 #(
		.INIT('h0009)
	) name666 (
		_w491_,
		_w501_,
		_w895_,
		_w896_,
		_w915_
	);
	LUT2 #(
		.INIT('h4)
	) name667 (
		_w900_,
		_w915_,
		_w916_
	);
	LUT3 #(
		.INIT('h04)
	) name668 (
		_w900_,
		_w895_,
		_w896_,
		_w917_
	);
	LUT3 #(
		.INIT('h80)
	) name669 (
		_w900_,
		_w895_,
		_w896_,
		_w918_
	);
	LUT4 #(
		.INIT('h3332)
	) name670 (
		_w914_,
		_w888_,
		_w918_,
		_w917_,
		_w919_
	);
	LUT4 #(
		.INIT('h00fe)
	) name671 (
		_w916_,
		_w913_,
		_w919_,
		_w887_,
		_w920_
	);
	LUT3 #(
		.INIT('h80)
	) name672 (
		_w888_,
		_w906_,
		_w907_,
		_w921_
	);
	LUT4 #(
		.INIT('h0666)
	) name673 (
		_w491_,
		_w501_,
		_w895_,
		_w896_,
		_w922_
	);
	LUT2 #(
		.INIT('h2)
	) name674 (
		_w900_,
		_w895_,
		_w923_
	);
	LUT3 #(
		.INIT('h0d)
	) name675 (
		_w900_,
		_w895_,
		_w888_,
		_w924_
	);
	LUT3 #(
		.INIT('he0)
	) name676 (
		_w895_,
		_w896_,
		_w887_,
		_w925_
	);
	LUT3 #(
		.INIT('h80)
	) name677 (
		_w924_,
		_w922_,
		_w925_,
		_w926_
	);
	LUT3 #(
		.INIT('h04)
	) name678 (
		_w900_,
		_w915_,
		_w888_,
		_w927_
	);
	LUT4 #(
		.INIT('hfb51)
	) name679 (
		_w900_,
		_w915_,
		_w888_,
		_w899_,
		_w928_
	);
	LUT3 #(
		.INIT('h10)
	) name680 (
		_w921_,
		_w926_,
		_w928_,
		_w929_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name681 (
		\data_i[50]_pad ,
		load_i_pad,
		\rd1_L_o_reg[9]/NET0131 ,
		_w250_,
		_w930_
	);
	LUT4 #(
		.INIT('h10ef)
	) name682 (
		_w920_,
		_w909_,
		_w929_,
		_w930_,
		_w931_
	);
	LUT3 #(
		.INIT('h56)
	) name683 (
		_w696_,
		_w726_,
		_w728_,
		_w932_
	);
	LUT4 #(
		.INIT('h470f)
	) name684 (
		\data_i[51]_pad ,
		load_i_pad,
		\rd1_R_o_reg[9]/NET0131 ,
		_w250_,
		_w933_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name685 (
		\data_i[51]_pad ,
		load_i_pad,
		\rd1_R_o_reg[9]/NET0131 ,
		_w250_,
		_w934_
	);
	LUT2 #(
		.INIT('h9)
	) name686 (
		_w342_,
		_w933_,
		_w935_
	);
	LUT3 #(
		.INIT('h1e)
	) name687 (
		_w631_,
		_w634_,
		_w685_,
		_w936_
	);
	LUT3 #(
		.INIT('h56)
	) name688 (
		_w270_,
		_w276_,
		_w286_,
		_w937_
	);
	LUT4 #(
		.INIT('h4080)
	) name689 (
		_w342_,
		_w936_,
		_w937_,
		_w933_,
		_w938_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		_w932_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		_w936_,
		_w932_,
		_w940_
	);
	LUT2 #(
		.INIT('h9)
	) name692 (
		_w936_,
		_w932_,
		_w941_
	);
	LUT3 #(
		.INIT('h90)
	) name693 (
		_w936_,
		_w932_,
		_w937_,
		_w942_
	);
	LUT4 #(
		.INIT('ha251)
	) name694 (
		_w342_,
		_w932_,
		_w937_,
		_w933_,
		_w943_
	);
	LUT3 #(
		.INIT('h1e)
	) name695 (
		_w382_,
		_w385_,
		_w716_,
		_w944_
	);
	LUT3 #(
		.INIT('h0b)
	) name696 (
		_w942_,
		_w943_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		_w936_,
		_w937_,
		_w946_
	);
	LUT4 #(
		.INIT('h1428)
	) name698 (
		_w342_,
		_w936_,
		_w937_,
		_w933_,
		_w947_
	);
	LUT3 #(
		.INIT('h48)
	) name699 (
		_w342_,
		_w932_,
		_w933_,
		_w948_
	);
	LUT4 #(
		.INIT('h00c4)
	) name700 (
		_w942_,
		_w944_,
		_w948_,
		_w947_,
		_w949_
	);
	LUT3 #(
		.INIT('h02)
	) name701 (
		_w936_,
		_w932_,
		_w937_,
		_w950_
	);
	LUT4 #(
		.INIT('h00f4)
	) name702 (
		_w939_,
		_w945_,
		_w949_,
		_w950_,
		_w951_
	);
	LUT4 #(
		.INIT('h3c36)
	) name703 (
		decrypt_i_pad,
		_w460_,
		_w731_,
		_w732_,
		_w952_
	);
	LUT3 #(
		.INIT('h01)
	) name704 (
		_w936_,
		_w932_,
		_w937_,
		_w953_
	);
	LUT4 #(
		.INIT('h2010)
	) name705 (
		_w342_,
		_w936_,
		_w932_,
		_w933_,
		_w954_
	);
	LUT3 #(
		.INIT('h20)
	) name706 (
		_w936_,
		_w932_,
		_w937_,
		_w955_
	);
	LUT4 #(
		.INIT('h0001)
	) name707 (
		_w938_,
		_w954_,
		_w955_,
		_w953_,
		_w956_
	);
	LUT4 #(
		.INIT('h0804)
	) name708 (
		_w342_,
		_w932_,
		_w937_,
		_w933_,
		_w957_
	);
	LUT4 #(
		.INIT('h8040)
	) name709 (
		_w342_,
		_w936_,
		_w932_,
		_w933_,
		_w958_
	);
	LUT3 #(
		.INIT('h10)
	) name710 (
		_w936_,
		_w932_,
		_w937_,
		_w959_
	);
	LUT3 #(
		.INIT('he3)
	) name711 (
		_w936_,
		_w932_,
		_w937_,
		_w960_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name712 (
		_w944_,
		_w957_,
		_w958_,
		_w960_,
		_w961_
	);
	LUT3 #(
		.INIT('h0d)
	) name713 (
		_w944_,
		_w956_,
		_w961_,
		_w962_
	);
	LUT3 #(
		.INIT('h12)
	) name714 (
		_w342_,
		_w937_,
		_w933_,
		_w963_
	);
	LUT3 #(
		.INIT('h10)
	) name715 (
		_w941_,
		_w944_,
		_w963_,
		_w964_
	);
	LUT4 #(
		.INIT('hdeed)
	) name716 (
		_w342_,
		_w936_,
		_w932_,
		_w933_,
		_w965_
	);
	LUT3 #(
		.INIT('h04)
	) name717 (
		_w937_,
		_w944_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w964_,
		_w966_,
		_w967_
	);
	LUT4 #(
		.INIT('he200)
	) name719 (
		_w951_,
		_w952_,
		_w962_,
		_w967_,
		_w968_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name720 (
		\data_i[32]_pad ,
		load_i_pad,
		\rd1_L_o_reg[3]/NET0131 ,
		_w250_,
		_w969_
	);
	LUT2 #(
		.INIT('h6)
	) name721 (
		_w968_,
		_w969_,
		_w970_
	);
	LUT4 #(
		.INIT('h9909)
	) name722 (
		_w491_,
		_w501_,
		_w895_,
		_w896_,
		_w971_
	);
	LUT4 #(
		.INIT('h9009)
	) name723 (
		_w491_,
		_w501_,
		_w895_,
		_w896_,
		_w972_
	);
	LUT2 #(
		.INIT('h4)
	) name724 (
		_w900_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h8)
	) name725 (
		_w889_,
		_w902_,
		_w974_
	);
	LUT4 #(
		.INIT('h6000)
	) name726 (
		_w491_,
		_w501_,
		_w900_,
		_w896_,
		_w975_
	);
	LUT4 #(
		.INIT('h0600)
	) name727 (
		_w491_,
		_w501_,
		_w895_,
		_w896_,
		_w976_
	);
	LUT3 #(
		.INIT('h01)
	) name728 (
		_w888_,
		_w976_,
		_w975_,
		_w977_
	);
	LUT4 #(
		.INIT('h0060)
	) name729 (
		_w491_,
		_w501_,
		_w900_,
		_w896_,
		_w978_
	);
	LUT4 #(
		.INIT('hdc00)
	) name730 (
		_w900_,
		_w895_,
		_w896_,
		_w888_,
		_w979_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		_w978_,
		_w979_,
		_w980_
	);
	LUT4 #(
		.INIT('h5510)
	) name732 (
		_w973_,
		_w974_,
		_w977_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h2)
	) name733 (
		_w887_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h8)
	) name734 (
		_w889_,
		_w918_,
		_w983_
	);
	LUT3 #(
		.INIT('h10)
	) name735 (
		_w900_,
		_w895_,
		_w896_,
		_w984_
	);
	LUT4 #(
		.INIT('h0060)
	) name736 (
		_w491_,
		_w501_,
		_w895_,
		_w896_,
		_w985_
	);
	LUT4 #(
		.INIT('h0006)
	) name737 (
		_w491_,
		_w501_,
		_w900_,
		_w896_,
		_w986_
	);
	LUT4 #(
		.INIT('h001b)
	) name738 (
		_w889_,
		_w901_,
		_w984_,
		_w986_,
		_w987_
	);
	LUT3 #(
		.INIT('h45)
	) name739 (
		_w888_,
		_w983_,
		_w987_,
		_w988_
	);
	LUT4 #(
		.INIT('h0090)
	) name740 (
		_w491_,
		_w501_,
		_w900_,
		_w896_,
		_w989_
	);
	LUT3 #(
		.INIT('ha8)
	) name741 (
		_w888_,
		_w976_,
		_w989_,
		_w990_
	);
	LUT3 #(
		.INIT('h09)
	) name742 (
		_w491_,
		_w501_,
		_w896_,
		_w991_
	);
	LUT4 #(
		.INIT('h0600)
	) name743 (
		_w491_,
		_w501_,
		_w900_,
		_w895_,
		_w992_
	);
	LUT3 #(
		.INIT('h07)
	) name744 (
		_w923_,
		_w991_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h4)
	) name745 (
		_w990_,
		_w993_,
		_w994_
	);
	LUT3 #(
		.INIT('he0)
	) name746 (
		_w915_,
		_w911_,
		_w888_,
		_w995_
	);
	LUT4 #(
		.INIT('h45ef)
	) name747 (
		_w900_,
		_w888_,
		_w985_,
		_w976_,
		_w996_
	);
	LUT2 #(
		.INIT('h4)
	) name748 (
		_w995_,
		_w996_,
		_w997_
	);
	LUT4 #(
		.INIT('hba00)
	) name749 (
		_w887_,
		_w988_,
		_w994_,
		_w997_,
		_w998_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name750 (
		\data_i[48]_pad ,
		load_i_pad,
		\rd1_L_o_reg[1]/NET0131 ,
		_w250_,
		_w999_
	);
	LUT3 #(
		.INIT('h4b)
	) name751 (
		_w982_,
		_w998_,
		_w999_,
		_w1000_
	);
	LUT3 #(
		.INIT('h04)
	) name752 (
		_w665_,
		_w666_,
		_w668_,
		_w1001_
	);
	LUT4 #(
		.INIT('h5551)
	) name753 (
		_w687_,
		_w665_,
		_w666_,
		_w668_,
		_w1002_
	);
	LUT4 #(
		.INIT('hc0af)
	) name754 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1003_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name755 (
		_w692_,
		_w1001_,
		_w1002_,
		_w1003_,
		_w1004_
	);
	LUT4 #(
		.INIT('h1000)
	) name756 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1005_
	);
	LUT3 #(
		.INIT('ha8)
	) name757 (
		_w698_,
		_w1004_,
		_w1005_,
		_w1006_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name758 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1007_
	);
	LUT4 #(
		.INIT('h0020)
	) name759 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1008_
	);
	LUT4 #(
		.INIT('h0200)
	) name760 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1009_
	);
	LUT4 #(
		.INIT('hfddf)
	) name761 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1010_
	);
	LUT4 #(
		.INIT('h02aa)
	) name762 (
		_w687_,
		_w698_,
		_w1007_,
		_w1010_,
		_w1011_
	);
	LUT3 #(
		.INIT('h01)
	) name763 (
		_w687_,
		_w665_,
		_w668_,
		_w1012_
	);
	LUT3 #(
		.INIT('h01)
	) name764 (
		_w693_,
		_w1012_,
		_w1008_,
		_w1013_
	);
	LUT4 #(
		.INIT('h4000)
	) name765 (
		_w687_,
		_w665_,
		_w666_,
		_w668_,
		_w1014_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		_w701_,
		_w1014_,
		_w1015_
	);
	LUT4 #(
		.INIT('h0100)
	) name767 (
		_w687_,
		_w665_,
		_w666_,
		_w676_,
		_w1016_
	);
	LUT4 #(
		.INIT('h00ea)
	) name768 (
		_w698_,
		_w1013_,
		_w1015_,
		_w1016_,
		_w1017_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name769 (
		\data_i[22]_pad ,
		load_i_pad,
		\rd1_L_o_reg[29]/NET0131 ,
		_w250_,
		_w1018_
	);
	LUT4 #(
		.INIT('h10ef)
	) name770 (
		_w1006_,
		_w1011_,
		_w1017_,
		_w1018_,
		_w1019_
	);
	LUT3 #(
		.INIT('ha2)
	) name771 (
		_w823_,
		_w824_,
		_w827_,
		_w1020_
	);
	LUT2 #(
		.INIT('h2)
	) name772 (
		_w854_,
		_w1020_,
		_w1021_
	);
	LUT3 #(
		.INIT('h2a)
	) name773 (
		_w822_,
		_w827_,
		_w840_,
		_w1022_
	);
	LUT3 #(
		.INIT('h06)
	) name774 (
		_w330_,
		_w460_,
		_w832_,
		_w1023_
	);
	LUT3 #(
		.INIT('h15)
	) name775 (
		_w833_,
		_w842_,
		_w1023_,
		_w1024_
	);
	LUT3 #(
		.INIT('h40)
	) name776 (
		_w1021_,
		_w1022_,
		_w1024_,
		_w1025_
	);
	LUT4 #(
		.INIT('hf690)
	) name777 (
		_w330_,
		_w460_,
		_w824_,
		_w832_,
		_w1026_
	);
	LUT3 #(
		.INIT('h15)
	) name778 (
		_w822_,
		_w1020_,
		_w1026_,
		_w1027_
	);
	LUT3 #(
		.INIT('h8a)
	) name779 (
		_w823_,
		_w838_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h4)
	) name780 (
		_w1025_,
		_w1028_,
		_w1029_
	);
	LUT4 #(
		.INIT('hf060)
	) name781 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w1030_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w1023_,
		_w1030_,
		_w1031_
	);
	LUT3 #(
		.INIT('h04)
	) name783 (
		_w1021_,
		_w1022_,
		_w1031_,
		_w1032_
	);
	LUT4 #(
		.INIT('h9009)
	) name784 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w1033_
	);
	LUT3 #(
		.INIT('h01)
	) name785 (
		_w853_,
		_w839_,
		_w1033_,
		_w1034_
	);
	LUT3 #(
		.INIT('h51)
	) name786 (
		_w823_,
		_w1027_,
		_w1034_,
		_w1035_
	);
	LUT4 #(
		.INIT('hff60)
	) name787 (
		_w330_,
		_w460_,
		_w823_,
		_w832_,
		_w1036_
	);
	LUT4 #(
		.INIT('h3f15)
	) name788 (
		_w841_,
		_w853_,
		_w858_,
		_w1036_,
		_w1037_
	);
	LUT3 #(
		.INIT('hb0)
	) name789 (
		_w1032_,
		_w1035_,
		_w1037_,
		_w1038_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name790 (
		\data_i[56]_pad ,
		load_i_pad,
		\rd1_L_o_reg[0]/NET0131 ,
		_w250_,
		_w1039_
	);
	LUT3 #(
		.INIT('h4b)
	) name791 (
		_w1029_,
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT4 #(
		.INIT('h0010)
	) name792 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1041_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name793 (
		_w687_,
		_w665_,
		_w666_,
		_w676_,
		_w1042_
	);
	LUT3 #(
		.INIT('h80)
	) name794 (
		_w665_,
		_w666_,
		_w676_,
		_w1043_
	);
	LUT4 #(
		.INIT('h1555)
	) name795 (
		_w687_,
		_w665_,
		_w666_,
		_w676_,
		_w1044_
	);
	LUT4 #(
		.INIT('h8acf)
	) name796 (
		_w1008_,
		_w1041_,
		_w1042_,
		_w1044_,
		_w1045_
	);
	LUT4 #(
		.INIT('hc200)
	) name797 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1046_
	);
	LUT3 #(
		.INIT('h01)
	) name798 (
		_w698_,
		_w1016_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h4)
	) name799 (
		_w1045_,
		_w1047_,
		_w1048_
	);
	LUT2 #(
		.INIT('h2)
	) name800 (
		_w698_,
		_w703_,
		_w1049_
	);
	LUT4 #(
		.INIT('h0200)
	) name801 (
		_w687_,
		_w665_,
		_w666_,
		_w676_,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		_w1014_,
		_w1050_,
		_w1051_
	);
	LUT3 #(
		.INIT('h74)
	) name803 (
		_w687_,
		_w668_,
		_w676_,
		_w1052_
	);
	LUT4 #(
		.INIT('hcf45)
	) name804 (
		_w667_,
		_w690_,
		_w1012_,
		_w1052_,
		_w1053_
	);
	LUT3 #(
		.INIT('h80)
	) name805 (
		_w1049_,
		_w1051_,
		_w1053_,
		_w1054_
	);
	LUT4 #(
		.INIT('haaa2)
	) name806 (
		_w687_,
		_w665_,
		_w668_,
		_w676_,
		_w1055_
	);
	LUT4 #(
		.INIT('h5545)
	) name807 (
		_w687_,
		_w665_,
		_w666_,
		_w676_,
		_w1056_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name808 (
		_w1005_,
		_w1009_,
		_w1055_,
		_w1056_,
		_w1057_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name809 (
		\data_i[62]_pad ,
		load_i_pad,
		\rd1_L_o_reg[24]/NET0131 ,
		_w250_,
		_w1058_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name810 (
		_w1048_,
		_w1054_,
		_w1057_,
		_w1058_,
		_w1059_
	);
	LUT4 #(
		.INIT('h0e02)
	) name811 (
		\rd1_Key_o_reg[51]/NET0131 ,
		_w250_,
		_w256_,
		_w428_,
		_w1060_
	);
	LUT3 #(
		.INIT('h54)
	) name812 (
		decrypt_i_pad,
		_w404_,
		_w1060_,
		_w1061_
	);
	LUT4 #(
		.INIT('he020)
	) name813 (
		\rd1_Key_o_reg[53]/NET0131 ,
		_w250_,
		_w263_,
		_w467_,
		_w1062_
	);
	LUT4 #(
		.INIT('h000d)
	) name814 (
		_w256_,
		_w465_,
		_w607_,
		_w1062_,
		_w1063_
	);
	LUT3 #(
		.INIT('hce)
	) name815 (
		decrypt_i_pad,
		_w1061_,
		_w1063_,
		_w1064_
	);
	LUT4 #(
		.INIT('h470f)
	) name816 (
		\data_i[21]_pad ,
		load_i_pad,
		\rd1_R_o_reg[21]/NET0131 ,
		_w250_,
		_w1065_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name817 (
		\data_i[21]_pad ,
		load_i_pad,
		\rd1_R_o_reg[21]/NET0131 ,
		_w250_,
		_w1066_
	);
	LUT4 #(
		.INIT('h31ce)
	) name818 (
		decrypt_i_pad,
		_w1061_,
		_w1063_,
		_w1065_,
		_w1067_
	);
	LUT3 #(
		.INIT('h1e)
	) name819 (
		_w346_,
		_w351_,
		_w594_,
		_w1068_
	);
	LUT2 #(
		.INIT('h4)
	) name820 (
		_w1067_,
		_w1068_,
		_w1069_
	);
	LUT3 #(
		.INIT('h1e)
	) name821 (
		_w372_,
		_w378_,
		_w764_,
		_w1070_
	);
	LUT4 #(
		.INIT('h0145)
	) name822 (
		decrypt_i_pad,
		_w256_,
		_w496_,
		_w571_,
		_w1071_
	);
	LUT4 #(
		.INIT('he020)
	) name823 (
		\rd1_Key_o_reg[45]/NET0131 ,
		_w250_,
		_w263_,
		_w472_,
		_w1072_
	);
	LUT4 #(
		.INIT('h000d)
	) name824 (
		_w256_,
		_w409_,
		_w476_,
		_w1072_,
		_w1073_
	);
	LUT3 #(
		.INIT('hce)
	) name825 (
		decrypt_i_pad,
		_w1071_,
		_w1073_,
		_w1074_
	);
	LUT4 #(
		.INIT('h470f)
	) name826 (
		\data_i[13]_pad ,
		load_i_pad,
		\rd1_R_o_reg[22]/NET0131 ,
		_w250_,
		_w1075_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name827 (
		\data_i[13]_pad ,
		load_i_pad,
		\rd1_R_o_reg[22]/NET0131 ,
		_w250_,
		_w1076_
	);
	LUT4 #(
		.INIT('h31ce)
	) name828 (
		decrypt_i_pad,
		_w1071_,
		_w1073_,
		_w1075_,
		_w1077_
	);
	LUT4 #(
		.INIT('h31ce)
	) name829 (
		decrypt_i_pad,
		_w484_,
		_w489_,
		_w734_,
		_w1078_
	);
	LUT3 #(
		.INIT('h56)
	) name830 (
		_w1070_,
		_w1077_,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('h2)
	) name831 (
		_w1069_,
		_w1079_,
		_w1080_
	);
	LUT4 #(
		.INIT('ha521)
	) name832 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1081_
	);
	LUT4 #(
		.INIT('h0313)
	) name833 (
		_w1067_,
		_w1068_,
		_w1070_,
		_w1077_,
		_w1082_
	);
	LUT2 #(
		.INIT('h4)
	) name834 (
		_w1081_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h2)
	) name835 (
		_w1067_,
		_w1070_,
		_w1084_
	);
	LUT4 #(
		.INIT('h0800)
	) name836 (
		_w1067_,
		_w1068_,
		_w1070_,
		_w1077_,
		_w1085_
	);
	LUT2 #(
		.INIT('h9)
	) name837 (
		_w411_,
		_w585_,
		_w1086_
	);
	LUT4 #(
		.INIT('h0200)
	) name838 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1087_
	);
	LUT3 #(
		.INIT('h02)
	) name839 (
		_w1086_,
		_w1087_,
		_w1085_,
		_w1088_
	);
	LUT2 #(
		.INIT('h6)
	) name840 (
		_w1070_,
		_w1077_,
		_w1089_
	);
	LUT2 #(
		.INIT('h8)
	) name841 (
		_w1070_,
		_w1078_,
		_w1090_
	);
	LUT4 #(
		.INIT('h9b1e)
	) name842 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1091_
	);
	LUT4 #(
		.INIT('h0008)
	) name843 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1092_
	);
	LUT4 #(
		.INIT('h0302)
	) name844 (
		_w1068_,
		_w1086_,
		_w1092_,
		_w1091_,
		_w1093_
	);
	LUT4 #(
		.INIT('h00ef)
	) name845 (
		_w1080_,
		_w1083_,
		_w1088_,
		_w1093_,
		_w1094_
	);
	LUT4 #(
		.INIT('heee1)
	) name846 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1095_
	);
	LUT3 #(
		.INIT('h0d)
	) name847 (
		_w1086_,
		_w1092_,
		_w1095_,
		_w1096_
	);
	LUT4 #(
		.INIT('h8000)
	) name848 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1097_
	);
	LUT2 #(
		.INIT('h2)
	) name849 (
		_w1068_,
		_w1097_,
		_w1098_
	);
	LUT4 #(
		.INIT('h4080)
	) name850 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1099_
	);
	LUT3 #(
		.INIT('h01)
	) name851 (
		_w1068_,
		_w1087_,
		_w1099_,
		_w1100_
	);
	LUT3 #(
		.INIT('h0b)
	) name852 (
		_w1096_,
		_w1098_,
		_w1100_,
		_w1101_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name853 (
		\data_i[58]_pad ,
		load_i_pad,
		\rd1_L_o_reg[8]/NET0131 ,
		_w250_,
		_w1102_
	);
	LUT3 #(
		.INIT('h1e)
	) name854 (
		_w1094_,
		_w1101_,
		_w1102_,
		_w1103_
	);
	LUT4 #(
		.INIT('h9a30)
	) name855 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1104_
	);
	LUT4 #(
		.INIT('h0004)
	) name856 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1105_
	);
	LUT3 #(
		.INIT('h01)
	) name857 (
		_w766_,
		_w1105_,
		_w1104_,
		_w1106_
	);
	LUT4 #(
		.INIT('hbf00)
	) name858 (
		_w738_,
		_w745_,
		_w737_,
		_w766_,
		_w1107_
	);
	LUT3 #(
		.INIT('h20)
	) name859 (
		_w754_,
		_w755_,
		_w1107_,
		_w1108_
	);
	LUT3 #(
		.INIT('ha8)
	) name860 (
		_w736_,
		_w1106_,
		_w1108_,
		_w1109_
	);
	LUT4 #(
		.INIT('h0150)
	) name861 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1110_
	);
	LUT4 #(
		.INIT('h00fd)
	) name862 (
		_w753_,
		_w745_,
		_w737_,
		_w766_,
		_w1111_
	);
	LUT3 #(
		.INIT('h04)
	) name863 (
		_w777_,
		_w1111_,
		_w1110_,
		_w1112_
	);
	LUT3 #(
		.INIT('h06)
	) name864 (
		_w753_,
		_w738_,
		_w745_,
		_w1113_
	);
	LUT4 #(
		.INIT('hfb00)
	) name865 (
		_w738_,
		_w745_,
		_w737_,
		_w766_,
		_w1114_
	);
	LUT2 #(
		.INIT('h4)
	) name866 (
		_w1113_,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h2)
	) name867 (
		_w753_,
		_w766_,
		_w1116_
	);
	LUT3 #(
		.INIT('h51)
	) name868 (
		_w736_,
		_w757_,
		_w1116_,
		_w1117_
	);
	LUT3 #(
		.INIT('he0)
	) name869 (
		_w1112_,
		_w1115_,
		_w1117_,
		_w1118_
	);
	LUT3 #(
		.INIT('h21)
	) name870 (
		_w738_,
		_w745_,
		_w737_,
		_w1119_
	);
	LUT4 #(
		.INIT('h0777)
	) name871 (
		_w738_,
		_w779_,
		_w1116_,
		_w1119_,
		_w1120_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name872 (
		\data_i[36]_pad ,
		load_i_pad,
		\rd1_L_o_reg[19]/NET0131 ,
		_w250_,
		_w1121_
	);
	LUT4 #(
		.INIT('h1fe0)
	) name873 (
		_w1109_,
		_w1118_,
		_w1120_,
		_w1121_,
		_w1122_
	);
	LUT4 #(
		.INIT('h0804)
	) name874 (
		_w342_,
		_w936_,
		_w937_,
		_w933_,
		_w1123_
	);
	LUT4 #(
		.INIT('h080c)
	) name875 (
		_w932_,
		_w944_,
		_w938_,
		_w1123_,
		_w1124_
	);
	LUT4 #(
		.INIT('h0408)
	) name876 (
		_w342_,
		_w936_,
		_w937_,
		_w933_,
		_w1125_
	);
	LUT3 #(
		.INIT('h08)
	) name877 (
		_w936_,
		_w932_,
		_w937_,
		_w1126_
	);
	LUT4 #(
		.INIT('h00f7)
	) name878 (
		_w936_,
		_w932_,
		_w937_,
		_w944_,
		_w1127_
	);
	LUT2 #(
		.INIT('h4)
	) name879 (
		_w1125_,
		_w1127_,
		_w1128_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name880 (
		_w937_,
		_w935_,
		_w965_,
		_w1126_,
		_w1129_
	);
	LUT4 #(
		.INIT('h0155)
	) name881 (
		_w952_,
		_w1124_,
		_w1128_,
		_w1129_,
		_w1130_
	);
	LUT3 #(
		.INIT('hda)
	) name882 (
		_w936_,
		_w932_,
		_w937_,
		_w1131_
	);
	LUT3 #(
		.INIT('h40)
	) name883 (
		_w936_,
		_w932_,
		_w937_,
		_w1132_
	);
	LUT4 #(
		.INIT('hdab7)
	) name884 (
		_w936_,
		_w932_,
		_w937_,
		_w935_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		_w944_,
		_w1133_,
		_w1134_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name886 (
		_w941_,
		_w944_,
		_w958_,
		_w963_,
		_w1135_
	);
	LUT4 #(
		.INIT('h0201)
	) name887 (
		_w342_,
		_w936_,
		_w932_,
		_w933_,
		_w1136_
	);
	LUT3 #(
		.INIT('h54)
	) name888 (
		_w944_,
		_w955_,
		_w1136_,
		_w1137_
	);
	LUT4 #(
		.INIT('h8040)
	) name889 (
		_w342_,
		_w936_,
		_w937_,
		_w933_,
		_w1138_
	);
	LUT3 #(
		.INIT('h07)
	) name890 (
		_w935_,
		_w953_,
		_w1138_,
		_w1139_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name891 (
		_w952_,
		_w1135_,
		_w1137_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h8)
	) name892 (
		_w937_,
		_w944_,
		_w1141_
	);
	LUT2 #(
		.INIT('h4)
	) name893 (
		_w965_,
		_w1141_,
		_w1142_
	);
	LUT4 #(
		.INIT('h0001)
	) name894 (
		_w1140_,
		_w1134_,
		_w1142_,
		_w1130_,
		_w1143_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name895 (
		\data_i[20]_pad ,
		load_i_pad,
		\rd1_L_o_reg[21]/NET0131 ,
		_w250_,
		_w1144_
	);
	LUT2 #(
		.INIT('h6)
	) name896 (
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT3 #(
		.INIT('hbe)
	) name897 (
		_w599_,
		_w587_,
		_w596_,
		_w1146_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name898 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1147_
	);
	LUT3 #(
		.INIT('h10)
	) name899 (
		_w581_,
		_w1147_,
		_w1146_,
		_w1148_
	);
	LUT4 #(
		.INIT('h0040)
	) name900 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1149_
	);
	LUT4 #(
		.INIT('h0015)
	) name901 (
		_w615_,
		_w624_,
		_w811_,
		_w1149_,
		_w1150_
	);
	LUT3 #(
		.INIT('hc4)
	) name902 (
		_w581_,
		_w615_,
		_w621_,
		_w1151_
	);
	LUT4 #(
		.INIT('h0820)
	) name903 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1152_
	);
	LUT4 #(
		.INIT('h0042)
	) name904 (
		_w584_,
		_w587_,
		_w596_,
		_w581_,
		_w1153_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		_w1152_,
		_w1153_,
		_w1154_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name906 (
		_w1148_,
		_w1150_,
		_w1151_,
		_w1154_,
		_w1155_
	);
	LUT4 #(
		.INIT('h02a0)
	) name907 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1156_
	);
	LUT4 #(
		.INIT('h0401)
	) name908 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1157_
	);
	LUT2 #(
		.INIT('h8)
	) name909 (
		_w599_,
		_w584_,
		_w1158_
	);
	LUT4 #(
		.INIT('hcf77)
	) name910 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1159_
	);
	LUT4 #(
		.INIT('h0032)
	) name911 (
		_w615_,
		_w1157_,
		_w1159_,
		_w1156_,
		_w1160_
	);
	LUT4 #(
		.INIT('hefeb)
	) name912 (
		_w599_,
		_w584_,
		_w596_,
		_w581_,
		_w1161_
	);
	LUT2 #(
		.INIT('h2)
	) name913 (
		_w587_,
		_w1161_,
		_w1162_
	);
	LUT3 #(
		.INIT('h0d)
	) name914 (
		_w581_,
		_w1160_,
		_w1162_,
		_w1163_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name915 (
		\data_i[26]_pad ,
		load_i_pad,
		\rd1_L_o_reg[12]/NET0131 ,
		_w250_,
		_w1164_
	);
	LUT3 #(
		.INIT('hb4)
	) name916 (
		_w1155_,
		_w1163_,
		_w1164_,
		_w1165_
	);
	LUT4 #(
		.INIT('h76fc)
	) name917 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1166_
	);
	LUT4 #(
		.INIT('h8020)
	) name918 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1167_
	);
	LUT4 #(
		.INIT('hfdc3)
	) name919 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1168_
	);
	LUT4 #(
		.INIT('h3120)
	) name920 (
		_w1068_,
		_w1167_,
		_w1168_,
		_w1166_,
		_w1169_
	);
	LUT4 #(
		.INIT('h1221)
	) name921 (
		_w1067_,
		_w1068_,
		_w1070_,
		_w1078_,
		_w1170_
	);
	LUT3 #(
		.INIT('h40)
	) name922 (
		_w1070_,
		_w1077_,
		_w1078_,
		_w1171_
	);
	LUT4 #(
		.INIT('h2000)
	) name923 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1172_
	);
	LUT4 #(
		.INIT('h0802)
	) name924 (
		_w1068_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1173_
	);
	LUT3 #(
		.INIT('h01)
	) name925 (
		_w1172_,
		_w1173_,
		_w1170_,
		_w1174_
	);
	LUT4 #(
		.INIT('h0040)
	) name926 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1175_
	);
	LUT3 #(
		.INIT('h40)
	) name927 (
		_w1067_,
		_w1068_,
		_w1078_,
		_w1176_
	);
	LUT3 #(
		.INIT('h13)
	) name928 (
		_w1089_,
		_w1175_,
		_w1176_,
		_w1177_
	);
	LUT4 #(
		.INIT('he400)
	) name929 (
		_w1086_,
		_w1169_,
		_w1174_,
		_w1177_,
		_w1178_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name930 (
		\data_i[60]_pad ,
		load_i_pad,
		\rd1_L_o_reg[16]/NET0131 ,
		_w250_,
		_w1179_
	);
	LUT2 #(
		.INIT('h9)
	) name931 (
		_w1178_,
		_w1179_,
		_w1180_
	);
	LUT4 #(
		.INIT('h0660)
	) name932 (
		_w306_,
		_w369_,
		_w508_,
		_w510_,
		_w1181_
	);
	LUT3 #(
		.INIT('hf2)
	) name933 (
		_w512_,
		_w520_,
		_w522_,
		_w1182_
	);
	LUT4 #(
		.INIT('h80cc)
	) name934 (
		_w520_,
		_w532_,
		_w533_,
		_w541_,
		_w1183_
	);
	LUT3 #(
		.INIT('h10)
	) name935 (
		_w520_,
		_w532_,
		_w533_,
		_w1184_
	);
	LUT4 #(
		.INIT('h6f0f)
	) name936 (
		_w306_,
		_w369_,
		_w520_,
		_w532_,
		_w1185_
	);
	LUT3 #(
		.INIT('h60)
	) name937 (
		_w508_,
		_w510_,
		_w541_,
		_w1186_
	);
	LUT3 #(
		.INIT('h8a)
	) name938 (
		_w555_,
		_w1185_,
		_w1186_,
		_w1187_
	);
	LUT4 #(
		.INIT('h4500)
	) name939 (
		_w1184_,
		_w1182_,
		_w1183_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w520_,
		_w541_,
		_w1189_
	);
	LUT3 #(
		.INIT('he0)
	) name941 (
		_w537_,
		_w539_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		_w532_,
		_w541_,
		_w1191_
	);
	LUT3 #(
		.INIT('h15)
	) name943 (
		_w555_,
		_w1181_,
		_w1191_,
		_w1192_
	);
	LUT3 #(
		.INIT('h20)
	) name944 (
		_w535_,
		_w1190_,
		_w1192_,
		_w1193_
	);
	LUT3 #(
		.INIT('h20)
	) name945 (
		_w521_,
		_w522_,
		_w532_,
		_w1194_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name946 (
		_w512_,
		_w520_,
		_w522_,
		_w532_,
		_w1195_
	);
	LUT3 #(
		.INIT('h70)
	) name947 (
		_w512_,
		_w536_,
		_w541_,
		_w1196_
	);
	LUT4 #(
		.INIT('h007b)
	) name948 (
		_w512_,
		_w522_,
		_w532_,
		_w541_,
		_w1197_
	);
	LUT3 #(
		.INIT('h10)
	) name949 (
		_w512_,
		_w532_,
		_w543_,
		_w1198_
	);
	LUT4 #(
		.INIT('h00f8)
	) name950 (
		_w1195_,
		_w1196_,
		_w1197_,
		_w1198_,
		_w1199_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name951 (
		\data_i[52]_pad ,
		load_i_pad,
		\rd1_L_o_reg[17]/NET0131 ,
		_w250_,
		_w1200_
	);
	LUT4 #(
		.INIT('he01f)
	) name952 (
		_w1188_,
		_w1193_,
		_w1199_,
		_w1200_,
		_w1201_
	);
	LUT4 #(
		.INIT('h0f06)
	) name953 (
		_w330_,
		_w460_,
		_w823_,
		_w832_,
		_w1202_
	);
	LUT3 #(
		.INIT('h8a)
	) name954 (
		_w822_,
		_w840_,
		_w1202_,
		_w1203_
	);
	LUT4 #(
		.INIT('h0123)
	) name955 (
		_w827_,
		_w852_,
		_w840_,
		_w836_,
		_w1204_
	);
	LUT2 #(
		.INIT('h4)
	) name956 (
		_w822_,
		_w823_,
		_w1205_
	);
	LUT3 #(
		.INIT('h0b)
	) name957 (
		_w832_,
		_w848_,
		_w1205_,
		_w1206_
	);
	LUT4 #(
		.INIT('h0f09)
	) name958 (
		_w330_,
		_w460_,
		_w822_,
		_w832_,
		_w1207_
	);
	LUT4 #(
		.INIT('h0069)
	) name959 (
		_w330_,
		_w460_,
		_w824_,
		_w827_,
		_w1208_
	);
	LUT3 #(
		.INIT('h0e)
	) name960 (
		_w823_,
		_w1207_,
		_w1208_,
		_w1209_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name961 (
		_w1203_,
		_w1204_,
		_w1206_,
		_w1209_,
		_w1210_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		_w823_,
		_w832_,
		_w1211_
	);
	LUT4 #(
		.INIT('h0040)
	) name963 (
		_w823_,
		_w824_,
		_w827_,
		_w832_,
		_w1212_
	);
	LUT3 #(
		.INIT('h07)
	) name964 (
		_w835_,
		_w1211_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h4)
	) name965 (
		_w880_,
		_w1213_,
		_w1214_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name966 (
		\data_i[28]_pad ,
		load_i_pad,
		\rd1_L_o_reg[20]/NET0131 ,
		_w250_,
		_w1215_
	);
	LUT3 #(
		.INIT('h4b)
	) name967 (
		_w1210_,
		_w1214_,
		_w1215_,
		_w1216_
	);
	LUT3 #(
		.INIT('h10)
	) name968 (
		_w917_,
		_w898_,
		_w924_,
		_w1217_
	);
	LUT4 #(
		.INIT('h004c)
	) name969 (
		_w900_,
		_w888_,
		_w985_,
		_w972_,
		_w1218_
	);
	LUT3 #(
		.INIT('ha8)
	) name970 (
		_w887_,
		_w1217_,
		_w1218_,
		_w1219_
	);
	LUT4 #(
		.INIT('h9000)
	) name971 (
		_w491_,
		_w501_,
		_w900_,
		_w895_,
		_w1220_
	);
	LUT3 #(
		.INIT('h32)
	) name972 (
		_w902_,
		_w888_,
		_w1220_,
		_w1221_
	);
	LUT3 #(
		.INIT('h07)
	) name973 (
		_w889_,
		_w902_,
		_w887_,
		_w1222_
	);
	LUT4 #(
		.INIT('h9ff0)
	) name974 (
		_w491_,
		_w501_,
		_w900_,
		_w888_,
		_w1223_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name975 (
		_w895_,
		_w888_,
		_w899_,
		_w1223_,
		_w1224_
	);
	LUT3 #(
		.INIT('h40)
	) name976 (
		_w1221_,
		_w1222_,
		_w1224_,
		_w1225_
	);
	LUT4 #(
		.INIT('h55df)
	) name977 (
		_w889_,
		_w896_,
		_w923_,
		_w984_,
		_w1226_
	);
	LUT2 #(
		.INIT('h4)
	) name978 (
		_w900_,
		_w888_,
		_w1227_
	);
	LUT3 #(
		.INIT('h10)
	) name979 (
		_w922_,
		_w971_,
		_w1227_,
		_w1228_
	);
	LUT3 #(
		.INIT('h0e)
	) name980 (
		_w888_,
		_w1226_,
		_w1228_,
		_w1229_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name981 (
		\data_i[4]_pad ,
		load_i_pad,
		\rd1_L_o_reg[23]/NET0131 ,
		_w250_,
		_w1230_
	);
	LUT4 #(
		.INIT('he01f)
	) name982 (
		_w1219_,
		_w1225_,
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT4 #(
		.INIT('h1020)
	) name983 (
		_w342_,
		_w936_,
		_w932_,
		_w933_,
		_w1232_
	);
	LUT4 #(
		.INIT('h5554)
	) name984 (
		_w944_,
		_w950_,
		_w958_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w935_,
		_w1131_,
		_w1234_
	);
	LUT3 #(
		.INIT('h20)
	) name986 (
		_w932_,
		_w937_,
		_w944_,
		_w1235_
	);
	LUT4 #(
		.INIT('h083f)
	) name987 (
		_w936_,
		_w935_,
		_w959_,
		_w1235_,
		_w1236_
	);
	LUT4 #(
		.INIT('h5455)
	) name988 (
		_w952_,
		_w1233_,
		_w1234_,
		_w1236_,
		_w1237_
	);
	LUT4 #(
		.INIT('hfd31)
	) name989 (
		_w941_,
		_w935_,
		_w946_,
		_w1131_,
		_w1238_
	);
	LUT2 #(
		.INIT('h4)
	) name990 (
		_w935_,
		_w950_,
		_w1239_
	);
	LUT4 #(
		.INIT('h5504)
	) name991 (
		_w944_,
		_w952_,
		_w1238_,
		_w1239_,
		_w1240_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		_w932_,
		_w937_,
		_w1241_
	);
	LUT3 #(
		.INIT('ha8)
	) name993 (
		_w944_,
		_w1123_,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		_w935_,
		_w1132_,
		_w1243_
	);
	LUT3 #(
		.INIT('h80)
	) name995 (
		_w936_,
		_w932_,
		_w937_,
		_w1244_
	);
	LUT4 #(
		.INIT('hc840)
	) name996 (
		_w935_,
		_w944_,
		_w946_,
		_w1244_,
		_w1245_
	);
	LUT4 #(
		.INIT('h0057)
	) name997 (
		_w952_,
		_w1242_,
		_w1243_,
		_w1245_,
		_w1246_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name998 (
		\data_i[30]_pad ,
		load_i_pad,
		\rd1_L_o_reg[28]/NET0131 ,
		_w250_,
		_w1247_
	);
	LUT4 #(
		.INIT('h10ef)
	) name999 (
		_w1240_,
		_w1237_,
		_w1246_,
		_w1247_,
		_w1248_
	);
	LUT3 #(
		.INIT('h54)
	) name1000 (
		_w888_,
		_w903_,
		_w986_,
		_w1249_
	);
	LUT4 #(
		.INIT('hb1f5)
	) name1001 (
		_w889_,
		_w897_,
		_w912_,
		_w888_,
		_w1250_
	);
	LUT3 #(
		.INIT('h45)
	) name1002 (
		_w887_,
		_w1249_,
		_w1250_,
		_w1251_
	);
	LUT4 #(
		.INIT('hf600)
	) name1003 (
		_w491_,
		_w501_,
		_w895_,
		_w888_,
		_w1252_
	);
	LUT3 #(
		.INIT('he0)
	) name1004 (
		_w889_,
		_w903_,
		_w1252_,
		_w1253_
	);
	LUT4 #(
		.INIT('h5d5f)
	) name1005 (
		_w900_,
		_w895_,
		_w985_,
		_w991_,
		_w1254_
	);
	LUT3 #(
		.INIT('h8a)
	) name1006 (
		_w887_,
		_w1253_,
		_w1254_,
		_w1255_
	);
	LUT4 #(
		.INIT('h9000)
	) name1007 (
		_w900_,
		_w895_,
		_w896_,
		_w887_,
		_w1256_
	);
	LUT4 #(
		.INIT('h3320)
	) name1008 (
		_w889_,
		_w888_,
		_w918_,
		_w1256_,
		_w1257_
	);
	LUT3 #(
		.INIT('hc8)
	) name1009 (
		_w902_,
		_w888_,
		_w989_,
		_w1258_
	);
	LUT4 #(
		.INIT('h6660)
	) name1010 (
		_w491_,
		_w501_,
		_w895_,
		_w896_,
		_w1259_
	);
	LUT3 #(
		.INIT('h04)
	) name1011 (
		_w991_,
		_w1227_,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('h0001)
	) name1012 (
		_w927_,
		_w1257_,
		_w1258_,
		_w1260_,
		_w1261_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1013 (
		\data_i[2]_pad ,
		load_i_pad,
		\rd1_L_o_reg[15]/NET0131 ,
		_w250_,
		_w1262_
	);
	LUT4 #(
		.INIT('h10ef)
	) name1014 (
		_w1255_,
		_w1251_,
		_w1261_,
		_w1262_,
		_w1263_
	);
	LUT4 #(
		.INIT('hf35a)
	) name1015 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1264_
	);
	LUT4 #(
		.INIT('ha400)
	) name1016 (
		_w753_,
		_w745_,
		_w737_,
		_w766_,
		_w1265_
	);
	LUT4 #(
		.INIT('h8400)
	) name1017 (
		_w753_,
		_w745_,
		_w737_,
		_w766_,
		_w1266_
	);
	LUT4 #(
		.INIT('h0032)
	) name1018 (
		_w766_,
		_w771_,
		_w1264_,
		_w1266_,
		_w1267_
	);
	LUT2 #(
		.INIT('h2)
	) name1019 (
		_w736_,
		_w1267_,
		_w1268_
	);
	LUT4 #(
		.INIT('h4a85)
	) name1020 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1269_
	);
	LUT2 #(
		.INIT('h2)
	) name1021 (
		_w766_,
		_w1269_,
		_w1270_
	);
	LUT3 #(
		.INIT('h10)
	) name1022 (
		_w753_,
		_w738_,
		_w737_,
		_w1271_
	);
	LUT4 #(
		.INIT('h2eff)
	) name1023 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1272_
	);
	LUT3 #(
		.INIT('h15)
	) name1024 (
		_w736_,
		_w1111_,
		_w1272_,
		_w1273_
	);
	LUT4 #(
		.INIT('h0020)
	) name1025 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1274_
	);
	LUT4 #(
		.INIT('hafdf)
	) name1026 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1275_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		_w766_,
		_w1275_,
		_w1276_
	);
	LUT3 #(
		.INIT('h23)
	) name1028 (
		_w738_,
		_w1105_,
		_w1265_,
		_w1277_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1029 (
		_w1270_,
		_w1273_,
		_w1276_,
		_w1277_,
		_w1278_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1030 (
		\data_i[24]_pad ,
		load_i_pad,
		\rd1_L_o_reg[4]/NET0131 ,
		_w250_,
		_w1279_
	);
	LUT3 #(
		.INIT('h4b)
	) name1031 (
		_w1268_,
		_w1278_,
		_w1279_,
		_w1280_
	);
	LUT2 #(
		.INIT('h4)
	) name1032 (
		_w700_,
		_w705_,
		_w1281_
	);
	LUT2 #(
		.INIT('h1)
	) name1033 (
		_w687_,
		_w668_,
		_w1282_
	);
	LUT4 #(
		.INIT('h1101)
	) name1034 (
		_w698_,
		_w1005_,
		_w1043_,
		_w1282_,
		_w1283_
	);
	LUT4 #(
		.INIT('hfd31)
	) name1035 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1284_
	);
	LUT2 #(
		.INIT('h2)
	) name1036 (
		_w687_,
		_w1284_,
		_w1285_
	);
	LUT4 #(
		.INIT('h1000)
	) name1037 (
		_w687_,
		_w665_,
		_w666_,
		_w676_,
		_w1286_
	);
	LUT4 #(
		.INIT('hf700)
	) name1038 (
		_w665_,
		_w666_,
		_w676_,
		_w698_,
		_w1287_
	);
	LUT3 #(
		.INIT('h10)
	) name1039 (
		_w1041_,
		_w1286_,
		_w1287_,
		_w1288_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1040 (
		_w1281_,
		_w1283_,
		_w1285_,
		_w1288_,
		_w1289_
	);
	LUT4 #(
		.INIT('hfbfe)
	) name1041 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1290_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		_w687_,
		_w1290_,
		_w1291_
	);
	LUT4 #(
		.INIT('hfd3d)
	) name1043 (
		_w665_,
		_w666_,
		_w668_,
		_w676_,
		_w1292_
	);
	LUT2 #(
		.INIT('h1)
	) name1044 (
		_w687_,
		_w698_,
		_w1293_
	);
	LUT2 #(
		.INIT('h4)
	) name1045 (
		_w1292_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h9)
	) name1046 (
		_w665_,
		_w666_,
		_w1295_
	);
	LUT2 #(
		.INIT('h8)
	) name1047 (
		_w705_,
		_w1295_,
		_w1296_
	);
	LUT3 #(
		.INIT('h07)
	) name1048 (
		_w709_,
		_w1001_,
		_w1009_,
		_w1297_
	);
	LUT4 #(
		.INIT('h0100)
	) name1049 (
		_w1291_,
		_w1296_,
		_w1294_,
		_w1297_,
		_w1298_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1050 (
		\data_i[0]_pad ,
		load_i_pad,
		\rd1_L_o_reg[7]/NET0131 ,
		_w250_,
		_w1299_
	);
	LUT3 #(
		.INIT('h4b)
	) name1051 (
		_w1289_,
		_w1298_,
		_w1299_,
		_w1300_
	);
	LUT3 #(
		.INIT('h96)
	) name1052 (
		_w1070_,
		_w1077_,
		_w1078_,
		_w1301_
	);
	LUT4 #(
		.INIT('hfddf)
	) name1053 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1302_
	);
	LUT4 #(
		.INIT('had00)
	) name1054 (
		_w1086_,
		_w1084_,
		_w1301_,
		_w1302_,
		_w1303_
	);
	LUT4 #(
		.INIT('h47bb)
	) name1055 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1304_
	);
	LUT4 #(
		.INIT('h0002)
	) name1056 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1305_
	);
	LUT4 #(
		.INIT('h3302)
	) name1057 (
		_w1068_,
		_w1086_,
		_w1304_,
		_w1305_,
		_w1306_
	);
	LUT4 #(
		.INIT('h0990)
	) name1058 (
		_w411_,
		_w585_,
		_w1067_,
		_w1078_,
		_w1307_
	);
	LUT3 #(
		.INIT('h23)
	) name1059 (
		_w1171_,
		_w1172_,
		_w1307_,
		_w1308_
	);
	LUT4 #(
		.INIT('h0e04)
	) name1060 (
		_w1068_,
		_w1303_,
		_w1306_,
		_w1308_,
		_w1309_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1061 (
		\data_i[46]_pad ,
		load_i_pad,
		\rd1_L_o_reg[26]/NET0131 ,
		_w250_,
		_w1310_
	);
	LUT2 #(
		.INIT('h9)
	) name1062 (
		_w1309_,
		_w1310_,
		_w1311_
	);
	LUT4 #(
		.INIT('h9dbc)
	) name1063 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1312_
	);
	LUT4 #(
		.INIT('h0800)
	) name1064 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1313_
	);
	LUT4 #(
		.INIT('h72c2)
	) name1065 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1314_
	);
	LUT4 #(
		.INIT('h3120)
	) name1066 (
		_w1068_,
		_w1313_,
		_w1314_,
		_w1312_,
		_w1315_
	);
	LUT2 #(
		.INIT('h2)
	) name1067 (
		_w1086_,
		_w1315_,
		_w1316_
	);
	LUT3 #(
		.INIT('h60)
	) name1068 (
		_w411_,
		_w585_,
		_w1067_,
		_w1317_
	);
	LUT3 #(
		.INIT('h10)
	) name1069 (
		_w1089_,
		_w1090_,
		_w1317_,
		_w1318_
	);
	LUT4 #(
		.INIT('h0c15)
	) name1070 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1319_
	);
	LUT2 #(
		.INIT('h2)
	) name1071 (
		_w1068_,
		_w1319_,
		_w1320_
	);
	LUT4 #(
		.INIT('h5ac7)
	) name1072 (
		_w1067_,
		_w1070_,
		_w1077_,
		_w1078_,
		_w1321_
	);
	LUT4 #(
		.INIT('h0504)
	) name1073 (
		_w1068_,
		_w1086_,
		_w1175_,
		_w1321_,
		_w1322_
	);
	LUT3 #(
		.INIT('h0b)
	) name1074 (
		_w1318_,
		_w1320_,
		_w1322_,
		_w1323_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1075 (
		\data_i[40]_pad ,
		load_i_pad,
		\rd1_L_o_reg[2]/NET0131 ,
		_w250_,
		_w1324_
	);
	LUT3 #(
		.INIT('h1e)
	) name1076 (
		_w1316_,
		_w1323_,
		_w1324_,
		_w1325_
	);
	LUT4 #(
		.INIT('h53fc)
	) name1077 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1326_
	);
	LUT3 #(
		.INIT('h10)
	) name1078 (
		_w766_,
		_w774_,
		_w1326_,
		_w1327_
	);
	LUT3 #(
		.INIT('h02)
	) name1079 (
		_w766_,
		_w770_,
		_w1271_,
		_w1328_
	);
	LUT4 #(
		.INIT('h0002)
	) name1080 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1329_
	);
	LUT4 #(
		.INIT('h8850)
	) name1081 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1330_
	);
	LUT3 #(
		.INIT('h02)
	) name1082 (
		_w736_,
		_w1330_,
		_w1329_,
		_w1331_
	);
	LUT3 #(
		.INIT('he0)
	) name1083 (
		_w1327_,
		_w1328_,
		_w1331_,
		_w1332_
	);
	LUT4 #(
		.INIT('ha0ac)
	) name1084 (
		_w753_,
		_w738_,
		_w745_,
		_w737_,
		_w1333_
	);
	LUT3 #(
		.INIT('h6e)
	) name1085 (
		_w738_,
		_w745_,
		_w737_,
		_w1334_
	);
	LUT4 #(
		.INIT('he4f5)
	) name1086 (
		_w766_,
		_w774_,
		_w1333_,
		_w1334_,
		_w1335_
	);
	LUT3 #(
		.INIT('h01)
	) name1087 (
		_w736_,
		_w779_,
		_w1274_,
		_w1336_
	);
	LUT2 #(
		.INIT('h4)
	) name1088 (
		_w1335_,
		_w1336_,
		_w1337_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1089 (
		\data_i[10]_pad ,
		load_i_pad,
		\rd1_L_o_reg[14]/NET0131 ,
		_w250_,
		_w1338_
	);
	LUT3 #(
		.INIT('he1)
	) name1090 (
		_w1332_,
		_w1337_,
		_w1338_,
		_w1339_
	);
	LUT4 #(
		.INIT('h6100)
	) name1091 (
		_w599_,
		_w587_,
		_w596_,
		_w581_,
		_w1340_
	);
	LUT4 #(
		.INIT('h0220)
	) name1092 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1341_
	);
	LUT4 #(
		.INIT('h7fc7)
	) name1093 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1342_
	);
	LUT4 #(
		.INIT('h0032)
	) name1094 (
		_w581_,
		_w1341_,
		_w1342_,
		_w1340_,
		_w1343_
	);
	LUT2 #(
		.INIT('h1)
	) name1095 (
		_w615_,
		_w1343_,
		_w1344_
	);
	LUT4 #(
		.INIT('ha3f8)
	) name1096 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1345_
	);
	LUT4 #(
		.INIT('h0302)
	) name1097 (
		_w581_,
		_w808_,
		_w809_,
		_w1345_,
		_w1346_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1098 (
		_w581_,
		_w794_,
		_w795_,
		_w1158_,
		_w1347_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1099 (
		_w599_,
		_w584_,
		_w587_,
		_w596_,
		_w1348_
	);
	LUT2 #(
		.INIT('h2)
	) name1100 (
		_w797_,
		_w1348_,
		_w1349_
	);
	LUT4 #(
		.INIT('h000d)
	) name1101 (
		_w615_,
		_w1346_,
		_w1347_,
		_w1349_,
		_w1350_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1102 (
		\data_i[6]_pad ,
		load_i_pad,
		\rd1_L_o_reg[31]/NET0131 ,
		_w250_,
		_w1351_
	);
	LUT3 #(
		.INIT('hb4)
	) name1103 (
		_w1344_,
		_w1350_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h8)
	) name1104 (
		_w541_,
		_w555_,
		_w1353_
	);
	LUT4 #(
		.INIT('hff96)
	) name1105 (
		_w306_,
		_w369_,
		_w520_,
		_w532_,
		_w1354_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		_w555_,
		_w1354_,
		_w1355_
	);
	LUT4 #(
		.INIT('h007b)
	) name1107 (
		_w512_,
		_w520_,
		_w522_,
		_w566_,
		_w1356_
	);
	LUT4 #(
		.INIT('h3032)
	) name1108 (
		_w541_,
		_w1353_,
		_w1355_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		_w512_,
		_w566_,
		_w1358_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1110 (
		_w520_,
		_w522_,
		_w537_,
		_w541_,
		_w1359_
	);
	LUT4 #(
		.INIT('hc480)
	) name1111 (
		_w512_,
		_w532_,
		_w536_,
		_w543_,
		_w1360_
	);
	LUT3 #(
		.INIT('h07)
	) name1112 (
		_w520_,
		_w533_,
		_w541_,
		_w1361_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1113 (
		_w1358_,
		_w1359_,
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT4 #(
		.INIT('he4be)
	) name1114 (
		_w512_,
		_w520_,
		_w522_,
		_w532_,
		_w1363_
	);
	LUT2 #(
		.INIT('h4)
	) name1115 (
		_w1363_,
		_w1353_,
		_w1364_
	);
	LUT4 #(
		.INIT('hbeb4)
	) name1116 (
		_w512_,
		_w520_,
		_w522_,
		_w532_,
		_w1365_
	);
	LUT2 #(
		.INIT('h1)
	) name1117 (
		_w541_,
		_w555_,
		_w1366_
	);
	LUT4 #(
		.INIT('h0080)
	) name1118 (
		_w520_,
		_w522_,
		_w537_,
		_w555_,
		_w1367_
	);
	LUT4 #(
		.INIT('h1011)
	) name1119 (
		_w1194_,
		_w1367_,
		_w1365_,
		_w1366_,
		_w1368_
	);
	LUT4 #(
		.INIT('h0100)
	) name1120 (
		_w1364_,
		_w1362_,
		_w1357_,
		_w1368_,
		_w1369_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1121 (
		\data_i[34]_pad ,
		load_i_pad,
		\rd1_L_o_reg[11]/NET0131 ,
		_w250_,
		_w1370_
	);
	LUT2 #(
		.INIT('h9)
	) name1122 (
		_w1369_,
		_w1370_,
		_w1371_
	);
	LUT4 #(
		.INIT('h7d00)
	) name1123 (
		_w521_,
		_w522_,
		_w532_,
		_w541_,
		_w1372_
	);
	LUT4 #(
		.INIT('hf7bf)
	) name1124 (
		_w512_,
		_w520_,
		_w522_,
		_w532_,
		_w1373_
	);
	LUT2 #(
		.INIT('h1)
	) name1125 (
		_w541_,
		_w566_,
		_w1374_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name1126 (
		_w1194_,
		_w1372_,
		_w1373_,
		_w1374_,
		_w1375_
	);
	LUT4 #(
		.INIT('h9fd3)
	) name1127 (
		_w512_,
		_w520_,
		_w522_,
		_w532_,
		_w1376_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w541_,
		_w1376_,
		_w1377_
	);
	LUT3 #(
		.INIT('h20)
	) name1129 (
		_w512_,
		_w536_,
		_w1191_,
		_w1378_
	);
	LUT3 #(
		.INIT('h13)
	) name1130 (
		_w512_,
		_w555_,
		_w566_,
		_w1379_
	);
	LUT3 #(
		.INIT('h20)
	) name1131 (
		_w1195_,
		_w1378_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h8)
	) name1132 (
		_w520_,
		_w532_,
		_w1381_
	);
	LUT3 #(
		.INIT('h2a)
	) name1133 (
		_w555_,
		_w1181_,
		_w1381_,
		_w1382_
	);
	LUT3 #(
		.INIT('h09)
	) name1134 (
		_w508_,
		_w510_,
		_w541_,
		_w1383_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1135 (
		_w306_,
		_w369_,
		_w520_,
		_w532_,
		_w1384_
	);
	LUT4 #(
		.INIT('h0900)
	) name1136 (
		_w306_,
		_w369_,
		_w520_,
		_w532_,
		_w1385_
	);
	LUT3 #(
		.INIT('h8d)
	) name1137 (
		_w1383_,
		_w1384_,
		_w1385_,
		_w1386_
	);
	LUT3 #(
		.INIT('h40)
	) name1138 (
		_w534_,
		_w1382_,
		_w1386_,
		_w1387_
	);
	LUT4 #(
		.INIT('h5510)
	) name1139 (
		_w1375_,
		_w1377_,
		_w1380_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1140 (
		\data_i[38]_pad ,
		load_i_pad,
		\rd1_L_o_reg[27]/NET0131 ,
		_w250_,
		_w1389_
	);
	LUT2 #(
		.INIT('h6)
	) name1141 (
		_w1388_,
		_w1389_,
		_w1390_
	);
	LUT3 #(
		.INIT('he7)
	) name1142 (
		_w936_,
		_w932_,
		_w937_,
		_w1391_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w935_,
		_w1391_,
		_w1392_
	);
	LUT3 #(
		.INIT('h0e)
	) name1144 (
		_w944_,
		_w965_,
		_w1235_,
		_w1393_
	);
	LUT3 #(
		.INIT('h45)
	) name1145 (
		_w952_,
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT3 #(
		.INIT('h54)
	) name1146 (
		_w944_,
		_w1232_,
		_w1244_,
		_w1395_
	);
	LUT4 #(
		.INIT('h4100)
	) name1147 (
		_w936_,
		_w932_,
		_w937_,
		_w944_,
		_w1396_
	);
	LUT4 #(
		.INIT('h001b)
	) name1148 (
		_w935_,
		_w950_,
		_w953_,
		_w1396_,
		_w1397_
	);
	LUT3 #(
		.INIT('h8a)
	) name1149 (
		_w952_,
		_w1395_,
		_w1397_,
		_w1398_
	);
	LUT3 #(
		.INIT('h90)
	) name1150 (
		_w342_,
		_w933_,
		_w944_,
		_w1399_
	);
	LUT2 #(
		.INIT('h4)
	) name1151 (
		_w1391_,
		_w1399_,
		_w1400_
	);
	LUT3 #(
		.INIT('h69)
	) name1152 (
		_w342_,
		_w933_,
		_w944_,
		_w1401_
	);
	LUT3 #(
		.INIT('he0)
	) name1153 (
		_w940_,
		_w1138_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h1)
	) name1154 (
		_w1400_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('hb8f0)
	) name1155 (
		\data_i[18]_pad ,
		load_i_pad,
		\rd1_L_o_reg[13]/NET0131 ,
		_w250_,
		_w1404_
	);
	LUT4 #(
		.INIT('h10ef)
	) name1156 (
		_w1398_,
		_w1394_,
		_w1403_,
		_w1404_,
		_w1405_
	);
	LUT4 #(
		.INIT('h000d)
	) name1157 (
		_w263_,
		_w338_,
		_w682_,
		_w721_,
		_w1406_
	);
	LUT4 #(
		.INIT('he020)
	) name1158 (
		\rd1_Key_o_reg[14]/NET0131 ,
		_w250_,
		_w263_,
		_w451_,
		_w1407_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1159 (
		decrypt_i_pad,
		_w434_,
		_w506_,
		_w1407_,
		_w1408_
	);
	LUT3 #(
		.INIT('hf1)
	) name1160 (
		decrypt_i_pad,
		_w1406_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('h0145)
	) name1161 (
		decrypt_i_pad,
		_w256_,
		_w313_,
		_w444_,
		_w1410_
	);
	LUT4 #(
		.INIT('he020)
	) name1162 (
		\rd1_Key_o_reg[22]/NET0131 ,
		_w250_,
		_w263_,
		_w321_,
		_w1411_
	);
	LUT4 #(
		.INIT('h0031)
	) name1163 (
		_w256_,
		_w309_,
		_w316_,
		_w1411_,
		_w1412_
	);
	LUT3 #(
		.INIT('hce)
	) name1164 (
		decrypt_i_pad,
		_w1410_,
		_w1412_,
		_w1413_
	);
	LUT4 #(
		.INIT('h0e02)
	) name1165 (
		\rd1_Key_o_reg[30]/NET0131 ,
		_w250_,
		_w256_,
		_w296_,
		_w1414_
	);
	LUT3 #(
		.INIT('h54)
	) name1166 (
		decrypt_i_pad,
		_w463_,
		_w1414_,
		_w1415_
	);
	LUT4 #(
		.INIT('he020)
	) name1167 (
		\rd1_Key_o_reg[32]/NET0131 ,
		_w250_,
		_w263_,
		_w348_,
		_w1416_
	);
	LUT4 #(
		.INIT('h0031)
	) name1168 (
		_w256_,
		_w302_,
		_w356_,
		_w1416_,
		_w1417_
	);
	LUT3 #(
		.INIT('hce)
	) name1169 (
		decrypt_i_pad,
		_w1415_,
		_w1417_,
		_w1418_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1170 (
		_w250_,
		_w263_,
		_w409_,
		_w578_,
		_w1419_
	);
	LUT4 #(
		.INIT('he020)
	) name1171 (
		\rd1_Key_o_reg[48]/NET0131 ,
		_w250_,
		_w263_,
		_w400_,
		_w1420_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1172 (
		decrypt_i_pad,
		_w408_,
		_w637_,
		_w1420_,
		_w1421_
	);
	LUT3 #(
		.INIT('hf1)
	) name1173 (
		decrypt_i_pad,
		_w1419_,
		_w1421_,
		_w1422_
	);
	LUT4 #(
		.INIT('h00cd)
	) name1174 (
		_w250_,
		_w267_,
		_w263_,
		_w633_,
		_w1423_
	);
	LUT4 #(
		.INIT('h000d)
	) name1175 (
		_w263_,
		_w272_,
		_w391_,
		_w515_,
		_w1424_
	);
	LUT3 #(
		.INIT('h1b)
	) name1176 (
		decrypt_i_pad,
		_w1423_,
		_w1424_,
		_w1425_
	);
	LUT4 #(
		.INIT('h0e02)
	) name1177 (
		\rd1_Key_o_reg[37]/NET0131 ,
		_w250_,
		_w256_,
		_w417_,
		_w1426_
	);
	LUT4 #(
		.INIT('he020)
	) name1178 (
		\rd1_Key_o_reg[36]/NET0131 ,
		_w250_,
		_w256_,
		_w420_,
		_w1427_
	);
	LUT3 #(
		.INIT('h54)
	) name1179 (
		decrypt_i_pad,
		_w1426_,
		_w1427_,
		_w1428_
	);
	LUT4 #(
		.INIT('he020)
	) name1180 (
		\rd1_Key_o_reg[39]/NET0131 ,
		_w250_,
		_w263_,
		_w485_,
		_w1429_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1181 (
		decrypt_i_pad,
		_w784_,
		_w890_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('he)
	) name1182 (
		_w1428_,
		_w1430_,
		_w1431_
	);
	LUT4 #(
		.INIT('h0031)
	) name1183 (
		_w263_,
		_w350_,
		_w356_,
		_w374_,
		_w1432_
	);
	LUT4 #(
		.INIT('he020)
	) name1184 (
		\rd1_Key_o_reg[35]/NET0131 ,
		_w250_,
		_w263_,
		_w375_,
		_w1433_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1185 (
		decrypt_i_pad,
		_w358_,
		_w1427_,
		_w1433_,
		_w1434_
	);
	LUT3 #(
		.INIT('hf1)
	) name1186 (
		decrypt_i_pad,
		_w1432_,
		_w1434_,
		_w1435_
	);
	LUT4 #(
		.INIT('h0e02)
	) name1187 (
		\rd1_Key_o_reg[17]/NET0131 ,
		_w250_,
		_w256_,
		_w442_,
		_w1436_
	);
	LUT3 #(
		.INIT('h54)
	) name1188 (
		decrypt_i_pad,
		_w504_,
		_w1436_,
		_w1437_
	);
	LUT4 #(
		.INIT('h0031)
	) name1189 (
		_w263_,
		_w314_,
		_w444_,
		_w440_,
		_w1438_
	);
	LUT3 #(
		.INIT('hce)
	) name1190 (
		decrypt_i_pad,
		_w1437_,
		_w1438_,
		_w1439_
	);
	LUT3 #(
		.INIT('h13)
	) name1191 (
		\data_ready_reg/NET0131 ,
		load_i_pad,
		\stage1_iter_reg[0]/NET0131 ,
		_w1440_
	);
	LUT4 #(
		.INIT('h5554)
	) name1192 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[1]/NET0131 ,
		\stage1_iter_reg[2]/NET0131 ,
		\stage1_iter_reg[3]/NET0131 ,
		_w1441_
	);
	LUT3 #(
		.INIT('hf2)
	) name1193 (
		_w250_,
		_w1440_,
		_w1441_,
		_w1442_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1194 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[1]/NET0131 ,
		\stage1_iter_reg[2]/NET0131 ,
		\stage1_iter_reg[3]/NET0131 ,
		_w1443_
	);
	LUT3 #(
		.INIT('h78)
	) name1195 (
		\stage1_iter_reg[0]/NET0131 ,
		\stage1_iter_reg[1]/NET0131 ,
		\stage1_iter_reg[2]/NET0131 ,
		_w1444_
	);
	LUT3 #(
		.INIT('h3a)
	) name1196 (
		\data_ready_reg/NET0131 ,
		load_i_pad,
		_w250_,
		_w1445_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g10087/_0_  = _w252_ ;
	assign \g10220/_1_  = _w253_ ;
	assign \g11117/_0_  = _w269_ ;
	assign \g11124/_0_  = _w271_ ;
	assign \g11125/_0_  = _w287_ ;
	assign \g11170/_0_  = _w305_ ;
	assign \g11182/_0_  = _w307_ ;
	assign \g11184/_0_  = _w324_ ;
	assign \g11378/_0_  = _w331_ ;
	assign \g11393/_0_  = _w343_ ;
	assign \g11415/_0_  = _w352_ ;
	assign \g11432/_0_  = _w362_ ;
	assign \g11433/_0_  = _w364_ ;
	assign \g11453/_0_  = _w370_ ;
	assign \g11500/_0_  = _w379_ ;
	assign \g11588/_0_  = _w386_ ;
	assign \g11607/_0_  = _w396_ ;
	assign \g11616/_0_  = _w412_ ;
	assign \g11625/_0_  = _w414_ ;
	assign \g11641_dup/_0_  = _w424_ ;
	assign \g11648/_0_  = _w432_ ;
	assign \g11655/_0_  = _w446_ ;
	assign \g11683/_0_  = _w448_ ;
	assign \g11689/_2_  = _w450_ ;
	assign \g11694/_0_  = _w459_ ;
	assign \g11748/_0_  = _w461_ ;
	assign \g11880/_0_  = _w471_ ;
	assign \g11962/_1_  = _w482_ ;
	assign \g12016/_0_  = _w490_ ;
	assign \g12038/_0_  = _w492_ ;
	assign \g12039/_0_  = _w502_ ;
	assign \g12094/_0_  = _w570_ ;
	assign \g12100/_0_  = _w509_ ;
	assign \g12132/_0_  = _w629_ ;
	assign \g12151/_0_  = _w635_ ;
	assign \g12251/_0_  = _w641_ ;
	assign \g12279/_0_  = _w646_ ;
	assign \g12288/_0_  = _w614_ ;
	assign \g12290/_0_  = _w652_ ;
	assign \g12311/_0_  = _w654_ ;
	assign \g12313/_0_  = _w658_ ;
	assign \g12356/_0_  = _w662_ ;
	assign \g12357/_0_  = _w664_ ;
	assign \g12427/_0_  = _w715_ ;
	assign \g12441/_0_  = _w717_ ;
	assign \g12442/_0_  = _w724_ ;
	assign \g12480/_0_  = _w684_ ;
	assign \g12485/_0_  = _w686_ ;
	assign \g12506/_0_  = _w598_ ;
	assign \g12544/_0_  = _w729_ ;
	assign \g12549/_2_  = _w733_ ;
	assign \g12614/_0_  = _w783_ ;
	assign \g12678/_0_  = _w675_ ;
	assign \g12680/_0_  = _w673_ ;
	assign \g12748/_0_  = _w789_ ;
	assign \g15/_0_  = _w793_ ;
	assign \g25/_0_  = _w763_ ;
	assign \g31/_0_  = _w817_ ;
	assign \g6843/_0_  = _w865_ ;
	assign \g6861/_0_  = _w886_ ;
	assign \g6863/_0_  = _w931_ ;
	assign \g6865/_0_  = _w970_ ;
	assign \g6887/_0_  = _w1000_ ;
	assign \g6888/_0_  = _w1019_ ;
	assign \g6889/_0_  = _w1040_ ;
	assign \g6890/_0_  = _w1059_ ;
	assign \g6891/_0_  = _w1103_ ;
	assign \g6892/_0_  = _w1122_ ;
	assign \g6893/_0_  = _w1145_ ;
	assign \g6894/_0_  = _w1165_ ;
	assign \g6922/_0_  = _w1180_ ;
	assign \g6923/_0_  = _w1201_ ;
	assign \g6924/_3_  = _w1216_ ;
	assign \g6926/_0_  = _w1231_ ;
	assign \g6927/_0_  = _w1248_ ;
	assign \g6928/_0_  = _w1263_ ;
	assign \g6931/_0_  = _w1280_ ;
	assign \g6933/_0_  = _w1300_ ;
	assign \g6967/_0_  = _w1311_ ;
	assign \g6968/_0_  = _w1325_ ;
	assign \g6969/_0_  = _w1339_ ;
	assign \g6974/_0_  = _w1352_ ;
	assign \g6975/_0_  = _w1371_ ;
	assign \g6976/_3_  = _w1390_ ;
	assign \g7006/_3_  = _w1405_ ;
	assign \g8882/_0_  = _w1064_ ;
	assign \g8883/_0_  = _w1409_ ;
	assign \g8884/_0_  = _w1413_ ;
	assign \g8895/_0_  = _w552_ ;
	assign \g8896/_0_  = _w1418_ ;
	assign \g8898/_0_  = _w517_ ;
	assign \g8900/_2_  = _w612_ ;
	assign \g8902/_0_  = _w1422_ ;
	assign \g8907/_0_  = _w742_ ;
	assign \g8911/_0_  = _w1425_ ;
	assign \g8924/_0_  = _w1431_ ;
	assign \g8927/_0_  = _w894_ ;
	assign \g8929/_2_  = _w821_ ;
	assign \g8967/_0_  = _w580_ ;
	assign \g8969/_0_  = _w1074_ ;
	assign \g8973/_2_  = _w529_ ;
	assign \g8987/_0_  = _w750_ ;
	assign \g8989/_0_  = _w1435_ ;
	assign \g8991/_0_  = _w593_ ;
	assign \g8996/_0_  = _w1439_ ;
	assign \g9099/_0_  = _w1442_ ;
	assign \g9543/_1_  = _w1443_ ;
	assign \g9751/_1_  = _w1444_ ;
	assign \g9755/_0_  = _w1445_ ;
	assign \g9786/_0_  = _w831_ ;
	assign \g9794/_0_  = _w595_ ;
	assign \g9817/_0_  = _w735_ ;
	assign \g9836/_0_  = _w697_ ;
	assign \g9859/_0_  = _w586_ ;
	assign \g9862/_0_  = _w531_ ;
	assign \g9867/_0_  = _w826_ ;
	assign \g9869/_0_  = _w1076_ ;
	assign \g9876/_0_  = _w765_ ;
	assign \g9887/_0_  = _w519_ ;
	assign \g9895/_0_  = _w554_ ;
	assign \g9897/_0_  = _w511_ ;
	assign \g9908/_0_  = _w752_ ;
	assign \g9910/_0_  = _w934_ ;
	assign \g9915/_0_  = _w744_ ;
	assign \g9938/_0_  = _w583_ ;
	assign \g9970/_0_  = _w1066_ ;
endmodule;